`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j+npTEkrOuoAYyMX9/wRnMYX5goQTEisG66YW+i1AlzpOzLle1lXgu4EgeH5FLw294DViS5wgySE
5m4qv4CG/g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gUZcfjlaOFMdX4kb0TbR60nJXJPsPe1GyqlMGQubcZlG9I4tJ/ZhHd1EMxwWjzpXAI7Q26CbWB5d
M0N6EdylvFtjmg1EUNKbV6Du+MfiD40m8//+pZe9DGyPJfpmuD4+Zj3hF5SrXabgZ6C1Xp1icJbQ
L5r4LZJ7J0joZtYvw4s=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m5BR7gQYyud1p/OTN3ItnmfZf+MrbBm5KEryxpppgQ4iwUC0k6E0EmeGOhQnOMR89C/Uz4vDj5vP
kR/7K+K3yLfHLs+S12FpPBZ3NyuY74QU5rOfBxCPg1sdBKjM7iwVGn/Ecb4QkpmrleGslFvuCXCG
V1QSO28mdm007Vi1l3E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B4L9p7tgqm98VIH/YFg16sVSk71xEJ5QzzMkqAXSOWwulHN1TAbp/Anvm0mHWyNUaf7zrkLBC1E3
DyXIIdN8sGBbSREiq3gWYd0NIbQUfdJZZYvs3uJPPU2+ALQYTUwHJ5s3WX/NzIzGuAAOCxw/hePs
QWaSntCuSjeJws9v8g1EGOV7yq5Osdtd8x2LUU5JN2WFDJuVRSHIv/ompQlok9q1EkqQ7S7sQz+i
a0PnTbVY7uVeCYr+SXmQ0ogUGteEgW6M1VHjoHTsYDuZz4WbwB51Vlt9WJ1soaYWFGDCJlDxH59G
F3endzqkQitpYnFk4ShPiMODHQv12VpfJYbHRg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hwYr4TS/aBHf+wunP3cLIe0CYKkGOTJ5Jld+NMc8xGN3F8TLtDkRxbVMutpF4XfSBJhLcHSU4iQL
iFpWN0M+yLVcuPEGASE+OmR037wzVwI4JbEmc01MfjDNWHEY5ss30fwhsdWHpqgsyV3rfWe51mO/
8TIpFsSC0FG+zpoqHyDwegAf/Lmf4zKpgFLLo+3OtJAc3YmnzL6aNZ5o46AbwYzVu/XN7Ak3E8lI
/q6Y4ANFXbA7iDszKKZ71HKX3ByW0rvpUTg5gri77obs5l7sIyfp4En11ig6Opv8IgX7A29qw9SP
SM2VCK7D7eVxqxbxDEPCIbcxsa+cEizeFb3ajA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fLcMKoU95J0rpQurE7HrpDJ+JK9crolX2l3JMVmKcpL0dY4KtTMeR9YZVRrUm6v6lYXi1gKv9VGR
rJoz1MY0q0spfAy5jHcnDVY24WoZRTIRmr1rwKTVmYW99Be9KcesnhPZ4WuQur2Sv45IkqlI47hK
jnLtqX84PKzW0ap4HnvRWci/sP2vA5n5UU1zybiOUtlCnJBxpHY65IfbMy3yrF80TfTrR26jC/co
4alM2f8ErqkNMnUr0tMjzecZ/pjdWFH5wg5jNvR9C2o/vcUC0kr2fnXRwsQXgxT9vAbEitKz9+8m
p1Mwc+il16beY7eojdApx4J9ojOFXIxI8G/fSg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1719712)
`protect data_block
VNYkwl0rEcKPMuF52+DMTsHR6VK3mFUVlRavY+1qMoEJd6RSiKV9iv+7wZi4qu/mtmdxWhWs69aM
tlQ+O1GubAIaI5VIDbUp99jEG13mVRFGqe/Bbtuc/vIDOwgv2SggkNsfbmbqOoKaK17awzcAh6jU
0qoJxdAzek1gXMw8FQAxKt+aD1HcpTF3wlB0jrzsc2nH4zkROYDGqroyE4zRLu8ZuQ8CqZ2G86EQ
8W4ptV1ZJbqWRuDcM+8x+0ishDPpwg03BFj78V14232FpWZB1ynMPYEFK52gjfAakIAI53D8FBig
Fc220JG1uT6DW3hxNgQuCp2RbkwB7Z+s7U9AC2/IW29diqCK6+BvopOWdJIsLUogSMw7fqqQ4IFU
ubtJ2OiQ9q0tqA5O/CQTXl2x2l3/Eeb/HwSWG5tGI+eFn8XhUgdSI4YZk4xGarJgdGThA1i3+cO8
VaB3Q4B/bBX+193Y7E0gLWwh8gKC+C5TKdY99+qAt5vjE8Tn+5DSnQzojKa5VAiuGZ4iNzfboAq6
ZpIY9OzDM55EGobnUYRxLOkNyMhaNRben9i3fJDac60dEQB1a1SJD11sFVs785zaXKCk9YBjiGLT
NxP1Nc8/VRMLgVaqTlVw+SHB8eObmp9mpz//z9kJd8FYh11lSZUz+qnM3o6ilMh/Poa/S6lVDHYz
MRZoJTimQfbxNN+/izG6zNVmrDdD8oi6QD7mF/0vIvAEoAhxh7rrxj0wvwYPD7AabaAO/URCJaZ0
4MvSY/lBNmdOWfyGXr8NCqARNMJaCJnw0RrqILSxQWZBqVZBaJRPsUFF/oFwK/QXQqskGEOgD11H
E5RswR8Iiz/3Nje4Ygv3RyTOURSiaOiAEvWlJ2xdlD1oofoKTGIDJr+gCwQdQ1hSI0m2oW3Q3+C3
wUjnPraDHCUdYuoZm+L1x2zpXClv3Tzdw0SpcdSkOpde8fQX81UrFC0osCOZ5o0vaibVIUkc/4CJ
A8iRMcUp1ImFsf2eJd8LAy0txsT0uEY4g/IOrHVh/c/rznijW7Um0UMxQwlzoEpVX/kfvT/crPoe
JNMmUXYlWgb1dw8GMW8xEyQ9nrEoM+ESDiNkx1pHjlpb9U72RX6yrFt9uYC06koYogmCrkT+GI/v
zFV8GXWHwRFQSB9pqf9F9JetP9ls+BAggKEEg41qwkNhRYgaTL4hxHpn1AaoF+f8nMhyc6/ygsV8
OSneO/JZu7zOS/PybaYejsl1I0jQvOr/bOEnW0upvG7RwMaf2FuGr2fNgX/geN7GG650etM8bmQh
OXt0ik4UFl6mUzUyOHuRI5DbBctKahNzZPjVlU3JHB9TNeUdJ/SfCWz5Xt15xbKSQfjm4YhxJqBd
ZuUfjSBLNw7j9QiEpFfi5b/d3l5yGIhbxqgjt04rhKQ1LEVGp/ghGSMzoY0yQ69kHH7UuTbuA6Ct
QpOq8EikujPIA5EcUzxFtpeKtGTunEihDckMNUK5AVv4bYcS2yemwbDeN9SRO2vuD6xsPNMa5+lE
SupunKxVDpLmB4aQpzCv4dDn0jHFGpXkp5/tZQhsTBRinDtDiaZh6LlYr1MoE/0jSx+qV7OknRVV
lEVjVoh9oaUeMAM3tJU6XHP1uuskBvUBylVLuP8yfDeEHoC8inS9d4m2hRQGCBKIEz8AgLZ29Fqx
of3PZ7CtCxOxBJ2d9z/iIo/3F2ocemaoN/61DBqJsrIG5rYk4sLRqBH8M8leKWspRn289yXhxN0k
GppzI92AZDP52wLCEJqPj/ZIi+edxsi+QVUpoRwo/mSACJRFq9LUCUdt4Kf4nf0X50ShwekXQiK+
UgitZVZY8OSDkmQ+qr5y9mIFN6YzM+vTDzNek//m8UlzE5U6Y02Lb3GY9rCH0qysgOideBhqLrui
I8mh7NFXf48ysyi+M3m8GfDsmVaowyLFT1AIhUIOyxtMhPEgjW6bClGfhSWQYHzzIyeyHFlM21gc
9WxtIZqsrb8Ps5hABaaeWvKdJLjgf8Vs4YN+wr1+GjGqJGn4TNAi3wqfORvmfuHPPBQmlwOWvDJe
JcmMsu8XlVEbpKQDD7YqgISC9Tws+ULJCkTZOeLWyRKxb4VrfbxfEntLylnXdD7NVuDJUCfUnr1k
/3JYdGfFahJSMFM59+FZ5ndT3kuvj3B6Jca0NcF5twppje67+z9A51NX7L9OBrKuaB9tHmyrNqdK
awDxV7mhI+8uLqltZaWgrbaTBpoXDNBWc7jb3tQOw3meJdpuAwnO5jFlihvZqHFN/+xOfHl8HTpP
CuxXJGWU6pfTjIJhPboWO1hdCxWKwbtvBiFu6thptZHPaB4+8gdXBrNm7JLVjA0qkPYUtSEbk5vJ
VnUoUeli0pxivkONDpbjiq3aGGvuUuf3+R3bmxYwLL9lyZtdKjlzduwJkpX1bmeYr8D5b/1APp28
yQCjH4O+XCt6ooMzf6iHRcuCQuMAESXY12oNLBp3iVFKgk6TuiildR1DmQr1Yy6FCrgOeC9R89hR
PFTyL2zGZeGbtELSZ+OauwTU9km2nC1WNHBGPw4j9Wt9QtaF5Trw1MpWxsRDHFmLg77q0vaknGQJ
0e8vomyhnwMv6P0itVs6Euxe1n5hb5knYdj+CN08d9R9rQTYGdaiHGS+Uu1+nRII7l6yJ0D1cThZ
Huo1rSN9J69sCelYx6VPOwIeneATO3WVtXYnm/adV4P/PT5QvWPHx/oTUa3qZrDeMLrBT7wQEhPK
/xkSvvNb3KUfgo4BkhQ0t2q6AIsM+SdOeY1IlQaPIZTzdwvfEaub9lw59kW7afBvc1sRYwQQhBJH
RsIywfmU4wLWczN9OL/xXFp5Gm0+72jQEJf9/3xab8mbUiKLGegksxcnqlFE1yhJOZ8yy/Tqe358
otctZUmy8rtRSbILS4pypzd1aEOf2JMjkqZfwDQPJADrCrL0Qqr2dMybn6dz+LagdDauMmkLC3CU
WwlI5vWMPxyHdJlo+g1XZWkAJNZkL2RBQHWm4GZoI9YpCcYNaMI+CNlh5MlYFthmP6lJJBtX23gz
zUJxHY4CWuWV9FQFUPD91+FRcBzQHvQWnEvNXTFm2BiiA7LPYp41UoYkEsGepD89OquNuMeu0D5+
4KhUFaRD6h1qgnhJRjpGI8ntcapsL8zfNuJ+ICjTk7RP13NwBd76Dj6ub2KAGC4TbcnCoWL9FF0l
Y0VDnioMpknUc1AgE/g4VR/+JyKuVjo6R9oYMc7hQPhOH3t+J8r3yuWyDfhSS7usxE5Ih2YSRxfy
wqBMVXunVAppcRJoNVyZpe1O7YE+MkuZE/PpXOa5IvIb4cv6R0ne1KrV86UAUwCDS7u3yPSGOrx5
Fvx66SptCn2bwodRk8tIg+GSCYrvtt07mZ/RiMqS0lN/DPA+YlB0vH2q1pOlMYf7x9iknUn6T3xh
Pd0JtLGNl/LlMmQaTKUEnJuEenGzromK3ntTJHcTdECxu6a+QcvOtoaPyW3+Hq9m5b1RY4gew/3H
caS2P6F7BsMTmlOTKfEnVP2zQuBakefYso8e1e7JJMQX8ZnO/put9UNR4vw4yWKu8BGlDGn6pBoE
I91nBRSZHBQlDU3usNQ3RWUHrNBMhwVkOZHfmxpx2P8skOvt2b2bn2OCpDq6U+k+5jkpxeaMrudN
KDQXhBfgOsdjpmTaoZFNCg3H/goaxAhb/eE1qxZsFXEOfNf9Q8ctLz7jnJrjZwCdsyIkJUtAEg7A
OwvEBjZ/DBlK9eDip/imR3Lv/B7G8cQVHQ83Ooq4EdOyhlGavpJUvxY5PecMcnvdTYQlz/9PcgDN
whKxjKfbqIoEQMTVUe1w3a08NCCUkOHiFvsCox3N/5D3mxkDEeAKiw033rztgBdkLBHaHHAKExsB
a0nymZn2AFcEWLYzsV7wpJOmkxyUHDNGBHiM0YnVMGIZOrsVe+/0YMN4ppb+9vtxvOHLK7b98ILP
sZCDngnuMPzFaz6x/kPpYTznEUp4BH06vRBF2WyO6WGbJxWL72Ed7bB0aKcT0WKkynCkGYSR1j4i
1DdT16a10Mj5y5llki6LoCWdQAgmnELM+xnq4UQbRc4I4vCJ5N0hq9xcORJLExtZ+7FYKP/dDYzb
ZOht4ruqBGxPeGXqg/9p0YegHNlFS+OQXmMmNmaWstCUy5RPkns9y9f+pF6v40dBihccFORWE5BW
FtUkBTkCggjT9GrBkWC2kyGSeVG+JdPYRYjD55Hl6eZgyQIHFLctQGiV/ZXYcAjHPRgEgVqdhKrm
SF+YXPKXDMDIiusLrD578BYCA1j0fQ0wuzWsy1gVC3RnJ6rTTjwi4i8IO2lcSLWiE5yEQbZlIhHa
0Eca9CmJmQeP0ffVnRE9HBXz+N0vONtomWx4ZF6wNGwwnntr1Vy0SgO0k2HMz3GqpWa+PK0JeyFN
tiwqOPtFH1HeVkil4JKDO4Gwhj9xfGBdio//CU/Uzwg+1QPBJBfpBlEzm9ZQLBRTJ6pLsbuiJOcN
NQfzRshm2Chg6mHnFujwaSENu3m7Gpwf7vhe4tEAFnMphCFCEvZIbvlkRsxWoKx+Sm8KlKu/EeHK
SDF8JaOH75DORCIKVts5nkmLu5JbELm/vTMw5bCQDtaYRGNi4Ajswcf2PClhnA7jQp3CZrqcWFZ4
6CVX4zpexuvv5jKXq/BpVx7kmI/E065XI5btYlmSGWK0YeMBD+y3T7NlAqpyn30ifO6kLGd/pHAb
AHQCREywh35rI6YwUYnB/uhbjH3RBtPRi9TbjY+T0HHjmI/yFv22Fh5M8DPJAk8f7KN6FXCUVcmv
NNfaPUyKjj2AOjpNgSzreYinq4f0T1mUWuhEvd8jfBrGJqXXcsu0PqHe4HlrN3ffGs+D0bXBFc5H
B3AN8HN9/UyWCA3dpYyIt8/wxkU4MRKmZWZJMY1HERRVl4nCQD0MWjmbCq+nVac/bwFOYq0HSbhu
EnCJuv5ri8JQ1AAsMJDgvsD+CIdIFK16AOHPEi1OT52bo7xyft1oiwTyxZwNhEIRDc2ui5aSpdEJ
eSXkhrwAIBcp8VsnefMc4nbsVKYQTupMTK49zs55dH2Se/2m+pqPxH95SgQOd0q8ONw/0eFa1pAi
ZWrn9hyIlt54JgvnG4lsKs/ydZyBYWrbSMVQoj24MrxyNTWted2N6g1hSx3NTy0BGJljqvNuOzng
UniuRvUCx1DtTogDHXpxHSOv6AVBu7ugp7CkgPDGZB1bSNi+rRbiju4TqR/7hJQjZ89mTQy/jcyR
X2mO9z+sjb0CNrcHs03+p2i8YClX1eub+1AZAVCcrXVzxLMZ/uGjJ1C7KKwZtifLiDiSCBbzlFFH
XfZqjtJUeP0j5EjatbCbgdwvl2J2trKGVRDx1XlPDKDFjrbtXJyGNvojEhXbuDXReMe+Dm+PsSAr
uXvLR3hOnvNLhtzvmsp8nC/PgRVx2rFSpSiaiSozteNhUrJ+BcE5KljqWBtRSnQqPZwB58qFSEyh
3kntaRbv/Nrc/wyCm6cyXVf86nZ6m9eYDhLY/tKTDr1PYLFWtDl33p2JnRb9zrKdRABt50XJRcGd
axHMxfSjOrj66HEAE6a7LmEs2mcI+FivNMU89CUIHNo6zAkGNocDpj5mXdtyYu8K2WbjBLLvUSH+
4+VOdh0r1dwBQ56CCiE2cd1FMUluJu5TG0Sq41rrccEG5FVOoCrcNdRYc8izKeF5n672fPK9HytU
pqfEyT2q+0xkN/vcWPiD3etgnZLZXgO/yUNJMGxWMEb6xrVxF3iHbmL9nlFzS0oVtdX5vXWvc+Y/
jyhA3tqhPo0acK0BqJ/EaPv5g+w4PSlhUtIT/qhixlNnjxw1otKh7GfKHFsu+0V5o1Zc6UFcfurd
9qhrhPLVvjclX9GEm+cdpQNrVVNG0MyfyZGIfWguqIy1+fsyPnxMlh348bChcTgOHpUC0ZDQz3+q
+7pAGEmuqamSOE9q2LTe2BpbvL1xo/FKUoxDWXUdgjLKd+ko1/MUtSd9OUN0v4ul11T15/iGq2/K
utIKdlsb/tpnJ1LSWRSGvjgZ/J/pmMgB6F03mzwsvGFJUsl/pLqKv7tdP/wy6CwPGzRg2ciKmP0s
A2+NNYe3zVXCcsl8yNN1EWtjeASj2hLKBEc1Jsof1SHJCj2T4o69CsxGoJYj0ncic/i6Stn5i9PV
TGSqKxWm80v48N5oLKxnvmr1bCKYq41CEYnKfcAMZAfcQoybzyxMI/od4V+Op2hwWD+9GyRb7855
fYFe/ChgWorgd/u2qsPtFo417pS1wmgo6VcX6ujOU6XEt93tDYLBkHeWv+T8B/X/QXQJ8iAwnXhf
DeN1SQwarjzM9di5EXzDI5eYNT//InDbaI5EZ4b0BRxJTHaeA1Av8UuR2aJK5rguRxIwmb15C+8/
lwuDwg249WWXNWzeNZW/h+xKV4IF6/FhCr2CY5+LaI1YtWxZDxKGuo/+DZ3VWsl6Jav0UYTMEjPm
ssRKkKCwBci5SPM+pSZHiYyUBC27W3+jcEp+S2zaLrnN0t5QDPKKxV6E+uSoMh/jvFPN+BXwXaNG
1hc46hUILPJLa/yGkWm50gSiWwcZFV6CANECa+3R9QA48RB1b5rjrlDEw8pJGe0WzYlsN5M+Ujho
S4B6b+xNh8aRUHMxThvnI+uXXBh2IUuHHqxH7/vBjcJraPjPIwAVGfQR7aZowWKf3/rJmZMJHTBR
kwECvll5mGthXxVdLPly7k0Yn8GawHfxEBqaoH5t/tQdA1Uab5ydKHs9/eCq3x0d2Xy7IF429D9c
mh967BAqyACNr3iczbI4DWFDM760+t8HF94vkx5PIvictip4awtL2E1yrNtfgh0UTyoaAbH9ekQC
TGSdcJfCzFwy60S9OE6LMbNicMoAXPaWv8eJTTT0b4nPVmUlu/+JufWpk1ezFpMFSwmeglRNC57p
QWq39l2WZYKm/S0EVdgYSUmL/lPRWLpejfium2ATcddvLjZQH1Y+cj8D8XNRbsdouCtHuFtOtx0d
tsRBnfRJCYn/eYW5sa5b2feFvKCum98Uwy1VnT5qLywL5vG8CINgKnVxDQXe60niDxeeYPDKB7XR
cdRDtaaoiJAMxbXaWmy565JGc3Yf8c/MZKdmLyltO5W7wCQ8tL5qPGzwMJ2XFqoZ7ohCOSctgTrg
C8dUG0d6+DXO3LpLY8lty6w9y2i3JrmeDykljziMLhuyNTr22ZhVav/Hll3AZsP8nM9pCJz1pGWE
P/QfstkLYy08Ts7LpGrUyYC4z9ivYK57bALD0ZQkVbnKhoNgALy2Zw+vyja8/l52d9AQQFeN5CMy
C05NE+kFnM3XOKHFhmKagf7KoQxVoBxRaWM8nhkxFReGWMAbuNRJfi09JpSY6sHQXARZ5bYE5FtA
2mXbDqRP8gwDHE4AbgtYF0+ONG5kOcsBSES6PRb+RBk0ad9Aown0pvqWcjd0c0hRJytwAc5St6J7
jIzNhfM2osA+7wUS60fvN28HoA38/m5VaPllH2ZlGpr5uKYDWdn5h1Xlq6SfvpV505vzmuE3mAqK
zQuU1P26j5wYSCEwGhnHmCF7mACQhG7PVJ0zsxpX4OSJI8K0xwqTGGD6IN8dwHW+I9SgwcV9RHga
a/v/qbG0etOUBsVPrqaG+oztYUheG4J4LlGDKM/uAr1S79lOi6Ra/rQy4Hnq+L1XVQ4seJw20fQJ
eqpUt9/9tUqpN1FGc8FgH+k+omiH4jqxLAaPzwgZ49xmIrZawGez/OUJo4kpElOy9u4ayIm5P+ea
ogzfuCK0WhTJgNxK4prJtYvhA7WlG9S6L0oJpS/6y88xRMk1j0rCJ9mbAPbbMpu3LI3n2PHlcIhk
BQ7HjGVK+4fdzoHWDGrPOUh/srbpaqGYvpGwt2D8t3TTmsi1ki0AE9B9r6l+PWTBWOU+YUYdstkm
DFtkT5a7MbxFncQoEPrxQDovt40dtD5twD0DvwdwN/xNfV8PsIOEg1l+PoFH0xozKLptZ9TO8MXQ
x2N8dLa6wPsxbYaTAPME3aCZbnl7Vy0nFo9Z5LZqvxL0wR9HaxhbRe16TeAdBfluK6hTvfcL/s6L
wphwiHRQt8rwFKxL+m3Or/F52Kh0fXlyMJkJrt02eIqn3gPw0QgwCgR5gU+N4LgFU6EvpUjTxtMA
9cMs5EOgq/IqcLfp2nuG/3OYxGiQtqe7Yk3tLTCbcUt3/QJE7sSlircvTnq568ltkfmIdxoJv+Cj
Ck/K/w2Onm72CNuE41zfct1Yvvb7R3SqtnUzPTYAMfUVkGi2a/fsgitFVZBsOTV/xHaf5UfxPwrN
NV2HBHRxWniuGETqru6/Cul1WPz7cUJvftB/3JxL09cw9283W4ykHNsNorBNrPMjXK09DYwqYmk4
nj/dcRJ2ARNFdpoFHbtSqmJmWQ8ZNMVoa+13KCfndmbe8RCHrKJ0C9v/anSdzi8rVv78C/CF2il1
w/FTnixzZfetwjSh4jeD5KX4yOzlIzCsE7hbJFpVUcRjTRcPP2InKlM0gAPwaj7r5PBFdMlS3qmC
PeRlWV+KkxTjMjohMGuUBPBm/2d0tScIYjjXJtrwR1LtZRFMYUFM+IFSQszHSKt29p983VSjddEG
bXkDZJ/H5VPYJxo7lX9q1HDmvfJ8xQznlTfTWJEF0ilhtYT04ffO3so4zN/DvbbqBM6k6QRgJX9g
IYgc+NP4divzu4PBPchpkbQLlN0uZMxguR6Ao04rZC4jSNkm+UIcpg3rCDZnyNY8H5FibzQ5G8ZS
e+39y1H1f0CdkmRStkMLU9DA0P/JwZanxzEFt67peeEvUzEdJ7kFDGfY2JbnSscK0RWQmDsBwDvu
OnPwsmH0zinRp6ry9fQOsRwoX4WFQJSlsC5F33BsYUyEqQhvflojUoV59guI5RhwPgFedOp7kHxW
LUw8ur9wrfPefkDap9FVZuhBE6Lz3ReM+FE04D2PLE0BHQsH+MPRE00AeqUme1OMH8xtoDrwmx/J
f3iBaYugjEbsj2Gh0PyGf2Bu6vmz9mFHlwJLQoIPFqkN0VGxFWUxvDRAkbgmpjYMIFBDedIFv1yj
aJtxSj3f8AD6/nI6HxHbTqkrJENFAch1A2dlGTcEYGIRj0IkpJxVn+DLcXNsQff/cTxbfgdOdHnz
IHJYgwQaITXC5UlhSMHx8UHca19OsSoPi97pymInbDJ3TrasT0/Ddh5+UNqut2MDDG0dT7033qjr
kpEfSBTj/8xclAUOuYpRksDM0DRAHBIR2BM1WEbYp9DsV7FPByTsAqUOpkTSMIy+L5ELo2cxUzzv
mojXF3wKswM5JEupK6R7DtlkVfAfq4XbfhNDS2O9fFNfaTRRqw/UiScRHyEhiOptY8fEsaKl/20Y
YFMtxJ6QJWReGPouq9ZiLq9Yxnq16JXVXqkeNQ37J4lhBz695pgvz69HJ2672smr1p/dCmMYNQxU
wnGw73CMKL0KfiYm6VO0nwMLYdVvrZKSM7T4jwuXcNzf/4eAMKM92xkfAOpR9OcSqs7RKETdKhD5
U5e9YagprZxFX+r31orFMHT4p8r7Ke4rZyKM6l9MvZ4Wd1XaICLlVPs+i2AhYPAuzvZ09Drr4+LP
9OaFHu0u76AaYXRUqo+lAToGFE9548DHudLMag9diyaz1ntFCKw1T8/hlIgJRu7tDM+IUQREokEn
/Xw0kfZZ6JPNc1XmMV1GsEoDN4njMjPZ41kfsHmegVbmcNmDxYu8Xq04xBo0jjfzzF8RApWItTTf
55Bo0BDYRmOERlQGO8AkPa85cDiDEbqhqunzRWRchNWAtVgbjWXCNvo6POW4Jpb8gzZTq3K/R8QU
YQzTuF8MHiMp484N3Hyii87+sMacIYYi0+SJE5WiR8fZdSs1UPQWlk8qD79lZ8QyHxXLM25/DMX8
IKPLKBxipzFsUy6owfgK5d6qkfFUeCnmP1pskyDB2ZhYIok5nvsPypjV22FM91wiocKWNVWs6Z2F
0Uw8XT0MunkNXlucI8WWKaysNuHlICFHJ+KmNf2vWcXBJuxbmr9sguwguif4rOsjCsDCqAyIMUyu
o0zyxjhGcOFYwC3VELXv+gNxyd3ZJb9oJAK61e1dlDz/QfRLo+1SZEjMVhcuijmaEFNVekDqCYWg
2BFt5UXgiT6E75SpSeIpTaVEKBrKGIsJsmfsIZ5PTuBlWJrSiwew6+PrBEPSJqM8IIa3TeqKma2Q
/pcZxgDxYMYPTAWh98eDgYYaAOMcu/uh4ZTX6PmdOR3EDGvR0eg9p73UDuUbN2oNEAE+JBmgE5ce
m9TS+LkDub6+nuU2vN6PmcdUcD1QkXn+nsbRfOazbuHHw8rKgSvZptoiSCqh/FIyJhfr1hnEcQjl
RbiKZYiMdzezhFqRikS3hHa0GElKl4n0Ls4JrmYrIx/rRjV+Q1OVAhnM3+QTLwWpzcATqKy49g3O
UHEKrDJRKnk28AhgzcXU9sWBJ8Qj5teY0fRL+RynP6clM3auRiXv0W20wkF3zwuItWD6hAz7MQFh
Wv+nESlK3boofatzEGkZlYRv+8f+nf4/qSOtLAzdbPcH4h5Ey06mGeAb+N5nExXOnpwreN18S+AE
YYsUcEoePS2c3iR7nrusXL31VZdJfhGJBRpDgUY3VRi/Cn4FhVUBF4QDiysiU2E/n8dCpYxNRKwF
mS1y7lj9xe9g7qc6XU3RCarLWEHGGHEyNcpfFxhBr103sLRwYFwYwIo5oOJSeBtR72WgGjxlKb4R
95ohCaiqHqujZKV+kvx46Y5uPbGX46Qm5cr3lSS+m5uzJIP61JD+RdGF+goP5j8gHaufKIZ1fyCw
GyI9Kw9zJ9xUDTFPpIqWwVzDUWv1gyZ95+luhZig2nrOMc5U1hn0u8RbuZ/2Uh2zZqdBp1rBVlsC
yz7v6TWEo/IFy1I5TVHbRIXowXeXpOr5eUl2JGq0/5ANL9Y7GrJJoc33HzwAI5fqoMQWrlGkMWJg
kIB4UgPmXAlcBV6O+tk1WxrN2ayvzF8TC/RX4R2h3pFV24mwazp3MnP+d91rnwGh/9bdiDp/1boC
ut3FMPWOYUiQfGVaeDSNWmXpINjbkvg6vzJw0WYViybItLw5JnVs2oXSXViUuUKrF2eWcVRIhIqI
9yByXIzeN70DiwFsJdl56y0r9A+1IleIyALrZPecYLz0SLz01sHEpiglWpTGTwFZ3kxeEZHh7/cN
a9sCtY0Uieh/agu4ZLy0DnP1xautrXHVqFbbqW60LUmd9Ddx8kFXSD8vlFfD42Xpx7NPv4mNWxGm
TtUitAEUhuq1ssXVFc0cjT9Ti35Qvsk8cHUp9eMyTxsHlm5go5rKxwqFMqBMGbSZo7r9KajVGrch
lrEPc4DFxH0QsVJBNoEclCsSZjgbwCoSnwFAFeKnEgHLCZfkmVCesAMPnoRQiVfXROsOCoNPrJ+4
EhtpSgWYZQfbaO9yVyjF8tvC8HKvFXrHhg/B2cDNlK87MuIK3OCvT4kJOwMCMrq/3Imo/w+KUXmB
lsZFsvHFoE4AMtOiWRr+YM/7K7Gvl1LDDLO//p5tqnX1NOxKvy2kgtOlqTentfrQXOCnhQtWk+di
h7hxCviRyOo2pcAfxlVejg19JGzykvM4lZSMWDCy36uR17r0aVGirx/G13vQPgx1yPXOSCZrQSnW
2bzvzVgnEkvfqArTR+GAKtI3O0oLWuITmJdAvri9FpWpAmeTxhnse1/rFpDtRh7FWzb3474VcIk8
J4FEde0sUgNpuJmhfmSk/WX/AxZ+gD4JmKdmPsqSUQruMMkMmcwucFKUDYVJkSXoDL3yjHbPwJcj
c0JdhnH0frtpWoIwPRyMs8CtB68RdSYiJanTO3uBT+6z2yjRWCzoKw9kEiqvU4qZapLqV33N00Q0
/R983Q1JeWm9VL3lq2lZJ9SSfVVxtlUpWKdkPVVA1XiRWGmeBmbFZVM7YkmCKkHZ127ItprhD9Rc
71TNrbL78YzxIg4WO07yTyOBZg8lRReQsk3eOqSyVSV0YTCFOL7MdtgIftre4nsia/Jqy4AK39g5
bI2RgMcgTLu1oMf/n0TJo0GxWLN1wdTCjA7OFwds5FOo/nfSJ1oxgK3TPdBK1f90/T67f6foJ7pF
gkpL2YYt6phatoolOiXwB1T4uf27B/RWQwUHJbVppD7Zu4PYgkvp0ejpDixfSqt2a/lA21061KQS
1KFNiA8VdxvYfRdur/WiPhiQJzN9erWd6WrtQjwUhDpAPBXacDdHLDTBRIzUA6D9tfRIKo4JIibC
1ZBXhhTX42tJh5x5hwCvEYY0T/jutqJZspX/wGwxhtp/Myjc1nIATBXaDhY9dthXQaMqlnl4Olde
dZvvtvAzcREjaFCzTqt0rzKUk4QOxma0rDJOIFXCFStTPqfesEtOCZhmsk9UuSQ21eQsEe9qE5Kp
MEqU2RpEIh6vd13IzrxpVUy/Qm75ZvktBCpwSUxp23lilt9K2wg8hX9a1GINVUhaIohRcGx4/Nvd
vKFMYx+x2kd5AOQCRZ+bZePH8ZcPMrDI0tHX8Uo2+zbXL83hHmUWBeh8/9GI+tN0hi2ZaESgV7Sm
YxYh/JeHsf/8BYmOvDlG/wMe2Q7BiyODvo5tR6plN9vjG8f40kyYjWyq//1O70PRyM1tqJOEyfgF
p4mS1uoVtBCa+c0GeT5/au7lCYVdyWaComgsOuRxE3QD4vudBg4zoTSFSqFTxJ+5lBOnhWD3y1on
CxBAi1qVkmMx89wGQok13UtNkio5kJORPHSnPyKRkX0bcTXxzL9gxjx+9pU9TPAUEnFNhN5a5Q86
aI2Y4H+afH7/YyJ3bTuM0xFXj1touxa9JVuJX62ziPfN0lnBzVIe/WOR5A1y4LQxfaV4Wu5Z1RcF
fm3xppNMxFTUWfeinAPbpl9ze9XVynZG7wHFBFthbDoEi334SYXe7NiSz366ZNxKPLI6zPupyL8f
op+vKOerlJ5uZV5zaUl6cLTP5Zd/db/EFIlkq89gn5QEiRo5L0bQWtK2yYozKODwKbwBA7MKHo13
2/kg3DYpxbFpXTjJ4JaOzXhaiVP2WfXkL9TcwQZ7uY0Ejs/x1hprtALzjD55GN0F/lC11SAAfPfL
e35DUNdzrwVcncRNxqsXUud89T6eXw5TVP3XkVJsAsH+mCCSI+PaFNr0rGr/azpMzvuWqy8YDBBx
ybei5ISo3PoKfw2o7ZLWrqWbHu1J4OvCLPwue55pgQ2uZxJ4qrc3fvQbHHVYdoEcYWQBxMv5L7Se
r69gU0JOVjrWhFawOOrGCjHSXbiE2mIlOmoeO5PCjYYg5Jafkecya3J9JWhKGKM7gO56+gyZ6Nft
Mm19mNOHO/00LTkz8eCDuehMSzNzMG0MpEXwSsUGpL+HO/t4EuPbGfARVL7HFIv9iU7CFL2+wLF9
TOyrqCNM1Zzv6OuufwS95Ox/HlW4D9GRTi4s+CTi+cP8caWonla4ZHfMzx2pHZzCcDVe7yiMKr0u
QWdjgwkDJsbVaoJiEs7l4aJfWmmiE695TrFkDmOHeuZAbLqWqOkLpX4ielbk2ltfiDQqFCHFFZOf
L89iCZEDsqnbR9Kj0EsKEKF+WusBok0EcC80yOyUdSC7SXOVov+pWO++HUgWL0pYtLbGA51kM1a5
yKHZn1gykGAcapHDHJBPW5Y68fX/Oh5OZWXyjnTzyroUWjdYNNS+QclnFQzc3TDxPnSHg2aAW0kp
ebIQQZ4PxlcnJnp1n/j9TQo1aDemCLWh5qEo1ooQXEqgAHkv4Mux/G+pizWc+bcH+JRrE60YWnTK
t4j2HEbVmQUadK8SUyXNaxZEIxxamnPP4k7b6ghCiVJ1/of4+MFO2oHQAFLSvm2MODyHtlsFQW0N
u4jLqWFYSX8FFP5QXtktB7/zzVQC38pl1663qfEQQIUDZcd8nkjS7qZ/H3JXoP1mc8ZUSBXNLZ6D
l4SCF3qrIDKu4ghWyeQt9EQGFcSxzt4P0KU1ChPuKVLcK/x4gKqSI+y9uzHUzpnYz4RF3KFMULAC
ANHtzeLXIkPU7OFW6RXDcnSFuJFXsDLgiMyzAqqA26FidC73DBIfPbS7DaxbvhDGIsqjH2JDo8yQ
yZc8vnwAglhDLgbUgKDcWJcueuwngPYXyOg+/UXDUtZRf5y8gv1gHO2Wuh59m4vvvFaC3Y45PcDz
BASfWSILBSyqu7j8Fs/+6anTaNYo7V6VpbJSt+NGFjC6sqpAnNewBfK1f9mdC9mmDOWDLfEJNKgJ
ueyVEXlniGNk2UMvtyUO5LYh5aaHNtVXV86MYGqdxnYFh5kAbuhjbXlfz9L5xkXdD4v+yxfVSuGw
mVIgx8fJYXt4LvzI32Yc8vEIeOp8dQnufZYuXrEyYaXYX2GzLfyd+XOmD00sawnFRUKaAtgoEQjH
agzQ0VMrIrCaDqbBfra9zWipkdWTwfsenbiM1ra3Vpxo33fftifFLTTpGnSrDposjvY/n8TUkP1X
xRWkYI89J7JqWY5ekKusgmXC/pfQmrTkpNPzkRARiVzcMd9ZWyKMB6yAg4I5Z1SIVDYTA9Gyk8eN
1vsWVGmuO/VYPfk3BFH/0XBbqrDWPpC6ceywkTXDo35MAVjtjfSklnc8HDvucpSYkiwPFmuJHknH
jTa1PMLrVJ12DeFLrvjUt99xr3p1KPrVsyt74FSQgDdy/h9QtWraNLI0Q+oSAcKKmcR33aGv5QlM
Q7P8opzRLUU5RFK8ueYCk3On49bjhjL4Z7gLAX2ngqsbPASJFHBxL/MGKwLJspHFV9n0ymQs1PJ9
li7KCc/4a+s8m6hyMM+Vpu9P0fb+GmHciYA3Ok1KNspM/3lcyR9wBSJphLGeFQ8Vc4oQF/XifCdD
CpLhGf7m1EKJEQDMVZNg83ENC3LD7HWZfdsWUEjWT2dQbh9y6IynOPVn716fn6DLAoSt8gIiAhqU
rwRRJlJsA7x7gMmLlIo9HpdkUpttTHbw84rUAVkSP3Vf2ghxGF6uXbxDVsoI2bnPVr92wrj6OtCU
tX1miZgrMlagA19PnGCWCprohq2FiYjBcbzWoPMY9dztOVWG2Qay6BIl4DRtyQC6VTmQS175VLcO
dbOYgxftJRJUIHe+B9sDvrtmOYMtwXdoO0Gqc3SVc3Hhq0acyYvMh1bWyQ5H5JPqo0GGFkUvQfN4
U0tKcjTi0JHqNZclkgnHEm/+tFdteUiD2ImtA22kiq3Y4pfwmzSfoEigH7TixHPwa/EGmIM++acT
MqFAeiMBAzpb2ImN6FiFHC6DCbt1F7wX6lE1HgjFmTuJhKp+NeN8mDgqDikSyu4VD/+gVen9oNW5
i0f5AJ1FbeMP5tQAbLFnrBdVzXjbISa5SvbqdlggDsImO8T2cQMkIBzunZFXl9kpRnO+AmHP2hWb
rhvf4NrwHe9oZUyHsF/M8ksL+zJovhdXDfro5JYwZn0tNSwgVnu9EUjU3RzWZyM8XE+IBVinobKK
XQMnbPHGr2MWd/ryd5yLyOI+ghnhB20p9YMWpOqkzgY0NbszZlH2xHUy7YTHLRCBt7xfwRpoMENg
esarb2Pr0w4HzedKgA8VX1ooM7+LBaoAhcTDARP0nn3YbumB9PS/dG8hY8o/t9dB2bmRgRGSUtmQ
Ozj5HKpgPuV+dnYmvJ/Mei2KYMBGtPxO6rU2iS6Ook6S3IA5RgFw4hOla6qflgpH8PVDHsJqbTdT
ZXlottgQPqMzAEjSTfgvMeqYyUOxWsfYRJweFxnfxi4ewhgQUZ0cQsY/9yJuaKWp7PP02XF/9bjz
TVROwjfU4RwGIAvNasXoC3HngRD9XDV81SL/ms3kdcJY5dyKNGyFw5+wnz5zEuUg9VtTLxQugxOe
sOF9Og38px/oR20aZDLa7UsSZSYfD5XkQ1vfjVXvZg1HqJ5DdY1etwRRpxUOnIt7DKyD1qxXDPpn
Qt++tyz25PwM2H3gJ6UCESux1px0qWU1s6uVLcQ354Y+yfOTSZXZoLDTnzU4Gw6NfoKOcoOrI4w7
WFNLODdmBMOBrl1hgIeOQcaACSBHKRIYsdYGx2yiABYK8sUIManhkyWyz5iMD6IiOiRYW/+dziAm
VGIJARoi1jaOcNzgXdpQZEx43i+f13E3QZ/28WEgYkH1y/n/tgFrRkqWyAinJRADU5kNGh48ZBN5
D4X1cQwbXOHE6S5TduVqhwqR/hZpR4xCP/tcl6G4PMAdiAy5ScJqEImtKZGSkXkzi+9Cs3lrYpH9
94E3jA/697bd60Qq3XF21kNmsSxQTG+iAHUQffe8i23RY2FrTh5p/xXiFwS4JFiumzx+ki9p1nIs
5yW5Rfi5kfyobMJHJTaq5RStcRj+9i+p9p1ftYFFf1/4vOxjiQb5bqK/9kshsPWC3Xfk1bluanHJ
3Dx/ImLziXBe9hAqa56oHl6h5fQces7ycd0wWWsxMAJBNtuEWpe4+AvSfRIHCMI0vxPBHW8AJ2U7
1Tf+/0iaRmMvO8gLwjwtHcl0WSAFOU5DkSyC0OgOY5Jew/kXHWj/6l9stpO5ZLJP6pLoFqQqKGOT
W/igAgqov4kabf7yS5TzmhcY8ccktQLITtrylgQigPgyV71Ky4qtXdUcRxDsC1j9w+dN4VLm5SzA
8VEMnB9vvsHKphaWMqb0EAYE+dKcQeaX3H0On/NgOkA67FubPSgMgIOyKuoVuK+C0rgnoBx/PgHz
UpEc/AluimHHZDUw6JIoFUgjmzFvYHMvDrbwB3rB17/ckfXa2zcnt6bGcjndxVzXFOMC7tP9x6sK
lMA0m+B8RXdO4DI4jxf3z4GP7djSo6ix0Y1cdZ3e2G1N5kLf4SmXXplePaIZhL/oZXvLsa+sX8Jk
6U2JBV3GwFNrLF7RhHTQYUusa/QmomBXsBio0s0bDogpT8+a5q2GlNd7hDbNXML4MB7nDtiqnC2q
tmiVoiiKxFByOrdfG98lk+ySEyhuoyVamho8PtUAU1tBb9mkh8nMqGkOrbh1vs3Nx54KhMHL+DSc
U/mjcpXW6Mk/+QzWmjJcB20oDLpGwvxvq4JdSZrWtHLHoLwR+h255dqt6cS3se5mtRlTD7rrom3Y
GVfMxBFs1cxWkHx5qkfQFtRbzEbpUwhxzAzeJF+j6xWnRXdS20UnwC5PXMcobaKjdO0JoJiHYg0h
dTGOn6xgdDjukN8TPgPOlhj+Bwm7pd6/QIGmJrGk36pSvBi5Cne8WckcD7DzQWSqzvros5cOXRrb
RVYP2TXC34p3D7BYRB1HEpwVxvH4xoYN9o+8TSFWUZjfFXK1utEGxuXbpwMReSztxaLmKEidfxZd
ANKU8gNlsj8VeIDk5ywthmJ9cIGbQ0VkpbqESuQiq+ClDwniDone5mAWiTq0oSv+9uPjqCxwHQi4
xL07FSwkUWN3nPjWh/8qcf/IjRVMWnDm919A8M+tnJeGP7Tg2tme2ROjCbvysNNCkO1KZxcUYmCZ
CQWQz3NcE2WNLZ3HCZ/zUG5VDKZlYqaiEswNfnQbWUo92eX4FuT3zzWoU17I4sNnz/TrMbV1uEO2
/BzHCcEsaKE5coVUfwoBbXCm0voqUsH3q9kPfzlFK0m3+o8A/I8lEj58Keg0Yr3XezLdbzVQzd/h
w0KCimc5WfHQ6e77rhaaDFfhSs6/WwdAzMQG6HN9BO7QxQWc8ZNnt66QBMZlwjlIdyssWfqsZYJF
6pGpy7+HOBqp0m8z3cOVrUhh12lAHWkNJo1LDTYQI6j/Xk3SWjmypexud+UvMruGtWtr9JJNiYad
/Xd4ilwK5YVgYVVEQuNvz9UzgjBb4kwWRrD0FRPFkoIUjtlBGda2rOlJ0j+PcX+3+HSBeDxgp8VO
RBBwZWt6Us9u8fepbVtQUhVXzXUIyNFqU89oJmvcUgxHxjvDt8OK583y8N8vw7edxEzhHpsLbN29
3M6LSDQ6CxAq7Px7//zJ1GEmWu1xq9SBfxsNlni2yNs5omG4zNt1PR0VmYeA3BZq4w4zPwWQTxgF
kHuFbzcjD5XGkWcBnEFiA5bs+5pOhxwYTwon1MWr0LWp2bt3A/jl5TI9Gjm9GdIALgZ2beLkfB8G
e6q7z8Axu2xTto7CdODm5xOSXs+UQgUiSzwC2M6+c6M+vMnPcmR3ROmYgLtfccm35071Qop96LCD
QtxVdB6FgHscCorXFfKB4bMRTjOYGNAbRX4KF2p65rRpWEUfpPExhLQx3kHd+JwH55+W2mqV9AN6
StI+PVMeSnOSbAf2vMusIU9ubEUQgZgnOsXjgSE0UX+bGm9l9Rp8iUfBoYZbEKWF7cOPa7JnVxGK
ML43lbqutHLCQGpxzaBpwa3v/DvNy8GPeqGn6s2+NBrOlfaEr6WVoXDcB0StS6Ht45wgfynyENNU
ogVQkOkNpXKohLOP5rPbfLlydYtVfoy6h/9KlhNE6RATQfEE8mi6VaL1NLSj04DGnPORjBhZjzoF
LOt5WhOf3/d5PFVhPlvNFvXkKsPzNA03hJHkCyw3hR18FxrUfYSXZoJ+oA7R4SnW8jzO1hM3e4YS
96AXcNrWkWOkZmdVzTeHxFEja6gHkVgLoZ+9C/rRSKdfjmjlPK8OR3qa4G5OryDf/yB78k+sDZLj
v0/a5OwmZdVWin/ifJVSraDfuJsLsPSyr84cfEvEqo/foDPb03sE7HeXkl/0unBIHIoVqISC8oLa
WLef6kAWCLEgnZi5IT1IIPHAaW+d2cKBD55xsnLXcsPuaSEhAxOfPRhurFn0EAAMdF1l7auSWqgv
1PqMw3sJpAEh03+ocISz7a72dWupEFnrMM3A1A4d18h/4UiA5qfegwBpyvEbNMZM3yPziWSE2lKq
ckWDOh/0FhnyMakPRuizKlnT9x/2Z5IyFNGlpRgerJXM8orkkENMrOS2+o2a+zMsLVHsvQDfbOSh
OPEBD4/n3hwynD1Jprgw0kqK2IHpmdAnVoccjs5k2erY5K6hxoWPT+okKeA0SYxEkbyLgioJiHxm
99d5I1TjEj3OpJbVXKu54xuWJDtj1pjl0ituzmSzhz3V7lE6qfkf5gAJoaXIteMSzKk7U6QJVwJt
FRqw48GuFWrSkVh4DY2UJljVWujzUBbsu86fMN6IDE6TmMw3EjtzOKBY0yk9AJeFnpLXgrNuBkXM
sHbVLn4A1C6jSsBRJIv6VbBGPVgCl8wWMT3bx3MzDKy1bzE1BHHt4IiTExX4nF/RYcu4sqUoq/Ri
Hhegos/G0EFtKVHPh8nZVRvzHcu+Fk+gXRinH18H1fm0nGFa/SIULdOLHpB+10gNaHG4/C/QCZO9
pAQ6gP6jGbS1hRMdjXj5ctTRKFYPW+gn3XEIlc83/7vmpVmnCKhqieFQr48hqAG4mKSJ7Xj3Nohw
tWmu/v9gZhHNbgBGBKEjQAcbomkmuHg7SQ6j0j1uayXrAJHGA2a/QZaXl7VT7eHjxBWXJ6vH5qGw
+IjeGbV68cPRdfKV/JkbEsduKceus7UHbt4FA0l8iCqtrMU2DHhZHUah4bq1naniQK/ggw6OV3rB
EguOfSMZmsn605L2mbow4r45SWKlbxriNkSBVyRR39b9cP/PR3GP0MVoeq8NNgNuzgjmk10QB2Mb
AtUh7pFt+6MuqyhfWZfA5PLOBBMAvpyCy+Agcj1gMq+0Nxxa5eVquJEmurEcV5U5gyztDJARgLti
+IlNRc+dDR+rOTb3d0q7sHpsRncQ44K7cWC8YKU1qJ4fuEjOwgLKsBPjGVvCLJ9dGB59G5UluU0z
IheJcOOSndzY3XgMFGmhs0I2cH4YUzX0AtkGBOkmDmA8ngHN8jcSUh41Z8W6qUfELoJgqKtOYA2G
iIEKprcxtoRyUO1yTjV3t98Vh3b+0mLffnYIs8TpIbCFLBIF/iPgPljd/zjqH2Y2g12kJrO8+ijg
uUsACy3WOuOvG504cFBIl3uO1sZYmm2d8AoGFLaSSsgtMjOHNIB9gvXEwsQgYU3oRsNgBcFTAaq6
KweuDe3upJpwP1/LWRIw0GHl73nsRmdv0bP+zeG7lZBsJTcLqETYCuub2KE3bPazmScHNaux0pVk
WZd3IJsyuVP7DcBc9ieR96zrt9lE2ls0J/rBPHtcJ9kRRXhn8sKPmleIf0MaAsOWBezOVvJa6c8f
eC3Gy4ShVO5+GYw7j2vapTIKG9jE9RdIDEzQYGdu1zFmPK553/12pTKEyFdsDizMn7vFBVGBsms5
LhaTO4I5RADa4hYkPGzQg7QRT/iUVDpMyvAVbmySpXedd4o2wEIxCfmRNNcqpy6VBAlJvvRqFppa
2vKGhKO5qg8RqW2vHMak+9lc1dA+xyc2117i6NXcqaP3bwFgIvRRWXPil0cxuGC9Dbb4eTOUZbRy
6s+nmjF3FtiN+swxnOsZUj6DdYNpmzO5FCBeebbsZU/uBpiQpPPj/d3DxTMBeegI3bDO2RmgdrnS
13IegEoLYsLhGqtqb/iTo+on8V79Z9lN9NbcZ99Yp5R/31tOO50ZsGyUR/YW1ziIpA7UC0wTywjL
ezkw4w/s5Io8bbk6qUYnc3cXk8Xbsef/ayIqfTag0JOzXpXtor4BSYgd8ePU0yZsoLbUkdDJabuC
k+3CjSEIoYeB4JtDbAIWILMbn95Kq4EZ9L1pA4VJpLK2J872k01UWIN7PpvoaWJCOv26ih2i5T2z
4UpdvZaY8CgFf6A7BUFa6/bsDJBJfJrLI2t94rJBvCS2JqcJnR7xWSD277aRHXZjMZR7HI3v6tBX
JznfHPPhAYJ8n5JYNHV0ZnFam5YE56kL3zjilgvRe9ZePKEEOkcDw+25yEkCj4pzM2orxoKlD2ef
/54MHFHcA6ZrUjavUCFrrJuPhSuza4WsDyWHSqYcJ8ABk+3ooI8Uf4f78ENlQriZ0BTzCy86gXnH
/Z54zpstnndjgrtKNBKwsVrt+xfeybRLdUUxvLTBAkG2JChRGTHRAunq0bQFh6ZwIyxA1SWLNmKW
SIR3NaJ9eAUOfyWnbxKQhs+T4rlLqaxU/cXreFJ6fsljTKw3blLPFQNkby1LWehi18ejy0Rl+TnZ
h1lATjtYk8BNMzIaMwHt5t1SUxfpp9Wd7Nf6gZlvIT1PWm8Fyg8ahpfgycMzzOF8JePhKVvbxdX1
f0K8TLKnjPTn/L7zcTf72FC86N02Dx0RrqVQpDo9gn48L7ilDGDlqkyQi+zSqLlwcm3whsJ4bGOR
Nz25ISow5SuvwW/UlrBVoSqWFuUTJ58072ORGyzXiJqgdC3B7FEl09KNPvA9scTA15RPGNASjJzN
KWhKE8mGITWuUTJhISvLUrYBLYM19OaHkHbM5jAr/k+TSdBshpYF2Wg/EDvwNzwBzTcex+Jm2wZG
IYaH4qi55XPd855BZyfjxZZZUuSXBvuJcAlFSdNBrr+A1Mi9zomCW5pGJZQcU9Cpo4Gqwp+s6O0B
GY6DVUJiboEbgprg+L4PkSPsUGtlPMTKLYGpuZc1IJdT0SQ6VVpoRXcyfCfRfy+Id2tFRxm1BmHc
272SsAlkGyamM+TkQzXD4E9zFTWqrRFTdJJrs894Oabtn6jLWP4Y1B1q+7NJTsdXjSIc5X5zHqK7
nUCpnN9mivj99MuEkLl/bwFyJxZR8PxRZ3Km4VdVFbiE+FBzC/knApw9ICvAivQctnLIeSGMTRwz
bNghvC5ExetjpD+c9YH/pl8Um+FrOeUPbjhTxnU2M4n0lUnsSPxBPJN5rQaHJhs73F8+gjTEE8i0
CGm4ufDMUFJjcY9uoOtg1e6MFtBUX/46uRK3iHwhyaP64EmBa72b6q1XDD+hFe/gPigeuAfVIJuO
wYrH1CMhH3LzNWsu3+rNV69xLtTi6WIK7WbFQprOXrVrYQaC3y5bxgreaciGyJ8yRqGrwlNoUcoQ
s1fTTW6YfNExatQuontOlIGtC0dUyhZeIBXq1Qv/h+kazFKFJrWWXlrRKWomeUXQfby7mKrzIBhb
4XtDh7L2idbcq7D3T4ZwORW1OG5IOwnDteR9JunxkA5PryMBhathG88Y2KdZbKQ8OQKAVMhKj0oK
/pj7a5kNFJfyfkPZJi69qxJcx6rJg2q7AGAKOKUkNEcrK5f45Lh78pM4TGvmmtdU8N5xaFWzkNok
OkhP3MYVwL48/FCuxC83QQIPU2Koi+kvlTlrk/Dcz0XbvJDXclywI8k275fVNSf6YTxfmnXXlvxM
US8Ju7VIGquEN5q7FjN7mKdZr9VOVYgpsueKf4sowxJxyuO5imDNF88g5FwfOnciAe4Vmwvmnpcr
bFBiYpo1jYpt5UNm9EBVDuYwuA1ogBQxQgNEnV5sxOsOV8PIsudvQAfe3o4jUrZYv3X/8DDLqENU
9dLBYJ+0M68V+DJjuRyJFjtnu6haw3UQ9PVtBKgPrX6qWidWFuk8yvRQf+PGqDKBDtNfevZWRoQB
JGJLQEHBM1VEMQHZvKXMc2gJhQzlK1yWSyNMpsZfQOzP+a2NO+yFKnbsuaSkfb6qJATv1LaPmC0P
QQEpX7n0mE13QVJShKN7bxjg1tttEcgeDOwm2ro2Cmm/Ep13p7/vh9jZyGIarrx8WXb91oeteU5I
8UmbsqNa/DZdYaZsyWE5Jr+yDz7RqtgCg2z3kBqCLkUJoURtsDNxc8TqfPxTBSIZnfuzetdg5qsm
5Am+7UTUGFPTd6YQKj37mBw3IuoBVQYz6ca9jefuxHklWHc2q1O4LvX6h5vGfTtCrFRUukXNsZ/w
hn1iaLho4raDJJR//xtLMzUTt75N9dtvTe4YtldUAYI3nJibNYLGap18Qn/k844AF98SJvYzCpzR
4e/th4v4i8VyLHBJpGtSXrAyR13Cu8uf9O2a+OatltjzExQE3g33pekC7fa/aCCfzQG5t4D0N9S+
hiM9s4/RVsJ36ctx1CYwZ4CCLMuSbSuMCtFeBoEmfFEio6Y88fu7++N9izNFJqVUJ6FrBx8axGXf
RGIiKysIyisIpFmMnV1YpTyTOicWUSOQObAkQXdHU5lVpF1/DYbtzBD4ETlhsanQCT+1juPsSRgi
YNHGd6osbkghzq3Ky7M61vkbwKpK60cjqt0uHonLFrwdLl488iFBq2IgiCYgjvKsKRKrPd6NlMeH
vnPTYnU9LGUQlnvvkjqILEAYAyV9GPo9vZ40hah2JRkn6+0Jf4/rt2FCAdXZdbbTEAzBhmadl8T0
NweslHmV9ACAVF4a84CDcFztA7KsL20XvMzTr1lVEYAGgXMdd0XnBBU2gR7kgE6BU2AMb0XOLATx
CjJiKMQa3TIeGnGeKbLkIbFI8msICFlWlYRzLmREgd5+pYQhXYCU+snOfxQJ925Zu+HP/eFfKRYS
egJKX2W+WF4niHcFZmiwEZ7tdwv0pESS+rxa7Qqt6cW46/JVfoxiW+LDc1aGT/ingcJTpK5Cuq+S
Cxx/FIZ2QsXHcQa19fwblmx4ubCVlwnGINjx4QWsCG8j+R4YVMaHSE1nk3qj5FX/yU4DvAc/Zkjk
OduN9iamIykhtLZ7TCEiC+oRu3PhB0gb8yLtyLfg76Ao1Ng9qeiQtiwTPSO7FiacjMz9XbMw35Vz
Zso7Fg7RlrqfHTVkBYudOLuIBIfktk7C+e3nv/7ep9FCzW/IA0f/i0W0sXkEKQWup31D2irkYyrw
z+vl+EzAcoaaIBWbvjrPWh6TAT8KZdSwK+7nTk7k7MhSEZDh39k4wl04raev3S46QTOBpbeQARXS
bktarjAclQGw31uZt+3e4AFpS/IrSyTnbU6QipEiH52aL1xwK9He0bwYIdJ8QQ5lPZY6Ji41J8Vm
QzeIOs3AqdirF6cqAtRN/mx1vqGl0lWYgP2mQUGqZ7OwdN6xJYG0uLVrtcIMmF4v2nt2DoGQuQxP
neFCsEnL1zNpvFDeABpGDxhXw8nnJ5QYeYoNOVhJrpk/xtbD0By7rKDeELeGdskADtPOC1L1FzT2
WpAxPH0tbJlPNrRwDhpPrR1LXN/QFiqZvScJaVMb+xXjHnG5B9zZRwt1ENI4RhtTWhpCYpCeW+RE
KBDxoN1x5IKooO5UapK85IpEubB6cqtEZ+NMVBhXzFhr2kz3gYZQuhmbg8UxoBJcOexlr4ZZwfuz
Ey2jgtFiZNH+dPNVovACPDVWGZWRtB9s3BV/GTFELpvTg6G2rjo7tu2zs91vmb+X76wI/3QLdjeu
PzhbsqVd5yRqOwYDJQNl6jV90cH7HFTHfqXCy4ucGcmC445Pq1SgzUjX8NA07HsZ4dgXuis5MA7i
JY7JWacVazYCW1lIiV+C7Ewic2H6Sm3R7H27YG20igpNiyS/cEdvdsRACYc2NnHUtVi/DDg7Y8qQ
JLyunDU2sL55bK6YeC9eaeWIbsRNdBKjAhk9R44a/2ipFHm1UJ3Fe0UamXZMW69d1Z6oa+atEFUN
71Rc3UIRRdh373TEG1BXlAdwuLiqH3o89oyPWsPu+x1IlYsSF5YOma4YleF69v9KQKW5PiD8TwFF
Z0qqrJfk/v4/AuUidCq8jUhG3zuNsAa4Iq4U7cNBEecy4busc0zDgsMETFSaWXBAGRQf+f65/3GS
U6Zgs/UazJgqVyOQZqsbRN+WrngIn3dlUwgXHswhUxATjGDPle+ouCvXAzYrwSDOhc3xkxTrM/lr
+VVV/r5mfoMTBikeBHqvEJuaI7QrjPIjVhKGKhNeqLYhNHIa65i9+k3YtzfDJIb+jTMB9cn55Fq+
e6i9oqMJpP4h4ax4IEJVHr1Pwerh9sxilYSV7yEXuXv37SSIf6tr/eqsLuib7EqjK2W55pJ8mmmw
n2Tw8v3V4Sew7h4OAOjqV/NN0TxmtPBQ9re2uQNDp+D/fMy6aDGRzsBTC0i+WtdVacXaKeGVrM8O
WxtNt8Ypr/giMLe/1A41pax8SpnlAjum226w35EwlsEfUX/VG/Z5ZRDaGjhPp4vozKelL9DWfZ1S
RreImNtk8OZckHnxLs4M1jPbP8cbBrq+KFp8Pe0dgb7oS4wYvobcrP7JQP40DKNJzXLhK9VSWvbH
6RXt41uJhr2xSQAfekL0rr2idv2MKylpjF3IsCR/55OlDkbEjtqMNIPEuRcCu7uKkaPYUueHsl20
amVFZTeiztL4hUqxsywUDfrae+Hu8iGGA/cdr4sxxkGrgbtRw7hdHPCKS29KaLOFUHpYqvsOwMHi
hmv9urQTVrJ4bGY81Vdml5+qzJwcROwdvUwevnwzKQF3JLlQW/uLJfQ3Up2QYCndZ1fWHZgCrujs
hTpmgPMMpXOqgxbhZG59OyKR4zBlxkb5PqUNQdOUH/KLaWW3iuofJNwtZnogtAK49m1ke4SuHm/z
ZhTY3vBT6xr0d6ALovtuamPgcgw3vxpbJ0f65uPfA/DQV0eyJ4D3iy6lzvRk5PNL9sI7wTa7YTwQ
bl+iAKa5gNJE7H2nZ3tQiiJgIK4anRI45uchms945QrjE1nw47JbB+ClnnKnqkRjOhbFgV30xLh6
861Kf+UVE7UcP/lUyDAKPllBc3aCBcYCx75YDA74peFDfIJQ/1yYtKh65gmT5uiNPm9zn/4wyOL0
fS3acwRQcOzvETeZEEDdsX5sHd4sDfKVhnqIOYtSOTqAcMTy0nYrkgjcYjGc+6ZiAqNHl/QeqBGK
blTaWFXg2Che2U7Fxny7nfXfeft9aVXsH8oMgV1T6Fjiq6G+6htUqaFH6i8CwT/ItUZRodUnkjXw
/xiA+gepco8fPSoJ9+GHsfWsBblTkjqyogkixXW2cSZE8BFVvyQzt1JlL+qPeiqQauTqCHvDhtBx
HH+C5Btd81Mf5nC+1LSpOpVUrqSbwHFi8w0z4ewmshc/5eSIH+bHslOLnGJTiRQy0TYMJ20Mc96U
4ip8tJoWIk1xTZJ1u+tuXbW5SQAVTbPTM0nAJq7HpnUCpOihn4SRv7V5v1kAeexYy7dzh2hNXO7N
BlVnWE0tO05Xa03POUyHQrM5zOSaVsYiA9M8C7VNzSG/YvNF/mt6KN6d32Ld8PmE1cklSyXQrXzT
8BJ2tJRu2SmwOCwYiwg36WRmACoucy477Stn2Kuf7usq/NtHmo8+1dixLevYnda2i50/4JqD7Un5
UAL7Puq/rMJV05o6lwzkVS1hzWYKOl63yws5vedDGUi5Xum1sXtU5RIyLkBPlo4JB38k+SaZIkXt
IO+3ZlXeElunZp+ja+zXNMDjYiuWXxIa1+2hdGVfQv3Y8Lf6NGXKTCnE7nUhRcZ1laf0kTkdEvzm
uk1KxJGnOCebGz8d3kYhnAF56TSbfDG0H3z0z5dXIc1JWyCOvGprQuMS3scgfRX5/8Yv+F8w9d2b
8OI/GpE8QYssWsffKK6wNW7h4hnmhELlnmb41Rr73yop9Y2P7lELTWF7lmgNeRyvkOQ+pEvS+ZSu
ynAxRRE0aPOBRhqyWVSlnxdrC+wRRkiwd4JqTm+PhnD6sI+7csVGz1iGvwQ9LEWtALo7OJLCj0FU
a/DHMqMXSrFYdaUhWfLbbP/BJg47FzGITKA8xrENgLU3S1y+S+bSxH/IjIhgVwzGdeYCCQIF9DFe
jXmt60oIWJtnlXZ1I/lw05ee05M5Qgr6E25Ws1NWZYB8QIOmrsvflXphL3PBt5R06lydxt4CnV4N
zaWe8gQdq4nyxKZ+n8Z1f4TG8T3GRb8uB97jcRNzGjXej6G8m+LnRekq+WCFaXQAXM29LZifxzNh
Mj9fstBn4wZaSnXJium9JzqownljuoLJa/QQu2kZqxbYfMGRfM456vXX9Unm3tMgnzNFxRDsnVOe
7nV+H13P5jXywYxNQAPm7bxh4Gl34cCmY9uuv1pYT8Kd5Q0X86II26EdfIb5ao80niOMgXL39rCf
MraJcOEc3Qx1KYg7bV6GrQqDsSjo1Jpm7o2KT1HS27sOYFdkAUjxkFbl4ywUOKqBTlnt8FnVouXE
hHtQjtzoKHaPqjaGe2DRDyMKvZpLDSB5yaw/54SQ6nbr+hkt4VXIiKAzPJq00WZwyc9DvzymO0Rg
4/2R56AW4FaX5S81mWfnF/xsb5pmSv7tJgo4Ylglqwmlv/y0ouDAGV1DXNkLTrhYsu97bNupDfMT
JTMSHwGCPL6INXaR6/yS36s3GlXTrZTamjc64YyfNmJXFMEagRZnfgCPYWdYvKdszONexavdFseS
lt290naxP6SU+WA/GF8rQUB0l3OMWUlmy0t4xfNaQIUxDYYGN8sXLu09S+wr2ea3fClevzPOO4/B
r6n9vQEaBBfxuqd56x9bz8t77SsfG3nPyElhPtjXOk/G05aYQjW/MvtRh/hvYQwRlYHZEufq5lhG
JGKWD1TrGFRh5ySZu/sDpOkXb4SWYqKDCnrjDsf9LRzY0OAUHFcit5+N8HMbKizG0TuIOKbNiPUb
NB5xvomySf6Bf4QBORXcihf2PX2/zCU2vFRnh/y4YiKqM8XrUBxFXaZzw9wjzWR83E8n5Bf8LYah
4tl0lYjnQX4znCuc4XAagzQp1xAdrqiBxYgm0pV17rodCVQHsdn3QTquPb14qgWhDMBgEi3akiot
+e4HlPrp1rxcjIlRLv9d/035ffALJ1D1B4JCvEIaC78X3tqpIg9LMta/cfLE+O8tOnIIcn51C36Z
yeVfWVxNGeIzzWQbig4vKXB0lCDJkK+R5ElHtME0qVa4gIpmHMyYMb1wrJtjydH8lu2ks6TL1PRH
iyAtnh+B6OY3opl1MtF3wqcmVjPY6qHhjWOy5XVFL9DpD7nacX35fqEPycJUTS3W4dG36bNjy/dr
RsgFehbUWHzrLP9Ufq7Drl8YoyPboo8WLwaj4XK3fii4U8RKWVNZkXQFQ3jesMWKUjElnxj4SMgf
3N2aWMD3joMoDtfpm7Sdna1352CI3cFi/DZq+5eBgZlhIYHdxRkJleCuBoQ26m/pdojqGMZdiPx3
O0t2dCtbSIEvDoZJcjVJELvK8KH+9Xjjbu6L2l/EFV6ztdF0Im/6xlaXGFu2wwFBwodgN0N8f3Mc
nvDdd1aOkTpdDTIkEAIkqQf9OSNZNi8V1lDF9pNRsETV4LNBzjeiK7z1nbXOhfFfVDCl4kusOdEh
kTXWy1SxHdi+8CRToT2Xz7Da/46yxPW5BYLkjqmCTfnLxM5X+FEYWwgbEOd6MmlqlCJE1nuh3icb
NEJRcCY+kIVRgemiBn0C0/qPsUQF0SCG2ypjNb4/VYwwmAVORPvRSnlzkQpt0rxAoLx5xYJgM7Pq
MMuEg2vo3mypwVDZAKdwq1aX/s2VLEJrgBvNQfqGQo3raUnFVYyLfwC7+6aksXd9IP1vgimX9EfD
Jg/lOKaOMCYiUQhlWHVaUaQItL2Py2QR9n/Rj4c9Vyp5UKk/HRprCgqq9fjX2mMhvzM9Wa7FFO5V
mAbEcOIAV3IF2NBUp2qGC3jeSw8K4ao+fsnnWwFr8fhJ15kHz2u6z5Hj2QTuLGgCOnul7+jc8nFQ
JAC5Wp7Zw2yuNJgi47EfyFzG8agkl+rxiHk/mpMT7x2tMPDXenhAr+Eo0FSwPADVZXpKY8asdqda
eWKIzf382cKd1lKuXFqeuEkrqANj09Jf/r6pn6LB3MR3PUvsW4IhDiQaSgpMo8tb+wxOTfyoeh8a
3NhavueLY7rTcJEzkYOfJtN1+QIqT/LXVWjaC+KPKC96TFBCjh5PcEc7IUA5RBiH0sn2UkRzmAA9
bhuWKQlwnSL+v6IfemKziJDyl+ql5iiLRST3EKhSJahLSJrvGevqw7414nWUCO2nY/dj+NSzmHqf
XNRGlVZp2w1Kl/A1oDC3GDJFWw+R66NUBZZhHDbX/tklZi9kBRz1JCSAHMGywzl2VFWYvdtwkgKd
/Lxm6EDHi7sBCaCtDlrueWqn00QEp8Qq/ASX3ib/rEjGqJuFu10jqMmRZK5wcDg3IORgTU0+gegG
f9IPKq1QkVHFwPJOjZSVSPVS47L24UG8XRQjNDGCzskj+MVFU+Q9zArILmLnVaFw6AFhXUSTOQQz
PNJVJzYel2+oiNBNwwQ/ZVZoLyCzPC9grOXZofqxL4CxV1IACS3TdiYzh//DVOe1qYEIXEC+qmul
JHYi7hKXrFGzqfsrM9B5GAfxSWW2IC4M2o7ekliZ1kI0EF5qOJAv7nz8CwIpXWPTlLhvxYAfFtlb
cSYybfp1Fy5Dx0r5m/Hw7i9gnSGCQasKFc4xO3H8wX+3DHAWtVv+1Juo8oDvzmfL/V5yCiTtrU0z
1JKc7+vBkwTlPRUcEw3B7VqDOuS2n90svXYDLX/G1wsPxIlRJpLqep+9YlWqxNNKeJ6X93Ww/ZOY
yxeEM43B1XEQ8qozJny5TRFCw3etF7F38W0FHq7Ncpr6TFVAvrv6VRbIDSpTtEXEAJ/jnbgskUuc
OGTAvvfxaI5Oa5OrZTuWZ4zgxV1gWn5xQ/DVjeBWYJGlTCPQXQ3Yb7bETJzpysmzBJPIBGEyUOVl
fhYTaBWRzz8RWqQq19x4c9JTFEepcUeicjNOdj3/8DBL4QhbFOuG7R6GwFW83eUdc5G0b0/14y9H
5/l8CR5DvjN5t+WkItnw5kdkWYEj0WF4hkWvdas+j/akRbpB5B3tfOiv6f1XsOWcF6llGxRTPG9T
NjRmyhfT0jfDYVIUXaJZRPYLV5gKVIuqGcj8BbfwTmQbgDAR7x6d6GDOoJZIBpRYeKUsgY7bSQnZ
PW2AErOaRrURcAu55IMb2rRSUcKeI45gmJ1/Y0O3WaAAQWDy3zEbQS0b3qlx9doHRajjt9Riejqe
cwU84kQJD6+6odihPwetGbxNepGk4TYrB1MkVn6vBLO7GXL16v1iTbk7bBfrLyBQY1bxJlzY+6V0
IJHinTwBmtRAdUf4dKIudyOPJoDDZmL2NumPsZ5RhThFriscdIxuf8wdVGY4b47wUX9KUiH9ocV1
SvrZEiIXMZ/zJivganODeUQ06PZDI/7tI5ojS7XpkyG2XZB2mGZHOxD7qeDOxNpI1W2RMpE6tBF0
8M6W9YCV+kRsfle35nHl84wTh+G4a3sZO1WMyxaKS/R2oLRdP3lonDd5DUrIXoN0BeJuB80zTvph
1detvv5kbzPU3hFAdfpNU9Klmoebc84YIv6XEaKEtZqDg8qQ0iqemUwAY7Jv7zIJd2iMejEQXv8l
X8q4O/YdYVkCcbLqXJBc29R547GocsuvQ66TnmkAHrxaMGh+HUFfKj0PWnVoD6oX362cP9oDmaIp
1LILTr27AzE8bj5z7pvNTJldSpVndI3RMZFZyBBbMtm7vdJmGOc4aa95D0cu1OFhrxme8dofrPx4
zy74a2YZjQU2tCWj2w8rHPAo1scO0uGjlPl/eScnGYYMswSBPhMeFaGadtiYpo2QMUT4TXxzm19u
0QRIWvFrrzsL48pf/ON0cbW7uju7TuZr84LuARrNtMCZZB46vBVL7uDP3Rl1ZzKUymJn1RpyX9gX
LIdX4XtfdNGp9LWBZfaQiK169ezs3NrrQ07fesJq8ywSjrWqr3Ip5KKCl/3SuxAnvblqzWBquOGD
HGUkrXCyFWJuMgroaAkyGhZkrvjK/A+m2iS3T8EkkYLbr/N1IiC10blzr26r/z7/jfmRocN4bX5E
6zCnQlQ5poggvtgmAwiPErPSGKZWiKrwTmTt2AMnK+FTiY6PfveR79I3RAbWARvd+wanrXBcjdts
REbrzHRuysgygncE3D7vDBKq5JMMeTi6Fyc+8s9l6M4RDo6JLz5XTQXzfl6jQQZDYT0VMOq877fD
iFk5XvMBL+jAnkrYEbJPdLlVolaNbpbISlEorlNOrF8nHhQZEWVc63yVQuvPs0uJYFKUpdEfzcmM
hHcREwS/UTKVRRpvSgrssfJQthxf/TscyTpAMCPX/cBTgEM6F8zCKFLx1xJPODAOuSxuSmEljFQh
BaKh9zriGRJCtaFsz26S16pB/uz92QlTjmtziaXZzHko9R3doyLJEiQ29vm560FT6q4icR3qhkgN
EAWqawCNFLOwcBqSQsK62etf29H+7CKDfKVNrl+QgjBYLF8tOgFcx7NDRDGv36uFDwLmvjuwBnvk
ckp2PxxcphY9d52bmbFekV3f99sa8/lqu2yh8aQAb/yiSe1gzL6CR0sfLvBd7oy/RRsd60V8k74C
Ap2l6n371ho7Zqn9za+T01IhB85BEfmAOglw10mFYXLB0fNFPmxB1l+JeugVwyeVAfifNWX6Q7ku
kAYujNsmffCfbmYo0ry+ho41B4Sp/adci1DtC4LmkvahonyfNMgtlUmx8OyFtxlEY2p2pAfN0GvQ
2ljHnHEbgwdtfIVxdcRqPjaW/9EPpmWwblXVmMRWKUQLOkwScJjMUdjzZ4HsDJd4DAJxYH1927pA
bj9WMZMH7bANXT1jtbvYtbAYF0w5TOTmejdO1MVrIQ1RNhZmhqPmWLfu4jXG5ccfzuub5kJa3CvV
H7Dq5W1CGSyADsGMyhsgizyJGf437SpLZ2ZZpGWp9KP2xQS0x3SoUINYDZm09w7cu+t2q3/4aT7E
o+FUnlPBv3v7IWOI4JMNDtgMuDCD5UOamJ7bkECTKB/y28HgFXYum72mdiz2j5n+9o++E53IIKEg
uLpV7rK3eMFsHJksi8gkKF6J36mvoWJXB4C4M09ubMpypT/xaRcs6ObmYbiht/MGS/JsaVkOiEn3
CsWLKhewurEtZ7COihNfy0EBI45pCkW9fTHls3CGOW10xwJ6nZHLam6mNu0/LXmjR0wrBG7TYzUC
ggCMkwYGWNEhsTr55CaK8NNIuPtq/awnpuUttMIbCmdFc6fOZq9ppDtu8bH8m6A+asfqJJW3EGoe
62TrlZycoI5ljV/QwcZXoSb5UsbH0S1Sz6z7BH5rWhDnQ9smtGNm9slOrVvSXxV0k0GxU9Tj1/1L
bfx4ySyoYlQ2PltYNmmRDPZVZlLaPOqHJ/IANoAdqFpo4OBhEp7Ab6OJGhCAPN9g45ykSPXz06aG
7fzkVMireLaTjBz60tC37js8iXJ0Z2fbuODmnZLd8H4BhabpCQEJ1lRkcTnG2B68CE0ttSD3Ndf9
LKh2uB3SueE8u6/zAbQ1j3lywCB1VIBWBytf0ZqjmBt/TXARQGPcX1yzDvbsvV9PlzAj55IvXLtI
VsLQ8W3qAr7/V0gTvezjCOAryc2lAH33Xz0vOmdCUEVhKNhIo9NT0apaOOC87qirJE8fNNZv6Wh7
lxzV/Pf/sLvXtwX+5z8AC+d+Yuckbi86fX94m0wXn6GfXICHKmpuC6XwWszizpeJYYDvRtHNmVWH
1EeCoYlMznN1u3ZG8LzIu0a6ZaSi0K36nej8lMIqjPz7CNUu9nBlnpwTfAwfGn/VOwE0ar/1yhli
HXNaDAo63H/0+/2CSxsCT2j7DNAiHyHH1h35VqajLZ2tzYLHDzlWc6RUi4qC/LUO0BBFz8gMo6nT
myfVG3sAibnfqp6+XUvgiZ2dPcBpWTfKMAGQisb7lFC+qSNoZFPdMTHSp3/h9UXirA/KiIu8lytB
1m7Bqxx7Kj5wuk1vkuSpFaA98m0NMpsL866mYd3FEBY72pp66IEECqc8+A6FkZ2ENeSIbr9No1Dc
v6AdwTdR1bjbjWtOe1bIYTgfZsTjySTuT9Y+UdEOyyicAaiS0REAfgJmgq9vdB4C/f6/aQhlSA+q
1J9bNhntUwLcTkTsu+VwuqQrX8LBzIzV4M4Bt8g4aqNP9DjsiAIX9Nh88uWI1jBkdiiz29jLORJ0
Vq3lgFL7/MEgB4UMViw7QiiRHh+nq23Vzt2L9q+r8TMP16WhWj06AdtRVClAhJOWx2z0b+P2TPsN
6ebWXAOrtIuC9EwjcSjxiTKyLbh10ESygLW8fkOK3A2VBnP1HWppxezw6OEfZdDCimRs+a5HS6KM
3doeJjv8mTHsrauL14DJca7oAs54zjoEvQ0I+M78ptbvyc6bZLYpiQ1deWk5Br0GKJ0C/chyBRwY
/iyfvVhtFw4WnkxSC6VQXWfV8QY6/apotuSBbDWDH0N2KF/KthP3JIMGktcEyKDNJIUf43TozlT0
hncXoLgvo6iO49/EjC+oRaMol/oWTFdXi/I3An85vHCzeU0Rh3onyfwAVSUlO9Qu4tntEKw6Jv9H
SAsxSNdoY9vz7GnHmTIPEVyeR6edOw/cD044Zq+X5whrDXp1BjLyGG3nh46G6tdLLDzIn0Kp03fq
MD2dQqUHc9eJgN/MN0BqvzBrlqDGfEAFfdOSzlaP55XDcNvCsl+eXPJZRtgLPcvmI9B2YxH6Bo3W
zFimadJ779yRpECab2/WD/+Js9U3ngSvYd/lHjGXDSLvalf2wPt/gY9R7mBwS/pbeb/ZnESkPCgy
Arn4s05mIKbeYVCn6RBqjtxu7jFuM/q8LotoOblrCBsl/b+sEhEh3be8X9UTf/6tdb4bGuhnK6W8
Ejt8QcLM6oUs4mei3lrhLzz5ViAhVfE31H8yR1W2tltRpY+Hvee59E84DPZMBxU53p43ovgrt7mL
g9SRIFD680xAhOO7YTgGD0wbbwAMkmkHFhDLj3uiHQCM5GvdwdDHXWREci3xzHNOUR6qGe7+gXGs
FIv/wwCId+xLyZwRsvbxNV4lu7DZ9A/NF4+ArSYLZPoFyouvzdmdSAMEvq0XUD/HbDaInLS5Lcw4
bfQX7TDWemq4D80EQqZs7uK5VL7wwcOc/rs4SjJFNSMIxhAFuUG3IThdo/hqRCDug3HQqoqFr7Gy
IyGCHawyzbefADMtdGzh/dvT2khhdkKFhGdYPe6m7C0J0JCcQS7vcvDpkYDwBbMtkztQEBYBk18b
jCv80z5BWmUbYnVOghmJ597X82HT8GS+NqNqVnYQSm78PQefj4TuUb43qIEX8MJ3ODARofoDMSPq
as3OkK9+ad0FqxKNBvy+3BJ4Fh3CLZy84g87x/+GvBjtKR8eoLKzJGclcjg/mzxGqmFIpyvZyHNZ
8ECklwC1A4Dy4osyrJAiMjNpx6TRL2jBP2gS5OfXufl//wJDuP757f8Hp8kBCY73c5j/Yw61BLgl
oQJIzdCe72Ur/6Ys0Ik+th3OGsJcCF71qAy3TV19o6yea0CQ2Z4YDOZ+nNonpSFo3mDqAQzgyRq8
T4XFnj9sD7DMdllit0DFk8VHpypaG5ptVfkRiDH9JjnOU2ahaw0wgTMYbcRFPsObGK0edDL4r4sz
y4NFQxYybhI0PATXc7qmN8LaouT84VKR7bZcT4HrIzg5PgXl3Hs8ZWX7LY14zF+gX/YyU7kSwU0p
fLg7ZVMpoceTO7h94CCIlo/5BpDCEWa6gCUBV0Vbunxr9ijZjRvssT2QTFFpwuCpq/u9nIY/fSSq
aaC/KE0oIEYvJbhI85mcC0Zbg+fYC1nSH62fhy85/sWmGPsAEDo/NpH9il2InthOvmwzbLdR0xvJ
cKoaeHIRlG0O49tWzHHexLE9s5sPeU3+tnvjTP/+VOBlx4u7jy8fu3CzPsXmXVxkJedc16NhXPwN
7Zk+pbCJ6yzd+volP4UWdH31tD8+PJAm50Ke6E14axizRXEM8IfTsvIzUKXZ4y/1RR+lWV1yenr7
LW2Jhcql6ebWPPV2c4s3Ix7UrzTMAVYnbbRfJMOv2pfuNcvYPUa/w439AYEl3EbLXrsMrPF6PGKN
WAC0f2MsP0Q1WpT778wGqpCGmT9V847XfCj5Hn3UKLMSK051HMMrTdiJwOpsrLYzZr54a95DR5yw
/YZFZH1aZZ7D4LCGWipmGE9SJGVJSiaew4qAcp/zyBLAGPYhLBn3yb1Awm5utH+g5B3YQs+Z4RT6
Br2YdhoqsiLi+caDpCHPrAK2AOrBlMqmbjQ4P77HR/TrPVc7QlZkGQaHn8aklEIIsQtBEqFEVdSo
5Z40EECcEGmdFy0TFT8wR096qzIIOQ0jZswkJbTmQk/jB9FGE3/dNap2yeLN3nnekRZzLukQzAXx
NvWGWXlHTRNzKCuYVNS2GCXZRQRMpImf1DhbTXyyUWubIinABedZ6UYsNsg7IvvELUdgX5xntfTc
0J/emzYF2kxWW3lxxCX7AbhaoXltqPBTFGCaqCDchH7rjgMM5HJCrVR6PrgtYvuolJGLRIj6Ob4y
aAiU+GcvIuaCumPrEnKjbdJK21Umti2WtKxlmKMqdGKBulpRaYzFW4GHXs8AFdpB5JjzHC82KAks
fYuixm05yk5GOR+Sj+3gdptbU7CXV/jr8PJGI/vXIdqZznQFw1Dj6lDdcf4ugS2/WqOlybSfwyET
pRyGVjq+42m74pFApVYTxiHa2HMLB0VvJ1Q/+XKnYQtkEgFrN8114MP2LI2xKdUjj16eZNElMvWp
rEaueqbzswidj7Ma79wPzxbR/hTVO7xN6fHF8BMWE2jjIajr05kjs5J8VqyGmwAUJQDIHjbLaBsW
ucZJW9slVUALGTdUdzJJlUHIWLWjFH62OySYbEdOGePsYCZWcECJcMX+c6rF8mp+cbo1rgECM4C8
fVhmfjRFD7ZZsuanU1UVQKBm1t9rxoihNMN9djpR8q87bV8hkyFe5n4eGQxzrQLCPybO5BzIR9HF
aYK2ZbqVZMHDvFdetV6ofPVelLKXUafbrNKH2MfQP9PwnHl/V2kdY9ye5GyeFYxaER0zhBcjtWDn
i1u1vC2AokRIu6+WTjZAzJHXwe/m9a6ZoASWTj1kyU2H7X5eqWU5yUT+rj7JZWXMGQCvMs2WVYRY
Jaobenl+6yALgtRTJ/I5JTDFIPD1TcZXavmHRm9+2mc6znHtPbaLvXHOE1I4w2zQegg3irUWsokT
UALlxaPqRQ0JA2mMdO/YrCL5LhHZK7Xp/Gdy+JtKJ2cM+010+q2KhhmhQt4TjXcbXLuymGQ/wCWZ
0huzIZNZZarPSfm98pJbxZD61iv2GRc4+PYVF4qaXOkNvN+UpZ9tDbvGJjuSo9p0a43EDJmnbHDT
sczQqyM+wxlECajZB9d8unQh2zxWQrjsA692VDvnG+CB4D87a5BfvBxr3jLjP8rC6JjnfvpNfyDR
Jf6CqcZy3e8cb102eIQU9kL1Jt+t7TnuPye1Hq+qNzLe2NAbFQDDs6tCku2BCbmBd/Vu17h7ht0P
Gr4DiLl6Tl95DkFIWadYyX5l9rLivNok6rSLrXEtX3XBcArpQwlS6o8JWYUy+EmggMH4ez233h5R
ill6pTn1i/x/7b0OnEHmKEKQX8l2h8NrpXn2v1G0dtmKoiAZizMFi4fTkme3uNjWZHhZafCJeXQr
9OtQY9hcRl/Rlu3fUDosQAw+rYQ7+hYCKKz8VRZF9JHIJr2o7ZK7FECkcFAu4nZ+P1yJBs9fSgUU
Vm3Wz/8il6YvFzJTHeifW7NHSk8AedZMTfSKLDofyiFbqOvm2a+vLhIjV1XgnNSjyxmm4ZT7pzFF
5J2FzAjNIertcuLZjvYUODNaUITxBqbEq2TFZWEMZFFzQ8tFMDnTIVNB/C8T4BEGhc6M0vbRuz4h
9OmU/eqK831gNTS84h5oIqcMqy556Jp9HR96iXyjeeYJICE7yD+DBWajKqJZn7D02ZqUr8E7a3XF
DTU3JnQowSdjvlx9+65MVu53GjSjQTwdXSoUK9pElK0bPaqYYJsOIOZpuvjnjwbk3f1pnJFFt9uz
2AdA+WddrRMY+XigNgQ/+IEqHNiAOCtu1+qdhfneJKv8gMOF/2EsdsoALdjNzWZlTtlDEbYhuSpx
QuTA40avXN05Y8U2gb1bf/YxAmkz2wLICo0X2pBe9OI42VNBxIQfvy/FTS6oC7Ai36BTPxDi+3kT
ddz5UvEdJ6WAmwBOOZ+/d6m6lBUkb0bncKkm9Dk84NrrstBjNWsaX/XZJYNdzO5vLpuMUPxba06s
GNK+ibbj50I+QyMsiP1xk9DVTdEantVNSLUrhJZpQi8p3ArHfSNDqdQqoYceHeWtdlFzoeWDubxF
2Pvv7LBxj+XBAYKi7PW/2lFx+yhpeeM3vEpCIQpwoN1hk2VyI3vUw17TToXcsfLuoU5EuQqXRGKR
FZQHWYBNtx12Brizt7gtW99KEL2olvK8nO0Fa99N1PyI7XWcJONN0p9JKKAx8MMUnHda9iu8JlmC
yw0ue3WclpteEfnJ31d0R25jyR94TgCaFEpyv0zTVvadusmmWHpxcHBWA7fyagtZCIFSEvLnGriv
/70KuZkIzzbssf6/E0vymjmwgYMiNoAYjQsAx8VkDEHzyWo9skr67cqWi/35lGoVgSGP7IKabDI9
favuWnfvYtZWktcPEk64xDRVTW/VxO8lphUsyRy8ESAwEgv0KdeZ10Z6fDdl93V7vPvmHemlqfxw
jbX+ITzhmjKbu7jZTLnfrYlaYCdOaBAWycQ23b9zqtzX8jWAMQt2XA4AV3bCJdphaSZP4zikxHtu
kjEUURsr5/gR5O/yCRdsVbHN9XuPTiKEQUKvdSNpL3tDGVx5XR1LyJY/7dB/tO1klIAm7cUo5uQ1
bmJcTnSrAWKtP9M8AnWPtquzGxMlqchAH9h9TTqqUdFgc+UhYyNHsccCGFUV8ut5vv1v4KQMxv6h
VJZHjeAWxmh03ofJjyttPr0fiyMR7zhXcJAXMYBfXc5xAs0SAhUSRG/qZXj4tsFIveNx7Bu34whU
aPETjaP3sXWx0MTd3eQuDHqT7PsCtePsHNWXmOR76m95Ref9d/2j7kpRwjuRIhmA2XcXT4aQ6ri1
cvn4nBJpYj33BtkKwBQ1YrXESflAwbNmfQpLVIglWM4H81bHZSWRWaw9Lh7a/GvVgvTmzZ73HFk0
gpVEFv1sA+UCTCItVpgq8AaBJrtsiMlJhF/WY0jAt81JYfgrGfShl77XisoPFx7/mQ0bYaztj7iX
/PwOjnXOiNLsVX4h2Gi34S42U6zUeb/rSOEtn+m57+l8zt2QFLNYvcVb8FbEHAZO/cJfx3GWCfGu
OptY9mkTlQ6h12adSbJKfL6gMxQbdEv+5gTapKKzJMRPGwrX9PPFFoorFZa5lrfOYLFATfugIT/s
86N4vWOT91oU8qH0mIXPJ0Ysa8gbWHzPoSRO5LBmdM2e9hnOXbnKKQ1th5HtO6Gl4AJeDvu1yR7v
sK96zj50X+c7osQl/PXW6UMEUAzj2qreRv+J991mkL7WHlyaUJR2WZ4kIfGORlaePhOBFAI/4ddu
TAhaS9A7X8uF9jGATQ+Pp4bDsWrRqsUG5oQmzNpcnK9a0u30XZ7yYvElahlh1Rp1REXa4xU0ksDD
HpHsKFKIjZPvgjx9Omx17D3mDJ/QL6Mk4jL1ZsUJ2abs1qKHMVN2qImVHUlnClb9SE8WteVREVpj
JSIUPiOv37G5pIblFqVKHDvS8bXJV1ZSEqULpUj6TXqcyQvpSBS88PwNuSl43ea+lvQkRYP3J6s1
2dh5c4tFhzrZa4OVGxtjH57WxHzSrmgOaPXqhBC3eoghQhtb/xlG8t7pBaZHAK8rRHPJwzCm72mR
eQQv7J8BkyP8DSdkWTlGK9UR91KhKQw4YEH+gKcIUTqrC9sUuVSzuvB+7VmiEID19MmBcE5wOrc+
J29V4BU1+ybygUtp5UsqEZ2Evyo2dLBDTObnQ6J+CdJMouR7YGNNIGITbloLLKjI9gFauklNZXKC
taLJlPURRT/LkBYwynDvF1mijTfyxQMSHT+KCcEcLKk1UpaPCdljXR/JvQGZJdsiOKFHVGR4YGGM
1vN390qiB8ab+Hj73OGp3u/WET5AUCe6NN+2vcO/Ov5HlJn1RkJMKnVn3eSx2AgVSJcuBK6kawLg
PB0ep6jwtoz4Y1YMLsyInG4PJn8JXTAC6dwKcdy15Xv2Ub6tl3Iwyyh1xmgZ3APV6Vj9gf7AtM4H
t6EzRG/xs/1S/gNnY9slPbBctE1fcFfvY59DYp/SFpa5XhqC/4gwgx9uCPAbUlfYqSKXd0J871Xv
2kt9/VvPHU4C4w3kz6O7L823Eq9pNCoq0llsXhTGWIR6MjiJswyRRqckciHJYmhQY67xAMIPang9
QMVc3nfxeMnMKfJ51movxOCkAUOmhVYX4PdY2FgVhoPNx+RHHmf0NXwVS6diQpjKEk9ti+LQz5XI
UVqBis6x/bCRnCl8lv9BZp8JyegTcJvjjCFCdUvGQeZO55FxaPjIXif8megXiUJusB5uvkYze1/v
YJWmayBQBAmyso6FTwUhGNNT0Gcz41HF76glonml94ed7+WeRnCufpwUzrPdplQ5nsnHtz3wfONI
0ouh2vSWMVOqYPaihBB+UhSnbRuObiO2Mf17C+Rzt98ucHpJP3td3r0yd95Or0H/H4todlab9Won
BsaEqb1b9/UcZoDksN7l5oSchbVFoY4445defV3CuolAOma8e7ISB4uDs5flxKQWyH/dHEOklFAh
q05ylHIlAvXS1d3vP3/nIny2YssP31vM1XvHySe60yKwnjO50oVvqkKKqFBMiSOQj9U1nyTPzbnB
Szgb+SIrK6algIjlx9VbwJAHum98ZpPcMPPom1Y0TzdgtCYCEJytF1a+AISWYd+pz03eqpBGx1Ag
IafYG1HjTViVPpXLSPfk/iLUfzock8+R0AfysV7ZsOup7NldtqPchTxn6TMtpoKwwTuOR7V9fP/L
POb5hD1x2UVFiCURE0bEW+jNdIdgdLSSpqr/FXs6f85Gh6Wx1pDPRxmWFOpfeed7R3bPKoHsPcAj
bC2ggfjvRF3Y0Adh9JT005GdXPmuODc+uS0riekk/2j+TkZePeY83giZn3nPR5TThOFelzdhMKHY
6srvtgIwe1NK/6qo4zM4uAg/yQTia+I8OHcanCcJbNcO33Mor24M2/O0pGQwSnwhuWXyyMr2bRtv
tniJ71mMVt9CUN23vTCU1HHbv3j81UfO9OYJ5iVhKxj4VaLAyJGSTbx6qy4+oV/lpvmOR0tQCVZ8
wh1kaOJRzl6qREh773p7j7CoFKYhuEhLD5jQCsfemKfoFmzjPACbroPmIPsZ5VxXwTOGrU3ofTIP
q9nZur45MQXaTL+1nuT7MoTlEgQoryZg5irBhvfT/nLRIFEDsWDp2XBHLvViYiCpjPeyQyUqGORx
SgSNIpUAa0113Bmh+vSdViBVt46GKeaHeqGMMTiTptDXzUanLoZX30OAvKx/W1Ns9iNmCuOTdFn/
WgMQSgVsw9RiGEzNpd6d1kwcujRDBA4NXiTFW26gPidHMIJMlPh57HRbmBLEwfKZ7aNVpD/6E4Oe
pz9NB345IFBmS3rmAflGi9UZB0317v1y7r80y/naSoA2HsS1dieVG+hCefksOh4xYptS9IFUS0Ug
Plwoib12fWaiUBkI6ma1UYDndsiL4TI8MGcEaN5qNu2q11gqtr6YMDEqoPmMVlJ5puR0zW+lFzce
Fn6+NMtljE2gDBLmxr3CnQwwZoJmyn5vhmbCcgeWPvgrJkeH6sIgRIG6kDag1Ob6kmeLJEaR2h4h
gVSmtno00a2cIOL95h5Ee/X9LORSR0Y6dRtYMBMvc5SL0j61gtpXuwgvPoAhzyKLYG2SBQf0yMI/
1Ovl+WyKlcCyqsoWyfp0xPrWZHsv2NUTl8fQC20cT5OhlYeFtxGamgKvyoTYdqi13mFtVSrmg/R4
yCuwzphdWwqs5vtShHYVKRJ8010+/6a6a/hs+FUzGbMet4nf8ktN8WJfDFEEn5WPacb+F61eEzXY
UGxXvM7ASMTvJZfQ+0st2XrhZwX+QpvSmLK+I7D/ZnOFajfvzDwQdw5pq15O07aw09Y3pJ//NYaV
2gSQitXfHcE1c5lyYQYTAGbgf3bTglDPWhh41fqCojwbtitFzp+gVbtodRn7JvBPDok1yn1uLpJ/
9SAFhhdiO4jWrlxR0zJxPZgADP0GudqykUkc5LeViUFfmiROeaJvOcFlB+fjd0CUtieoFVzNlA5i
iEzx6B93xridbFgUllwN+woa21akmxwFNSm+tQqfZd2BNlAgySLkI0ajHNbEvy2ClxdV+d/juteV
HU5gK9U7fIeDvFB3qKfYzmL8wdKNNH0lY+VNou3HZWT7XwKxe15+yCvlhPpIuNP1I9GKGmBozhJS
/7+KDwfGhmzm3GPz6J5mMPvzA++NbSzcJIRu7UIr554zdX18JOcQuWseQyYrVNQVeW4DhDPykPMs
6MvBFBF63cUtN22pn/67ilmZDGGDXrzE9frSNOz1YjtCyGIrlvQ89tUiYp+ddNpGmB7A+Je+sdny
OIeWPCir5bm3vhzaGWxpUD7GZeSQzDJLu66OOeKQ8e7Uolcb+YR7xuUEhJSPLXRRZ4LnrAELz6IK
kPu9vqGC/nmQJUSF3i3TqD+IOF82jXu43tSRIY9Nvd+grZz85xCMBFWJpeyb8D01Pex/8gJFXZO+
fOMEFhNZQNB5hpTdkS+CY3lW7zSZI5+7fMhFs6LGCn7NDoFzmScMwAzbw8Z6j62ScAjjJM0sU+dM
FJdr4x51gCREFhumwiIAuFgkGT848dTzuzd4iFdLrHvFDezezfzr5wjvJFDX1K8PCaC42aATNn+o
EA8jCIPM4kUVKDF91D0tz2haBdlNahbCqEdcfbq3PiHJhANXHPJZiM9RlsrAAomMe4gUDWtRO5Hk
Gis8QeSEy+SnzK0hgfn5GDXg3k1twDPpBXvSPJy5ZH9KwDW3mc+QdyOrE8krCl1w5YDPjGfeFhos
G1ef5TXKr2T9cWtKk9s3TWVCQCrcLRBu+KwUrux6ALejQkmTAVbGuLvFw+9gFjCIjMTuv3+p7moT
JyopQDurGbXhffD39HawcTwcFhRhdGj1XoxgzhliIANYZYqSyK6IWGiymb+c1+7RyDD4G7gwtcAz
39UcE64ybGMysJjonIe+NiCJPNgYcaHjSwr56SE3xg/Ta+dlOZJ8b9nSITAyqr2RK1HBer09H+eQ
JyqAJ0FH5JB0kJBq//s9rHCqh8HapYgnitWx1cNRVk0uxx7U8j9C42XTuSbFaE23RoyEpc/6HjTf
5FrgDcXbjs5M4shzzbXip82IQoWNgmLpowDjaY9OiwkwT0eYA3L73sbnc7ZIrQlgpxQvyWNj0W/N
A80h7+6MLUgK2N/uH2rS5TG7B1R5CO7kgQu3iiBI4a5mS8QQqVvBp1sn3DEgB10jH+SIHH7NqyeP
X3wYdu0dcpADpAfNWpRj58yTzN9n6bcascM11qxcZUH8vwqu6qa+MixIEeYhPiZ0/Ee59rvonx89
C3mX3tI9lTioicxZDygvRcubK/Lh9D8zLjMyCLPv39W3dsVf2JZSj+UJHtwTy7oVcU0hKeL3vI6R
2SGKTqyb+9c7SZeU9FuUgYw7tG3QDk+h6vWsz7d84TP31MBRkWXv45UpgRHvqy3OxqMqlFONZOgs
j8DC4ey8pwSC03NGWwe43khEv6m6Qi1g7C+KKxqG9kdaon1G3xOzDLfc1d43g/qkCKimLK/wO1c2
p8tDlszbGXoG/Ga/haodE4vPF4QMIeZX62YtSxVM4vOsBpjdStKzQNYOg3f2N8FwPFPPLks5aKwu
M5CEGiK5QuEtb9E3LKLCyqQvHZKTXMEVO++m8rAL/un8525uNj4eLtPez0b2PiVO6OmLrfiE3S6x
vm11Z5VCnIR6n8b7+U7j8AlLprsKFbtVq879vwSCBDv91z4hMDp69jDKz8BpvG2NJlpu0/wCpn3R
6QAjuYpfWtL/boAspDhNmzDAQMoH2ssSA+9HcTcrbG/nZxeTKtHh26w4+Se3GKeIDa9hUT4gopwb
dvlkeYStBFkh1BbYahmjjfNBiWkNCy2i/sDsrgoZskeVJI2wyEZS2ZKE9hTo2r+OV4TXgHHgO44s
MiuzcYGa7fAcMBSAzGQZGjzGmmlHS3uSgOUcv0Lli2PZh4i0WH60G2s8WtjzfQO9vFIUk9Za6RkP
G6oHC4cGnGiS1puOQDkcFcPPOFds5ZKDrOgxTVvHChIXuJzS61MquFuhNFRVobVglOtU85qFbsVA
SPGL9/Tbe/SCsqjlAVT7Z6ht+zv0gs+vhC6nTUUJFK2keEFqjfhoFRT9zwEJJaLnjSqIfgei0bKp
10grGjnLscSChtr8TdI3FVLMKeAZ84++Rz0xXlHbYKN3dm9KxpR6Pu4KYN8IrR7W7H43yEvOTPmc
VSVI/vQUpBrmtNHRqBsamcm2JHzfrmhYxqQbSy3US3jMpBZxZpZMoI3muOhF2ucN7aFbPwVJQpdh
hX328/g/H5IODPfhyVT1TwZnar3l6A6mp/3L1ECFtmu1NU5wrQW5K80UcX4cLbRMvTd8hKvIkPxi
fEyIINj82VNZmv0oCdw2/08rcoEixoxu88EX6jGka1lD1DHfsYtaZ/k4GPwbv2P5vQyVew8zrPIS
YIXM8nJhm21gdd2/Pf3orbjuoSkmCBdzSWAk87qhB23QXTI0XwpJiYcgLoUaA2jU/srq5f5LUZAk
Ncyeaq7xuuNOB9+Fh4SwFbswtZAP6GzfAmGUmKVjEVkV3zwU8mUL6WLoFAUnlhZFsrLHbu9p85Sb
zmAXcVVeQoeQspH3leH5MhjUxD/KGjwVMhhjrLygVFLvEz8d8JpoQ6g/5lXxTULpdC1RRastThxx
pFsmyg+TtZLIIE/RyMEA3fYB/hohNJbSN1168op0zUex+a+xh77ig3VN6DWehvlE6NPUR9sDyz07
KA3yZqO8lx6G2UdozoL0Kug6CYS9XpteNVq9tZXTtgfGb7HPlp9byFTp96kiNmT4YVnnst5nq6Rn
EtKFz/st0vf2nnatoe+4KgF+Ko05nkfHI1nZQvoOiHepYRu21/nOP857r/jICP3TX/63Kh6TfZLr
n8cm1yJU/c0vLCY6oHcWmmuYetd4M7BzUQqIzmzBKdJb9FR0Os+NVaTY+br3B7wvqQE0HQCUFkg1
9f9afh/nVTgXFJnlSmlwni8my1UkNEk8vHqcpXdPwvwkL+mXcR2FCazeYVCITKq2A/pjioJ3d9ZL
PD3dAiPN5nguZ8t1+O7ovBHwXrTNWFNrpWY5kZSfXhC8IUA1ZjLkVHJlFwwId48nOsdhnnpbHUoT
k8Bktgvf1gb8ph5r+qiPSn8iDXDK+KmMO4b0n2HF+3Ui+X27LU2kDYcaU8dOVJmqedpb4w91nYy/
dCHg4dezuW+iYWPSMQMYU3YbHuW8u2pEc2gTuwRahEr4qxlV61WdHst3ugZm9kM7TU2AXiTC9vRb
NJKeRSOkELHA6txvW29KLvbd3EdqkQ7Ng0uanpHSnooKYj6GG+6g5Bkon7rCKttXasMd3HVCkQ+Q
v0bnOxFuxMSxw9uj8EmTnTum/gWfQr8c/UF9ZMgd1J/emych1/5zmTM1An1b+qxcLuHYpnsoupTp
MC6VN2/QYQ+qBxpmyfeXw1X+WRn48ngObSMsQz7QmB08bG6zmRqQ2611wA7Y0Xk29H5o19TyXLAQ
Ildxb0cw1GYU+HtgyOeBrtFJ+MUwBeya7BIdDAB3CD47tKb5BPSHEi4pNa2u8EQePw4/gF2cJ7zb
wtRXaR982KUcN4AupjTdkUEcfSYwPv51JJK6I8zSNHBtat1EZmT25Dl5ThTJyPmTnRRsejehmlBr
z1HUqU7C5mRh/a7jHQ0YMJA+Pv8w28l4XGcqeja8TJnSPQ+EkCCX/TYPhuG9MxwVKOMyALxEyjg2
HUY6eZ/a5g8qaD2dqmRZ771H5XkQq3Xk50TiNTNCwm44x2l2zuwcddXnBSuw6AUMy1aQIwZR2LMd
P/y/ACw7FwgTeMGwrUm8l93gkYrnTj25Bi8+9wsO4By8ZY+ihJ+znzVlMwrKsXU762vHcFIREx6Y
4HHuWbbLkgGOycpKuFCqjZ2ByvH9f/uvHghrt8JpvS0JTB7z6fvCQ64o+S6xH7vTnID0ANXYx0yy
yMDbBY2UTNrlXEwDfCI7TlUWUuY6IT92GY162ardgLZK1Uyt5Xs0nlnLnOyZnudC8TYPMpcKCPRt
oevwFNH9AiRQ4j+5W6RUlbR3V103oid11P8s+3z9fOkQ537M5INldBSSRunZkEFWKFOinZav+App
sS8cSLZrKd2kP7bewxEAZ4rG8tgZiQmNdFi28liaMDOqoAGXlV2oG1acIj1SwpzSlzRicQ1IgLHL
gmpODkMjo6q9AVgi86mMLuhgHf8/eq81+pV4CoqejQNHbXW2cF8tXM/25OIvjjSR0q+azw1LVPfq
iVs0fIYlttCKx9uc7h2QU/sA2VitbFNdF2ooLiiaiGHTIJYBllVeCa9Uvk9meNF8Y3ac4Dp3acUh
mBazbHfehdfqxdWC8wkBTMZjykXhn8Z8mj2inbvCJ9UASHCgbN4oulXAHu1dAuMHJZI/3b2Hv/F3
7XkE0/MLtF+ucXhmknodABBNZ9Xc1X+6X2TILAuurMnzIEoGbkU4w9p9b2tBwNaA1BLRa31sDe5Q
x0+JV08gWcpTG9MO6fDMJzfM8Gf00g+X4cH/AO+kr8srvwDsMXns/S6AChjKo4NECLfh6tExSRAt
senqBMy32tzstDKQRTBy5xjGmJ8OF7wiiUqpmZ6S+KJiAqDB8BtlNoWfHa7rBB3JBbHtDXGP4VIT
0Rf3juwZ/h7NrcfH9rdNNRKHezdtjMik/SyQ44nBdfIWn+bQHK1aoZo0nZFrjPAg4XMGWdwzhmJp
fVJ/+ck7sVeUtnzK4kXgi5n+dw+c4k9uEV2WneqxhTEbtsMAfaKZ3zobDrgiXgdfUy11nkzHDWUP
WywmDjQ5StInD6Rz+ULfPo5CCzDzqtaqbmSlPJL/VAKtUVEIzChsGkPX6q+44W25tGi4xzdwZNER
rCOLLatb651GO12uuGHrOpUU8RA8zcurPiCbtr7o3cOvMB14Wfsp/GjZQlvdB598TPV3TEtCaREZ
YDOZ2cVxrvQZ210ure4L4q6kbR78sEoKKy67ba6K8sfIHVfx4N9FGEa2HPUyccfJEcRCj9JQjwx2
k2ZXMcYoZOOeVmXuafWcOmkxq4Tg3Th2p2oxrj9RC/0MMueAdREBbc1nT75cfn3feSh+X6nVBcLB
lTZhfMhg2/Dr4BzXdX5VMCVwDb6FVR4hsY/SAD+fGY3IueYIC9HGEiJtsVJlRvqsDrKg5kOZnFOS
JNHlaTiS7Gxb6xTo7OD2iXdFB8M2ArQYt50oaim90LoxojWcy6Xd449gnoFAcOpZpXwT+ByTbSV0
IVGA9bHhpnPa/RSyJp4zfTJDhRW8e+weZM0Z2KkTw2iQbNEfIEYcvqyiKWkZkRtUlgyewNE2os9k
WjA/DxibHjtWU4lFOqA+67mig54ZvFjCpBW8RLu5NFRhxnHjNTguDnBI5hCbaFau0lqY0kiw0Mlb
Aw+eYszq+s6Fq2p1rpMETNFRZTw6WmmfloPdv9mVuZ/i/V1I2d+T8pR/RSnbs48Sk0286C1So+cP
6lNN18HIxqEGDrUF0F9JDWd/lWSzq//ZXTtooOW52bMut7VmGq9gkpD4/4SKEY9ekFS6UJYblWfI
hvuwmwjx4DTnUuE1HQw9ppkcR1OdQnXhqUR2aZbuittmxnElseyHlbcurYw2YaNKeWzcfN/8RvD2
1JZXsOV97UXEVHMk94mt/qL+fNg7vHQzpGCZ2dRb8/HuPEr2cB+yOgy9RLQ6Vc9eNrIgf3xuwSfm
8ticISoBVX4mwiU6AUM7Ds/p5D5dTXkeVcSEfNEJdub7Rgncy375RvZyQa6uJ2SnIcDVgDSZ5ZnG
hX2+3UaH1AOpaPUmumzmxMaln3ihzzIe8Znp1MOIFUmReKQwFirjRRm5GFNEVEC5mhfR1tpzoefu
+xuwPP/sh28ZPFu86LY4CTHNtNsqjBd4KQoGotZm/aCtSIrUwnWww6LIpz9XkmCBaMiRv+WdoS1D
LN4GUDLecpltkc0v0n3GykDXYWZUbvEkL9+LpLrzey3VJuLX250ubrMuaQpT1zOmgvtvuTTOcIu3
Mk/Asj36ph7D4f0YEUg/d47yPXdUydIqI94rmB63I2FafbLBHUpR53n+sL1IuEwMLBSJKI4dagtN
B+7YPSXbhp/VvvVFSL8fDrp+NdRq1H7PfRTk0Flyo2tms2uCPSIfx13QHigTxjUtTGoNKJsHq3JV
u+yHLbJ6dBH0LNo5SC1E9XjCQfDopMMn7fphObp+nQChGmtDKD94az8OHnJjyK+EXkQp/TgjxRPC
Z1HLZ3Q0cr7Uny1s+zR9S/sBCchqVGjIvmkVO4wRH9HlgF1p8T5Y+Fgp1Ln2OHsoY7VUkQN0JP4d
nwQs3DQP7fDOvq0w5sagVx2UVfffb7W/hlZNZ1/Sef3R0CNae6lHlVKjBXz0p7lT7vUfvBTHaXMg
5Wu3HrzDuOtdPyq4a19A/VqlbXs8ZN3q//QOec0zT9XkQneqQlWJTz+Xtj+wC8GAVJ06IVQGQa/3
rxYp8llUx2bPC/+dDuCCSiYidnL/nO9Z+HO+EHl8D2/l7uzl0kH2r/fTEwLsso5xdVOE+tyBXrDv
biiKzVdl3FVzAngi4GgAxHKfufvbt1pQfBdmk3ZGzRZ8Ak6QaJZNlm5VvwLHsKqD0caEW8xU6CQJ
kYgALc6nConolNhhid1ZBH5+fy2WUS4HUHIjX9ZqXZTvc3kttlgEBP7qCDLqRrD2ZpT1gdrdPNry
1921yAWL4Bf7/qJtF6rKvbhPJhuGVw8FgswpM2NefbYxhud4uUYgtfj2AmqgzvGDLoTFmQPRXg/+
xmjuQN5owDdiH3S4Ce4f4EeCkU0NQQBYdDPi0eP59I3/6y3g/o0IrJsGS67MsD6DTcTU7DRMTp8+
m4O8y6Kwh/u202+6zV1cOIVM+dQsJxPtnG9aKnbbMdL827HDYim2XH80Ymq/ym4bw2eq+vtxwFdx
AP/qii29P692R+jQeqfd1b6Sum9JlDbfF6eE/zl/vhxHfM0itZ/rjQu9l2Q6q+a+wflT+RNj6AgK
sWb3ALl2l+z5Xo8lRphbjstcDLFKZwHTUNSHsRW5JpONCWnd0szPF//b6qXd3Q+9ELtsRwKmrua4
TNS5I6cOOX7PtR6Lv/jV89aYJINnDecC9Uf7RcM3o7AhVGwiR+jxqm7cAKdoyf4imKD9/lhH5CcW
PZGhsiwbgX310jAUFXsbCNSYamJIY9U2+wgFT0qs/UXVlsREcL5KtVhMR2kR+4QkYV+9icVmIAdq
DxyPrPl9qhEydxL0Ds803GtzxkdetQWNEAk5t6H8/CwSFcF5iiF3AIZVKnmtMjcw2fzoB/Y25GNs
twlbOLUocRmZ6znQEzlAAp+AVC4OzyrR2reXi5ZT6wVuURF/46Mo/+Fe3pZGhgFJ1Cr/b17FV+w4
/EPOYKtm7mFHWjCRikQLVhjsdhpIkM0uctkBBwE+8MixclT94UAjprDVgwVY0GgdncDKXXYDyn+A
UnPSauXZAFdgdr5y1pIWOpthL8VpAadMeOsVKH8EEgyO51L3BW3TYWtGX+Xun17l9g9wgQN88tzC
3+Z8tgV0aQFnLNbYjwi8TwwkfZf9tZLh4hCTHIOtNKBRlqIVfneAR5VUl3GjkFkTCbjcVRzag5x/
Tp0wxGBuKASDJ/0yuKRhy+NA2YrLth359dzFQzms7M5FxJNyxWZEs/TP1xgVdF3XDNKB/ONorr9u
NmMWraaQPAL1Q4SH+D33FgmmQjKs5FzRGBk7XSxxUmMFZOAAzCdvp6aLNSCBkMGNMYCHxEOFfBSO
cJec3FkYb6XejdJ6aWzX50qWVnGK6USZElU9NBT3NF73HkJwXfG79Hj46fqsoA3OY+f3esqWmtFO
CT/+yExYa2d1/OAvADdTjlgmslkIQC3q8DI/qfZiJxp+v/bDE1YvZLrTpoyl41/GSwU9dz9hDITJ
fNlVXsdltokc/Q4U3U8EuaZSzDd9vXAYkZXOBROmQEu5ExrK6eOkGEejKCRPcLy4t7ENmSoRI612
93wGO0AsZPqXYaXJOBQ9ImPQqiDnj4+3ltcft85pD5bhmdHFPmx/QtBTkupz24sboe6VdITWHs/q
8AqDoGeMnJeVe6PwKzrBPVaLvBoj+46BKUO+3pIavY2PdrCDBy/og5cuov7YmQPLqYSFdWKQN/TA
6ALYUAIKVxR4diWunePTlIWjqnmbWq0hBD50wykNWkaXjolXrwDKmFmfhWu4JQoz/FWT7qht5zRc
YjswuBjWTpuABQqnU7XysM/ErWHNVT/CB/TteU/OlGF174S+xHrtsJGOI1kqxUbhxv9Le/PXSSOS
+WCP/n+atmy4tZmDQugBYPJ66B9R7POldgSshPS1h8KJPhLMCHFqXTzBB5IR2yG66eyuiU6viF3V
tSO2xhw9q7xyE+COYdQMbpFcJs8Zbi8usoPfuLX1toVYBHsiRo+ROtaWnLmK5KPW5Q6IFcabF6dK
5nB990fq40mmUZBoTf3byHnnqAeffBAyMD6Q1ila5KMQKBMMkysHNGvkeb0rTHY9o+j350a2pMEr
b+3nJeZImQBVIWM80IAkh7DFllLzzJtGExtbTRHTpYe/Teu9Uvxz/8Ks8wzcdPDahB/dUo3xa5WP
Ho9XFSD7JyBw8oI9p0rXNMqMYGIJI7VHeRkc/gIYRotUSzZ26yAHBzrWUIRvW0E09DUqSjXzO7jU
g2dH4XSMo4vuQJCge97g/wkP5p+Q4i5nPIKbvi/p1fH11i/Gd+dpuGgj4Wpg+Pau8uXepcZDYwMu
QZSyzgy4jxPyuTDUDMwkWN6ptVIzbybbIu7EgcRz2Nu3FGtzKrV67bstD7P0BTZ2GdEEhUdsgqzi
OltLCZlkSKa0fomizk/URzoODdfHLCHxxa8UiggT5+6kl1pzFDhQZM5plV9zTvsJFo3HWeNZk2rB
w4kP9PTx+VLS5+g2DUtiekKaidOssYKyyJ8RUK9hq0ynqJp5BMGaQSJhZsEVkNY4va5AQ+dXrSDa
SqGJ+JXPKU2iniPEBqFlkUc48DmeN4S8KposB1hqCKS4A1WNLEg4WIcFgbzZjt3/zw+tYqhA41er
0P3Z+p8mCH2p/unvjoEv1gfbhL+ingtSjJG5nFyxT1GRbUetYyeeE83XmadO44euVJLnzgjvvBdz
0+W1ZPIbAPdArFXoTUVoRxZAXmOYThCmssGaYQ4f/TC3R4bycwCCmQeqEk3XP1AYFS/PikrOTs9J
hw9h7Gi3RSoVXBOq3ekiJJPZw/+9PJs9TND90AvM7o+9nPcFtD77E5FuYj4hzgTRBcV4huilAQDT
E915EoI00W8p1It/UZXoBiUKsfZWzhHaP2woTmdJHI1r5svJXrUYhfYEveXinXr84JaCJEoktAnV
FGoUH8dR/8AG0qI/l2nwRzmPb1VBBv9MkeuDT19qyVb56HZ+JH9CPZEP5lJp6xFG9jg4hmAjJb8A
WrbnXJQa6B4l2Xjq+KrTV4sKcVj0FQl7egv6Dcf3VZPyxNspiKko3NnOwIm34NyLY77Jho88oom8
PSCVcHk5BMTUhnWCbQMPhQ7ZhmPzx1vXMQrFVE3KsBK/Nz5LkWWa6Ij1R4TyQNRlbaxI2cqgapc3
xI4/2VR9hMjeAVd2ya85E2EbU+WDP0e7JumZruIkO7+xoDaq0mRGLJ9B09B5SU5iU4tGd9wWhDMZ
3k78zyD+XVenY+2+N3h5W+nsPR+rQ5Haj/1woARj4b9aF3hrmkAulkn0gpQwiSIniwVUerPHPPYC
2usL4nZMJ0Fx88khFHDq8FKhUNbJlHBiB6MsWNyFqA5JQoWMKOXR117HHIgpWvTPv8hATAnVU1oZ
JW3G7arMOjX6Guxf47vQ3C+xCd7cpg7nM7UFbFIDqXdvbwde6w5xzJTORoLu0mx41STbAUS5n4pi
atb/TLUJQMlHwrLVT5g6KMGSmUuPCNutZ3g3/3PqExWRwp/P4xAQgYIyvZmBlw3uZc2VFKmSz2A8
U59gpI43gEkeqyh/MXkPyZ3xtliL0WqzV2JLD08t0vdn3rvwSc1XJhHaXGERAh+v6AmLxd8S/8uj
vO9CpwVvParRhSn2a8zHPmt1zAOilLCfpn1Bo3O2NA26dIm9Rn4WLQ22pNSFEIDJNMEXMzDb1Wwp
KBvRE2YXK/NCatvfaQQKGcdxxqBT77b+dC9TvcBlC9jag9JN/vYA++PLJOOKdMGx1D/lK2iMgdsg
kuv2wcMr4K7qFrCdKEJK6aFr7qsDqqk6YAWPLwfORkp4EKEmXh1y0cvqOxHqLPtCwveYFLoQ6J64
RoHvkXyLXWVDN9Ld4VF1Ks2l1XsUNfPkv71E3H6BCzKv4GakkH+18Pw9/qJ/cpEEt31yeHGURGcz
y6abmHwcSJs8KE+aKmWEbMHziCfxTbozXTPJkn7VK+VRkzO7dUaO5hdYD0YQPQAJAqKysnGo/EgW
NRYqW9ooI45Hvw9vitQ68/HY19n/7COWUqHRPugPiXCoqrcW7Prc6u7JhyXxUtn/sbjBDHDNl+FW
4iGYC8nD+eapJ4DR8dMWpgKmuv6F+HRz/QM862fjf4Xb7ajTJ9SfyEd5TtABO98RJCL6Pir8a+Cc
JDVr5lmCj7dxPgT4UtJXnsOyCOelR4IvAXy7rzkFsiOQsllmCNQp+As/3yliS6zGtRyJAMNKfen6
41tmuRW3AUZyAq3du84C5P1Q/BPc3UiZBhi1J8XiMFz/BRv713nr8GN9P4DkWyxQubxP8xhSXWZK
YcIGHEeoBV2A2bDbdqD97HEsnfoPv6rZYyvc8FYbeNu0VS36MZRp56cu/d0SEoHYcPTQJFl2WFMB
4Zd6UmHUvPhovIrkUAQA4r2bXjBccLE7GZYzVBYewyEst/RbYy/kyPvZSicFnLNHc+163oeHSrjJ
Rn05Tn51NSkhx1vXWbIPm/rYNc81bOFUMCbTyr3ThKF6JKSitPhXQBr0Rm3PV8wHBP+Q+5xmWMqe
vkNVVihAXklvXVInQO9c2przMbJbO/1BEN37scOwlZiRshbsXWpEkWBmjLlfBu6LJD1nYF4eSUWg
FX5xEgLpnto9+Z9fy2UMH1aciZ1PqrssidfL1O51TV2FH4nDYONZeQ+49ct7NnkWa/W0l/VfjJUQ
FzV4d44ZZeuhC7Sq9KTGMbpUY7JUZ+9bidpzbgoED3Y7+U5SxYFvlMvutIFIRibnKbbYFnqPXatF
1tC0Xa4OSjH21/Gi0iY2TR8fPcewTMqenpLgu5Sklk+tp7fdfiGFHfXYZj7WHsOQRQqf3PTNSHX5
h45Io36YlaLtfXC9VRljZFGsd6FDgGGp3bT8ePIWMYhkcm7w6tTBmIYDIyHNe24siqTPfRvZU7M6
adwojtkZXln/t03nJLZCFZ1whPJq27hItRmNlcc17N5enCYed//CfCxeImSSYiUK36uLJ9hTMdCw
OMujrvwAqnFwMP0hDWbso2oJ4Jy7ClMxngKWhrHebbIexUMcIwtUkn5uPM1sQ6GVnr4eEvKV8dS+
b9bw6xVasQWkQFrpUv4+xxClE3jagTSrXRVZwyjyeoa3fEA+zlNXBvCIJIqAAmT8fFhoUucD7+cF
HvcOs8MXgW3/Fh/t++bBFiOmPAbE+s+lrgWCRGGmawn4Yw7YkTilo2x8cvGLe6ZqxiayR94myvrX
tb38lk9mkCW6lLn6okhmDkoVQuBP7ySJnzfFbPxAH07CPHNph6u9AYFTsXYDwJqGg9dQhRiFjdhO
oJ1liFXqyl07C5fbceSIlL4cMLPZQ/ie+z2R9NNR4BdhO3JwxJjwxG1IUK4qxURNZyIxsfq0SGvC
37+Jm3qnoFGREHdWInI5LzPleL0BOXdJHXV8oZ6Jk6NlXPLlwym00E4+04KT1xPPxTE8i27F/dFH
QHJI1DV5TJWkUxK9W9vhP3oPayB+7Hv+DfjRs6qDCgQLtbOItl8rDGfP6fvRSOILkJ6HBevAr7Qq
fouLZXi9DBViLNR9Z63DWW7U6RifeeqPgd4vgpVCGC2H/PaIUcrWhC8QSu5rVyqu2N4fjnhVP4a6
Laml0YPCb2B7+VPPBtUl/ddenRqehunwDgUzAIP1MBw/nRtHlR2cUZUfLF7qd9vU83I15wXD/K3j
o4IzCo2CxoEV/bqgB1iJ1mBiIx4AsbvHDCm9Nn6sVL9PgSaViIRZph3NBlz0oOHmQTk/RtB0RnDY
IOTSlbtrjEDKk09f2Oefeu08E3d95vKdHOOdnz0Gu5bITJMjaWZdgCRT9U6Egtp2Q3XzBy/5jeha
d+QYptHHnvX1M+DaS1fqR0/o6KnmkcPQWBIsnTv0lLd6/0JJXhdg6I0XQnvPFzyAp9q9eN6eBKhR
ealSfT5cq4vE7Tia6iA0teSyiwOBHyVRQAgQJE4t0KPhvVhzDOtFAT6Yy7xpL7Em11Rtfo2mnbjR
RXfweTq3ZWpGIl9MCr6Xqb79VdOMj4XqwIP2dON/QzBUgsc/u8gSF7Js+R3UBJyQwPyvJHIyU/MF
aN0K7GdznVVrEclnVDczigofQflNzz7CXGwiQjwo3tqMcUtSkMykQ4kXaxcCKuLJG9evRyD6XTIg
bKYT9l3xaJPwFE10rm2ochqrLJrHRzHFQYce6YcnxGKzdgy4jWOwaTD/MhHBiWhZyl90jCGCutl/
ZvxIu/NrH1+wYhsVZ114zgfUoTKaLEwFpZPBbPGldRXNuN6PTAJx1aTb/R8FlWSXJyjX1P7zF6Ik
Y41uia8iEMc3n14hcjrjnGK8GEaUmE9tVAkcRxUwvM2c1+lxzHW9l6AvAmlCs4TWIiZSCZLufU56
WR9vN6iS5Ez9v7TKHbMKnM3RtZPIZtygw36IXGSrgHserc0d4S23JfxiUtkd9j+gfUU6VQ3xc01e
0T5x8ybqm4S2VLepuHmD+MlUQiqNfw5hLGHO0SjoW5BQVRSHNQadQZCPdt8R4SoeorNKl2IrXCOE
dq6WyP6zBSjQ+ubDzvqJGJ2y362Qb72RyWThVUY/WtnRztdnh0PIU0jsmx7k+rMVdX+2Avx6QZTF
ZcErKGvG7Nv+kTRqiMCOliz4CtpFOH85vYyUQIRRUlEsr2vwjy89K0vOcf60t8bEHsuKVZozfnFb
sOuxbQr/AIPnZvbJNT7OWxnD9ct/6RFtKSOuBLuuh1E7GvtRTFCgRBQkJNazn3dpa4rshKlgRoE3
lPXx/4tsBVIC0hldkuPlnFwLTDvohiG2ouySMRUQnS0vo2rK/K72yKczzvSIIcrRMbBsCzCzIghX
JL6m1Tc0j+jykkyyiIS/9GQepCazZonIHMrRT/V9HNVhmYebpi3OcA6q4p3GOUJG0+AdlueYhM9T
gvNkmTQdYINm2I7Shw7cZrsTnBBJYmEV2npnzkTgoUHesqAZuPPD1iHUxqnZzAhE/YSby7YUxCOS
53L8iiHHZS/YgybXCpYQX/+Wbt6JOr/zJOznwsHvIUWAyy6vsiGCkqI5l8xmseiMqronpzd5YGko
Gkre8y4sMZB0y27z+VMBPtZs2us4aVgaX2hL39gGb643IYoNVeY/xP4hqw8PEZLoHWhMnjvX8vtd
qPJaVa/o/b4BkzahWATciHAPdqNkdWnicDa/A7rpbjbOWePcsiBHFwi60WmNwnvjteXCAhEVCcz2
VrN/qMUQy4ZCke8Emyv89J2nLFmvEx26yCr/4cENmPykpEIBSG1ub1HEKbRtqKKvihBRqDbYOMPX
MVS37FlaKatDpzZeKrJwXZPuyJ2NM8JsvimWCypY/66uVgWcJk/KKQx79Oc8EbfVeOgskiDNufgg
cH62WrO8aCQoLYktKz7WOK2dcKgOZxqBgTq/PiY2edYUxlTmpAs8Wy6HTnpKSoIjfN2wDuWCIYnu
5EAHPbPuHCAZOZqTySVj4vrpbfZeu/OouY+BUTMU3PEFc2DSlxFIKlxytok2/Ofq22pLXC7FPoki
w9aI0YD7Hel4CULYDYzyRm98VVH/RATVmbkpYXrL8VaRuS1TKQp2u+l1CqUnfHszviQd+MV1VmQd
6rKgISjUIJpwOJrX0gb2Jb4DAHvcauPuMoUTlVREUspLQCr6EkjRe4xqYxIVZlCoBmMUEy0hqpZp
g0lZWOsK5HsxdAtsNADFBYMAi1MRNN7c47rCxv0OTd4xmLP0s1vjQzGnCykoc0wVG6NNaHtYijkP
V3keFdU1A7HVthZp03nHuYJjxl7MT5vSYCw3eYe7RrpSykSXvqax9uIQRsZTKcEIBZzKJBlIp7X1
KRey8BQVklPmUueh/LZWwhp4HsKUBytpmE76DfECDhYGlVg+Mh9fcBfmn28ED/4/80zgflF/+ip2
Tik5qOA0VFJTmGRTb5LRyuXBX8ArG0+6nzICXEt9Vi/tJ/kU8TDN6tPVY0v5+4nOr2FqhsLQAizZ
MVVugurkPrbYml9rszspLsqQ8BcSLRhlidkh2WtadV2DnFgx9YtC7DiwlIzC3OD55ilv5TIJp2oR
OTiLKwAChrNAV4FFVIPK38clpfI/PvgeES7XAHjIpOyQrWIz8xwtFNVG/uMKIAfHT+zgFLz3HLpe
mXwJcEn79eJ9OZHtx+S/dbEWmHTEVTYrrCTSNS/ovTnJMz4xv8qn9DIyWxUloj2VThSPU5nDFDTw
56CabSqrcZmlgjCvrETv8Ax26vtxKTE9DJxCCr58hgvDdGsSNR5Bi0MO6DTklkWkMlgiUWDT04bb
29BcvmEnti/dY8aS0ytKxARQEC3lUeCja4MkRmpx8igO2zzbmAYlDfxOtNc/Vp91N7/NHTtNaLkc
LUvXvmbUw4TbnjFSwhJQYoCuT/WY1zwLsxTwvHVVmXIv3faHeMo1q5qNh8jemOHJwkwiG/ME8ipE
pkYqmitpMZygUmPCyAcdANV0bQWtXgOJkSYeLuh8wT4ENjR4rTQ/8sfk35B9JfSeksOOJYLwFfQI
Hphv4t5Kyib+D2onM/7v8OHY8HhA+f2DnVTAO8XubegrcCmldZVKQ+fRSmh95hiXIRx24S0Eawpr
2y2LXORbiSC2fxB7EqjfZCV0D7V8DYKGxQ6lXKopQA8IWEgdh3EDkRo9xpxtA4tw0OWBWFV5VNlx
oOor3AkmDx/GMHdV2AUPr+ndwGPbbY+4eIlJdeJ0+25iej6Tzj/VvNX5anD6qBcv/rDthwSdaDVz
dOmBCPKxqxDvpj7VNI5G0NdxMpJvcZbLpAJXNo7Mbhdds10IaGShMBrjWMkzj1/gK/P+dhCN8Z4V
yOEa4IvqiFcutF6qe/76U2DqjFvpJTicImjaOwTgVozr/Rptukt12cNadstf5EZmLKUtWm25zi0A
VvO9GJXVc+Spc5kQ4F6MLhPJB6W0KKHzm09vm5TjDhtBuAwFC0UXsr2aK2hxeJgWLRAD0Gv0EF0D
27Xha+h077XyEYDdrvPnjmfD8Smj7rdDUcFfJgPsjyJXVzlxtTaaF5c4cyTIkafyAf8od8SNOfh1
nGWcZ7Ls+d6irz6+BoKMzSXLt0j9RPyjBoKHv9J8PMMHQEToa1KGq8xfmT1Bz1aPu59AghhXJcHr
hbgKUPZVlgXcMzCNx/GR30g7WtFPqqOMVV9vImaYj86n244QbFnp0xGKcq0w4kBFhKRy1fmZBjTW
rDeN8IR59/z2OW32UpRigu/I0j6SpylrAv1LME+atNHVMWv+TlixngOqN7FdCkXWgJWrC14x6FjV
u1C0eg89vhdCWcNomfWpuVEkRxhRNs4rlhHHZhGmbU7i8mfDF808/rtGbJUoUmo3dQnA3LnxfgOh
BN6SupelHpgWpxCdskx19CtDQjWRPOhP7UB8oFn5MOP+XaSflnaFFFqbmuhMAxJSW0yBO5hull/8
9F4Bee6nrbMHqxGNaKo0wU6Pg0Wb6v96FnsfsV9kAIOrAF/ytQBGIOqR7cqLgnD3Os2kHyWZn5CV
k3U0oD56k8hMH+ecHZx4KGr0IPmKQFrk/me9xVdVuC+S1P/4rrdqiqDvc8690PgL3Ol3lN28Q2Io
2ofUwwHIjaXyCdmS+U3A/6Mu1uVp5nW9P5uS8O87Ur2aIYJe5DS8cnq/5pamknf7by0LrUfdxVDJ
7IESfdqb7RD384dQuQvca6umKhdoBuSBkkvdFlA3yGVg+xHgBm0D5IDCHV7js6i5Vka52hcQ/Cfm
6tagQgDIvt1g2IgCH2q7qUMdxC7GqRY4d4z0rmpIqadrNYCW6T9MXi/Q4qRgKSwG2m/+Q26jkTZh
++JoPvg4voVUoH7Wucin0epirObk9+0O6PQKmz4x7zn3U/nP98cf91/zWBc5m6uqkT3GsevXw1kW
Vk+Dq0o2+Mv2De8iCxxo+Mqn3ED2j/ZJP7XUaGYnI29KnTlfokv/nrzBKco0nKwpJMiX17xM2J6p
+u6MgBY/crPOGUtbBIjjNA/3Mg6a4O4ZWekLD31iUP82D1QO/Xei7rXQ7jkRPCWce3S8Qc1SfTwt
MGHwWBUB5t7+0lBqVLHNZCpsjmOsENgumQEvRemeBMBoXEJjJPauxyqgkzCCS8hiUoc0QakYhd8D
q/2Byo86DxtfxBA150vxkLd16cPdWP8mOdaLj7hzyawt4oFMTs72R3L/lpIT19AgM1VnDk4AfHEG
/x8lkm3fZTRk8PhZKQgvU4KcMzJltld/uTA3VLxmpkZTG6UYfAzSycqPiNDQI7H1vVjR7waK7864
5rKsTO1hwXhAaRABksVel82BsAKiBtY0PQqch+pFc2YrRE6472u4F7I4jOKLu7ELWEGAzRf0ZbEX
2m5IVj991MgT51IE6IjWwB+4ONzDkWNEyKLMIN6p7br7vqdJKr19eRwGt+rsbHBlSLnseNZ7WST+
VvuDOy91zXZwRsJC0aQr1EBxQJQrgttc+t8UwlL4zM29IQa0zGv0yl/T72RSSreAN6nQR0T+IYLp
Oo2LNl/4hZ928CDvUZyrnCTWVXg8KNL++pL1qR8UCpPYvJ7OwU8qCvLdfVjcYzfumNnH9tYsmiwL
XYnBG9lgsTtu6RMzgNI+06KsKmcuNYpDr+axRVJmyeg5NKPg25nstS1U9kuimOJ41ZJKNNuLYm2y
emCCawS6E5BwUcvW8R46q0CPkRsxrcjZvk5sv92trK2UptzGgkwzuVzdwXeiFm34Y4BigvQfaKZB
QjEJD6+lc/fA4T+Vt2PtZ0VKPqu5ywfxO1voPNsE9l8fygEwxN/WYuJVDn74+Ke4WnEmthrGrQI/
xnXsBkfdjk/crl8S8IKWKwov0oMDCFr+lmQFYJhyniqf0VVYLQQROJEo06OG41coi6+2piaQIv8z
4EU7+d3nEZV59s1rAkyVjd+7v/iaxBdIhYlz9sJlyp7aGejT1XrZ/Ri1W5Gcnube6qs+G95buaRu
eMHxDDkS5J2+o1dSEkJ7jRpxwrh0heYltZjUwIHLGMHPkDKO3dYqxTQe2oxSt95xb20f4Q4XIz00
szLj8eUjT6K7ymFLOE/Gov27caBg6eYuAgYYq2cNDdYh6dloAgV2KQnhg7loJiD12rlxN7dPpM+z
odoJ3re2xCgjEqzwsSGwrUSuyOTVr9fpnUFwb8F6MdGmZHIUvzuhXJ5Y7vN5ANIPgOjRXDSojgNN
SZUwVGMWbnhEFLSSZMrgpIk6po/9DvP48jRmBRp/WYVoSw9VlaFyOwgyF+7ctFn6O2pCBrDIdGYn
6ZLNJXjKNmh/K9yFTB/sPZheRGzAmpB32n6SqRf88E/m0BiDXuf74N1o/9Mo3yKbL5O1opYRPHZj
lpLTPQLl9vmkGn+N48rnpar/cbFxk/fgVIul2P6MXJvIRnFVeMvvph+epL6ZG4StNq0VPbYbncFp
A2UU9ST3VT4ARu+rDfpCu9cIxM7TJP+rdvfAJ64RfWgynAyq++NEAzD93oZH/FWKaNMeMHwcoTpb
OsTggUFA1w7JezNsNl/PRuJ2JSuk0vJsxdnKH/+7QotSLj11Y+gni0/Aef0hWGVvhgeT481FgEqd
VK6LJYgVMn4CziJ9DyYTE80K+or6PjRUgHufKX7+KdlsW8MfPZFcLasaikn/z+EzlGbNXivW/9/h
vcvS8/Jxt6LccTSZrvpBPvEOOzCfDPEuIlu1DI6WYO2vpQpfVXNKgBpHngeVgheac33DCwfFmlmF
nhsT37ab2zXuvfqqPVnbV1MxyVj2WECYaPGSvTxo28FLwOSyIUDyyS1Rb+b2N6C4V+KJAUaS5Z4j
HahUbBgMFD8IJE9kW4Ueg/VhJABjYzpdysR/OBdEWC5CMllVCU6foFZd9NYy5yutpsMUVGbSfgA2
30nOw0bMfxvIYVlBXkuOs6oKed/SeEUZ17eYj6c1ONnRnSglCxVDBN24zCgqJnMu3kVA0w9CvkhQ
nugtKytb0kshQugF8adqK3XC1I/o3pT28G5XGVXZAdMachjVPkUrBHlIUxvwhYnDkDNrLfYJIGe3
HQNgN5E3eWk80dUrKvFC9gKWd1W5WC/tvwNucCa1QYh32a6nkkcmEBqiJ7jEp2WfBRf755hcxwC2
F5sI1WhN7PdG/9YmWKkoUMM3XeqE7Eq8Y0qYuuntnTU5yvKTpWx4grgUWSHeC7131IgayIxwVWZu
vptLhld/WDTXU86w2PSEXt9nqVmD+f9QYqD86OEJ/KhWH8xXq6MwmrReGLHFBYqEPv3b/Cxrkp9y
ScPWtiNDRiltAOmyZVgKMhtBKrXSLXs9ZfOfyrcnvlsfGbIUbSXh75sCqs8ZhzznZpwHX7RP1IOC
ciz393D5fhCl9XyngPvPC8JGv57uOKGPRrFj5rTqAgC2QLjaJ7cVNa445I1NeRmOZrdDriNU1xEg
j7cNsSYv1fHq5kbi54usVzwOTmJWubcYZwC3Agszn3IXMdoch1RPf60j90Li8M2lSAOSzUsI6LoN
L+yt7WkbhbV3X5s7lAoOrgRJPQqdtG6gunLZ1g64Yelc7eS8BfksJ2CCU6Ka7VBT5l4FYVyICl5m
ZUNBYxwd74KtF6iUATs2BeeNBVFsKLsV9KVlMUb04fDhSval3G5F/3QvMyoYRrllcVioiecyxkvr
a2M0RByK7alKVYWjQvJIz4isw8EYPsF8LeeYiBiopzmAorvXVY0yoXhRkQ10eHlAcwrk02lHE8A1
dzdkeUUJxxptFSmncoHMOFpk+Dp0c6vd/9MqRWrvP5TFnRpvk2Ch8Y5XUnmKx7gliSfzE3H0uObJ
1lSGB996MnqckF12Bve7H1qumhlq8bqF2zu/BrvsMcFCT9Eg7rgmX7r5jMMQ9MGAE12NTXc5cVIt
8eVZVu61rLNn7sUnJ6+M88JIaTkcXUeHvxykrcDYwgB8JTjyTK7phVy4s9R7TL18R6MHr5WajBxW
zHRXuHKww8iUx/CZoEivnUOXk2Gcw8dn/9D/1/6UUpnmzxOToGw0HS6cj4QTxYwEyTsNH8jtWFof
SHu4Wbo/8M/IIgBoFi+xzC1G4DHoJ07/ahlO9+zUokaEjyqUb6U/J8Wa9GbxPpOlHjtFwdWolgQO
7FUfd05CnzJmVsseY+osx0LkzEh0ldNJFAUesrqIgfS5oz3pK+TSqNwuGzzJwttDL2wyvizAAwAI
XlLlWKk9T5PNqYMj/XW3Vqz5ZthNMVt/f5oV95A+X9lCpUOVJGl41OjBDW/Wvmj2aqkxHaktcKjk
oXF4ZtRoz9m0m5rhcRpe46KCofSZSlHjyi90ZrwIuaUPdYBIfvpQxSjvrPGXLDfrdUo4Gk/FrI0i
P4yWTEZbtNycPiuCyriW7Proy8vkG8iZ8eaKsk8sSBEmeRj+lk4xj3aV9yDkxtNNtjmgrQ4ECO3j
ZswFjvMu+lZ+60clnUbkKLWsgvfqYTWLCAQVVntbIu7z9jEPa/0TK3EJye9FH9OWy8B9sodn+wDp
J9TRrcJ0yLfhzkaXJiKzEUze5osBPYsWL6vLBJO0/7ohUe+KYAuz3rTPhh0y3YAq6bKGLZEuKlcf
cKI+Q3MrFge0D5CjAlAmDkHbpxL7Y8INn2CU/wUQwAuIqZWvXoUlr1wVhv83/aVXpSp0dCD0Ebhj
VOmbMgtcSNU2x7yLzdGWDfujs6AL3oql4Nf7f6j/QgVMj09sEQCPmfQ57zrCTkLSBWFQ71An78Ys
oqpOBv0nvDuIs64qCkHHEUa+yoFowVw3Te8Hf37V7t3CU7rjEQ45RG71tuvC63TTJW012UQhzCPw
srFCIIZWXIGv1e+sJ51QWwxzNQhzP2RNG9IKPHlS/KEe1L4TltTacCtA1RLeBNZM2VRXh8fPb3uF
AUCR6sfMTj4fbg5qcDNQirrtDhayUeMxNPR0+KYtHoSGPXqKYExHlOqXughSOdDXqoThjiPf6Yfz
jUnLlyt3zf5IfbIMy29zk4lFmk5T+n5UMkmRwWaXPzcuVro/PtVkCxXSuJQtyPlSCXxNyE6fhZq0
JpMNMXwmN2uc1+PDEtiPu0EdeCSqJ14YT8TmUNNB3+M3peW9UVP5LUAouBZZBaArtT09FdN8Fa9h
BhrmGkw+czgGxzrKOQroDOhyoSz99uaPYjFMSAoRBd5T0VlJq+i3qRYcsaEjubg2enhT13wjPin+
BZOD0snBs8lmDd3AgO8tY9LYrdxOsmR0XG8iiMT/uc9kMSuP7Q6D+nbb829oSrbWIM5cztlPfk7x
X/TBYOl/4fVzZSlolDTXd5z+Zx1QxtYSZSJcGz33JpMZlmk+SXtEp1WIDWj96VWvYtsYJ9NhNBLJ
mWN/EFiOhy8qM+krzYZ6RIyqUs50myZmiddaYeGcBzfTcbDRyS0fzjNdJwYVNYxmJ8M7j/B/EkBz
3AHc0iVDB+D8Xx4CwDAypiOr9uoChA97l4KrzIs4r3fFmG1xQZvUNHQZavgSaO8VrCTeDH6YjEr9
GnZfOBlQupM53oeLtZ0FZCgqLFH6NWGBQWSXTxLAHBKydzCeljE6ZXASYJQQH8dCkOJrF9BAHrzk
5AM9MJqOYLETkL4bDY6RzCg1t9XGmsRi/f1G9AjJjkjAqfFbq6rNl0UiTk5bDMJw1hHvkx/+8waZ
aEiZDDxvC1+NfqNaH2+32YweRTa/70lCVk6N++ZknpfA0y1LcwOowycp3Xpakgad2KDUuLAm7wzK
M5NFTBzvhQYDhLW2HsG3ijGiXwvm7CmnYZ3R02VJmWWgxvcNSUJp+q+PSQTmtEHMiMiTt0x4ZTIF
wlPeEiCIt0NhFLuvYDWfbMzotyta2yFHYRyNzNqjXprU/jrqJVKPUh7WylCP6dF/wVeZ17MNXwPh
Ze4zep40Kd0Inls8dUhcTNRItWVcDf8pXHVzwP0rhmXB39ftdoOOjjzXIBNv2QxjseCGrm1wQ8d5
x3C3EwHjW6PG2cZpP4iH2noDVzIO01k1Ta8ThIJoydFZxEr4fiBcxoZJGgqFLaTC0RskecYIE0GW
DBcu1NGhu+T1Wn4NrTMVa4LF5jqIiBRAZttGVd5G4na9Qkk2s38007eHP5ERyMQSWuka6DWxMLsl
M1LdHXUO6Kyg+MsGeO14HTaMZ8Li6YKZmT3df7BqwifcVTkc+lBDJmk6XT09Lne/ePVslQFgGokD
lpgNUESC9PmIBrexscyXx1VySn4KNLbdSDR1zohNbYCgGSedUebJ94JScGUDyXBe1AJKtQvsmGlx
gfn7+0CetqJtvHC2ep2upt1gOP8P2rlRjm7cixA4NzmIGCB/RjaTu+tFNX2sM7LJzR/BmfcLt2h+
GJwFbCcBXi5LMx/RwUTGo1DzZm3OoJo7ICWbVDHbfPm8NUNNcftQqu+2TBOTqiZ8g4xKD6kOVYG/
yZduYnF/gM8k4gmhgXqPWJQ1kPQAi3Gcw0MB4eODbpGHoBdmvJVBHx7x46oR7fVxMRX121ve9EYn
tCGu6vqpEo/WjLwRZrm54bhztUVvkzrFA1Oq9EyNSCC8uDQZdjhr6+pbcUCkh9rgWqDlX7utuunN
LcefqvLYt/LXAOj8aS8fQy9oM4ABwtqK0Gp/RugMO4YT0sb2YikLOajydozhdmzFpIFoxUCt1uyK
yVu4BnigX4W9Fpu4qtcsUvG7+x57+RagcVYfoXMUDNcYg549PIrmNgPfG8vdvSkIpK73UyCK2/Mu
azRp+Bj0xfZqOMWkKfxk/ZCt6m4q153GowHNSWh59VWBTaO/qobmgxdr7UJA9sDKwI825Ud7YnHg
HPW7DqUJXQw9M7pEdKEqO0iKKNBsRWaNPGRNm6fFS8qdVlEiO1BhiEBiIxTGL1yBZrhAhmTiKFrK
tj9pht+M90TrWasG90a2ZvJD8IHIwIGz661E6t/MFh4cr38P01GdYvxDH2v64LRWBf9kOLRMN1ku
csBRTo+pHC/QbWVkk+r/BRCt59cBBnnDcgtbyLefaHjEbdRr8mlHeUiBMmxgQ6hkvwfKA6hnxdUe
3ctJWMSbYcrxv1L9ppZXMP0ZAO6vgRzjMiL+nlu8ES/efHxxjJgus1cS86HsrHTWSnnIWwjv1zXO
bZEUrJ3/r4G0KNzvbvV8J3tlKwcSplqMnU1zzxR1RTSbJtCf4CSrbWs6EpsFET1TNGGe8k+GCBml
5PGBmNTnGBG5TyoTjvbHhsZsUJuoshU+2tzkIvx531EkJzD40nFdcxi5++VqbNUIAJPF0lxvXz5y
cD4hzo8RKlcmxU8UZFTt/a9d5wmYqSY6kb7r0CVffeWocWIt6xRipYnDFUlVs3G9mK71KS5eOq7w
Xr+KvbJ60iu8mphODMWMCxTWpwGvEGoMkrOgx37/SpFRzQeNizwepEapxHk196Fbgtfsvm1VgVQ1
2pfneonnO+3Ca1XjgkZHpO5mSATjhUlPnBTijiyWbBKSFxLGc0wup9N+zjSHk1X0wYDOBCQAQswS
I7xLQTlsYjCRFm9jW3QveqIj1CK2eKaPiPaPfQ8WevgKoNgIe9DyR9y9/81MvwFB/eUr377AxW8J
W4aT8W8fOpH+WHkecu0YdMiaCZXN6/QsRdNyhA9oeaAK1MvTLuC2NjdBA9TX2Qef9Tcj/RvYdAn7
bEoIAJkF0kAGMmoGxQxISNIlaO+XmjVu0A/3Tl72/yRmFyoODFbXcf8kafx3FhyoowGW5lODewaN
a/2TRmxKIoEwW5vpvAxpzYQhLmXo7R/a6lzqhqzRxDVzDkoufRygXjib3LuVvj8yKfAlvjNJikx0
VHt9qQ0nnoGUal7DT9TYCdnkYBij+hOQH0P1v7+JNMneKm+GsqPv69zJccl+5q5Cq3tpBuAfCf/a
Cq9eay9GxXZrz/6uER1Q50rlcIxqNrkakms0t7N4m6gMtsGN2B/6E2Q46vaOPu16mdo6yI8chxdl
wWLTMebk7XqJFKBnbfVkAvPQEbZ3bf+tEkHLDkMszOHfZv9EjbU/ZPTaHOO38NGvkPLvUd7cJ/ZX
dU+o88VXgAScKqi8PkUZyRUS6AyxQWDTfnSFbJQ7Sg9CuA99URLLmu5QOU1R1ZvAi7Zf4Z49jrZV
i8UF8dYTvB6DkmcTdTQIJYdcOZ8ZblX5cbPbtqBDRZ9msaNGPNxqPn9s4512yiUfDlKftvJFVXHz
mJWPjGvpIFz4WsYX4wUZJG5IwhsPci67XPEg5PEJg8G1S2ID52CmQQ6/ncSPTtPygNBg2mthMpge
nn+KxVi+/tYx6L3PmXtgVKcXkVm7YOCm2JuU98SvQZaUytpQkfu/9w8o1qSbxKC8Jcr18FVsp9Pv
1NY0jgcUxPiMfRgURcgeDsOcYYJpytCBgPvebN7XUdNLww0pjre/qpEDCMCiwanA5ASVG2FfiA14
7ZmcfwCHYOAgGQpri8UJly0CVobJkw1v8r0bRdhDQMqGBhD5oLOgQYOoJUvNbdsnoTdBnmJ63qt3
+n5vVowD5dOAtFzMdNyBzntnjq+j4knwwFkDLeilbeREojnfUu3XXhULMLpn6rvsG4Mad9nHkFfw
ApRPuZOnoDuP2kxmvUOt1SI0YK9sJ+6b4xUDXTvXFMS+vjBnNvCtRLyXhZaC9p5KRmr2adqGNsfa
EG7H3NrcYjcEca3x/pHjm5+lX0sEO9z2/a1DMhN+tO2DXBRX+w7nIexWRunOBtMPxcWJN93O7lKJ
fbwWVjsM3m5lS2mWXlSCdhHDKj5QxdjjDQgvBvQcWBKe8Snnl6cEl0TgGyP1xNASKdU/NOOYKi7o
RCWdU+0r3bYuAEHujUVIbkv5li9d9q+vgbZRLRiK2Gy3eDpKudYscrgtnbe8RAfHECO5xOpC6qQ4
fjqFQf/B4847rrXnpuUSfk6n0CxSEP71ZRhKaFu1KMCW6F1U55kcbL3fCkgGvVWcR2q7VTxgPWJU
/VRisXVBhVebOdGSA3O0JXpNqfag5yYDBb30B0yGUodH7F2tfPRgP2eISfKsoYx1hIIY/G4lhbBS
jbUYtfPNl1GsbV1b1jqClyDFSUUPm+ve8bs6WgKqlVVmFKrDy52aj/XOLgKATf2gywBf3cQSMnwP
LcctyZCWK9C8qiw1i0t55w6wRahKF/6W4A0fNhHEo3Raq8jgzYUoK8rnJ2p3g/hpJ3emjYW8/srP
p+et/9m+Ajuq9+iPbeT3Z2a9BEbnpNLekJPsE7EtcZjuvfl+QlPIsNyd5fLlv7EhENog9xeY4CUC
bIT7UhikyqyDbBRggxy5dekcc27/HlKTcmwPcU3P7zf7Gp+uN8XlwMo5aV+efAUhqMRpdENij9vB
rWyFVKVrkjC6si5SYqP72TGApHqO6XX6246Pc4HhlI2Fpjbw7MAkDMnuQp5Zntgr/lWwJbeJfXsR
t8xOh+n6Qw+5uatrlpUO+NPs1GI8KGxnlR8D0qYROFzk5PdYiRrs/9kC4Mzk4FVenC4Xqe7nIhnH
U0nYe+VIljEuu+8fZljHHwqKn1V22CAPmEybF0f4gPr5Pl42H566db6U3KOhwwGFqGLstrvrn4x2
aBf+83vWjJYEU3s70cdHCP4/zXbdnCY4QceyZxJcrMk/x7JtRhPn4vrwkGaEq06Lwcyz8eb+P+TF
OuIHrY3FDdaOEQW5G1MEsD16yu2pzp22K+oP/gkMRd56eAgL0KAVkoy1dZXDc8IEEKzAr4B7j8Dm
EuEUh4BuyEc+Ds1sVMeuYsBJewEVowcvm+BbWFi1+bluOi5IUiSzR4vQ4nQ37jy6aPjnKkMdL4Am
d4h8lrMZ/QU7lEfa9kNvI0431PJ5wwj1PRhM1vbnGMzt2+BvI7T4h10zrnhZbi2pYXAGmoDHuNvi
d0Od8JeOvRgbHqMe3ds4lZNz4rKzcv16sKid6I8UHMT6auSyvom88TV28GsPQCT0Xu+JlPgJ5Xu/
wmd8BLfMyPILEfeuH1YryMK7FuG6MWDs4t10x70UDSq5ubdwlQSsDzHGdwtVnHB7TxrOdMFVupMP
rFnlSIIsMwak+7SfdtexIsgHVBEvzQ4tBHZODHydXHzobqsXaKNQLyP+ZYfuPmHohmldMSB9z6O1
00erSXZSKja4h0iR9bY1yyv1SNff+asl34U9OeMi2hlZb6v9AhgOY699bWroJfZvM3iPV4bM+EQ0
In9JCammWMvTdGo3pCMOD0RmGczWHE/IkG1vCvZ/b4Vi6oCmKgEyDtM61NIlnlLBP0icpC99Ak5+
ujmC+bvo5ygCYeNjyJxxJoI2gWSfwQnpxQapkblGltziIYjhEDZYsqT1pdtSV6gDR7WwLZNBIrcH
b63pfS7kn2l/tYXzWN7Vqm9BZVp0hMlvawfpP4K+mPV75hJBG5rhYegra24ips9HZH9kJqjpMIFH
zdDjbg53n3iHrrjLcqXFPxTwlEE36RWhKYQfXzXDnvPgB0kVP2GZNPpzV5WJei1fLuKR6N2z9QDQ
5rn7Acui5OVSvCBhb3nHh3RF/aKCimV43KFQ8jx5QkIEV1rwfDhksAsSF0iLoBXGPfEOOt94hG2G
wnSLhCqxDiFjGKE7PlUS6wxUnw+zJwjP6X7wKw7iOZzLQixAt6uGKYiYz4VXN7XGa6sXH0tHD3LL
CCUzE6gLAcnMRvszzYoCNNkyfpGM8YsK5hyn0gqlNn0aVTttTykqULRz11dz1XOwsOpKV27ANJFk
T0HYP90apPAaJf3ZchWA0hOvUi6N46876g4kch0m5T/DI/mrgx8orzeu0qOWnARxNEOeb7xxBbaC
Chd52Tt9Jo/dnmdLcyotOHcHYFz9LQcgiPexDe4RUv/XfMhDhK+IyVFGWP4N0ElJWq0YqPnLUgCo
CkRm3z4EkEFBJifs7ZEzg+WwQ/N6Gied0n4oymLb7sw/4Z/odqHRso5fOIKaVhNILacmvdSLiZci
dn8IutE/v1RQSiKB6uFzbsp4Iowua/irm0WCTCjUHi3entZQN6wCFrPKxmcYfXWiMsSWeaAAnaid
A1x72TxYk2FDV/jUf2vwbzI21YdOictT48MbxB0rylRE8tPtJAhabRVrarb+HLaX3/sfXgaKSiSq
uEf/tinPwt/uJvDm74+gZUKZVvO6iniRatXr5T2+NLxO2XZOfSu2itCFtVTMcdtHvgd7pLAZPxbj
kaG7LOO339wN3lT8j4/qRJ5EDkDHZbsK2nq5yLPEb49uMVbGvDGVS+EIVTznFSTDRLpKXCyjfquY
DQRdbB80T13EU3Sev7lCqJUXYjebmHBWXI195KLdVwhZxcuqItoS9+dL5FpEuyOJ/d8kh57VNnNX
RzBlWi/9nis4bq6MCZ7Vm87OyDNqNYWsEYy3AETpmZM7rQq7NbOyMlX7OwlbyqjHDsZBPAokVpu/
dhSJ64BTrFijKL1TIb2lkMyoo4QF2hEccjb1VEhr1bIvGtX/QfL50dxdSgRGij8DCDKuExG3lq24
q2cq4jpFyuJ2XNXUilcBk14EtmrF0FUH7UxzMt3j9rNe87PhxSeNT0hkyxoemuAC79BkZVvatE1B
ONL7vFyqvMiO7JkkMCbJiLDe286s0Cg8gk/785M6gnukd+6RW4e0cEAm9xmu2FSFfjC2lagXFq0/
ok0ra5FPTdHWriB7oaElIntNseCPaJXgKwskv80OAXFYym4sD4LF8NgQYoyC/Vhcx7xQ/fG1gfn8
6ptKHBdq+5fbKBAGmNPdTSWzHwVTuj9xQwcensPcOkC19YjMMBV6yCvjESFGeoNqgfdLlSmfEFQc
U1uk6A8Y4h+IdmoyB56oqNra3xL222Z4wCwQKcxVvZkzVhgqNHYSdVUXtmpuSpBBurLedKY8IVG3
O9NG4hdGvgv0OHMx60xer0qSCaiwHTyM022P88Ohg0Ql5CSP8GgOi5qvOYVqyNUvJOMtP9CGI2GY
/FclfbfS//9MNGHZKqS8rgYrXPi1LrHuhYcUKzE5LZEznwyozL364h5BIP4rOOYPmB2xX64Qx5OC
M3+OkCVoGRCzoutNY07h2aI2ZEIi/tXrPkimAyCQH4mzrz7/+dRSigdBnGabKw0a4Fhp+EqFAFzI
GCmyb7ZdGpl9ShkrSE6PkgzPtUNW+YayRdchxn/DIIjva7xujFwEFWhyvkryOj5VyyMmQxj6hLRZ
rvxY2B4AwGkaBFmKIAjaWMqTX6ygkScc1IvBXSXVtmlz87Ltha5HzBq1I6GFLdEv4yl8cWONRPAS
hRGO/b7D4DFUyeMuMaLLK/SAMMP3cFf4ufV+zTC8JyxsURvJmX5gd12VrPXawifVpMfVU6bjMYiH
9FsLHh3qH/ME12zVDb5JkinEi3lnpg2IM55nOmC6cu5D0VHF52qycBPr3xIDf9Jh9cp4P0+uADMe
F2SVKh3yNrXO+k9wxT7M5JXdRZV66WeRGO/FqsNF+BxKKa7ptzYg4M1wCmKHnS4cKiXH9YHjeBUb
qxy/jMLuej+OwMJnOB9KhrGEWJbP6FzC07gWdB6Lz/j5s4Toi5x00nZjp7GpJTvcjNNLvIsxZsJY
CHq0caJxFs1Tq9piCXHaiwsdZC+/mFYco/FKGCESVLKKD+UzeLYgiZCJUUlfigRbmTN4bb24EHHI
UmpaeX27VM7cDbz4w2U3J4MR7KeFCXRi+a/Ajy88XZ+ty2+IylhVAugjF/WD7JdwF1oRsAHc6KML
OFCJyPJcxmH6Yj76p+Km5uUWyALPmxIae2LvuR68UQR8TRN4+1L5Lm/LxtRvnZ3+fr8bx+9Ea2qF
BaSuhMH3uZpCeMEr5MJ9tmhZVDNJ9yUzbKuc9rSWiXsngKMRnJBM/l0F59IhWSvOwwgX8a5/xY6Y
lIuCocbkJ5FtB0mBV1neHYVlUUMxQ4R2p/TYAhW5Gwpmt5QOyTZfswqWX915PQNLlNTVyIAe+XoJ
SsxkzNnBSb4f+VZIjL9EcTnR816SKDiF384mu9FlDtf2LqOb9swkfarr+WfuXWnH6/lOFMZefo1T
zDVfcg9WcSpdHK57+XCLs50mLZqQIk7vbYIIRsC99dH8R3rNUbrW7N9n56sBwZGaCFF3ihpfpP0G
MfGfyspJl6QRtAJ3aItg4iU66/R6FrXkC0ewzAXYuW+wvHfrxh1hncu+1XL+Df307mIAOc67m4ZG
j9TbiIQnENtkFxZRyub2pLnuS6GwzPHKhG2Oy7F4w5L7lzVjlmsG12qh4TcVaRHanchHf2c/2PHs
7DqQHglB0Sgin5rqWSzf2CrVBPHiD/gQ4I/TpCjzgXzMM9lOD5DxmVLhrNPY3QoE+VVT5WcFJorZ
+2UjcDEIib1sNLuiIw0MGU2uplJVRdIj6EEGVJgLRR4uTpd8ThXl+yLC3coguLVbdoBtlOwtJpsp
di4vDneov+5jUHJWGtyL75ZldmHo9yD4d68G4jVkqPlGNrBoFNTEme8fS8xo+Qblzqaoc6CrqysZ
z395FYgk7QhIaLJQvv3qdkVPQGw/bl4l5aYAKNN1JSh5/Pl2GS34swTDFJTJ0BmA1H4af9OHHaSd
Fz83/rtqZ+rHzVd8PdzpUpCcBwlwtucjkOCCdURdHT4pa3ERwMJySbG0DtC2kFiduZGis9O5kMCU
yMxUfpjZmzxlWEn0YOMGBjJX8O4UZodohMhHE6hGxVSs3hX74pi9aTTVjb6zI5KEFqXQaRWdDYTp
5AdFziwV++7P39WZAg8DSoLK84tzGvN2wtTQs+7ObsifXYBkyq7PJIm39F7Qy9JGFuIsYyA71yHZ
vLRZ5QZSaCubgWx5FD2iOAmkdjn1mQ5wxJua29cHqq1zd3vElMVfT59b3OPSpvwltaprS7YVHgAz
sT6RXI0ZhsA0ZE1/xGK9buuTsjdADZ34UM+JExXQcLpIdtzjdgmdgVGu787RyYZXPH/oqB7hujZ+
Y+cd96/74XjedXKfnY9SB5HbNLMIb9Zw0gGxVOfz07NJl+o4ogxJV8GKMgNejMd414mheGFo7oda
dn+FSfGaP4E8CX0ZW8gzLTZJ16MxhmQ4Oxzc26+kgyDrar+BSyvOzQusWqOf/oE0eDOWbjbQoH7b
o9E/OdGKUwO45GJZCHgzLi0wtznF2xJRD2Ep0iquHkMpq0+jKkU1e+RzW4USOsyT3AWuykvHqawv
zgnPCc7L9D41aJJsMW8zVLt5wAVyVJHfEV1hM8fz6yR1HSwnGRDKphFX40rqtHCBMpPsLRYgFgIx
7i8P9IvYqLKg5WtbgcioIGYWBxHMfBjB19Q/WUGOb7RoAVaB31da1Rzk1JS/ygJLB2Yj/q6Vfwb/
zYE97FuKkkpuuvMEgyxpUOXUy4HsirDq51Qe0CoHefAIzl67ObToR1SeHhm9LhUqHUg9+3oia2ud
NNiOYHC9RKGOG3VR2Q/VX9jyXpPfe0R0mryHrS0T049/0uAvwUEhN+0KIzlbFdUpRDSNQqHMJq+c
y0YLw5C/SfyyeHWlmDJ5kw0kGqCy66cnU8VJEa31VpgrMnI/3SDSUCH6jIy5h48Z01TEX+Vjx1CU
RSfeGSpu6iP7mGjhovlR5SP++7149Bbnfyey2oK3WrQO4wdmdOV7DMdHBzDqWBJ3oNecZHmcH875
M9mksousgN6myGSnovUOklTk/WwlnlE+zikZ3CetJEbRE81A+qRjnTLATVrJJ0cTqcBe4q47QdVP
gRBd1goinwGLe1aH5AFMCa0mz3mf7kVj2erTeFabrBEQtZESyL5FdB/FZI/FCIEeSecOM34jnzZK
Szpx7WFWBCk+kM3/nWPVqpI6FRtZtCpQC6oGkNs39pYFpVZF3I3a5A4n9Elubhzc4bJ3ymL+SAqj
OtfAhttDUjWtJTZ8cHMTin0QpJzWGdSvvX+BNMgfNoHaL5e+XzRLXqHLWfpiaTjBDjITr2yzPBBj
4h03u3GsUVTfFChi8LSqX3YUIAGck8zjWCUhHLX/9tvPLLnBSXY3gQpvB4zD4ATwsYr0rLaJsPcU
rFAMtJ1XHzFzHWbs47yuXvMrrinLLvRU9pxn1W/xKvLrPM/lMAj0ujBE9ASdPkkpSH8B7SNhc6Bg
W8gPiRwZk7Jx7OSMu8CjrQq2FoJ++YTE7b7+M/0kdB6vCLJowhFyJw/QBPH21SiuTmo/+ZYeu1vy
DTtX2dk6X2Om/oJQUKSnJNRAlXEmgvXIyFB3QrKPP1JeZBUy+im6CDZqk5JapZ12Fuq5jyqcKv6K
yiq6cxC8U9/D2lIMC9UOrdEgfnW9aRICZ/ggVzMY2bT78XveQwfwyXJ/bX80VzwJV2/wQAhbsHFD
+NwqVgdfnXPcBhnQ6VEIVTJxdP5uz211siXIzCOGJNhXkmejYXXcydz8Ef3VrlwMlewGg7QiFUd3
Vq5AQWJP/krCF9d002zkTtBKyFK3BGpygfcI80a1GX3GRnyX3fI9YHeQexpLcBxEMEpxX8g15mjd
NsF6T0OvxzdQnb6TAHTQe/xpy+kULpxxO32FXuypomS9cuaIAEz1xpoE5VLjYtVyMc2VBhWDTkxb
j8QeHVcAGh1JgBftMMrfFSbCXnv6NuEMmHJHfZ+u+6JVr7VKggGfjGKER7GdPbCgfJYpvJiLvtVl
yz6mV4t26NVWiwP5bPpLe0FpgR3xRvXiCobSLNbt0tup5mj6qfEPC9gh8pr3GQsUnGC4pG0OjSSO
3dgE5Kst1D28FaotIinchGOBOszg0DvULBjgjQ4pgTosTVMxYRK3C7dOELv7Nw7HDnTPhlqD+iBq
My61iZsRb/C9vx0b7r6MJkB8A8+XJ2KrspN6Y6q9oCu+pUbQpfU0cpuA6YdaDjmNKuGjunQCFsae
6kSF6fbYI1QTZwCxGCIT31LCEciCDNeN4o8Z0/hncOOSodPbEEizV5oslx4C/UyEdQIbFRL7EXnC
hdwToBWsXh05LdCbAlaOuET7cTv6z4J4wieh+2zNQaHvKVEgN9HVOl+MSrF98TuzC+NnZKgbJlNe
gVNgv9iZdrWLeF1QyvuRK+w4qdaanDII2R3TfTklZwjIzVd+51DQFT77FP6c3KFsLlBqQnYie5nw
bFrlA45tJldGqmtLwHxrtPL9q0RVCpIFxJ9YTunLvMKOyuI8HDKwpMdbR4GU//cvAGI+kyHu4I4T
iu4YfHw1z3vZEjXA6n+p835tTqzPYDZEiA/fhW+FCKawMXafRiG0cMnbzcyGikPFeWcldaepxEtD
GsXsTWpHtKydp3e4Qr7CLzVdtQNgiYNFRrHKeljv2NpJyyl0P+S7nHwsaY3NjyYPUfSWvSDtCjin
wGNU7By+cT4Npf8Z/XY2+dhTRACt0eKjSNGlzy3WiYOIh+9d8yeRwU65Y1TSSouzt3uRo3MEg3bq
yEl8Zz8RNQhoUB1vs7ck9QIbVwvmha4rThIDJwKX+1/n444WsX7cnWvwdjofX9w9vIjK8Ym1KDsi
cvw8AxQf6JqnNRZoFhyjM6eGya2/xdBXhLSWmlYC6JFDKKUxB8XJZh/mDN8CNF8yHOw8QV72Znkl
TmKMq2KcJHMAlqUiAMMgaD6hbqsuASHGpSF0mWcnbEB24mD8Cv2NdFjbm1cnLBHRuNCK9/3PBWFs
XWFARosAqvAX/GwZWokD2PS1NU3DHL6QTkpbLI34nmMFPyVg8kc2J1Rm3cREKG/7rGYV7e5eImzE
u+rJordhDOAT6UauSmD/bUlDTIlGVDSDnltbI1AvCExTPcRsRP4upIZ8Mm3YiFBb3wCo3kduF21A
dTPsf4zKwUjPn2xmwddJqwz8wWrmULRA3zha77OjRosPL5wBEaAMrxVlxSfSuQgBw7tcYGJmMd8Q
n8RTnBNCWoTWah0GwXdv2RiYNbdJe4qPXC3hFk2FaolpDyRutQxTaYV47DJzIwkZ6pv9/bXAQoYs
wIc48biS/gvcdMOHNXTpdovprSAJEB+NXaFTjCBFLSv5lMtuozYI8whXwjJcK59TIvBkJEk/oujS
+Jq2sqH6Qa8rEIY5FwzyZblrw/s2qERIlui/ulO1Ha1BmVxo1GbJDgZ4fujyJBUH1lQrxAln2Hbt
Ablqpgwawp8MOwDsLOh9lVL27VNgvuSFjcnSLPvb0Wa1+c0tgSEiMiCN/Y9BOMqDqgsB3o2z87dK
JDkFoIse3jA82LXUJn8/WUhs+V22XqooRbCCQcz9SH6w2a7c4CvZt0P3Gm15yDBKWWTa6w3Q7lha
vwFp6i/JPP9tuYTv9iVi6M4k1rVCUw93lpAit3E1DGoPaf4xOAC78Q9a2eIbAqSZqz3IaegLhKPo
vVAOs5pnwSuL/HkZuflI+sEDe+UKUSCJAiNcV9EJtcPQ1Zmi5aNVSRjARitewk544jLTeJDmJ8dT
FK95KmQbs5ldO0yvozPeKU0HCNcFZZ6LaBZDzfEQBrjbzyT060GFr9N+Yr6L11+OFJGwR5rKbKt3
MdxTTyBbepwmS+Ew1O/JYxaxRKUH+gz3kXBvyK0vePkkRsBLnlQKooAWPuFrLzNJGOk1047bQjE9
Zj47D1olZyP4F+nI7k3R8GcmobwJ7sWS9uwdtyhlwBh2v7docGFFbll1SlCe0AGMGftYClOFkWla
qYcfN5yiTAbtWtgfwV3S6AiJQhbedv2h3yZeSFjky85nIBdbaPwZQAcB6ZbIScKJmKJAobmNxKQj
qg1c94Qgns8nsT1n/YK+raFuJiO1Q29IoVOWnnnnWOXGxbv+XOFV3FinxySISFu9qPGLp68PWENp
+6XUVAojLGyndMsVb12M0dWvviMcHjFgp0ck5uvTT1d9OrJMG8dAaBKiyVdD4kWvExb/Y4ZvSaSU
nwFor9j4JM/x1tvppiW5ThvM/hsUk+JUrUIDYmS4O+k0arYQLE/Yz6PGybe0h8UqKo57BX/fxdCG
+0j9A3Rcg8tNFf+6p037muNQNTsZoZ7v7sqQ2qnS+fO/GPQtTdanckKxeAztYsnYBUOqwBHBTfUb
iAjNETw/X/xyft7eOCk2YSxA3Urk7ZyFxS9cANBOX0eV0JKSCRDSrbALgeOZPWeI2dUO2Tayd/ec
R8ihn4f1wXjb1bQYsdTkb5RDcTzAQt5UkLjixteye+EFyyb1PVOtasV9UA7gpm+Ou57AhOJS1o08
k9Kt0asWkSho7aotjK1E9QdvUekUt9Z0ZSYtp+zvbFUnvHjuTZIF5Qb9+lHzdyDfGeY0mwC/A7cM
gCiDIq6vhM3FBWlUwyFMKb7JUJg7RJYXyDOcztH3EeRS7R+dSga6xb90ERd0h7VJXH/AEC1A2S6o
1zQuQlxPLjhdEZ7Rg9Fk/EluTFjezlgmz3BaplMZwxoR3ozvhZRqSdI3Hn6HUa94uRNCTLsX4YuF
BMMjVKdBFxaJhH8zMeT6+AXBZJZFKB5Jf1GWY4eK8cF4S/e6oXMCnBQdD2dwiQA3vWEN7HR4bEHm
vaspLVhwpfUSsRthGW5Js4KxcQqP0wUj22+H26WY23RD+v0wx/Diw2DdZ+PCzWlPvBGtSu0BB9r3
VO9hTjo1w5IgkBgGsSkwpYeKT8gR5FOByTujzEbEOABqWcVLBiCGxvXfPiysjFzridoUBRg+bGxy
fbr7Y05/lBWqS6tVBvlbcHQqhiaFSQnifT8uzfWg+zqzorZ7CrEwvlZk2dvkDM4yr4Gk3sox/nI0
WlboS+wgXuchbHXosBk2NU0TbBIYyABbbPWsBubKOZwI2r4ojlneDIAj2ilCBvTAnCy3JQQbvkHq
5M6leNw37Y94iTEL3RveJCivokrXZ0b0+bCEdebuJ381wTesumde2WzdQuzF0Bbk7OmpASYKNgx7
ogX5BFoGDCX6YVx42WjKldDby0p1VB1HsA9wzy4VknMri02i9Wk8UCBn/MxRKgqrJbWGMWSk2Wk2
kpxiunmlJ+xaTqU+mzKfj+hpVxcDvnqrx8J4hQZtaS4LSg9xzmchDCXss4FA+THk3JUyHVNtUydE
QS03ul+p1CdDrw+Rf6vgd2RiUoEmYs6GYJFyb+ZadOZ/pDF7J35eOec6+jYFC2dtak8kxZQrO8yT
79KD+KDg057h1PSwY1NtDpx8qY5XkRvGZ+Rou7TL1LRzuRj/puHey269bkm56uJiHH7sdDH07YB7
dFtq3xvb3jn0pJma14Lyo/zRZtiqBEml+3qh5glXEqYfpyFNDUx/sUvEY4RC+4y3jVC9Ic+O5UsL
xafkyioUxX4lad+fmpiFSI9x1TPRTjgArQdYcaoq5i1BdAW84iCq65lfhFLNeIwUUGNcZd3ZZZ5t
uqaEx2QRHQNXjw7QDG7cYCpbQhmuwPlg9KvNFmozhv6iUZNguOURbAn09llTU2dWoREqpxlg0bHa
yujDWvrFD94j9mYhHoh6pLFgWST0JqR7phy910tKmjhGI7YHGke+sHNUgHmyqITmoZXn2JvLX4wr
UtbyLM5f4B4YgWKcih99gynPXOr4LdwFpyr74SR8KB9FmILeOKqrKnq8W0R+YbPl0Yjuu+0DdGI8
2k5YZ9hjYfqTDC5/hJ4XAnQIgd2ScaC2zpoap3NWJuu3bg4hvGaT8PXqRLe17g0tFUaS1oUaoasL
JvRqS7zqz02iWFxkxf3KuP0MPeojewdWBK08rMRSDXHSFEOy2qWyvUhjeBTq9B3BtAsyRIQSvUvC
+J6dGCHGykzKbaHpEFBON7ia/rBAPgh0ZUSGuQYraOILiXc7joN2c3PKiig5/NOfRoCJ1vq/+OYF
mULdP0m++4xScpDGbCohqSJPAGPjEVUdj6Cpmy8Xflju6HgZ+gYMu23EO5OsEGrOovAc6aLf//bJ
Nv+W5ucR9SYMNLxZdNZ+KLLr+uneo1BCeHVWaEERLWiqNT7WYt+xM+v+UrfRx0w0t4GdHhQf30SI
0eLWzB4AVLRtvXzTJs8EwWH7mqFRHuQTyw6CmC3SupkJf371mLhRQnRq7sK9jit91HmjMEu0agn7
rgAO1wbMyR5LcVcSbZweDc2cxYE+dBNmtAHMUFXCYEiMfJTmsSaae+R5lkVA1XKdr7OFbn+usBev
lnV4bURQOltECNFFxP/0K7GC2QgiZGwEdRnJIt5REJtzEkaW+1hryxjidQWfxdV+YRzKzSMLEXqB
uLf2krOpdi058ADNWqphBl4O8sRd0Cf9c1xQErO5EJmivVO7owUaKf+ZiLpHJmoZBjYdANbmFj0t
6f2jqKvkEu1r/GmNDi4hh3DxyhGrJY8KQQDv7ulNYRnuznfHMQ1ZbuS3sz8jhj4D0K1/mzvEnvWi
QL3nE+nCBBLE1yQGpWoI9dX/CX56KDvRF/VEM+ZRi6y+F2CwH0YRPIsbE/jO+iQ5yzK2Uiuesx54
svA8oQpE4Ez8cAbSskIO8wXwhcKM941RmcwOy9PjmctX9nhwhcLVtg44Frw8L3kzuyBfZ/MbGYBR
YW36BmiveVpwXS5hfcyu0OVUYFa2F+v+JKayLyGfWbNuqbJPCA5ldQVVIzf97B5axZhrPnT4DJtn
IMx6CiO1Mgt998xI0FvXWKNn2S+ytfQAZMKhVxTXe8fw6VO/LK/kqz8thymgiJcJbxATS+81uimt
5itmBoaGfVeNkrxgOf37Yucph7HKQPEAxdW/yoOH6lRDsEtrw0jc1H1KawCphtuOpFacQ5wBZx/n
/0SpfUdc/Rk0HeMqNW9REp9Saa2fUCUNCzZe6fxOkp5Q+38djiSifl3CRPjVd2hizjVgdP2lJGv/
Yoedw0BBvDk4N4CRXSGN2ptdsG/y2TG5+/3xEDE4pkmmTYM4PLBn53b7T4cKty0le5fYbsdDrZml
ekkqKzjcw1TVxokUtNZsfRMgFa93zvz+X6Un6pITWyXPF52rtkPdfLYQqLioFYNYemm22BXUOFww
U/RgH0SfcUHT6oKZpBGsB3MraI6joZHv52zwOPS/EaevJmgcUADInFJKqVgjkKtxl4tnjvEqVQUx
0RbIvXWocAVL45O6+o1pyNm/t3cwfMtze+sTADKZSVFFss6dziNTA544nfGa88sxr8R9i/mCgkhb
FHOJM94UeNU93WBhLHC17NlrJVJ7uGjHnX/XXWgPZ/EyaFMjbwjscF5a54r1pHlSQkSV3ZPSVRQi
EAbpcrfdRXDNYik0SithXz9Oa8WrLbG9pu/Of4VRWSF2YBNEUF8/Ah5snr5hfvXQ6NYJMiFIzyaN
/co2RJpvUBsZNxxLhFckVHlWRmzimWMgg6JSEFV1ZbqTyUwrPgMt+r6zVTNVuCfAVtynWoTJIaFL
nhJMsPalQkWdhn+qUWm+Mb7aMmJDOEvno+Q0ps2xwsUEgZfcKPk7x9KMJF04GwRJ+sXvTczGRS30
G+XXB4SPSyHV3vqmLHULem/PdXJ4kEaYdWlc7UpkziyJEbdOzko/Jg3ysVu1rnPYy5k1GWt3Gj4L
ADW6h65zqP/OUG8p5zV9Iylh1cDdpwp8ZhL4YCx08RRN0JAPNRh4pgdMaf4/5k8sXnrTHLLnkePR
9uQiC4QgXPlMKvKYtgXnhm7p6XM7Etxnwfx9SBAIWNVTkU03B0tfp6ZN5H/fVQPV3DyylqB2yM/e
CyuHiiIMubww0gy++nT5Fbu1hRb+lKIfIYBh63XG5OOqrHjiuWSfmLGUpNa8EzQ9jAvLBMqm1TMp
Alqtup6tFP3OEaCn69k41tsukEbmj6eYvCk8sJQG+e0chgsgA6j1DBM/yey1A2H1NqjGm2c8FXLv
FpAjRlxr3+YYjw2E0SBgz+yoWCIuh4BfmymjlYI4LJ127kgTzdo97FUxMnHa5Nb/XusTtiOQaNzv
Y2H8sJbwnXltlhndB/Aq2KUArSKTVcqMt7u0HzpZGBRxmISAMGaISx6DmHy1lOzAVmH4tc++pgaa
N+e5bTtj9CGZkXjfHLrAISKPcUCrcwiZhvjJMgcq3z2fEA9t3752VoKq2BR8/NauVasVwdhQwoQT
ISWA+gpfmdykKT74Ixe+S8MjFSa0pXGG2BcUwMtujJ3k7ESl0DC4eiwVYycuNuQQ56cWOgVKtZZ9
d4xy8Yx8xIRYAr/Vi2ar3INs4x9VJIFBe6WiXbBo//rJspYq3eSnHwPulUhTvAl6Dn0PqvphUrTJ
1wZo4zKZT68YN/KVhYObJjJgjD5fWlU+GP36uWrezwl9L8XMikzwAIV5+GmbL0L+UcRVGT2pEIs1
Nzc8RZgOlU7aS+S/n4Nj7dI5vikMbb9CE1QzCY60o0ywSwwFZdY40d0x/rRp2XT8QccpCso6FcSf
2xqGXQFFLGBl638UfC6oUfFgysGLlPCFcSrqDemubAjtNZ1I4J95a4W7omdK9fMPebsdC5YQxwL0
8ZCdVCfhFqmyLhhEPBQIlZbC+k2ROAAyvVlEw3eHWdEzOyVOURJ0dDOMk/8cPwpKAax+eAaKLiHN
w25OuSBp13QU1xYS8OhXpnG+fonKecU5FCUmvbJv6P0mutZXFAfVHQmle3YPWgxJbvxS0v34ICnS
9JlRfy6OL935BtNShLiybb91yXU7aXwwzewNuHWYLYu8wi8m34CZDnVR48hLgH15ly/CDUAayb/E
VdlYgqaQc+bpzA/TssIMl6P7B5PXqCDgTfMtplq7gqjI/GPmjXpPUExieFdEF08yCI6/LjAHc886
2s/RX1ftGbICQKhTcEQOGEOqpmA3heceN+iuFVrXS2n7yJGsjyYySVLnTL9yeePhb9pLjQqrE1+V
m8YC8E32s7Ygjec/Ygc8TzHMm872gSJfLeKQ3H+miqLaW+MdQ14BVt/5GaSuSoSeP2n/cKwgeVRc
9B4sXxP5fLyvmEaCet6gdEYFL9e3pIX3qlDW0WoGTTrSE3qZF0qh9gdaBfrj9hj/FGFaL0SoTO+w
rP7nto+3x4d8Y7CYs01lAIWVGlI70jKVjX7JImutpL1DS7xDXGQs40OlK4GmN4g43h7KkelBsYKB
skI9W2+NFnsfSG0f/VDWupF5aW+CAT+cUN9Lv8CxtM5NFFlC+fhB0wHHux2FRnZGC0baWCeNw3iw
RjggfEW9LeXe5T8UzfVqKFlJyUY2jsixNxwF4getiNvpemfaMCB/Y4jDQxnCbqcWUPBqodUNt3tM
QyKJcGvwvbOQBY6K1lTZddGZKnmWf+JL9SDI6TpInFy5P/XqeFu2sN9D1h6haTKk1TiVyCGHvq8H
5Ey41jlbX7OmEO5p2yMF1JJlRurexM71z2reNSgG8a7cHOUAAVr0fRtGXhFbZZaBMZ4I9Svu44Wm
Vcn+TzsoQ72kaWP9EHjPFOt5YEa/AH1sw0pYalMLUGmaDrCMSeY9ZmYcB66oeQqbskbqijcsaxoR
SU675SxVdl1u0s+K9EhCr8uQB3TEaORNFiA+9oRJAHEMg7PX887W12S0uOFw8ZR5h1rVyKop7OCh
zxiTnxwKVdkB25JlYwY2zxNwvmNFb0YtwDFUJ8EM64XbUDTN97GU9bIYlWc95hUREFz0iFaw+MDQ
Al3jF/NFPPtasfxwh6WYNB6WrHRte1zV+enannTDLxPsZarl8UhIl+3QuvhyXveMs5t7RE9qTGvs
YYWkyLKw4QIUbL9VmZNwmIJV1AkDq6mUOnvO5dUnSFtGJpLGwKB9m4HuYaoUDSo+IO0rHStGs7BJ
3mEpKqw4EwnPMXLjy+Vleb2DkOblXONKLd7Jf4c50p99rAnfMQIFX4o2puBu7kBMHEg9mgj3KCg7
PnrcBS6PpSnlWJCX/E/YDkPxT5CvsWpzXLNXE/+G28reVLTPKqxs7sfHuWOXrIItGTYICvNr+nHI
j8/H9BgvPJCT7RewFcMmpFMbJEWPtZ3EdAISemEPCjsJR+FlhG5WHuw//7gZZS3DzVFZyhP3bqur
NF8DpT4s7R3YGWLK0jmaoR/DNH+MerOpuvq6nNtJRGvFaZzDWQnZi7q5gptWJwVSSJ2A0ynBcziv
WoyWR5cGrWtkRip5Hu0IWfz+SaMDnehgdEc9D9eR6NudDnn8mS48vnLlDVmKm28OrAX1sKK96BLq
Og3x53ABQ3ssPVMvKUMPC6UNCQ7leVexqq7cuTIsx5sLotORDBOHSb238q3U0yDfGq2zwZsB/Mz/
qbCiqdonO4Qok2tNnbZGFzB6NibNsoayqJve+vCtNaCfUEjYGhmHjdNEudSXmJebkKXrNwmIcLV1
32waLUpVus8OrHFPb2J4T+/J6dOF0ojGU+VJEMuFQHQzpa1MvuhUM0mUEGFMTwsOiAJuPR1UaP02
y/oBrFy02JGfXVm5UbJpYm/AqqGjZviDycPclXyAV7VxrNS5YcBgtMucPwBv0pWBIUThaJH7FyNA
fvvwQ+kxJYka5t9YnYzJ16HiZAYIU3vYqNgLgZAU8pPVp1/f2SDZrWQBiDCtdbDVLGC923lXZf53
LEmJQjviHGDhU6RL0tDnSeLASva6D3dsrQAuLpwpZUgOvMvyUNh5qxkb6ejDuvzdovt2VTALqQdT
baCcdPPrFB/32gADi1MPYSfPTI3bFogHkT2bNTVtAcO70mGSbA7QzZLApubgcfgxskF0pxxMXzhL
iT5doUNn4+mEuugrZsnQxHDEe8J8J1SswrAZyjg7LiRwO/AI7ESoR+02ssYNEw2uyTacHmgGbKMq
EKnlusjKEfH2Gg/IdmX7yACVnJzwZ/exZOek44u6MKWdEPvN9jKk21tzUIlxGc0tksyWJdl539fN
KzFEBy9R7G03cBYnn0VAzmcjbgvDU3nxkdMMhKouWgaxJ4ZX02BaNIMJbqs2306KwhAq5SPdfkuY
2Iwsfc0rsJ+YhH7QNMLVRbxnQcscxGrucNlVNuXGVU5pJJG/skumk9rmDGkFUFlLEx/tGc3tocWl
iB3swwZ1gTRssGcsKPi+hzXG/hXAo4JTdSDb9Mmjt3NhwKj5eqMpp4gETsAuTklBSL1nSBd+z5HO
sMNxpDmn8OavQVeHsiENEnnU85JUPGfrCwIb7q711oh59g5TsoDEwGeHeV6dlxWB4Wg8uvb1ZyML
pawEj+1N8lKSOq6cuI7iIr35Rtyw8QD1XtqbSwoec9EAWH9CDf9vaxXLnhy6z4vs0qOQsoBCFU4i
ZGEMUX8SKoy1M/9MiCuNaJZkvdPEMogIcNDjorgdFGzsYjQ5MFl4skdTL1qoaziLTPCQ13LOqx4n
VW4wzH2wAXFwfbkgTY08+ZuP/9HVQ+sn2oINsDdXukmFGZUSaUZNqVrNr+lh4dH2oS+G4fiTYQgm
a3dFdHxdoRAX0vi4ReDiDB0CfQUQcZ75ySBUcaYyUrBSr+GYKMaCHK21rTZIXNQBw2L2hQ43CgDK
OWbRJYsTI7NQKOho13ttddFCWPcyKgCq+LOf3Bn2ZrhsmpNanXpAop12DDmtG2uu239Glxi+vQtQ
Hk+xbNXz4IcEVSSRKU7y0clMXZ8glCdNfSJUwKrlUpW8SbX/CWel4eW4cVFLwMvUV5DmzviBVdsg
/nODHMhIEWQoX1mYG6LVCIVXTO+PJ8bkruCwsUaxFcHenCqbxjIX7kpN0wTOpRsqj8VMct1CG2Un
j2AsE9i6nTIKXfuTrztkNABJc0a0wq/uplLqH1lcnMLHStmRLHjp1jBJwGcpqkp7wNZ+fxa1aaz1
JPTBzKePoZgg6mHGcRZpl3UllEb7eFQ25ekphGAQAuEgIZ617lhP/31QRWZv+3foOs56CIov3FBj
d7btLf/cffr2ANe8ipw3MpjrPRS3tPh2Wbp90KN5pXaZ2HE6dxDmDJbOl2zIa7HblqIUbNEY23do
6UNY0GvsydCYRGFYDB40OepRkCe5oHk6kCwrBrFJZo6SZerKOD30yIxBpbF3tkYi0n5mzEXEEzFG
BlIdiX4naU/W0Bjf/S16lhmxg4PMo/hFPGQVjzO09fnNTX5PeE8OElAxUgGi+eR2N4f1kipaz/uW
V6++dTTber7wO7zh+vhgmB5l5YP6W/QUHcfgQ5o/gzc3mGvDPMhiNq/Sh6mZck+C4kyemEeDFMy9
6z0raR7bEL21BuiCeXuRLhg0faWYGhRWVwQuss08EiRf09i0nXE6BCpDdptw1dakJ90hLRSgFYxU
GjLIgsu3nLKq7QTbE9WMb+wv5mm2EUaPWNKA1m4IgLXcEh4OeIt5MTxbDyLIMMlka6QTl1W0oOpR
ofEXiAtBv2KTr5D1y39VyuwuzAHnD1HPwkTHhNPAZiPfq4hUwIdcBaLBpmucDaEpDRkN4qkrE01v
kMA7QX/ZIltrvTrTs3KPWSZ8S5nu3xQt45zfKRaNJHcZbye8hkRhqkw9U6SQExo03VDjseKa9rVJ
wPZZYtlAHFSLzjSLWpUprmwiu6GJrH1CywkuwvtT8u+jwofwRWwBdthAWiEkMtUTvo08EtJp/OGO
q0wByXp4bTtED4tWLJc4gqBklvC55HMkNZmP3GELnf79Qw9WdFSkGJe/+he4Gy9HSbBr/5c3Tblp
B7L//I+pQStfNtGqesbhCGh4gxYQu9PAbY7/hY3Yk4jkYprPrdT/53Ve/Xb0EbIdNY3yLnuPkwjI
OufPqplVPSdzNgpfmF7Rx3xJ6JGkrTQ5+RhT25FQ5YBxe2uvDAs9P1E0jpgxwsh958KQJ4RWlmKU
+rmoQHguoYTCycnhhL/Ohtt//C3l4TfO6nA1g9aUB2csvViwTbyWU8hJsul0QUUDKcXRVybum5vG
8TrBZZxI//c9KzXJZLKZ6X6do3VdkJifJiVPdNktqTlAw+gLJJ8zb/c1ObHH3KbngwClxCb+6j6T
1A4mXNyD953ckT3nhBuynT+FGxDKfZiMxwollmpFYNqoTA68U1Ixp5huIhStwfWNxQ2FeSShq+rC
dzmMppstJQrKbFvXP98Yw0Wy4+7jR6FnvuyaXpY1Wy+sU0PLAlj4z1gP2jsRI0u6jkhYchsPE/aV
wF/TNbdmp1gmESRvRoEj4VUSZ++yN29TtjcXJnGMe+WOx7zZNlXq4Ek8kls3EMUlCO3TCfdT5z7P
iQ/A8NQnq2cRgm6S7ywMfyS0KVR5rHpVDGGZBI0hSVKpLEYxUxAUdlgP6ZLkhoPEN7+0hh03zdbF
lCAWiZ41KaTLTLvk8kw5ahB+7DbOI9gljP5b7G8UiQnsyW5u84gedbBYgjcpSY+UV0wWzaqWyrr3
Uaog78zwFY5h/fyJnWeU6JCiAn2hqlwVVQfB8bZGYDS0gWiPOXAyv9Pdsv9ptyeK4NuEDHsTdZ33
hg80EkL7RyDnI+qxmJnL94x6nWYfv7cK/oLXTenz8JqDAKJG21ZcPCSohR0+cY68F3f4IhM78p9x
oQpFMQlenH0gU55S9pxadbAbzKz0O4Br0F/faABV8+PhwbRE5Oozqre3V4JX6uSO/IQHU8hKqwig
oJZMgB3f99PIoZAroSGu2O1Cn8sQp6cmBEeFfqke9JDxEK91x3h9C3j/hu+alaMEDV0awHKKMqUG
ZHfn5g6jtJ9i4u9nwS0I58fpbOnhB/Ds+cLWprCGphq6BUMYU1HHDd3he89dNPJii2UF/6XAeGig
TQcl0tNIGe1Iqk8IepgmV/ynOHbbyfeumk/DmcOSHjyXdvPbO5lspoXS1R0Kkq9mOTGqp9O2XYP3
v6PqLXl3bZnPHzmyYKOytsyWqHIWHZ+XBcm8DWvGalfd02E0K0V+EFzvt3KFpgviOuqUjSdrxmDK
3n/4Ewt0OV3uqUgpHzei7vWBIeni4LtP1duajxxmbKmIxVA3upBk4Zpf908dCF37ZB4xRJ1jVSfB
yRIzIEIgjJSP0JcWYh/o7dojFys/nWywngPozTE7PvxEjodE9CApDrhtwoHql3Zdezm00+bjfBUv
5c46xWcew77Pwcc0ptmJraKQqYddZr7MwrygAf7jXo3bF8Bo0jrm8gEYkNg2R6EQslDNmEHK9uGs
3efV0pDb1QYQn5FIXQMWuWAkS5h22DD/+J07hN+yhawqnyM2ZaaqeiHUMz9jUeNeJqP1hx6itfwJ
RWtTfKMvGCCQgNFmbo7e2ogvZ7fjzZvI9hnd3S8oJp4IFZ/d2uZizMPBNbv4w0c8L2AQ3m3A8Bft
ewQ6pbJdThzaDoMxPJ5+zJpqyyzZPR/WmfQXd9wtUOPnXcxtLuiJ8bxwznfYyw5lAycDnzLzyRbj
kCesgZ1rrO5hbSBXBtzwnR/2TOXzNhu6iff3BufpJuYG77reKI0KY2XMXV3hbum+w/2M6aZeWgCS
DMKFQbWWCDTDFR80Kwxqka7U2oPzBj5Mw120UGzYY8fusmlp9Fb3sGFK/aWOGbwoh1N/GbFiCD0e
0Fj/ms+Ic6/BEq+k+ljo5HSnJ7RW7LYGwgoU6IWX4vhgqvTnb59jXAVu/YsUqCnYurfOE5G3pR8C
vsRYw659qL6wleHhuqQQH9UqOTt9/slhLRQ0L+/PnKS3RNfjahdmeGARaYR65ujmg/X8ORfS+gP6
wvOlIbR12fHY1tujGHgUHo01/Pdyt6tEMVhr4n+LeMqjOtYj9LG6pAtvcmMJzDLJ5TtSJyELKcjm
tqEoKHpPMTSbLL00U7jj2tPOXI3XkWjJXmLhLrfozXAbLBbvoHZkQmot+o6a6ipkSUYF9zCvQMXQ
q2IVc8CACVlyFTi/i2YixUjwGO8iZMzb6buKn8cmLxlQ79VQBxAVDsioMsJ85kETMiIkCOqSYSTC
+2jOFVcaZdqHizaROIa9o6H+euzUSXPTq+85Z+D1xZyQzw6OStyBKaxLgJHhdUgtfvS0DFcIHVkx
+QappQZl38t/1uiFkpZjhsemrg7mBN7CGT3SKwJdx6mjxZsl91tIzDxAcWa1TdmudqdTru2fqVUI
BKlZ4UVl1NSeY/UZbUsdpy3Yvsu/5Tb1LjdCbg0XFuDhsgfy4VDpnn64mMCRMHdnD11TB7TOpLZS
2jLc6Xuf1wL58kOfKqbA4CTtaGhfI0nEu/V4y+7HZLxvz6THxf/m86v1cUBgMN7WTNC52k5CkbXN
g2Oomo7fwl69JMXTOT9bvOu6e20PRRB7ziAoZT9YKxo0IOHHB5/i1zblvc6a92u5HzwvIjaDtCnW
TcSr+jADHbNaOnMc6L4ckPbIX+/nwq08RGa4wxE/bKsFC1ewEk99hYA3ooKt/YOc5fQPrO+xnsS9
MPvY1Fl4oD4S43l+Sv/UL0naxGNbKkGEdkfRN6ZM03/yYEwiCbDSc9B+fXXxHHQjAkn0jMaeT8vI
J5JJWT/BMxmOYQvPjX8+8JYYIP9EyqW/vNjO//ThhYWpaJQ3fBqWugsR69CM/3S7da75ZnUE6XnW
q0I+ID1F7atOHu+mIbIe7leG9+O9QlsOWvN+W7GQpICSjM51s20ovIofaRMc5k6N4NFKDIAPVWYb
FlVZUqRNtWLkmOfU5Lu7fLvcaL66Ol9y+NBj+BaZEfTBo8+rS618dCj7fDPVw4DLF7RT6/eDK6Y2
ueDA3WuO+lqSTN2XYjqhnNSERUcu6ngSOdPUDipqdCLXC8ga17ULYHAxh7UYwBLOx7qYWRyCaHsu
GgwDkcECqU8dFBbSN8jn0bvObf35ZGP8VictISzI2oJvEC/rSKtqcpTq1iG3Y17VKjjIsBvmbbhI
8wBh4+XgDYEusiYqqxrpj3zilqEOTAiV0q2vzl5EpUcZiAVbOKQi/BjD+fCK1XqD2JHb7OEs+Iyr
58Ra6hxncYhLZ/6HKdtdHC3bOgstWhvaFhlCOZP44vaUW0QGUpWvB2FeYujXV/kYjnMfJbXJcUgR
Fv2entxFZrvoYukN8Ng/ejIeCtdOndyhbIToL/IoF8znlkAq6IsZZMYkuIAEY9NHYjiK3lV87cYB
ESCnJzci2Uyxjag/0KGRBboKbtqHAYM3zXGLPg6pDgM7FPns7ksjxYoG7wIi6IFS8lT/x7hR56rT
hWTzVi6zln1jw6S1b/J0xDX/QCMgqP8bPw6IKYy40kL2b86xTrM4BcTQtPYqZOAHd/mgaViLH1Y/
h2GJz6/1DOSiA9tD2BBS5ferugRQG5u6iLglgV/rqTgMP6KMQZMsUandH48KPlQ+3u2tHIw6Jwtk
FErRx45Okvpxok/TIGLGkXN+FBM/pFK1LSn4cYqDisc4cFy2dJbHlpyWkmkhFoDM9PoPnnc+sAmR
839DoTDBzeFTTvVPSPcSAcdcEFvLvmnjAQH8ticdSnHqzde/FmzTD81REeozXx1LZkrkO8yivzKB
V5lH76lgI77D1ZHTkmi32NQhiYYTphxKo8YFTaUFeYUc0zDxlp/3kX0xX8sEfrSstas0J/OJe9KU
SkPdI5LlBKfhEcQgGSdfEHUZskS/JZ7QzQ3GvJLmysn28hDDx5/Ja0iPint/x/dYzDiyAuKURTuN
9OSXgPP6rT0jszqrTbgzD7vvysje+Ar8mPqcE4cXqh2ueESnY9xRmO2lTozVze06JVsrM4YujV51
kA2IQ6qeQr/QXE+fs8FZtNzmFaj882CgTgYPIpdwgl87owmbm9dbIURY6bi+tp6DDGtYcii9JAZf
qGnAKomJpJ0kau+c7EPwn0h6CMT6AociTIKt1Y5eJ/FDMb8ykuI38OB9wUlziePBNuYwg5GdyFai
dyqlv0WR35YfWr/wu5OgKDSbuOoSQa5hU9t/MPYXiDXGmL3Lr9gf1kY63RnK5Ym0SSwqP8YK6Yor
gNdZ494BpQqqHU75u1rqWd68S6htU/vU/H+T//Hi4pVrEouUfPtRI2GtkMWdDVT5bpt9ju2zsF5I
92zJs5BP3Snl88hLRD6UEkuNA7bPLzikzn805jWiweG6fDXFisUj34gWqczvN/RtFjOo6ShuiQwe
tylP6RSf78Z5R2ggPFVmLamukfMPdxrUdTgjeuagZPcHJihKMZdpXplF7lxHWI7V5Z5r9xhzDFUb
mh4MMcbQfCt9qy9i32FDN6UUyp3WwTqMzBEn2SPd3eefzkxTaobpbU93ZgXaGGammHA+R0cnTIMK
xgCKcxQZhsAqlYZU1r5PNhpWhy6BuFr9AURLjKJQBP2DzbgkUIo9VOpmeZLJkEnyGGsK0F41rXtM
VOqk58XwEoAxv+Z6Gq+secopifweCgaFvcEiSfQQwPv0RrAXoSckv46RfUF4gBsageYd0MftrJbJ
7/lgCVoVLcUPH4r+SqIMHCtXed+z1UHkjGmlp6l/8riij3nBj/v/3hLTwBnajueFbvCA7hegq+JF
2cPHqQNCzXiLni3oH+lPYFqMy6+OmSjS9iM6WnPu78R8sAw4vpRj3KarUT+rjgea3Syv/u8Cfkq8
SPcL6fMZ3mtKwTj2aj2NLy1ZNLORyzLMD8RIHGmFTvTjaRUxKh8i31CrAot1fiGPn9pZyK8nTpZ2
eGquw8+BUIJeGCdhYlmP4oVYso6zXMMTc4/Qmsyk9oRkn3xpjVG5QGGNjjFAglmzPc3xoGIp9wCz
R9kc8xgx3lt6j3PxqcntFEVGDaIFFd8Zm3bdl9vkKqVuCsfR50cH7taiLuVf+gdnjSN/gQKdL2nQ
mO+RDOP8t1O6NzELSCLM4SRPCeySYB9cCXXYHi4ykjf1ej2LdlhEB1W1mRGzhedKGYGUKMtVZSb1
Ct6tIhLN/wLUHvHGGkcv0npRzocmhVwjfm7iPYmQKIZvSE8w++5aL3gUX0OMq36yCj9dLhVIZbx7
Xjwgv6HsEcMadeoPkDc7A+axu0D7NUrP5hrQMn3xI6LM9uxk9JDoUjLxK4Cbq0WmAg6KBk40p71W
6PBToZuz7CZc544fRFjZMQdOtvZMteizlalIFUkmkYE9jyNxW9SkHWNSwTsfIaDYU9E2bsMOkjFk
jtj0Tmc+2eg5nuUABIE30mMMoTXYJi2f7+OmS8aWyVczzVSMMUZsjBeNhIW30R0x3PO7f/CjspBa
GOUFdhYDtaYUdhJAimmvVZO8DAVApz/He7YGWpK4bvvHapF4IpjTsxrxUdNqrSB+bKPDkPGWySg0
CuUKqFUxeKAVQyzriKM/4mBYvvLhAc4Q7zPDQWrIaW5TwKNIEr/QSF2+uaClnmyusjw1BOiDqUbZ
aSyTrqHYnvQ4JkDgo0AQ1wEf96Cq+fiszyVcrBXBCnN3tew6QOq1ioFAFDYkIGK1U73j0JRuOJfC
mTZdgBvuFHAuQsxo/1mUH0igqT4h63uowBlYauW+uIz84RoRCEvW4gQwQsZxWD6U+m+v510/ghjP
ar6eVUnXA2N33vRiGOgf693xGpn2qdT9iaC73GyP3q4S9t+aWIowaOfoNPidmwfnbbsOwLv8RzOT
3YO98E2mFqvURi/yALOQ73lfDns89ES98cTLeVeEheTQoTUIPjF3ufmULKicwCpqdX7IsewgBeGg
7mvLd3Ri4O2pyIBjKnCxRNKzBDldYoyhtTHA/NKHpr8+AGxEgwormmLgq4WVr/RueEYfLe6qnX8S
LpoTvQZe22BbTOxC1ztusATQpnn7oPnqKjLF13pAy9aKf5iGXmFIwwWXzx2Q4m9J36nB780FF8zd
vaFqoMqlGQkimMDJaexsv05lBg7P0pNkQ+fNra94mysOG0c0d5E3saj5YK82GRThe9ldhMHgbygz
M+gUZbgBNXZYxXX9m22UK1LeWy6Ok8LnDmGzfbL+w3d0MRxJGxBA1dGgh8epP0w4NiTD1IdhDhAM
W9FG5lC/B9eqaS8uDC1Cqcqaa/uiyYE6adzNBZWz62RWBx4xxlS5LsHCjNT46GFDlr2+FtK+zVyT
ENLHL7ls1SsBJdRMf67wQetNQlJm760bYpxSagkKuEq0+xCg2gHpyMHMpds9N7QX43GiN88fQQcU
r66aOOKIjjkelYAtbhlUOICIPiR3NaFVu/ABj0zMNsCFCuN4WVB3OLxCkQCwmlP4nNdA2DGB8PJ6
TIzrmYrcX0WtY7PVdVDfd8mYx6EIbCquWJFkLx50kRxpN9qVxQ2v6grsOUsAJ2XMYtTPdbMVFdt3
tUxT0xUvcHM25sWASVc1NJWycO8GWIqnSYOQyrAQB7zyvKMCdgLoc5iZIg8yaqf1H3hyAYDWEeN6
s/NS9jmD00rUW/o1ISlh8Jp428Qsy90QIREHiJXbaErwIDmvcKB9vDlYNOzN5m0aqKdPAofEmUQj
CV5AhlJJwJxOA++eZOA1UYaWGNTO9LRXuSGVa49d3LLEaERR2cyjXsu3pDzlSuPrrVGmQHy04O1K
zUGkdtt5F8leZjx/C+wDM+hQFTScb98Bze6X55Yy2H0/WKl0q5Cc/ClAns5o5UAVJMa5gptFYMoT
JM2rM7azxmbxX5/q0KCr3q6GEvtqThJPO+2pg7C9SScx/pdIklZV72vikwM8GD6A+xhg9vT4UoCs
/x5flYgfMnEC1Z81l9axj+DzhHa+7OWxxVxHwsG8lZQwbe8+Bqa6CCMccfGVfiaBx/YDCzLxWq6R
GZGzN4dq1XiXfqsxEyI5Egll30kLeDENooQ8qUKuzpZR3VJCmAS/H0JUC2lMyIYDhQEyRBFUGM+c
mv+6r4IMGl0f1eYqBdBgzyWNeeyTa9o1VFCc+IEnP4vPdJO+LuQn4zrZqKMjI+9eDGPee8ayvkhO
HM6kzWjaDM4cpSz+W3emZLLWmqZrbeKTjIBWFhWqgV0XLlKtjoXLPE5ZUPOTuR8egOIRo3HgqlME
rALaxaw4dYwHXiKzeWTJuzCSHpHG/Ucuq6Vw6yov8OYCZk8JeZuaAdL0LrRRPz2lPxu2TkssKXH7
AgJ5sxnjA96aGbdFHWbEIsrhV+cfRFzX+b/3DJHS3FcY/v8kgLPVn0TZYBqzlUL9qkxTZUpBHJdE
Gj7xhYlmA++P2tfaPgHNPJZMl/+HilmMLqzef8cE7uZWOClKmLAMu/Yu7b4Ix5oe1SqK2+jOdVtC
QIgW/kimErvsLzSIvn3X9QnBpZEgw1BOiZFaku+/irXVV2d7EFXXA/xLbvbmPNxdl5S1AdKecbci
svS2jYI+/DzO3WUQBeSwyalSGi5PTn+SCmdaAs5G6FSatMFFftu1Gqg7iRFFxtl5UnrqxXmycYRO
A5Y+PxYJMYLA2X0wOJY1436xpLUU79vt2fQ5Z9gmZUAjZFgnciA0cK8X2AdX1Xg9G336N/DdSG6V
Nbwe7Oj4LtmlkVHOklRh/wsBqZ72Ux0QLLxngRzy5+mVRkzLmldhawU3lgm5W/wnd07OGRgp1LlR
fwk6MiXPZ0LpXZhoj/syMktxCHxlPFmbYBof5fQZOGjXKnp0AJF6eTm1crpVLbns/LYq+5djHHQg
LOc4onQA3kYiNbh3Q+V1qWftogKxzvJxkuXk/Q/EAta66tO8v7T2/l9RvNWKLYTo1WJzLePK0lAI
vRWya8Vi8Sg3oR3QtNFxY4VN100GFpGAedNIanu9Xc34Ly98B+aVz+AFLsIFEFYtz/BFbUni2rbG
GeV8f4gT6xfEA4gA6uNG61pB7h1C1RV6KSMJENd4iKoRJ8uc26Lupi+DWsZaSUFzKz2vA4ZGb/ga
1wqqjktta5SlK2/ziE9zJ4LvQ9k0VWn+uoeYMLoeNR1lGZbbYugx0H6IA8c1lzvEhQmsLni7sMvZ
taAtEpwxhKbBvERw5LSQiaEbK5+0S9t/8EpNfVk1g7vHBEDJdpkxjy/116gOnUU3KNVyQnXPisib
osP8xSWwl3vuFYZR1EapEiC25MgIQhQUgG0zgmGElii9r/Z277FfUKV/ECZQr20U8if7ENv/0FXp
70vGV/7trIjlLBi2nwrzvWTJjiO/PpPur5g9dzshOE9vWKWNfwtge5bWi0kY4WNgmZhdxX+NrMrn
rX6hH/wptOWfr26pSz8GGLmc+EI3gmlI3mZHZ2hTm4JuTfPvzEq91OH5a6UnM/0OAADwsW55WfuI
pk49Xjnn1cxivNlwMuAlf7wOhELv2ctcak5A3RVWqmBAHjp56Svs+Knz+q4BqWtb8xY0wHUCz7GW
91dBh7Osq9vd/odXyqXPbpC3GOKrqlM4kjfM7Tl78bVU9+1DSnanrUWiuZxD2/NHhRV+o7PnseYR
pUTRAuuBdogRHOaCN7AnfdfEu48c7qWGdUcLgZRi48w+GGpUesjeSXERpxsbZZQGBOcS2aPxMyOL
/t0GaW9uSwYitQkzZxFaF60g9zYe0drcI7wRW9DvJe0mg7kLrbGFphuvQ0UjPczot/XFstPmqtSf
ysQZZhKg5hf56WGej2+8ZF1Zs/vgSGaX6fABYmVwlQPbDWx7pMVdu4zHjn5MRK7evdHLOpTMEuxJ
0Uf4KcXkkYZ2DPHEP0Esv6n2ZJup+vd7Rhz8nmS9s6gffYrNJVYr6DUQ/Kba3otlq1fJqmcGKzt1
oVE0U4f/ElD7bOwS0GyZ83WUjuBjpaYIVSrh3iGObnT9xpHzwbnhobOPWPVbmPWwHtfpGDWmY1n+
doLbtCjH+7u3dtxzd/s4YbpQIJXCogoU/wq6NUU/zADwIf2tflqpUMh+VA/yl1w3I4ti2jNN7Art
C/RbN2kGcJD+XDoeksP6lE73j6oZPJ4GcnTEUCHVSr/KciDXRjoRRlaKkZcAXmTpFQwAPR73iOyb
mripvbKRSmC+wo7rIEnvIJK89dQANv1cFjw8IWm3fbxXNcd2ePs+nlD9eJbapDDloQBd7gdJwZ6G
aqRhn7tjfPRWLohe67ckQ2n7z9EPaNRVh1HIp2Y2JaNhbOdkNT+jHvSXb5AKJE9DuLz2T+P4jbH4
fgCPIufBs+Ngztp6x4ZA2pvC13n6yjGw8PLQERWeOQrHTKyKtSPhnT7pBfXFgeQ+aGH0Bj7NdXKj
e+9051rGdwD52WJSqokn9hrkw5tOS6rRBXRgbdzGMRPPNI2RiVEpR6gQTpkLiCp+ENXN0yZgo/Y3
yizv6XGgGzvGQjh4JDMsBODRfB+hp4k8EX+Hif+c6jAt/AU4I5Gbir/Z+fmyWoQSLixtC2JVQaZL
ABh0DNyvIG4QZwYpoUM+VsGQSbr9LLaWf+un2RVsckVXUhGj/qYEvAf4QHMXSgZddfpS7CQ7uQmj
KO8mH1HiDLEK3t/rp29TC98G23QKl0FJzbWjwGt/jqyHy3gBfMwTEAM47ukc6A23iMMgyBObKyyh
Ue2Qf1AQSdCToQOdizE/ZUf1+h3t4/JT0xbP4Keo3KQZtQytRaSAbutQPpTJLZ6FwUO/qxk+2bw1
/p6/hu/4vdEGzxFP+oQiLzYjr/TjmRB+H7ZDwlCjReUhOe0mpy8R19842ZNmH/TyymVxD2iF1SBP
xBmFoDcG6zVhgy5psfH7T1EgEUV/Tm7+CRXwcCNVbvDCVcB3tL9xqajXGWEuwHox43AWEK5oyvCk
IYkWFQbbiIJwdZle0cq5AGKrcZy7ZXntOnk4dzB5ENfr/YmvOHZR7QsEvjTEzSF+Y0HbNU3jeNSG
qYKb17KVp1APzCGkRW366qyjecLQkJMveKKJLiwi56zZ1EE9A0HRI4T4NmQu/Ygk4grduP6kG4Jg
2EyMplnUnF8ZAD0yyciOdHdJC5nErCbWa0n/Ay6MvuHrAutwaaLUyop69ENUctqLj6cOSZryLiHi
n2q6dXu5IUooNhhMCDCsb1RxL/4GDhGU6jhLToPn6q/XxfO2nVRgRl2sE0H+HyA71xYWZuxU15xf
XaN1SaDUuTcvGarUEjZz64zk8ayPO/IGjZ+jJylpqWo7R26hn/+1aglhKNtfBURCUX0hXPZSVFi2
9ASf90Tg+08CNn+PnzCeN0owgXruqDAiirZ3vYaMo3zDzSe2uAyI9wThTbYGKwV5Ytv99YWqsHKJ
JJ5Y2JnS/oYsGIn+sGYBODSK5xVAj0XPRU8ML3QBzqB5wURhFFkMOfFaOTOMrqtzZ9W4n94e7bJ1
NQLld/2XiBTrgzcsyFKTC6vf9hWbxbBn+yDjlM0vfQ3Ks1F94Iu7BvlpsmXcNWXNyyerMy7EJre7
Um7gBny1cgyzY7aXU/x+1YzCJ958oBMc8aLHhHHnmdBot2PlmbOWsTCPq+H6AbfFM1wDlbDu4th6
fO4csoS5jPBivxCwBqOstW2J9xaffwKd9cCi8SijmuN+7+ovMKnkarriEW+XcTM3C3TuxA3T7wrr
lZISmLpOr9oqoWj+NkW7d1DDaUANwUA5jpZ3pQ2tn2y58FXmw9U0zLrJPnz70nJoRmxbB1Ock9Zh
MF+ZFMGLNaOmp/16Zfw2DacdKUBHZs3Z1c0XAPJjLm9kFZUNmXSF1vCKRPdeqTaxivGTYDDWNdcJ
UOX+Lc/uTGxNl+nDHakEBNzPys40a+mA0cVq5rnMm1ichihtU4Dd7LkVgXvUIda24hU8iRReIcdE
gSnVdeC9soj8PeEcivXeVMjpvdvEUFequE1z0wPuDOWn59asWxJmbEBqCKkVDqd0P4Sy20MAqRL6
AAa/IXovl2qDr+dJYg9SHg0MamHJsB22e9WuthzGYlZw2GTbskMO1uHdRf/HivpVFjS1ImOMeO0T
ZOaB91GkwaOxjVmBa0KhEXjOUQ11KT63/AlzimL6nllQCT8rm5WB/jZdc9H9drjDarQAxKGofYBY
s6eGqEsKa5sGRkYm0xCpl5i43hdHIcUv/Ex0eZook5lsUSXXkFVEcPZXjmLKD5cXoLGz0a6yDjTy
+If/I/4YTjuiOHvBWqJqJkWtDGrOqtipc+7amZVmUU4QStukxVniorusFKEQSBlChhrOOK7D+MIu
80HzJDK/7wrjyP0Ea2WjrLaJ24gBUPLS5K+oijG0lyF+2a8eDkmMZ38PvIgSIX5nrBkhUKGtdrT4
3isDKS7aN4FJmGwp50dNA00q7OgmsdSooEcfbxXPnHdTLQkziCLruFMyn3p7DazwO0rmUqk8rIw0
qIxSOLiXSPtMMEDaSUhJTZPy2X8VW0HFZOFrgLz1rCCqD7j5pY2mFEmDbEOR5uMDyfdEm+NPOoMy
SQyLvf0UjM7JpmX49GK/R62dWZLvFZ2a07Blc4ajgjq+1xMIdRC2T6b7yXU9JToq4BDH8kPHp9Wm
SWeD1WRPQIKueeTMGsg2FWOsaOCSqdLbLdn/qISeTaAwvTEMXBM71NvNyFpz1/hvY8iQtaBRYf1y
qX9KpPrpGw2IdeAYqPsFA6hSmk5CZWcnfd7IJSqNsoyAllEhG4LHMl8wD/rIEIV7GyZSejGo09lo
NPQAE/VhJUKITRsUlK6AWm3sXU0O9PSjbgynCBJLfiHzK8g6Z3e273hNSyW2DohL5FSoBczKUJ5L
Q67yUDImIPnGKZ8IWMQs6jHOemMU/Nf6ha/18XCkili1+bhYbjdNpcWAy/1U8FylZKthGhKkcT44
yOa7hm+viW1gzI5q/zzpOa1vP+tweW3eMlAx0pmOT4ZDTC0IwAba0Zn5j1+Be8cRLH9Iye58NUMb
MxWYjcNQV+glG3OKU2tesPTOW4WYTsvpiCRXry1ofcTPdE9/idH0PYdtEUGrpHSsOMnkmrw/0PCn
6idlYaEQ/wmr+yGWz/HjpXWbrvcPggpdKkypVTo82dX2ChjoX8iqblSXvO2yrV8pPGkA92BGxwka
Mi7vWnumB5TMjR5Nqn5h5vgY4ObO3jqTrp84E6O19OsPFCtmOe0nJnSUO4vIXIe2Wo9JC0GCfYiF
gC1tjodGePLRsdneBrOxX6BEZmP9/ZGqguHcER7Rm86DAyO6X9RCddccGq46iITt6ExbQxXQrhzp
3fyt2CBs61g17BpuBgHJZZYOcBChnZ5XoxCMxUmQe6YMMN/iZnyY6aUAA035vC8qlnl7N21iAFWu
TTIY6W0+WwKgfbPq7PR6VlVJ3/bHAYjZJ1Z6frf5g2QNZ1RluPKDGUrdYifV2IDGbX07bT3/MFHc
MqsxeMpVN8/NpGVlavZpE4NRHmSr0YA6KfMejao/Bak7dvAtvQD0frwhSKzQaJ6JlpKQFctXzp2m
xQDvnfjjh8hGou09xaVmmKw/p9nbJmQ0K1iV5JJRk2j94DFuPEAZu+7dyzmJDCkKPp8TIKZPZvDZ
UQ7DNExGPKVTseCIochRO+Vc3E7Uho7nIC42ObzC5S12GYzANN+llnfVYqLTs4X+F+rZ95WQJDG/
OuH+34X6Kgiw6Sp/49I7+zdw+ENLbKW27DnqrL6pA6YJlTfp4Ru0BEfLTetLKnnqx5PAkXGvKQAS
idjWLrsdqnB+wy3iPsEYyWTbmPubwrweC9iC1tdP6X7Q7v3BBqLGr2azZcHU2NnsTyKCw2i6OqXc
pHQ2XRPJRCnmmMS2O8Wq2Gyr9kB+lUNGiqwE8zFD1X27iTq2WJG24P3bdci1GoO6SBC19jRkiBxc
MjZzdlaEvjoKU2x54ARMO/VcPlkg1UZDpDzSZ3NIuEIp7Ik0O82KO/a02PDGHEQZFDwvMqmHhFdf
J8QlBvzF/8hwf2eWu5p9rjr1jWF5w0/LQy+LuwGpL+ghznFZ0bXN7nG34e9Tez04FIqPY+pDajIw
qXEI3RVxEXlcrh53RWEzQ/9uzw8U9u8EWipy4CofJ2YQdg3U++UHuA3wvX6LuEbcvUBCghFi0EN5
3iMbFKfR6is2I5/Bq/stj8Ns9QVu1xhD2aNIqwFEeMr9VjHvhX7czMzuwncUxWQ3x1c+OvfH2G0a
nnLPu9EVzV4nReH9kfE2KzZaj8GR6J9hhWYW5w+5EtcZGNpLi3Wjv3sigVKXtDzUfROaMl3XyLY1
TQrZZj1x9NwGd9TBjBoEa9hlNg5pjqVx63/oKHgWqRmaJqu9bhA/55km5IjEWQot3z4Ml8QnhhJD
wwcIdt4ih3aKk5LyNhsQbrh9j5pT9YOfAILhkGS4JnctIici05T7DTw3eEHdxa1TyFs2cHXxo8Fv
m0zRzPe7s4ucDgju126ln+l1U2/ZdXCsX1ciq5WH2mnUtfH7Thz4YYpXpr/S3ObKVoJHyUhx+PKO
tf1T7M5u0j3RTh1oj5aYlbLdZMBbS4XgN2M6yy5yMzTRQLwfNeDH8BOssiqJtwFJXKBHDBnC5Deu
OTL41G7pLOIbBy6GRObxn0c/kHMDtfqI1aaJ5fgKmD5CZ63mY3R6lvTVjOrD6ixdvR0jfn9e3Qfw
xdSDhBh2n15M4LmJXldE6CK0FKX8Fn8+yXYDdgJVq7n2Yk9tt8LhEpX01ERwyhqU2DDFcJh3sEU9
6lQ/sGQ3W0gfPzuCbWBniXUVrL8UkoGzRcsEzKn8dp6rNt+UuBWlRT2yCgopCw784Eair8bVgH/S
UDKImWX9DJ50qlSvprZQZ3TDqOrCW507U0AC95kOndrWgv3o+NYRAq4i4CTKky75NuuoxG1lCxN1
JWxe2Gh8Halcz583yg3Nkxzz7xTM1lSrTuhVNPp4BzLnydzUKjCTojmlyxAoXkcbu3rlvLFZ0cVo
3HCgUS52hZ+E3CIGflcOS+836FOdPyQYph53Tn8iIRAsHVXmM8uVd3wo4jnK/dawW664NID/AybJ
xvXxwG3gXU8c9ga/LpNQCTTcakVdTVvdEJSSWthqukQNNIW6737VRcnQVWPsse4ivcPrNg3T9lQr
98JuzOCTK/VaGvO9xvl7mwVwtF1hRVbIZtHXcjofJDVQC0CgrWl3f/MjfFC3wTOkIme9tXkeXzYE
4ZCYnM+6AVCJX0u3wjdN23fkHjaIZlfgeJrghewWkb/WvFnJc/a3JqEwknevBH8sfxkGKLw3M0Mq
XItgGVKZc0xLI+HnTogEk8cN/1weDCXWMBNjLtwLLeaJkaxof5Nxxfyl+LnBtEflXHqvNmqp2IiS
XnSyY03sUAhIeo2hJ+7FdruC71ru8/3mVapimVsUXXoPnGl0NQJTgvGVw3dl2WjMd/2muxIB1pb1
qCqp9UUwq/IWzCG3LT852xfa3FPHTno112vXP+Pn7js83A6R6JAJvoHEuOYUdtkfi0gvt+bwDuzn
7bpEPbVtnLOZ/bgm8RYSHU7H7KhhwPKo7xpc/9Qrwfge9SsB1lqrA8ZigvM0BfMmZ8k5+t/GRtDO
uhsW3TOEQSZbOd9eST6kwhZGt1Mcq1zMYnxA4p+OpHkrAg7tp/jRE8Ee4LoCC78uQ/+3WbHma9X4
oZjB3oFIQEZjUEF9xADNHzE7FQmuUm8TTCAAo5oRh61U0US9iJsqFrTAC0RM/rciTt1x1xA2QpAu
F9vd8OH/dDWSpMU/Ipy3V+DTNb3TFvmOwsfVwlcwqiywVy9Pv5o3+M7NjtQcGBSCJPkCK4UyT7Fv
UX3VYBsiy0x7WDzEAw6nOxZUKRZ15OYtqEGJeq0IvlOThrfu5KtdiOdPAmByEY+JodCM366Fh8EC
FKabYA/S0cIVq5JpydQDe9Loh/N4wBHWx1kM22FZOlJgGYe3wD2RKYRjlJFd0BEQ2A9CGD3FbK6T
pFp4CpPTK5vhcfFgcyXCmxciri4oanQdBGRAldg1NSGa/1T7Dd4Ce2rnzRwCUPUb2M3rbjPbBIGa
NLFCG1RnWhrgs8Uctd5PaUVsq71F60I5yXw8hgLC3K7HUOjp/PQujfknqD0xE2cEXNnlMCtS6l03
EPKGtM60l72mnwF4EsR4Jy08J5x9IbuWrshnU6svKHIUVNNkk53+jQBqHs5KmTwJD4mgQlI0MmIo
BGYqiFWk6PXAEeRJZfvvVTdNPsZZtpm0JqWOgq+2cTRsNnBaZ5FAbdLDVMP6Q9Z18BuIG1Dfir7v
sq7O1m5Y+QJraZyEWj1/tQaBO3hgGaoPTQ1XJstRkRwf+RJ+xlAG47aItTYFbii3D4xNQY4lEDil
aPAIkFDSj3ZupLHnTeFQxh6HdR1d6iy6n8+vyh3DCXhYkjqp0tzxS7BIQnw/9Q5ZiCPbaphCSXF9
BQUc4JPn9N0zBB2EztvG4EXTYg2NluzlSewDaHX++Sj6+/w2/0N84eEEAiZOFLU4K9KjDKFz4M/E
PcV1THRK7h4wV0JznWQKx9fbvL0XzQmnNU6GulTLG7kSGSnApVqjrTtwmdXfJIXmSSYbMsArKE14
EvRoRMHlVvehAhEeEJ4/+vzzz+eDRqZ4yDigGZoId/L94ZznBxVvcLi4tQkrKLyX2FQehAEioWB+
gSIdLKsC/5Wq2TQw8+Hm2I4LgPOIxMsdwozcWBYJ5LxgY/+mprKon5K9wPzpO+564PXLW31iwItU
I3D6HcewhheIapqBlc7VRjNErjKfvY3QOmeFyBklPp9GkzNRxAmO3Of80N9JGE7NB5AyVlbuje+r
VhaHKpIQgCP15RAghO7uzRCG2hfESKIf+ieNkeOMKYxdcOln4KFsP4nnh1kSxzv1B3IxjA1SWHT+
1/E8QERmQL5W/CjJ19GsZFcawV291mhNdkIhdYUDXeQAyou+i14LhrVekw0KdYzoPLKBZ41pY4jd
P+YSDV/aSWAdpeHMtBVYoxiMBMvtveEgoz3UkS+z1n0KU5GBrzkKgRR88PnWJb52G5ZvFFT7/BpC
DKGH7kXMa6zrHJ0k7aXqzlybE/PaZdkw8HvNqnEuQqANHe++51jijav8wbpPk/NSNh6hqKwTU2IG
IZeaxQ7KUEZ7+aKnooUTWZT10umHRKDDR2tiyxMkNckPdOpdqHb9Vz1DgiBGF92x6VFyik7YC07a
dIvCDe8/H8AayJgQrHOMV8sUlUU0NZ140aWYTejuNZl8+Hp3gAzU9/3VBAJgRHQ9oWIU4D2C5ZGJ
mQ75Rrg5gcp6WGo+GwWR2sE1QbY76k2nYsL7c+XHbpzjzb6xnbcmCsWiMAxD7Y1iDxpWO4Vdyz1M
r9oDdxfo9cJNo3Z0OzqlmS9zjyd0Mg64QuupcmS4WSkr8mDQ2Pg+oXpuS59pKBzB7hFKWHEvQLOx
OL7BbaS3W6hao3hB8PJ8hkct3P4xcHIb8ZGO0RIsiTHRSCSk0yfi8iILx9wqXuki5gftnAIVoxyG
M9GkuwUXfEkcHlHU7K+4NwyUw8ptdKZ8kE9/ALPHlFs2a2xrKulWlqoY9JUe3M9wSHRO/K4gJYlH
PeeYN/M9B1khRFZaPFxfylvwCX4qTN9AixcBhasiDjEaWbUB9RF2Uv3/Xy98Vxrp6wreQSbiPv5r
zlchSmeXqQ92b7nt/0i0+u9twOrSlCrRUC7e6RFyr8twleu7AMJffHGAyY3O5IhhNp8PokNiXkXr
aPSxVANnLIzDCpLfA6K9OekIQ4vfUY/WIcD93DXRo2/uPlBS2ZKN+4+mJQzXrUQLUXCpRRd5rQft
6R/Uidkp/CX0L5CtUSq+afqVIONG8s07oBHu7Wl55EY/FToI5rPrRlHjH4EN2sdTOnV3gMhfQTsy
tEYuOwkSNER83ot27SH/G+I8eXuLBoctjWWowxOlhxSbyypU/+r4B9t5mq+grGiaMvfNBQIICkCk
VcQXgEg+O8OXrsUGUbkTP/eIz6+GVt+KaJ2Ys5Orgfx5bGLsOMC2jz24UOriAf5R0/jJXK5217Rf
XZT7b1gZzCHb2PdBT5iusgV2B3teOI9Cyu2QBCIhHmJrUv/sZ83G6MnDcAmbrncEXdGr2Z0G76qw
IHmVlqdxuwYsQJsEzmb1xtBrwLEPCK0OI1CT5kFmFyBKQUUZBDq+dydimeajCAolMYMucMcDvGA1
btRO8Xc5+hr7LUyp1VFTwCM+UKPFoxx8xsGDjaPQdIC9J+N6zPbh3/HSeXevrldUXS7FXTP8yefS
LRXKIeXplLuNFLEydN6KEztsNPByacHt023pHjcGlC8yuvpNPSa9a+ttoowlVcmZGXdAWPYkaBT1
Ty8DOJQQx6qD7ZERN0gHK4+vcHFN+mXhgIqdMhCgRC2hh2Fk5ngRdH0NKkc7y/tzBEWeh0slKa7G
emjqVFgfsGXIs09IQJ1AFRLufzYYA4xoJyDOChP0R2FNvWtQM+D8Y+AIxiT2TH9xVFZofuvE3hxc
YZe1kCEZXwbqmYM9E+3jbRsoPc17gZ9vX7Qj5f3xj7QuRdlOYFJHZGaMr/3w9XwJnoq+wSwA0TGJ
iMI1P2PPgvTeW+5KF4yEAlFQGDwL2Ax1uN4merclaRt0NC8WeFAD71kCMBESHFEahl2mRQ1wdRCW
r0EefO8IyVX6+CfVjZQd5ROiCWOy35f0teKXp285M5f+XItKWuY1P5JESc3gtETmCy/vxJlmlahY
XspQ3fYJALO4h5SbM59T8Hd+rKQ/zAiQzObiGAbxhG93jdY1xJts96OAdoodxxOnqYzEdnPi1UaI
dfjEcwQflRAfGuO8FUvZFJ1JcK8I/wsp9vrYjz1YMgk3rrT6v8HFy4dE3Wpr0FJfHEESjf51kdBP
Z4u7p/tVkvSRTOA8imR2Cy42bwNLZ+H8F48lNtaJyVwKOWEaXrsP2yrQPfarYJT5OR/gkmW2iX/N
DKjxwdV0ZN5/AzPA+387/57PUemWqg7TdF0Iv2PfSEP9Chk7etK4N4/+ZLIpJRvKtghohNxYKB+x
UeNcJdvMi2+qfFQkyWUq4Jpz4hbl2r2QKQahM5SgriYMDhn91wPjnveNJE+SUBr0WZjgVP0gHaoY
SX7NDdBknOF2A2EPYMgGbELplFAyfu+yHyLMqvh7T5U3goPBKmZ5WnlLD2vTQsyeEEjQQ0zP+B7j
3T7afRT/uQQhq+CqqCEN3j5viDORFIMRGveOKM2GUqtaBCgqIc0yYrnLmlbhxXAVXs5PUnS4f3mn
saezUSxF6s+kDPN4uRwyvo5oBblmOXadK2KZj2/C01jNyXNi+YK4zdKbYSH2KWovDg8YXZFM4Cb5
rP4EWtp5VtlDMznbOSETPgC1fiJ3lZkt0kZgSWufMTm08BRfNvJtKkHOuJsPLYATK25FAdQ72T/8
egn1Pc4efAm1RtKaXiPRhXyl49qOckNm/svBQLziNDZ1wpgjMoSRtvCY/kt0ZqwVLV1t3PZPeyuT
rgkOv3Hq4Fxl0QUUryBNGtBjcb1LWf9iw/tsOpRb3bHoQb1RkR/DKHDOOHdZiZmDHeR7KZP4tQmR
2npNtQvQyIg5wvy39EWXKPuN6rQcNds4p1zeYclnHwpZpCjdKEM6OAlNVB+QB/d0mGQrMLsCjNxx
TTMxsIHk10UTznwSg1eNcanyokIRqSZ8RGr5nUlRwcr38etqhE6aa2XfCfSunUlROzS9+SR6t1G5
tE/Mi1BfKeNDzLy5jK1+7zuPANCphLHUA9VCWwxLbm+CV8b+TIPRJnY2/QZN84SQErvCfrVGSVhg
SaA8FgJZr5ReOYISjPlX2dLBL43Q4CHNqqUTOQG9ME2kUTF45Z/ovtbVHGbKwSAIzPaH65+0CJk0
sa+/AqDHoMLBo8N8e3xAJFluXXNlPp2lCiTn33Amd8oo3XzmLchruIRThES2Le09c5SEabV5H8Hc
2ady243QAI52fff/W3skDI6U3rdR6MMy4HKT7WZntgJEFj3YWyWgdGXMa25MjEzMws2iy3oFT/JA
gIqtocYAzdbWpGrt57gOC0w7qxL21fskdjZNXlVugPVNHDTKaASKJZHDkVdw8RoLwXEtWHJAbc86
ogpF/5eJ0Ao9YG70i6oBUSA16XmNqoYyLatlmm7d09Hi/fKJJYCQUapwwNAkD9ayochFTLakCOGW
vf4Xgjpzb0eNUkt9NCCi+ZE/ZzKIRo9tzf/G0wXJ7jPlKqKPyPAePHtqprHfFxfVolA4SbX1f3/l
UEyWgh6mIBMJGmHjx9T6hd74vJsKWfEmtK57jbLIYhXkCiiawbHbqTpS63pVRhTFmCOTY6H7x6gc
neKG1QOafMlliNWd4o11POTAQWKnfnEeVPElcJHz4XHDQEcMAsmvsvD8fIqhPpFFuWxfE92Eh26r
tNHBXrJDcrSZ9TK20g+YkNBXbCZyKVgWvaK2kepRcJy/J3xsaQieag8g1v0POqzPkradA5SsJ7Og
2Wym+XfVHH9jCKriiVygEJvqXNjd/g0wzo4Z6cSd+Kp6fGGfcMCAA27fPcRm50aUhvv4rGPP+Q80
soqhLS3Kl/WLVvtFzxP/HxaEGLgo2rCkbfxeOjddT99SvHEjnT/YSqzOnlgDX+zQQfMefRUsZHDd
6tESae9m4AJRwVU95zZAecM3LvSpdplUkAfShs+C3y4Lr9eOtNE9R3WVJ3waVTB7PlbeKRk4G58M
o79mhEV0y7ofD9UVs3PE0M5G5NjRbe7SNagrqbOm6Ow/lO0DGy4CtnjWOTZaz1WZL+DDHtdOM4CF
alfqfgpGyIUnfq8Z04sVpnw+t/NVBOQwbPQhN0k5qkkCU7s4c04vC6wdSDtrod9S3RFBWZJfQj+T
lOd0/pG62Q4UT+XEcMWAXR5rb/s9sXGGEdtbF3tO4df7er9mG6alLfNvQk3N8aNDj0o3TB1UhWoW
qXkeNISMpO3cRwz1EkGqMrp5kpw+o/N6Mc3vcHOaYT830tSv1VEHxrpq6+hxAHnXCBtE9kCNVht3
gtnpNLS5bbSPqhNRQYvENzr+qlW8H2V9gkDoiZkf8LhBNEAX5Zb+zBD3p2pa3ULSF/34RkjBytax
U4eW5jkIpZ3SCKgJISLV7EU73hk9ggKOpdv2fZ/ScdQu5I2d7OY9I7HZ8MqKsRN3z6TdO9Dnno9/
wKRnYwwVbM8Z45WtIXr6D9o1tvWCiYHl4E5tRGv4R/nSBy7Z4BpTUYz/ciWcQSdrB55ioqrRGFmS
gC5RiBXmGbIvFIRtf0AcoOJGESed26Vj2D2yyL9HCT2oPDdIq+bmkL0PrJL97+wlcLZTR7tiw3Wn
2EZxlYcFbre1BrlmRZTlvDBqvtCVg3Y43CEHFLYL0idBpr2ZV4WPW8dj0jXDrAYq4wXuP0ofYkif
FBvOIF2VYl3gcPSadnLImltqYE6YUJACGHpkW+CXPrG/0n+Bk+ydpDg2+JqgTojgyK1PKpjHsZlg
Leq1n++xLBSdLYk8l80TGnTr1lVHalgieBaDV2P9W55Lyo+l5qWqlfq8t8NePnm2WnbQePZYavkl
xOLmZZqEvcmvfeSEwWi2caotLC5rb8u+XTEIj3GVJ2Ay/sIDo67/k29rwgjyna4nkD3f0YsVpaid
e3HRvGwHo5g9NC+8Kh+vAawJiy3XN4rC7uCEMoxXltsPIASzT0oaQW4qPP3SHvrltYnNJZyZQmET
LPysesfttY3nYfWvKa75BmJWegfiIy86/sgBN+4rF4sU0NAVM0BBB+oHzOPFLYRICPhHuJj2sO8y
Q01MngMuGvXPlqcZRtJiQ5V/4FggWXfq7XKcYjS6MxedJI/WZHLi+W/t1RpUORpRqkalKDcF53v8
QbS+Db4xBhZ+dJHjE0MWrCvyIzMudzKG2Gfc1KE5ikit+KcB1RhOu3O1q3a5zW5Tqzu5polUQoqS
kW8JmW4kJrWwPZqA3QwvmwRDnkaF80knDpJ67wDXf9RUZHf6tXYt/Ah0iIdlPGRmeXaoa1rjeAC4
wLZBkmW7TgWXC+tq9bpAZ9eRkB1uuQeqTGMkz+ztG6+r7rZjy27uyiSy8Vsi1aVR7b/iVCQxwLjS
PuRVJLWmfGcP1SIlxtkcszgs72h1kywd0Zv+F4JqdLngReRcxA1t2AOXoZRPDVeg273Glsf+Bxmr
nX1gxzeySrZEHRTQ1Jvpip7eucJY+d4b1uPclyQxlV6WBRTtwSDLRBO5tkJpRxmnxV6Q2x0Y5eAq
J+z0gsrJ84Y5n7vsdKPt8ZfydFMMNWBskUWFqCLjobIqOZdAzw2BoQXUH5kHa2ay/j4jRQI7i+qP
pGl1sLcqRZuPd8++X/FLzlHrUjPxmjcxEyqizVrs8QfQflB2Q6Ha6Wo10tScBrBpxSNyzPQzgYx+
Dd45b/R+8Rz3NWVw7ZOYydR1HfYnvT1TkYhRtuOP5o8q/Lt5LTCZ6XZpE6aSnmm1OFRXopqHHHkF
VN9X4u9XTHTkkBESTGHDDe27gKnc8aeXZ+QMJhXfilHzbeebNjna8p/W3hBPuH+Hl5gEnU/Wh//i
Y1JsCctgrZBZA7/4yzE0tiAT/IZEEKqvuEyFjvOkhgOl58oj7nT6KNvfRnOpT6noogwIozsMU9yu
BG5kLa5zcpNC4iiSXFYxI3SSkF5FPPehvTVkf4AevBl399tzH2FwpPkcinX4R7bi/BmXGmQPihzU
Yifn2ZbpD6gFR5Nhc2w0P36dji0r0DW+X1mRboKHvbbo5ig3rIylr+UF0nc1n9pq93qtj3mfAhBM
T0bRCf6yeyyx0Swm74/SDG17eDOnxBZf46iYp8wKw2J1kvHUiruzbgB62fJryLBqAWsAC+LtCUtU
gCIYuyxqihU6JxYzV5kBbpPCswc2wsUVb6Y2Qz2eCGAFdv4wUOzACiVa4f1Vl3fdHfqS8g8H6gNr
t3q6XnuxvXKs3m4qmLuyn2C4FvuH3ki1PL9lEFnUloJY6EhJD1s0bj667KUYPAvQoXTHwppkRFnx
daFVeJQHUDQETfvpjjC5MG1cjQPvdZq8xMXyv3ygS6ETD7azQofC8kClmCpbRklRLLfeTRzWMYzA
qfeUS1tFyPouSs5FU02SnGSHnhJ/R/1frM30xhEn8VpSPsiZQNhN+0wSkPsAoPrGJsvXgGBhpS9t
tjzpCUs3As6g062vxIHjunC3vvHlUyfZQ92UviclYXOgAN5jc0txRp1Z5xYsxEAZxNTDhLHEMbm7
Rjmi6xR0lj81LLsRR50pzjQ554bFkJqBQg0nV+DUtlu+O+JL2I9kz+kxiutYag1WWxGNC+KF5O/F
bLt/ZO40kOY4kk10tntnIYRCf4e7Tj5pTiFIh8TNSW/f3IZQJf3yhJfOFPJuqNeiEmF8bOGM2mJ2
MSzM+PzYOgOHzq3dsaWDLDEk6zco2iQFQzQQtytF3S1jwzVAZ2bTu9iPEzQWdMX1iR0sHiPKPSZC
whWoE9IMrEcLyDqBzaMRvzsM85jYRtCoE+CukV5FDTmPjWxgThOPLghOeNBYuzJIiWaSjXHcz+0L
x/INZBfuf4e40U+wIKAWWO54H1I4YhJufqhYmsFhlB+SHHmRDcT5BoVGaXzfzdhPZCUM5i8We2Dp
yQn5SoPUQ4piP26D+3PGjfb4e6zoMos9cLhll4jSitaZjVJUb+kPk6sBezXn1fEJxyQA/5zh6NKD
g9R9FGMoGLBjt5k7WWhIXcQ5kVfQllirLvQW4NQN7Jr3uu2cMcPkuzIPC3yXCIfT4W6BzCQd8pZ7
5uYrdKh9PSCiYP57DmpBYNEgPY6HmpdatODZBdyfzbbsOJRUePlEz9uaW3fV2iMFGWpOH8PQonSh
TSZxuSiK1Uh2QxE1cTlqreRMKviWVxLCddd+GK4e5b/vYwBBrdnbYSfcPTF3+eOV/eVokxfY9I+O
dx4rcudgWz/Ssnkctia/ZOpTr1bM5ZFVHcjxD0O0DIgZ3KCEgJ1ar2CCXX1m6x8IOLxc4Kc6RV45
68lp7+WautN5trOlw1q4ltf1/ozV3KBM0ZPtkd/pv6/v61Ntbx9NqKCWZdSIcTJ0RlOiJM29oT9w
7wXqHe9goIX+5H/I+1QsCEcoC0VnDkWIa/rOUi7X10Z0/eNi5HvGu+FOXy+XDTA2bwv6MIooRcYl
E80PbjhYP9r5aKwveT3zTUmljHT3Nj0WuHBocTUYpRCCCEVyvlynK7jbg0mdIV51bhMGU3Cm1tAH
K+V71O78eq03hfLIBqZgyBjR7jOudUY1i1MJ+EtMF02n+jFkxhOB8zZpwIOkJVf2quQ0MayKT3VN
oXQY3q+MZiVUZsxLNOtMPSH3Y/dd+hQSPqTI1F+82BER2CC0mV44QGwlwWQnUOi7bSJiu35qWeCQ
9K87s7a4rOO86DKZ7jsuX2e7Dskrh1nFdTZiWAMmC3TCe13XIZ/wGwRh6zsg02WUMDIQ63TaoSvK
4ZsuU1/jdEc3G50bVnWOrtplp3xcgZJY7H47oPfhb6skyvKYEbXxlYnH0XwMyxRpRPfA0IZaVJdI
rDe2PELG5eXGUPetQD42AtvSVsXItqhd9avEJy2v8kz/E9HZOhJHwNIhqYpzM7YcLmzKzh0e4Z9+
+2TKDa62O05g4RN1UvOy3ZQBgHslq6ak589CSeL+LfK4WjImWiMDRdDLdwyhNTwDsX4gJaZaybfa
+lG+nYWnjIOa90EcVZMAf5oNE3Yb8WEaiAN362GiM0+4u4vIKTByFZRRcbDpXtKyu3QmoxcR8ehN
0c1wmd+T62mNfHjeKhNtHVWhBN1WEXjlSKXerw5QcCIyTQ2fAKhtYSq9EhSOvsNjs9XmO9qu1B/n
FxLWBzHE32us8lmTDfSUfkLoItLQYRU1h3P8tmwMbhR+34l6Kas2km2Ft9j43HjT9WVdUgjYePte
keQ3K5HIbQNHK4i9tp7vaNXW15Xd9izFBBRXD/pk4rSZNgJh2lkafu5uxFiJEBET3CxFgg+7KbUo
TbDzkJcSZQkbhoo5gocusblcOjRa9PJMYe15635aPnAQqJYYKbOYn9zo1OsTIv2FNmDMFxlVVfCU
/mmDrprBPK7/BroX3MS7DWv8RF+cH+TxjfXh86Is8V3unB0IZciHviNhLtEjw9p8nxS0kjfd0Kuv
crETpw1PeEf7FCHhvibO+QSHI2l3RzmWRUEejdEHmTVcGXozbP56Ua/DVV0FenEhcwKgOcsHa7iu
+GGvwA2a6SPZIpbPLHmdn9/0EkdQiavgMDwLBXEJCAXQgpu90XZC7U6xf9HZQiD/YV3ab7g0E7wa
LJFfSVL8ZI82V7N29a04Mys8qaG2mf7zISWdNNOxpflP2Xuf96+t2CqrRVqrnY4oAZVEQDXEGe6a
PJs2DNEutqmTnEhXPNKR1o+lK7m/BO09x8nEhaQ0czBZUFL/UFQ75wXnsjL+7MUmj0uY986Vpp6T
e5I6cwZ3aWCDvl9JfQrYWIRPJdHuaBalhbFPHeI7LqhZ2Rpxo/99qYI7PT5kokt7e9tqVOXF5r1a
9Ltf4R+S0UAD6FSNpJC1OG4xKMPaNf3qTUEf445reOwBlgXE/9HhdtYcd5Tl+oSr95uKMV0EfpPH
qbEkQl8riJbfuHn/h0MPFnmQKZkfNVRasU+jH7KYszuHjSB+6d6P3prQlMa1Z5IETdzox/bELavW
xYmLhJnxI1fp6B7mJn3XsDNwabGKchGKt5OhFz1+Bu66y37/H/mccPqrvIatFsV6UMvpbI0kkNb9
qN79sHXRnF+ib0RV+ozN3yFwXTgzDdQVsKUUJb99Tiuun5KQXaNC38aAWCEyLchvtUG2IaVGR4kj
bRUjazwz91Qi2HoDUtvB+vyMpSD4chkdE8SemfFaDf4SF+8QSIChvFIvXti6xNb0YDgtIrVGQj9n
CSSauuUz/B8ah1uO9GBdIx+6ScXfRuUAE24FQGwmLLUW+p2kt45b32bZc4UZvTg6Ar4GRyErufIB
7KRL8QY/PLoS2xkBAGMicpqg8DeHo0MKx+ht1YkiVi61l2s7nBMTuROCe0vzEuDmdsGtIduCAnAx
jfZF6iL0xtVVTwEvhLfNQuBAUGLhflhNcsfRNVvbpnChWfBr7Di+BLx3E76b1Bank4bPtMceyZ00
kyDtq0/DN/xCARB136kYGFP4LvFAr2VuyVk68Rcr28MCPZx17i0p9DevIr7wbk+V9dx3MRy1/6nn
KinYCWLAFXxZWz0VQJ8UPLB/+fi427svr9IM56vYphuTNBsOFtb3Pm6EPGRK/ZTIHbr3nWl5jAe7
o4gb3onRgcPM4yR3thi93oJXLyEAAeqoJdkCQOPhuEWoVO2iqt9NX4aIa3CAVTbOvrIT82SdEmI2
Y4GB2yJulrelk334xuT118J7IGSQiU6BADI17ngM1DwKUojpjF366mzC3u//cg3y2x+omFjv+m9e
nA2kjJFCxd2TMfkobCU2qICFvjpzOFOTuOCKC4psKLCc7E3BWdg6IrRoHH+NOwnxFXKhp4oC+xiH
1u+iICoSJa/iBLmyRJEO7f8negK1R7U0wje2jFktqewREugSsXxNjPvUGThHA7/uOZ09ErmdOft/
6KdLsKxzSxP2Ezj8tGzJ8d8/BUabk6ewUXMkFbzF4rKehtNSfMeUjXCfFKzbTrhMFK6uzPoUvjZ7
OSe+lVVrvTjDTJnUnyeZPG75US8TlKxlqJP7JpXkyMyGyQIHaLfkZWhgtYRBkQKvg8cUXsMsmT1/
WZEaKq7v2DgTHncikDoNYmyYWc3oU5y0FtwS+6biLhay58h00jGlFT/v7hvrsv6EKm2AACxVHLJt
pWifMB8OzJFb88spFuYOBDmYHCbEFkmfgSZWQ5QHp1QFnzwIh5MhDCbNBM9kyO5AfIKQDD4XvREX
lBZAJ4iby3Nacsq07Qb5sofBlTetA5gN6wUCO4hhAdJiOPrngW1U2N5NrahTVlaSmIiujE7ad2m+
R6JBLqKy6PuVYaVqn0D8jq5SAZfiAKlTLYH32AioY4eV/YRTxNWkXrrInjFYfNFLLE60G6ZV+wNH
6l44PfU6YIOHbzxpAUL88yr6udJX6uqYwRc7UCxLi0SM7PBGRj25I10UJKs66g15ksFocSZhaPv7
R2ZCaYAHIyBGYc/x1X5xQ7K7AMeygppbBeZ0ZjgRaAYPFgpX680fJUgMXZCW6xIlcuBU8ECbp48/
g4b+kb7pS2K72lXQU1/E7H/5fsZZ8/YwFH8qF7sCHwV/yGNFsPArYlEVaQJdeR/DATP+w/hRRBt/
44ZFjabG8jyJXCCHKSIFb/QqWzDZmqvsXGrArA5z1vTURx8BrtX7P5IAvQ35K0AcICaKlF0L3W5W
Gym5rWh+aw1Tew1kBWOMl6uQAybh0GNcg95ByhA/SUYRVWshrgnn/Kk2FnzBiyFSLduYLmkcBthN
z44RsF6zdSacUQuMNgwYrqr7xsDRLget2Xw1H0QJoSg2DtIokV4axXeolPH+soUkddVmZlH/P3xW
DH9YLO287Tzq//7fazYn8NiYIpBuf01rOxhWquqg935PfuNJ/Eoxe0KvqyyWo519e7wA8G/5Z6IC
d+oACH8BMYC1U2ffOWz9gTuvFnOw27HtiXQ9zmd7i3GpZ0uenQSMeulsC9gpg3HX261sD6wW8bCi
+ggMfOQ+TWE1MWwvEe2obqjb2jXdror94HbiNrFdzL8QSKiakMe/9HQc/Zg6syEbzNHwKJ8dc3Yd
vm4rNXhz6Rwj7aqC55S+kKvPZcqJt9P2FC9dNL7cau3h0yVx/mZRGZ2xQoA+EwyXpj54Y831jeQ9
NAWabWHlX+Q6HtBmNYcmiGSRBU1q4BkUPqO3eLwrlhZFCqYZMrMIIDViPL48h37L5VvuCkTciFXV
0Zwu4YTPh6PE+sTL51y2MsVLEhUOUmYGaeYrkUdeEFqk0awwNx/IDERmM4G5eGD5XlosgNnpbSgF
tAREaYYVYyyDQbQBpFa8aQiJOyqtpcX6e7pBPNMAPuYxPwxPuYR1dWPbTo7+HBs0QqWZg77zYi8l
ep/BVCdRE+rTZwyBaBCPF9ugOI1wPA06izJFwoAh1T3avbXjqsuVsztTuxxf0IwT1UXH2VUTIj6G
DlF70WKXxVuwvP/1B95GmQFTr9YZ2atcLsOmDTr0s1T1r6zjEGDe5fRiJUPVbUTpURfjnD6LvARx
Rzwfae9MMtkc6l25YXVmQSvr958GIOrnmOKZjtf/75LDbDTZ6lWmqGH5B2ps+EGEGsoPqVz/R3t+
gCL57tNFEZkDCRjOJ7v/MtwVXWA1/ypowqqOpmfYIqT/CwrRvRYfu9Nm+wRf3g3fQSNBg+ERjePA
5AVyuvFmtm9n9e0YBB7ewN5cHkS/RbIAp6IXwS2H92H+5n9V2CQvYR7OiCJ/Wwt/g935IjAYwIpo
LM2mDxy5lnvlgBYuze8f6zxutbDcYw4SMT+6UpgWQxCaNNNbHNIzBd2HU/4LyLLlUsmYCirFiOt8
P74El7ayQXK+Ev8RveE0R/tTbczRTxZLFOnIREh13/hBDda7QM3i0+PBSJJ/YrzmkpyPsypUgriK
+aJrL5C4whT5c1EZ+kIUjtRo3DcK3ZUuqnCbrkvMUE2TvctExosnLS5z66ZGuxFeMXXxuSRL4ijq
yCbfO4IEiO9+OaeOh1VpnBxFKJHkhcMgmjICtnLCXrh5DT6YME1AKDaNl1zLhdif8LQuqS05evY7
Lfy4UQrLENyEkGF3MuL7+l0Zx+bR5mvpazH/SrvgsGcKLOCIaOj+OtVIEDhBwlETK0cXz2Dhjo5j
JgoH3X6WHMjFUNERlRyDXXJxa8vpmKibRcA3a0dbrAi7e7CfKKYTWtp4V/es3qUbLH6wzgBrb2U9
RW6Pw43qrQgbofS0HGzWWhugr18uvyT/iO0WQiloNvuEV0B7jjRFFR70uhmk5k8v/Cd1aJwTBTRM
B9ZGW/FkEahwgKv5HR/Q5a5gsaC0kHdYWxHM98tt5bHxPMfzcjvFyqCd+w7V6gqh6RUE+DVNSavP
tzwY+jlXWtnKMH0DxfGEd9Hrx9mpq+0TXvQrJDtDg634vUtH803D80WVFkwZGa05ZCCFMnopTSw8
en/I7Xw06xsHOioH16/S7ccPIkmrl9MWEMNj+hyO45svZpbO1+oCoBPPwZ4IUMVU9zf/tYqxGfjQ
SyA93oAD5oDxvI1Yjl+3glo9SzNKM1f3zAlKyno1cXrAzKGDV38ZvxUkVKZ9HNvKcMrhmGQAA3Th
1Wo4Sv/MsGeUenPAC5XUUMKL78dkLzL3O8YGj4WL7bI8qx+e+/HFuFzviuoV96LBg/MVuyoe11R6
2PA9jb7CkCrjWfOte6X3eb3+xxP3jlW2+nXUhTfRKs7cK0yCw+lxgnI4Bk+vFeojKEez7+caqCEp
UcQJhY7JNGpzx4LRF9qedeR5nVRC7G42gqUuOhHmUk9nOiK+u6VsRMOd+nvWLYvyVr4iFZUF1c69
SRPayPKmF0P+pqHstIdHFKx3gsYcdkhiHQzqhq8mqyWbqQS0WxUFYCZHBiawcuPdwwM9Db+44+Kp
j0n0hUrXVjYVjibt+RRhRRCqjz0336mJUlaSm491QHP+bgbN2E6ZvpI4a705w3cFx0G2EA1OoA62
doJRn+0tyaPOcrcW5zfZn7B4P+prsmduH4JxDZnvcE9xaIrTTitCQm6nngsUuWSVzzqG2QJx/HJW
u3nq5CgqUFHhdSMf+2t9nqDDizaHpf92c0rsOkesAK0HL3+MFKQh1frVyap/d0Au6UVxeCM6GqDd
COXPITxiT0UKp4SEzs36712CzSl/qk0szSc/dL0cEZf7w7pUyGlwNBVpjmcV8+FyBoUezmCftuim
vvXFvNY/wKau2D6kIj3D3SALUJL89GgkAilB+DS08H3ovjSPq3hRqOCNZtSMfQGw9zOFkUFKSBoP
Ybc/y/038b6pBz8FDgm2Mcy5pLCl4rPu0hQq4jeob2NBNmRXlyZfQ+ounBEbQ+m04HPTdUrq9lsC
szldF5KJA3jdRP510RbtwaZ9R/F0CN7WAlhkn9bRzEVy15aKKbKuVGe7WdLLc12yKnQHX6xhluZ0
nBcl+WBCaF5+ygs1kBDG5UPtwjC7/UvdUyRhMhm0FM3Tau4iqmeTzplpoyL6ikjzwgDyvfZHPam4
Xsh8UYCWT6AifXUCsDTB4H816vThWcnyhDFTmcAjgTAXUzA5vCPZJ8AmjmPIhd2HxbKOT0Iwt0ZR
tOpNQ3EFbHcww9pPVyridedDY4OIJUaVubHNKv9MyuSW/kNuar40CJtiX1BFiFVg/pw83WGYZBtd
Dd4SUNpY6lAIdes+gxQZWoCI3WvVrovYnvkfrbesyhnfo3A3ORAy9WNGh05h3ydAlDn8Oix7o6Qn
yVAQeg+ryMZmry2gKFOFPldhN9c8DIf+j+Z8j/gpSMws/S22yLMB9ezc5g5536uCubRCGVs1i/o/
iu5MX2pHdf8Upu6Up+niZ9Ys4EVuoDxt6V8mrdY8lV+A7gp4xrUndZTfuia/8RWhxnOFHG8fKwJg
nc3mCxLZbwuJnxdlez8KYy6p7lcLyJ1knajUhAfaiTdPe6LibIfhbGWLq+52JXaIUTGILfLLjIxB
TB1oKrj4X+6cwozqaV93acKGl9QpXws4zIyEWPwFV2kXs4qcDK1mT7vgFrwaN1JqD3WkkJL5Er8c
H9b+IluxUEZLs3UHEoz9NBIaipadqF+Xk1jnaAGax0uctThIzThC8ksTVFRlKVbLBkff9DHc7oO5
jOcEkmAOeY7cbUetNaRlzjFQ4XgYop2L35C4WycoEwBzQlyVCnzIUFTcHwe7+pBzyGYhCc4zaqnZ
t//cLR11LSfL2vkUZw3XPBzn/fcPWRHEUShm+v3UsLfaYuwpxWBkMshMBEbfCwsZTT20RD8bcPsg
5FO3aWfrn2mxE3UQNk4s8Y8EkqfrUzjqYZrTwSHJZcFjW31fOqEn75ejvfzymj+wolhzSleFaLRQ
8+Ndv6A/QNB3jCngNvwP79rX/iqqcysvLx28f6MByTS6I5BAqo+QYgwzQXKiEdXYDXuS/rF13LsB
UEgYXWOMYvUL6p+BABngwudH3v/3oMtyywdFoxTxz479w96Z74r5KYlxaYkGTuBQmc8kLohz+7Nm
Gq1bNjnTOeKCRKkD9I1z5LvjvVgPHfG6Lgc36REh2zBqIMMiqQFEfHCJJXKRyINjVMU8HfudS8Wh
VoKtUdB+XAIf2Pd9fEPoRW9pTJwUK+UYevewx6ZZRa4ha97AOm/TExHwQOU3mTXSIwW4jJX/Tz4Y
7E0QkfN2BBRSvTS3Q1wCto+Zq1bxntNpPSA8DlXLTCXC3ElDYSb4hxpfrQw1xG5LqNE7dPQPdu1Q
R9HTWkMtbL53HPni4UY7rg5xefXoQ50d7Dyq7DUx1GGkOa6ot6VqdfxRzmoENBsjEuhZ9Dsuex5w
cqLU+dQh5rjJTz3n9v4z2AQqiwQv2sDgyetoXz4kh/rWy3equMv8GR5e/Ji5RNLtBTjWVWIphtKV
xpwU5tcGXYfbCoHhitNUP8LhRE+Qk4QdOHIVvxfccvhhmurueuK2o/WvX1KWILHq1y1QAMlmUjhM
G9YfCWPiRMGx8WDKNCN9OCLKAH2kkBg3iw6BQQJmy95scVc7grp/olgDGO39CfGz7Dk4Uih53NXJ
1LJxi8Cq5+W2TjyHTMcQtK3Yc0X+Acb3eC6iBPhSkiPcJ7hrnXs8cbmzKYCQHk+fLqEfT2cnaRrf
kUUaiJDfjPTx8oVpGZSwOS/SrXXByczAvxm/c0mI2phsb8KTmDpOFYC81i6fopfW2roy8COhai7C
LAJUrWknl9pHJq0RSQ/QGibjWcIW9o0Xo9/KBWicHAIeC50dOcYnlrcHiBwaLZjFe4ZewGeBk3g4
JbOi461Fw/Lj4754ZIOMNFcQdy1Jl2xbYYTgKtFHWm79rDKKp0u50ukAbF76zINMM2Hm+oUHd7d0
sQ1CgKL6hS5CMVyt5C55BBvG/tNKhb5PwAt1ZzbCC1kjZtLgFqRz/sOOohsbgluQdEhHBA0F87dL
sXcbrctUaXcxtLu6WgReIqrDTzl8chFrVqwFAwK+P/Dv2JO2JwmuCVe9y8XRNky4uUfJNvqKvOJV
RIHdWBU/09AuIH6bUWFCi5zayU35aq7uv9zKiwXEg8KGM65mtAQdW1ypZ+13F2GWiAFy6oqtW1Gc
MQurwk80UT/7Y0UI/KhxcOXGUwagccVZQWDGnCu+V5tSNWo5PSE3kLxNJ5WjqnFxEmfPOnKZXs2k
TOCbNa7F2Zus9GxNh2NEay18HOTeOE0X2uW15o6bpAQ88CT/xPWq2NrTyU7R3WQ+cvAT9Fct0gtn
pd9tBUtsXFiXV1l4JcWCi6E/KmT21MXRrvPxOzjqtwFlj54LeuCd7HU36pRU57ce8MxKy/9RllwL
z/ic4SplXEhDnrV+5H2u2B4sJGrl5rEa9KpuUg88xutKF9Rc3998ZZrrjVSXXzDz+3G8LZhFNfOL
SUIx/HpXDxtZ2Upig5lA1CNtHed0hrAAYH7Jz+BAy9SvWKmjvLMuG7A7p1O3RTQgt77QIVpyVYVz
8kJU8Xbx455QRGBxUDW525lyf8hgrqGYpmfGaTrzboREAH03Gkh0qrUmpUxC2mr2D6ZmQCXJTNmr
+ThykYZSMH7VX0utXM/6+DjOv3b+ajC7ohNx3iGdS9i98C39iIRwLN+QiPpBho1EGGMhUSPKWY21
8xr4yqsTS38qwImhBc/X9QGKFzMFPTIfRRuJqTED0p1KUE81ErCrttF5z2sed3TbRcnRlyA9Dqt+
xhaCbonggiRTG/3WqDs7xrB3ZE4KkVDvl+SxnnNP0rzAyr7hD64bY/J4HIJjxrnJCH+nLpBQ/LfM
HzFAVSlsFD7lnzS0lB+EtiReNOx4ui3rYO0Mpzg4gEticoFp68uZWG8MF/y3z1nGHptmmoEdJxrr
zEd1+JjDOvtdcO3Shsdui8h0g6yr63KxPGv2DwgtC17ZrQbq9NNdQOLn6WesBTIV//2rT8Z/2oCi
aK7DIPx5GKa2Tubhz26CfqzpciIhEDiHIY7DsDaMZJLE9owRA2NI3bo4dNw9cpix/EqTG7VW4Zz8
gdAFuBID5t+k/AgQSvuXlLo7aevqcCJBFPM1CyBsWHPw/xhiaFgIuLUnsmclqVVf9QTNzg3V6mjx
iuasafnLM9GD9whgSRXK3GzWY1PYtfXFZs4ALNkSOyiQtesCQ46RYTQKHGQcC7aqvavl3lsz0cr3
Gl13zI44O3GCkrTxzrwH4WScEDNUSzzNOeBAKXlQumzY/SyGVSV+Xo/GPOJmtto9oLfeuP93Xpdd
mlAqsXKSbj4JlHGIccmQqQapG3DSzLNkJxl6epqsPzxZgJu8C2NFktUjQCAER3yZsQlFJGBRCrRD
Ntr6a7PdOCvhxR6DjRDASeSyVIQME3nNq496hzDnOhihA6NmWnuu4qDlpgD97CNvhz7Ro6bDI54M
jlCSfOWaC+Yq/JpMZ3xAaT/LG8OwM4eThvoHFOei+Nb15/8mXGh01R7rC1Ls1kxBeTBHhJDIII9z
W98iLJy8p0DQkhOULpb3s8ffdlTT9Iox/Vxm+JvACnM+KWgzPqmRbe3JOJwreQdHsuiUYxPzk/Aq
ti47n3g6sUaKW/V+PxIL305wU6NqFPQceUtWrfRQV7Wo30RGnSLKsnyeMryBCLqCpL5M2CZQQQb+
3QJ95yd+frFF5vW5qKS4GXJH96iT9CpJcjZTbJiwoXCLokp/cJG7WfCq/k/5i3velv4NUtWegV4e
85qD20Jp/cE3vGrA6HDlPGfQfpOJGaHllmlorWO5gC2P6CM39utJjj6YIzy2o3JG4QNyQRPhPhwk
cwlCwF6X2EweqTL9NNDM52mWp4GMYgrYlynALhxcCDKqvWhVQ/kjWNZbSGfl1dx8pAGkJrdvOgax
YYBqWoC3YSb7l5ZT0mu5LqYpNDZtJTWZ9ZTwPxVB8uwAA524KSrRcVsCaciw8SCqBu2yJTskFcWi
k80Peq1P7i8TXTZ+yFpNzbOsK6OwUq7ueigun+vrFKXsIh+Zh06a+hTPnkD0RYH8r8TT/42+6era
y8DFdPwdhRNTA3Effjydezztb005Xeso2C+gjUbCcvoa1e7uSYbFHJm1nCD91xAY+oo6FGRA16cg
DlVNO12rnm/l01/zLHizEWBNVT8lL+H4USuRu1roolYdB9/PGw6AsW9Ueopdlbrj6v4jpoS/P40f
CG+0LtqwcQUedQ06IDk3zxXGzozfgJenJ1Rl4uwqxGWaEui6Hy92NUbqgAB7256LBANrhE2cl5my
NGTZbSy1CQ0Zqj6tB3Cv9E5NIbNikuCbFNqjBFnKddyuvRJN178XnTo49fNunOqQm04UbMJBQEro
laF9dPPaeVB3ptIxzEXnXVSjyoDI66DIMapcP3PS3ALdpVQwb8Yhw7naF5ropBQpq4lmLGokgOGy
2yCl2rB9jQtdCV4o38GKTWVk5Sy4x3gqQS6D2+UHOKC6baUI53yyp8AcDwVDc2aa1TTDUtjNS5j2
XAu98VJ5Tt9KKglkhds6Ov4AcnHDqjuun0HC9uJ364sSwUCBEddGiZNxnRhu7iEoSLDSkwV3KVm+
76xXV4JoV07gBBo8r8aqAlXS9VLYtPlk9Fiqf2MeYX8F3Epob3j7tN1tBBAEp7b1P0PgfCCdJumB
GswUpD+gU4pze/BOrqO8ZOSAiuIPf3dnJj90tG++ZIFkTX4ZGB3JwTd+NjJ1uDTgxea37TsNFWE/
feaU76Ip4y6B3qYaY2T2Lo30OBfKlqzcVrau+eFOh6jtJTClXY1LbuBC0xZjSY+nI+nngFMwz2d4
zP8/tTjvdl6OGHvE3ygYQaZQspKWEkPPs6kcqMcwm3Me+Du46upG4hAojmtWLNgNF2pzvvlgTA1a
Mgv/TyVZ5tbbzzpOP/RnsXQqzyhfjmqrQZpx/mc53TEHu3FbGx8mCN8DtqK91pbKxypMETZp55hw
KR5w1+QTDQHcKYxiRDjFC/JaNaMffv793iC0G5F9gHBG/1Tb/9KBhQP1b24ytIXzsR97PZ2JL3vF
9Vfay9eAUpiwfgVrC/XDbn6hdPCoDODZI363q/GHcJ1YhnG8vieHGJGdHov86IZawCgC9Yq1NaRr
BpL6XFvzpV2KrEREgZprUuGXxUl9UG/NChFzBsdooMtDU9xok3qAbHZzJrjRqBpIr2thscboTmqR
N/53fQpBC57qQ9r0tfu/ouTgWR+2Sbu9rqc5fWv82UMWOOd3sdrRibgUuKVMEQNCnmjcev7/MG/e
iWuVo4C18u4zU+WxrazMePGAXY3ZUE4xc2KFqAAIWx0kbHQOgBMS542bCu+NsYfPQis5Bnak7Uyv
Slf9o3o8YwvRF1gvI+fCbvOjMa+lXsJUF5eCABsFGfISVojkDZxy558QPbh7FI2NMyI2Iozow2hc
7zZnpB7I4RcrJ7xBtqgKYU0/LQ85zCD6+DUNOlwHdgF7N3RKPXhr1EEP20WOJ7VDGGi4edm38HI3
Wqfzo/dfREe5z46LJOXvW7RvmpbDl5BUzAdfl66NAiF2AmNFJZcpnu7Q00KcdntPzcdIi0baNoO8
PNGm6IymO43ATXtnwJy/+IewX51ACXc0jR4Cl4ojGPnTFFCkR9s8+k50hDMTaS89suypTOBjEl8z
rSdgFj9vU6Gg5h8EtUJK7prFU2q1mQT19oFITFbYJhs+omESF74rEP3wXnjyAkaFlvCgVip2SdnJ
BeOK6EpgG5oNdlJifxWnmPkZ4IsFhCB9BwfTtim1yL9+Df4Mrzjv7ItnOiB3O/vbMtoz2VtReamT
sbWNK9Q14mnY1P2xv7RmZMdEHkKz7G8LrGjuPH3FJ05XoDbiAdS4bVgbQKKYVv35cUU7QWNOrYgm
4WYd4H/dPti/EjcMHhNWk0Rm0saMdePQmiUBvXdLQJpKN8ajMB05BygpwD8Gqn5BoOskBSDBrq76
qRMI2laMvs7LGnmHlfLW+G/oXdKbQEaUCPjOA/mAUUJwZCx1ldUKzbXDyDT4F7rb5TjAzBg+kjw/
2DcRL32S1QR5nQHdvR7khHtnNGangxTl5VYGC1VRCHHESJOxsTDyokDvmiQL2bCZCv8zVOsLFgC0
wE4pgHpa6M1SMSVOPwC85thhIvHP4W4Mi1Xok+rOIYakZbAjid4A8KAZTLqGCRGP8G6ptgYev0h8
c4lltewxm0qDQeNp1oS/gFN3gnN2lmJz1KkeR6a4T16Z7OR1ZA/0bRTpOv6z+iy56ZRloYlS94mV
ye68JF8yuJx9lQ+IGF1a+p5ZFCXmzs7rYoivXMl64zSrAQ1W4bNzq6YeMejWA2u94V4nkpVXcsEl
O2YoohrINZLOaaMB6pUTfFVTqmCLLQJ4B+mdcjiPMHfLQq5vpvSvmAxi9yCe77AzW1/1MffgSieS
gl5zHFRQHUyXRPuF9jd43Ka+WreiIj4yZDGRjXVTCJyG9yfZ4AhxvcAvPS7LKSLjkaF0S+NI1hyK
qbkZWY8F3IKplrti1fEhpB3WK1hv/DQBKWuh0daYeRwmYIBalNvf75nly4ZldTlp86GiRXy9sJbV
6Kk9QaI26d/U6NHQK0H34+XiTRaEygGJ8HGSJh/Cp5JtEEmLUxKovImuwgBaBPktBCShCNBZWJuk
puFXPh9J5wUtPYDVbk2UYhvXFdtm22o8W6zVJTluUMw/c/oBxb2mfy5FLK7LjkNW+6RHj8kv/vP8
ecLmTPWNE0yHbOkrRjyyM7+4ORn539ce07Idi6tKy6aOqP5sZqQovVEfc679YcRpWwPMvez4VGI7
6Dbyvb+zoUJ+sG3LzLaj2Lj28hHmfekbPMabKx+o/JleAv6G0mNqG3ljZt3rHKaruMnwekwli6Vl
pVUaDy2vLfjbveV147105kULliihg1EPPPHlwSO9pB8TwCBQ9ujaWDEiXGogRFKzKDFoHlq7NlRG
t+gbdeJFN2ifbv8quO/oO4HwNHr85e95lyqdk2AlIAayaXlWK7JbFQECldq+VUmYFhLhGMXzAEqS
P8Qp13UJcC1ZigR47OhmR2mKU+bMo0QTr7tnIByExbq5X8+aT4e2bv3A5odWKn+eOxkZiQZ3OpS8
8XuHCYGMq1GW/wp/ETjmyrPMwRbltfr2TNKaY1gwQRGb10efSiQeC3dpmVodY8/e9Vt5VNLNzQmS
ciLyzjg1tRKprDt3v4X0DlvKWBoUORFfrJ1cueAVUZl35Fc0piT2uVCdbE4kdEgtq7Z4QEFL+usQ
huQgsKZKJhM2HgPkuJWcnIFUtq13eR6njVQxVHXfVFoy5H1zdTE5A9vh49NwplkfPqHNDq16esiZ
WP23t4IO8PyH5oaJnDYZBmlJCKfn7576dpzHO2TEsBUSbyRHxjbrBrtsp2Qpj0fNUuVHuDGYue7I
Vo9Z7MVv2WQwjAhw5cf2pE3rymu3J9Y0OE8q6sDnqVXUfWliHAIM4PdQuURVQmvtWWuVVdJtr0IQ
aGYuZYf81JjCgcx1Vp3E1CSK/xT7X2v/UXR1PJtm5+fIU/uz+UPozVZn1IbB71JUA3mraH+RNkz4
3uNjrsAdLpIRgCUg06E4ZoGD7MGCcT1e90ZKroyNg9x0SdpLt4LVe/FjONaJca7lWx1aubCXyXps
3gjbCd1E0JF5rZQ+gIpKEpPUvRM+49CJsCXMg+gTJPQ0UVLJapizMsAILP9m+aIm0t1ve65pKpEB
Rkk0beha3E+bkcvUQkLD2nn02SXn4IUGD10NqgEGoGTyap5Ow+khL97CXxCCjUMdIRY7flejMYIx
OwCcIYxFxa4YdDGhmTuwPQmWYxtjF88sf9CTkk/Ho9lV4XkauTaRY2hiwvovdqEe5xMTEH3wXYjg
r3zzLipb6eXXabXj8dhWrQZVmTPSTdWh+W1gzBjgqTPaLADZG246MvRv8QPqTwiE4YmRNfiyLGYV
mW5gi1U7p9CR5LR6LbFw6xGNaQ/xkRYJ+PU1ucGA3qDu+aBSf0PPsXFG9KmnCk+FnLoE56k3mIiY
cz3PdclIIaCL80VimWM7Nnsrqe5Ff9yY7jYTJx99au+1KIuZKVD0rB3Y0whrDuy1exbwVkyCu+j+
vn+DoJ6nABuzAm8/0yuebYl9Gn53oteYDk3Fe0Z9fqK3ruA3+2wWd+wqANqfphcD3HXf/Rs6R3Au
9AvmlP/Ipy+z1qYPBWqwnS1MqeHbHamxLsQKRw/eUdAy8sd6egs5Ei7PpOIkAE0lopW5QdcoZFK9
k+3Cups5syucZSzhOPZu+QJsF9i3JAbTUsKDa/glCdYxSKBJ56vtnoACQAU99Bbvu7gphDtqtbpE
ZS1Bf5ZpZQHTKw5bAjn0OxzLcui2bB8TvAn2+55y2rUW9zXwn8YStOsvx8tEQ3Nllb606zBuRnN9
rKQ54mEKuOY7QsA6kZn4rBufiWHTA6DpIuK30GHAGKfBI+18q5yct+uMKOnTeLeug4Ny5KDehbvl
Fno6bPasHBGzaWVHff4bYCGTWMe+EPxVzmedsOmeHByTzFpJcmqxG47YaOv2Ig8BmOxQrX4LhuLy
lGmslNcmhPZqMvfSNWuxXezI3PSR97OULDGYiJqcMe5xnaigOVij0cli9b8G//AY6KqBT3Qlx9Px
HzHWKNh+DQDdpEaAUe+8owHL4Nak+Pou4BF2wFwnfJLJHj/Ea4O1Z6h/rvegWeWXBVb4KlX3iuAk
ejr9IPoasRBa4wv7GQ4BwmjFksQbBJ5fY9vPfX5KeyRgmM7IeAfRd64nVrFBGJW6BahYcjqZepkS
yTpH/1zNfft/62sW+OHprgFb683tIP80fMcU+MjjK3Ksejlgkzyrf/CmVN4IoyLiOFaEF6Y1VVLR
Wp1qkvaXz1rpDadCUKLoDAjd/fdrP+tgHH2h1XJkv6TVLPyxtRsLg00GssKTVzJYR2nVbSA9fTv5
IeSwHTRA453MJHu9hTR59PVNN6+NM2y/K81ugrJMTfvcW3Gml5unaat2cXQ2yzuMp008DWSQQvXV
tMHs8kq/DLkQcWaS0w+OGqMbph8OsYsv7b28vWoIKaC9egRGfA0MYdU8UA+IJ+jFRdBlGE6MNVcW
PzOt0grXbmh5wqk8pi1BLTrzatRI3g1n8EVUEANR9+6xZFnIs+p82XW16iXJTTpFxVvDPElpIK4E
eZ9HtS9f6jTEJ2TRDcUxemq0JWUIn7/jSWKC2IxmeLCy9PRy1tl48STe2XSLIPf4hp811siue62m
bQCFLnbAB/o2ANC6YVU/Oq+AeHDPTS5YI7+ZOhltMrSvFdAl5nZYg6eQdyN3wmT8nMnbFuEXPtie
ijppxTLTMxBHN6u97Di1yilWbJXngTZ+eXdCqMp3pikfBSv0uu2ntmaIBn1toKfzSTkIzcRq+39A
FsZAF+yDgJvoaEWIAztLVcC+BcEqHack9+/cVHZiGyP/5WWouDzF2WQ0I2YbE0x/Bdh1IEIuB/FK
BymMMHJEkEpkMCzCJTq/fBrxY6JR+WwjOEhPyh2vmKQprfYcseHiNnhiArGkZIdgYtw9FG169MSM
9IoUJ0LzezB5TIJ06uHN7yyt6Hvdnjgfh3qvmuuKItTBuKrODvtAes0lzNnSn1wJ55oNFPsvneF6
/T4licRsDsWq7lCxCQZAaRGrdqPWKq/qKu+n4CqEHSl+tBbwhhPvutdxLuW62eeyljG1upEdzOT+
iBVOvOLqEEV40fYkD5oi40ejumirfLB2HPyQ7wXSvmpggYVN1iHsniJ94ZGY0Vw8gx8ue7V+/lBE
orrLv50TxxIkgF3KgOsNISVgEgbBdWgglbeOGtYMNDaZzi5GsGVhjRUsDcMf0myl0HPtcA/w3ol+
8orLpnej0cJc3Y7qbNBDALiEwdqtoFORRfJTMd+3zesZZqCThTGasYlzt199PCwYXB2emaqdvCc1
nZGWLQB8sdeOPEYXeQ6yQQAwVJwdwkZkJsNgintjHXmg1ToX+S1cCvZgtxJdjujFHn3vNoK7kg3J
sTpd8z4UgR/4AhDmFCC1UpvOaLnP3j+T0qG4TwfOhsa8fVjCw3Jm1ObKbGffVUo1WHnSY9PIriTF
FkucuGwK3j8KPf633ErlixL1bbBQNFQcfnl6nsrPLydsWZWQhFtPILDkhIFd/d3u6qZuu2oSZPP0
Prx9EafxI67Sw+PyUY44d0FQ28rSOCoEf53NgH07lvXJwJqrj3/+EbHG+YFiTGHkmwb7Yg9at6/y
y1XDl9ZNEmz3s7eSxqygfCxFtQkzo575/FySsfwS0UpiZCgM6MsS+CAx1/JJOLSlYeOPjgB6+k5a
1WC/oBwzoFyokLKaQIkMVMudhFwoMbOu4yt9ldt18oVcNDalw1du9cyVC+/E3X/jLR1YzbZdaGjB
bCeEV/bqmIRtblR5chuUXhDjf/A6Vn+UeTwUtxuOzRraZT9N8E4u8zxHbSuM+m7P3pyZIQI6yDKG
1H0uZfb2gL1IUwxdNbVVh1dKqOw7PBK8WLYs9uLcstORdYTrVI2/RyzJISAunh0RquSjhIE7Lfud
gAYstcV8pN0DGQUdCqwwn01ujwwzBl9aC9+Xhs+fWj6zGl62HPQggRmck8OoYnkstCm3crZJ2vxd
6FlrZ0X3xPdDnTGuurPjwmpk1XRbIb0/nq4L27kixrG1RJOLyzEshHSYu6BYsDAv8yu8Gbdvc48a
z1rMT8YHC/wkkSUl36JcpZgnmV29LQHhE3iZrqUZdLZmzZJlGOlf4wTTTdsb0qUbLveylxitGpCS
pKmw0NacrZG+T0tjH9JFQ3rrO8UNdXAej+zsdz4wYx+dCNukZfkT1nJEd+iaxJhISITuYTtHgqIZ
e5MV/FcPuLcDJ1Rm/HXMJ11Iu61ONkGKcoc/Gw4eI23ZcwORD14x1DzOUmL68Ok9NVwdHHtx3rpL
VxOUAjaiIfXLhV9rS4cpZckgxBIAFtHCJZb0tHae4WAbQYB+DtDYASkJrBBcNvNSvb3vDnXV5io9
ziTb9+bGgrN32v9sUOg71yVeRpUkP3owaqmIAb9Uj76fzO7/WFajmhaA3TOfmO40U6ICAlz6i4fz
V7ylnLnU02p4QZpXvToTXpIBMev85/BjXYMo/qgCKbULCF+VxQLu2d1MVU7g2MBkNYXfif9cz1hG
nGlHe6mosuWUc0+tmk4NUvuhmYkETI34pu0bFmEVHUwGYxA4st+SFdXz0wzHdwjXAfwVQ+Cumc4A
c59e2hlbba/+4vtGvWfE1v+4SlrGtOcXQFsniBWnXLu6eTLMqYnwc6Ps/gn+M4WgEMQmH+7kbiZT
gplp0o9PuRzGqZ/9JrLaztNCxd3UnMqymUv5INi6l4TM7UCyrLIXyqvwih9Y9DeHGlL/Pvx2sbU5
4ndp0iU4MqQg6NUYZ86flS4aE+CYNs0XaZj9D58mybu44sNiHvI5fWWlyTrV/psLuNQT14KB/XpU
h85+AhE0Cjr0as0p20fcDgA5O47HHRA9mUkQuMmTemhkUd7xdCJ5T6ZjItm7sky23+P5NPm9TIfz
TVM9OEywKQq0yZYt0v/Z/XOzTGUNVXs4mHMuBYPbZ4Uvwd24CU0UlDnyTKLDWba1S+frr9To1bm3
MiEC0w0ZcXc/i0FLoGDUZIf6/s9fkOCT1ntn80Xoep0QlZkaJn+a/8QNPJtnNEQznFPvA0EEbDJN
Lz5ESva/d/wT5kpnxOw9Q6peuk71xyloVt/T+z8hl31NgscBvRnO3lZfvOuxIf9axd0MKadmkuJK
BebNohzxWcF898cLfhu/VlRcW0nxPqK/kBZtpejm56uNpUd08DNJuXwvYuJy7YQ1cn2rKyhFncFK
IHk3fXvvGRvWxwWw7s5nPo0ZwxZ6pOnaF6qgUxg6eAo7VoNQcRCmunMXv8lhgDXm+FUUkNLHigs7
AdASNX+vbIMRRdnc/DbKoGlJl22k079XTPQwTxAEL+/kCcb/6fQGezgrgDLnsD/v4guRRDLZaQhW
FYfs1B/JObkedKhj9bqJTbxpu/WU1m81JQaI0N/kcB/3t11mUnqGpKooE8FfvG5aDlfxK+UIu/5B
9WMHBO4nRWC7o5m6Ip1g6o2wD4TUu56Rw6+sVw1f6eDyIyOueoZvF3qbTa1Q6Ocf/ekH88hS/Wvv
S1rlSUNYvgePQrGlaEdgyD71YzL6DfkkzC4Sux4FqqDWZ0WeawYiZ8JISkyojztTbZFytsbtkmn/
olyh2VRhmJs9SH0ag91aYs5KApnuJWduWQH0FlvPvkEaosWEvU1yX5DIDX2KbFeTLVg0vSRNk16i
mYEaMQJlcm2X3yUckiOELMu67oziatKEBQQNjuH/xu6fy2/Xx+d90H/GTLVIV/b736R8rdVZ3nBG
nhsr7gp1PW2X48V2wYY5dAbILkVt5btUlnPfL/B4C6CGNgvD+uA0wOK0S35fIoXYBLItcl7tEsWW
nhkfVLHBr5QnfiIYgvIMYkOkFtdycVYxP8G+utmVUNkaDdCxCJGjYQqH4psQFTXLaYQhVpzWOenl
gBI/Jd/R7oqNsH5zN99/VOOZydpFUIg8c5JxCKMEi+oJT9RTIn6S2diWLQMX8DfKOWEw1ogz2Ob5
A8eGhO9kVJDsGe+v4/xUBt2YSL+EaODHZVVtvGb53W2UMAUHwkeeDxJPSpzQRbS9ZDdmNMV6T7e6
D37GFDrkGYjb4hrCviWlRkEgtsfma43pewrIxfaXRvDQLnYAWiYbnlDANPF+cs2Nzvu90QlkHgHM
pkuSyIkElwXb9BiYx2Fy+vuejBrxApOL+/NDuIU/nWLuIlXvdc2qTkhP0pwyMPzhLzzW1sIpbjMx
tb5u7tlkJ2aluXjm3PT8UIyFb9srRGgf1GVBblLNUFJimfpaiPIeltSKfjt7Rwr+UBWjn7wBCtXb
QlLbMODTeRXBRQivZ8PTW4a8i0LyF1ivD4LSnVYRYmejMjhjJ9lL8Y6cZKQQFnKK7dT9kEqcC0XT
a8wKsBoGE8yEot4eecrJuqLYP5sbBDVFoweSGSxTFjM4kxTsun7IPxw+BravdRiALyGEWG95c5GO
8yF/VLoi4VKAJrlpRzuD/kXnn5OreRQn9GC5do+PldRbCwc71+VsMYficZACBOXdDfiIemD06PqH
JH+G/Gn22nc9oz9j54FAZJAWNRIhvuyNpVrB9COWv9TDjUeQFMLgTpgIYx0BXkybudQiTDIrdMwr
JN5IZz8pE1B58ns3iyOAg8OjC+Y1G9kyjrIpDlmdlop+cZkrPxs6BXGbK4gdWsoEVdeoKMcXEh8m
+mihVa5r0a56/k3uBhfRQIsCs0qTh17Q4wd5Q7p4VdokeHE+dtxivpMCZk3yoxJAUtW7tOHys3zV
52nnRI5xch6SpfCNAvXpOXQiPqmIdyuMDSWL1CtHKa//Yd7lfrG/Rv9zi6yKb8H8Dm78+XNu/iiN
tFiuKBZmw6bHREbAL/r+XYbhAfkMrv4UVX7GSTop/TeWP31NfwtUnI88nQ9+b6N0hBmr9yrW0oz8
mzN9kj/a0tHoxMVdXW2cYImB7is3pZHFgBAjRuosdiVsmooblyE3NFL0Ua00OQlVAtHtO4EHvSLx
UPkot//qIbsg08IMe2QEGhexMpkCDj7fG+hDpw1IjRUtfpXhJGXTWYDbSLczxuJEIyR95njt74Dn
F8OtPJwgccA2gHfZd7XxLuk8amsA1DRTNnsiOJ2tL53fMjFxdyiNp55ZFDS0vwY+jf+E2cUmzhhX
R3TD4wEsRJyfiTUyJmIB6nU4xD2ZXDX/e1GPF6jtbIz2NjDyY0jlIqDb/IYVeGn2V4J2pTg5mroH
pgZhW41kP4dqgKOcfqRmrXbdFtqOiIPA/tD7d5u2RR6oOY6HQ/HELKgALOyFTyRMBS5hjR9r+jkF
Q1SisJZeiJIlYTp4dkXqia/5J3Yu7Hj+mVtUZErbs8czVTlpt5Ia6UBvYiryVV5VoOvyAY0r7QoC
2T5gholvm/FTxJvT8r5RIPddNhnBGV4PdZAGMbu6i+kHp0jDtydNCS1gUMmIzA3w04legn/2NpZJ
NmaBIhin50sUis73rUYie5ZQxSIXHMRegJYs/9a4KL3cHteNWUDZD1v+P1NPBbyK3R5N7ldBgkWc
27StaUn4ZgSBpv54BzymIpUilECtQRoWgG69ra0PBjZlAEj44lwx3j4Ltx+NcNHmcFeiKKTJHTf7
LfjxRsesGFB5+BGO4og5DGHSgct99nnMCS52IeKdQQu0ZlfJcLfGzNhpVCWxq3V+w3OThe9YAQ2x
Fq2QGMTNgd0DNRzuKObPzVWCuY9CW/0x2mgTHu50Pq3QBrRTS5AKIu5bzfLMjHwjQOMDDqUKqS8F
VVolALvmQvMWhRgeHNpNwb/wkTs7MvSsa13Glb1KJAxew5YIcAC9MFrHyvNX09A1ReD61cH5czZO
672rzHZIB8zPCk0q9K6+LRfFWo9xF8bzLYRHCIcXLaPS1nlsLiDKxZAI/7nLRVL405phtgSRehCr
1RV+Xd6iN+XoBLahfOG0qFUwjgNFuIusnwxFa3WnC+yMwyCKR0fkLoq1LR5Qfi2eUU8iJFOF78l+
zPS28RWL/Av470QooxliujYJrDyJ6vc+WcQ3ZX0/ZuraoppOl5WYmA1L5CjHwRqoRpImFMl0LNGg
LiyGHdZrNkJp2hMp8iboMCbXaA1+0Ft4PWOeBvV9pnuxQd2L7pQ9S9VUtYhsDvxNKdstjmZr9W/3
l5zw5Ub+ls+sV/W9w3iie38Jb+j60rLPfx7z2Oe/n9dRp+nY/FxInk2l65hBZeEZh5ztPM3i8TOM
khtG1MhhEkDGC6drp2/qPb+VEaC334SiAoiwNT0lRE4PYL0GgkJtEWu5qY1XMqokIFP3xp0gCMy8
saFH/Rh9WacJD87TCfZw434UruDIuMHYJZwbep47eu4bWBduLSfElzE0whTKpmya67DvTrG4s+oy
qZZTDpXfZHLpwLV4wjsVZZKm51snDjXBzI7wRd/Rp+Q6irbHmre2XP3XbLHfsEoRVwiKETeEb5w4
DS6DZ9HLXrLgjU9qIVkIeT59p5gR4toSeIeAUVFZE2q1Xnr9V/D4HwmzT0Uum+/vOjeKg7hIs8GZ
AOZJiuxExYWOCmNSaWXSFrimHRDqrZ/yrQlq4zy8UpoAMdqooyQFYaH7nstAd65AnlazsVK8u0wD
dxjEyQr0vl0UKtQhE+gtGVLmugA2IIRXr1gEEVzigWjUI6BC8wsZEyV/kK66jOQ2wCOsem6LK3i0
FXckTDtA8g84oe0wuqVm1nOX5DWm50NiO1ltDr4gpc6vHX0CfcxqiMGN3WZcjGjakR41FK02WzdA
VjhWRpkVm2t/t/jFacc8YHz1XTzLwDaQOl1YGkqmL7hp4WFa9Ttg+QQsilmqeVZ8hyjKTvghuVYg
Xs0oLy2aRvlahzcoiYRJY8MuYoSJa+1AD/UM6VhHXJfosHfYWlSBmkdsoZbEJmz2uMTvU1PSTffe
KDG4UCQ+l+bQi8ZdUR+xl5+iEzoFiC1Rgou5A8ntxsRx97vkKDy5/98aLdYCyfpprlA5CHvjg7fZ
jM4hv9WyAx1KJLzQUfclzaA0yvy+SuEKBLxwQFCpaX908VSMmV7CPoo5EE1ofuDHnHk5aVIHIH4P
C+R2eHfa8uROdV8EPf5y6LPaxBu+xqytwdufE1JrPL6sVR29ZQibPqbA577zFNsDR5CK05vPztLS
Z4b8Ba8AIfWRZ3q5AzaY5Ey0UY7l3TYUsQnQnhBowq5MZjECTZwN1E+I5LDKEgzexIlOv+zbprk8
Sg2XzGQEbVnxd4iLKWzjSTzucB2N2x4P22+NEmU+OlpakC3b/nJmk5kIzv9LMeJYQbIQ/M56wcU5
Lz3jVmlvSJ1D6Sciv7HYyVUNac7ibsxXjaUbubzSQQmEfs8LYM7xV3dleqbROEhBZU0HU3K5rxLK
93Xurz57s0V/SVotktX7CPLp5K29xMC6bB96S4buslT5YHOsX2iI78616cNZZ1Urf/EbxbCwpOMK
S8ynQRZ6ql7CAYAAzEhqGBaUIWehbshW1JEeZFmnTSj+4ANizEtwMx2yliHEy94LlRPwNDoqtzwP
MWRrrJJ6YMP5brcoW9L/+AlNElz/8LJj5Os7Sm9oaN0Zn8A7UFCaK49mIa8U4qnU199jkxRWxeh1
5R6qo49Iv0y3Mtc9IT8nAx9YWg6w1/aOxb9eGw6Q35OntwQ5muRvx86RKFIV3QoKiozn+YI5BtAV
oeqVSFUDWN/Q8OgWoQaBV2vb9qFtnddOQ4UeU0qw7Z0FnWRUmkzKkZBIHXXsk+Gnq7qLPAFSPkcP
k9MXOPK0Mmbfb9QIviSltVitNtQoYPoHh7QGjg6aVIpYYD2DV5uOlg2urN6yn4aXHDircBDClAoL
JVqgEuRFX8YIZVS7zWHHbx6fJCZ40ebNI6D322uqjEQEXJrYLFblcKf40GuNAzie3S9+Wrag24PM
nJGYhQC6iV3vvQe98aSlORcdszDtDLftVJrqCY82VGqWIqRrWTTSSyUQ8vstetnfzhl0LjwQTHco
XEWKTMk130Q+L93YOC8VaZqnjzLYZrLNhEhP11H2GnmYEroTnCeQ5/yDEtAQJkoelBoTMZHXKe6O
cPnLNMaVrCeYaLT1TXTaX7NeSBlxvAaOGz3lsMqinZdD5yPk2BVbVINM+OeSI3C7wN4JkXBMtcD/
8vEbM1/qO5x+QTCr3uhB8NmMC6qzje/qeWu7CjJtdlUcSy33dJQSSOBDjgG63Y0LK/szuJKG/Xv4
E2eDlbjrdN4fgWERKL6uZKep8GKhUBlbv/fQNokLn5wle+mgwNH+Bi6OxzGDNCdh9T+exJqIoLBR
xcWPeHoLtF8odhcyXEWt78jxseswub6EDaS2oWII8HxxxUp4pf8CCGcVHqVlppKQGiN1K+hn/Q6K
x8VQ3ROiCTkACF/xebgE2840nKEGhEckkIYwlRMs8ZC45iGdaM/3ZhpsA35NwT8vUBA3AQMdqhYT
9yTDHCyRTihHatRPl9RvMPAaCbQG+2ApXxfQltyZtXiv6tfM0d4bXyWKV+O8m5h3duW7hKmYBbqN
72Wu77i5RdEKX/zAKahwE/M0nTRgl9m8hhlq/qgL0QO5fuHNGc0s8oFNi/8BQPng4WwKtQICXkCg
DUHj7aK18BzBX3lRfdW+zIeJRq4ybkTxMNWk5ZE/l40nnzC5X33HIu6wHR8w/XoCQQuiKLEZv2Sx
JBwlm12K6PlyASlVrsNYqVAwqTEtVdtVCr2qIAjF8mg2t/XqCrsYPbbl267x5E83ig8Z7Q0PkL1X
DqJfwih56WCnTt0jOJ5hABjci6PdUFJrmDFKl73+CCpu5hoIjbEiVHcGVVDaXxJmd3UTN0gGAobo
rjwJvLd+b3H8jue6VQW1zhM4+gkm1oSu274Ej2uiWh2sYfVzn69yn/VNoy3Pl6xf8PCjVGPyXyCw
8DlCxjL7l2vIWYJulMxmmWQ++ZylIE1KdDVSVgTr0X+WWW/j2RqztXq+bWIjDKFCfLVhQIRPOaHI
++zOwS0kUQgt3knCOE7QSEmkvYhE6m9NotJtbxcX/vT8q+redHwVNf2WzM5JqAaS1lk3BiVQNfJ6
jSWNL8rjk5HAr+vsuArbFW0JhAyt8Qc2j4x4DyHIAjfmgNDLfnxLerb+8J0t7HZ+t4JYmMEwW0q+
V+fNCjhP0uxxeVRnALOJCk7l6ePdTA8mfY9fjKWTRAB/hJ+63UZbbf1OvbaS6Nr0V6Iz93mWckOK
jCMR5XDrur4pri9yya8nbWbJTkk2tl62b2HQ2gHm6PnV4yrok2p0U0aPICWF9xGICQ5NqqCssBiF
19uP8MtzLGCvvf9R8Wn8y87uJOTm136I39z//TztCL9VPF9v7eEww6cqJ24Wi+iFiFDNi1R2dwWf
7Xrd10qyahGBEw7bimvQQRV5k/QCrXJJm/GlRs1fgoek0z34E+adv6Ke+SK3MSdZiax78fE2OWc9
yxmMOE78FhWZFQaUVUkrUm7cKRf10S1Ltkv08lM6oTcdVesfBH3QH889CLBJzWVkzf8Jmj/kdBru
qTc7csuKmoSyrLyRureUsKAZBRf4jL5HiO1pR9FscCK2BKkgDOoZqN2Ong9BnmhZ3ozrVB7tiJCj
rDKjxUAXjkLeiILHXsG7swowcJb3QcXqe5x5y4aPNk9zLCb7g9w6QRN+U3iRWCEBw1EME1ccsNcb
RDRQlaMkh+ZMFaOYdwqTgp2lu2LH1Owookp6+dpRa1I/wQ/PQrtlLB4jmzJU649bKtpEyxe95Ms/
v/VGBBErIMQbdrMOQ4iqbq8oZ9k6mILBi2/ewGXznjWL9D7GhoizXbTAVwjcNQy3P8bGE1rAjUe/
+bpVwpa8hRGpMsqh22kl72IjeDtEC3zHRMq4pX3QCsm/FTV2x+KgzulUp6Ju89XwdmghO7VGj99D
YNDrJFaqU8BUeAAXEACsIHC9VYYYre6DHiZrn0pq6hWrV0zPHDtiAVWa/alNgjSJyrN0QIBkeuSp
GZxTkvBrpwUWYgAuYvlKCIxU2Jo82PH6zuOYp4uCzUz69aRs7LabPV1FiTNY1Vzf83v681Q2CFk8
PjDAliFCJEOB35Eci9+ucbcTrT9umKU4ZsiGWUEgws1Uhh0QvJB5Y47WCUlrSHsOzpvrgrKkaWE+
AYUriDQoKje/5yM2TSX4+/A7ZZ2KbCXHT15k2x0HMThA96zuToHDNBpCs0pAXL9P+ahnWJmtrLIc
rY920wrf9bS8LpGmbh4Wz49p5ru+vSIcktcpeoXF3ts/akYO+2I/NCgiw2W4TMbPN2OkFGpYZLcE
XavTghs3827Asz0dYOGMEfC4I18SGm0sa5FPAKYz+S/jY1UT6AmCblG63amalYc9Ed9mbg3ikYDq
wv+vfjB63w8l6KL9CdEW5z2MjWUF2DijNAQi5VtB6iXwRoNC6AL5vUj3BPdYY4dE45NJPB03jfDb
wUo7rDuZW1zc3POp7QXC5Xw0X4ryYLoM4lwYcrAF5HKexQumOD56S7CXMvQ16jqS5P5czELKAQfv
rBsHvU5e0kk9+Bz49nJlR20Xfb/tQfzp/krBBV5cGO5X5iFGWw22/HUAMVHzosc+cVENq1V3cmpD
yLLyBpqzF/upfVvETnUl8S2LeXveMDXTdEFfoBic36tXMY+X64DN9SstDhwLDr8gIw9GAX+StVbE
j1R1oOIElJSnnHgb1074mUce34R16KZcqN6jM0NFNtVD0bgkqYtnZdbGqsYJNLOdsJAE5itGXUPF
xOshmIH/LgdYu77JvvIAtGBuIog+xyXb2eg6QCEBfpHWiE9ukJMagCnKXcLb/NhaAX6bOXoy4qqk
zk+CyIu+lbSoSObfcoOeJVg80fqq1WMpoCh/4e6SIExCo0U8J7hTZEAFwNky2R4kSpqtMDDVkbOJ
Pkdvy3r0r6lPODsvKlXWA4KJdXu4Zx6oooB104ydeKbltXaZEj/fl+G2esapg/Dxf68Li/4d5jJT
jazSaijGHEiEvZzgcClY5E/UcD1ZiEf1/uFUEdzpp3dLy4JcO69MvvsXWbc2DDbA+jl5LZm9fCcH
3++68SLLI7KJeBJyHZYARFMjr68OYXWHu3KE3EwlgKcKLArUxfwqHoGKDez4Mqo/rwr0z56bO3y0
NhKrGYIEdgjw4y7SLqaK2VcyiStRDOH2IvKCZP7AQoWRMgwkCsW6hj5WSEYpnV69OQsqlw4WHfhI
2NtOSKadyPFQYv+PWEhMrCXdAJOhW1hdzs0u+7L2X3kKKh+ECB1cryZgIn12G3M6kBy3CH+QfsZk
7EYdVfZEy4hFH2nbom6ESPp4qHcDexW92LqZFgwsTgZv2iawov9OqGzVcBP9uYIOpaTnbAswSPL7
LtTc9qxsGHDr8FfSoOOtDtKSUSJp4EaNeea9InZ+wHkYAOgr4UoXBEELhkbDkGo0MZdYErH7Xf4r
K8hcjjXakLO6bZgql2mBj+lCLOvrAsonVaDV1Gj37TKXaQ9oy2bVbpJWTxOAGeJXG4eZrzy11B7W
1Zo8C0+8/36RvQCcpcUTtsNGZWTLkAZbatLM+9VJhsoiw8Ls0CGzj/Yb++6iddU3CZxkzWYzZqFl
XfHqmO1RLWMQueoQcmSbI1wAB473+TodH9EufFsU8NX34aGwbv0Ukoq0LiEvCtU10+HlbOWYQam3
JkZ2o+f5WtWtwAmmKaG/yRhs/cUuRboeYsaW32+amT18/o3arLEIIdUyfxcgFbHUXCr/yY+Fwn6k
v/WZFCChYAaJ+DSpdxxQOSwScnZqadPl8IPnV+qxDg4AEOlTZWzn9jXgHNmTuFqT9ma8Q6av86EI
K8og+3YHJogoGonuG8cqRNtZYgfkjZMS2PTPfy/kGn1LaC7uiizOm4Lgdp+gOkc+dPIM7qEXump9
UaH7o6HXg65OnPZXrtLmCA9T+oFDAySuqkI9YK2QmDEld4iKJdHdQQOWB15AhPPpjzIGj4HGVrfu
p+WvdwdWmnQxb+RYnV1vtGoTUt68ma+ik+rRO+Rk2FjzvedPQQbu+jhw9f+hdvfyFEmfl5t1/Ivq
VpqPIMdTtyhF+w15OdU/x1XPz03Wiechg2DSP7MiK1HyiPX8d3pCN3toDOgSxoW9OwW+DLvaDu6L
2PpeHjpmlj6jP7G7JxHYQK02C7QfE8Ka2OiU3X8QRVoXJOMcbAZ/vR2FTPSG6B0vxKruic/Goj9c
6MZMqLhZSLerUxuKFgCZXZh8rPr3xaD+CXU9XCazxPO459YBsoMIpALog7cILCrk/A0Drb56AGuS
ae9uBI8v+su1uXm8alPdmGVLWbSCAPufnEuELs92E6iWyPFGUE+l4RA9Ou1G0YIAzBPZOrAuuqD/
v7X6tgRJLHL7LHOWyW6bqFbkh2CkZG4gGrTynF2Y+DDBHAJMzJh98bDTMng3BTOZuy9pi7ysbWu2
Gn0ZPYXPdh7i7SXyc0PG5KPH1jEqKXLi3gk3RQRioNsgPevC3gCIMfrsALo1PKCdwGzMsD023dAH
tm+Xb/R3r/KINZlLYMpCW6zQaWzUJDjhYc1IbFgl7CiG2C8HscyTYxxnXkRaWGPuwcqHFu4UH5Ui
k5hoES5XqGaRIu/qhY4+Z3Xpx0pZbjmpKeNeN18/tUbr2v2zeEYq1n0IqR3bmRpwOkAmga1HL65p
y+LvqadNnVd3IrBfZX4K19vPRqiL3Ud8jGF3y4w9UIn5fkXf+iSacWRCynOny7fIr9FPUMtiFqAG
OVEI50wmAsKR5AVIHiqlNvbFqSqlX4CNQbw5uwgfOKB+Oq0gU46eCeAnLj05kNiKl/Mda25QSFiN
yeDDtBUv8Cn58nEDSNsyy/AHSQ+WQ/GVPICuZOCUTNKo0uLWhXgSyt0XVWCCKG0l80cBcbw9+zGe
Nxz7eMZ6p1o45EBoAzKckj4snkJ/7TUAh3nZBaO8M8LxUqdEnw07/YVpGz7qjMCCuFyhdhRFou7Q
NY53Gn6zu4zAyCulhbfhnfxwgGC/w8TT4xyGKwf1KX0c8O8vC1dXshLTMdiZD9LGIFy50AwdbWW0
N4mzaSgA5WRYpEfl2b1o0R0PKuLK6SHOG3Dc1E25tNfsrHtG1eY7rAsnDlcy8bK2UqwUAacjiML8
WCGCsjfAAoKqj49918rtGOKCldCu8u5LlObDFK9gogbVVvsLuJ5adkZO2Ea9gmZGjK0P8jVvhW7o
yZBUy9Tm9pyrxluPRD/IWsEAf8z+r7dwUgbWXKorXX6VIIHetBia/zwwT8ez+3jzL+lOqZWK3dv4
PUFCmxWV5NVyC7pFDSrDz8lQl92F+19N2K4Bw0ojW5H9nHoPQ+cku1hR/K8pOIuBrDCfush14pyq
JEaFgJ8pHfeNRFL+BBsbksNRH+0PbxgXHPB2ACvlSIcbQk9KyWcMmFRvcj83mAgnfq3rijr5YATh
KiIXUFnEpFWJQGf84XWtxituWOxHYodLlFgvCioDjxw/ijDev0cc86HgbnHZgUZsJzoOfWVWjhwz
SBZj1UoJwLr9WBB4ENMvWy1NCBd71Y7gm4TQ4fPl0/nwH7Wwim4D6ZB9VkQPcTrDcrQ9IsQBnn4H
32UXrBODNAGcWuRDyz9RFVOhTfhmxTlegR1Z+s8eAc11nUdMLJiez+2sPECQvM2uD73f4NOgv79R
v1dmKCygW1XqRQdAbyCe7MmiqhyJ7l5VQAymu3GrhVte8ufVR1sQ+lBgXxl01pbi0qIW+yGIpRsR
t+0hLpQ6jv+ipQelukguUl5xWqds8O0DotqDcq0stucIWuhIfG5ZMCEpyzW//BUvrA46dU0Su6VL
Mh+qGxMMX8CWwnEFuOixedk7EMxnl19bBB18pFotyI0wGIgnJ/UP3Hv7crPhAqdJH5TZy6i/rsW7
oYigJ04lx5NdoB6ddjwwUZ+hZ1s66SF4d+f9ZSQIs6IBztlmYJLLYQxduKHnms+gjxGdreWmGNqS
gxnLRAUb+N8zlBaZXKzhzwkBoYkzls8j0r2QEJQfyc/zbDFDHLHD0rdKGAB1UJtVfiB3Uah2aNEK
xQUHjwcnYADkod9QZPFoMynom248X80etAmUEJfTWaPpwpmc9NfEea07hK7ySWmlY6gVRfht4su2
nW8uUNwNODKnIsbafWDI/LFUv99DTFzB0zJY55Z6SseXoLYkVWEWRsih92WP9CRxM2fe46Dq+tuW
8cj7sBbFJjDxOohxuQc5fyK0XVTR+CnqKs9SOiZ0lZAKWnmHYKYAEF7Un1c8ov9xWagS3PAdD8J4
68BkELLrJtcPWHPyscR+8/RIQfZIHh1G/4kKtbZtfuVT3gOLL6W9bDhsHnT5BK8e7/+b/E5PpAET
KLlyekIKfPAJi1y4Wql/u/pNCcXBiI5tSyF7CD83m5oWCOX+fgCmcjjKcD7qiHYvlek66go81vWv
iYgJTA/2nGf+JrHvnIfNzF6u5WAbmDj321VLBLZ/nq+rJ/xRTSp40obqm796pyZ5eeAPHHv22Vtd
4n/OMjifnHr7XYulON3BS28QqQaXv0FrwhJU0CQNMbRiWX55l8w2syz6fyIXp39v+jM1aRC26DvD
jxDs0PheKCii7xJB3T15mXJ+VdxMtUfyJeJ700/Sqt19AIyMgiBkSfH+wd2c9wIULunG9CGK1mCV
CJamdz8kerpnsUllu5tVl5zW4qILng73gcXgkVWu0rzX2zc4AqHwiU2hMoJXUSoLVCDb+HGDQT5W
i+sE3ae0KIOqRwlXBb4OcTPSSTduGi0ogZV2jmMzeMOvFeAuafGvN5ONcuRlYaCl8CerqKd+V1F7
4iPCXxwBTKDLp328t7rdz8FzripvGpA2Kmm6u1jBjoTYI3ew9BcV4gCHqC2hZQqAve1s1TuDub+g
hG/KL2aDbcfEP6FZLtF/D3HPiIR9SnycoSbceJ7CxPpIG0A6vi85jbIaHLOXP/0J4SbOc338DGM3
qWeqmWe0O0ARdDMee8pfZPSvv7FEaIyOuw0/0Z5z5HzJloFoaBsNKtbdDwUqD5XXx+b0YWV2Zqe/
uJDjFb4HqZlZAEElNxhneAkKE5l+o5FV3G2yiFdN7RR2lZaO1ft+YFGICYvnB3KHN9iRjNTue8eX
XZuuXz8xtb5/1g9nybwdLJrpghC5PCrpG8z6/IHikyRsKPuIdOlgURZ3HsyZIbDljUNdB8EiOwBU
q8kLt88YCTBioH90VUL9h6dkSi5NJlMIwICHQp9+gw4eoyjBdYkDBKgbJpPOqQqOvZcwdRPIT+Gf
7MROyOSsoDWFQEgvll8eKZdohGKUuB4v9K6+DgtxHZB78mnlLe84FB6+FgC4ZWKlU9RCfxW9mV+a
KFnHCTpLaA6unz6BljJwHM8oPzLdGoWas+KOAFD8OFQtSxCS8VM54i/C976K8uQ8tqh5cZXl30cf
iCYK5qbLGRy9st3FHRxf+kP6sAbC1nHzw37HsoKkQV3SxAearH+X1BJ12KOu9KqSHFgOqsuUETf5
Rl7ooLqA2tf26QnpkPyywHW2tubx/o9VBBud0e23AMHdeeFz6kyCdk6Vfm0oxoTptM8C/K/Ac9vH
GlhYF5BD9pnj29kFAQyMgQYJ7km1dqtbgEwmvrI+xTUjfyR2Gye0vaORrAJ6YlK377j5QTxE4RiE
V3j3Von+FnxaGHwduLib0/rOqe6AbnCtWAiU/xh8CSZjXOdnCbYCW2rY05qfjuPKB5c/YaCYd1PL
Wy14BUrZ0iTzhANP4AEF6EYkr2+n0FPDYJPSHNL5fUN9lxY0HtXI/ITjpDB0n1uw07ufd0oPkv+U
aGN3ZDPeaWA+UhkkebLR9yJ6q3o4tXJ39QSaVPkgrHkNd5o4O1DtgExvhguRoFVHIB3hxezfLjws
VnM2aqJa0e2N0durA9uvezAqTRcethwLScm6pwfIJGUT3CVcSq6dmU/2ikuvM5sVPflV3yN9lGu9
7G4VnkRDnj0kLcMu+APkTchcdZ2KApS7T5pe3k8P4EZbAr/DYHDoRuYnSlpF+mUz8VozTZtsdRCM
min+g//yZubjBtGq7IRQFpUMk1dR6+QBlfeOWgmOrLR8dux+745AaRz8aVRTRNUX3j6y3Sjb34ag
+aOqWGg29b9HkMMiU8tUbGL6KM0KPARrWfdiko5uG6w0bjBrxx5E/ItetsoM0dHBob94aip82XWX
BWCwyI+sbnaFwaJ1dE5TYZ150FHmTO08xFfrhOROn8O9O6LwugqSIu2BDEH9vKiN6rPB2TRNHFhm
DLgdED+h/ZMS6pv1CRbjyetBS2mjuyU0OaYdEXD8OCxp+6XFLyNSe8N8aEQLk1ZJR4ztT/HwyDW7
xJGMMmDpyYsffTtm6SK3QHxF/IOT7oA1YAsdF0oSHonKUtqLuz0aXH+25FR53gc3YyejBIdM5dcy
6tD+4CEnlW05M8nhmWeO6fLCHO2fkJV2MWLSrY8niuYy+Ioe88P9eTXWpulStYnOosDFY0e0cABX
Po5TRwr9qG2+rU6E5OstNasEKycisT+Y66stT1GCYXp8GeGpZcyX/eeyQSo30kTzem7dnHe6K3yU
gWN22y6GqvngA4FK8x06MGedBrd8XVRKEcpMVFtkrxBUTdkWH5yxP6oel/6rzPCuSYNP5bLtjGR7
g2OeFkptWo9iqJUhSY/URq6SkEx+Gll2Y/qOgCNqVXrxVQGuRrZt/CTBaQa1jap5h+0J35Ob81UC
dBPF+YeXchpgv0fHngKcTZvT4G8pZUo706uGoFeLVQDPfxWXXKkSmPhi970bDrEWRLR0NophI+pg
ogly9ccjpZ6KwYdoaV7OHCvHranpkROd1D/PpBr8BzijZ4BY9NZCep/zsndDcVLQeAvySt7/eyWj
4b7tuy/qkXVSJDpt9Qx8KD1BRDyj0fWCLWeWRo6mWC1s/8B8kFllpeDvRPG9ncKjYsA3iQEBjkwK
47vTPRy4o+0nyse2aoo3aYo9Hrhch1sBfdUxhyfh02uLGTZpRgyS4mSi95N2TaDqWR8Mo2q5dQvs
YFBX0godI/a6gvQSjKw56O6ITXpYhBQKPMptuqEj1quoV1LPNCuXhEZP7nldCuDsClrL90kOki2x
b05z1YrPLCqpbG6TJYZ0pwKP5BEC9Q3NO6JQRHnwfkBEoM4kTN+Or2X7r6fsCLzViRhJX2vZkwLL
QwtHitliyv5KsStWHL6Sohaf6+5ti8gEEC+1Kjb3HI9do1vAkStjf0VBrlSKVwu6scKs+VDxGyML
E29+69KdJLxphH9Tbsz556+vNFZp8May958ox31tKvc7kIJm8OOrAdJHfk1bEV7ecnpYhxLTs9FS
cKSbj0F6oA9J9AURaj6KyvdJ2qKYcuE9LsTHEvti+N8/07mPOWrCCkifBCXv2K+kQwDjZJmMPkHr
XrgwnT7uMuAIIAsvcjWs/UM1xHIug7vLTecqBqecdehyxXjAusV/NA7ocOxEij6prCQ6ULomLk6m
MtK3HBDNiVEVyxhi6qGjUOoOzDwhmv9XoXRR7GvoZh402A4MfF35akpGpFG/piCPF2Fnj/nFVwKr
wJWFbP4o8NoiTdu9wlD4izeI2C69v5Rr1Sz5TcoZi4MFdmOMW3Yk6rRyPQmbyyl4/beDETOZoJ06
Q8DPAzBoJpDP1SkI/v2JXQh0/d5fS1QwgyobkK9gh7t3MFuHUMJ+qZpC0bltGVHNlkO1SB7KkYsw
WUQYUqvhNL20xj38BHqFBm/i8tsbKLv7TR21Th8UOPYWcdCKIvnzwjxtj0sQRcJnplc0gNuLbc/y
gC/GgExECSYycOeWj1TKghkv54jDdil89qDz53rHsdr2e7rv+i7wWuxZSR4MPGZNirWpHdMlxqRK
384E1ZnskeE9nYE3Ugx1iS/VtMfgP5yLFn8NGgilwxJwZozYhPyYHukNle4NAVm3tI6AHI3PWFhG
BnLYCcu5zPtJeDT7XkzMF1V/YQZRqpl5Aw3nrvAURCD4A0/IiQEB5WZDUQ1h4Q2Jav1w+KN0WnBU
TD5SvPkCESJ2JiPEznCOPMqbbW3LNOgWav8H9ssMtS61tR6ZI6G3RL11n+a1y/OkdnYyVJPut7vb
ljE6VCnKg9J6CTOlAml7cvzVAxyLBryc1xHmWRXFI/bQ5uUjNYp15PzgmPx+og3Y7Nosz6TFxfd0
Uw/+3fH+0Rwg4IcJ5dM/ubCaeQidgjMM6DcyCoYhYXIyYfurK9h8OhCyCK4M/zegYbtZtsXyKkkz
q3T8rFPWlYv4mubvjYDUVuLjdvuCaVtQqjtA4Sby5yjT8qAI2D7ZVq/DIzHdJxz1V24ZNx8/T/4t
ajV6drZWacCQaEPMpQ51kvO/+FlkBoNfOv7TWqNYO2OAMGAOam80/xiiLBgyYGYqqEvUMlgXZwcc
JO/Uk3AQLvKXc/9Jq8lfmPkU3sHnljUr2FTqeBj1/9i7qw8gJAFJdAJGHIkt3TNrvY2Zt+F9ZiC6
kr2nfIkWBZMVsp/mUIM8Qq5bf/O62io0iHgIs0ydybVVlmP1TSM48Qgt37lvK3el1qDXdnF0gRjn
bMCI0FBVS1bBt/dbzFt8bKIhJMTYP6qfG3obeJhUj6Hm5BlvlPW93bwE5ZKnK4RnWikT2HuI//9L
nkDIcqpvmJM1BiKfP1BdIUPyBdaEb0gLLmkogrF2cyNxjv0N8mhv6XRxJMzZqEAbruTsW17gkHzD
7SMihtJs+M56jJ0cCD+7vWhneQVLtq36wJC8UpMsVb276OKotQ8yLjhvP/cOTn7x9pAlhFkSqQ0v
MIQwtBekXs32Wc+5oIez9QGmHsQSFVy5wm4YwfMG2Xj/SU8a+bUu9BCFknnMBe/Zdq7quF8apdbe
g5tmsSeVBKfSIKtzB6qqQvvYKkQ3VIcxnc0WzNiUjTfmf1+u6I7yfAXH9ZPAU5vsnGwBWG/smf+L
2AMKCbapJ7xeP+Ae4lIpGD6T9Z21CELyud8SXNqf5lfAs/0/MKffy0PQPHs649nrmhq0MsckOp3l
qBvnSudCEXbOOYRfu6ur8s0ryjW2olzM87x3r4JwmXLAj7uIJCeseuZjxoffDquYI0njC874U4ko
lIPVeEHRBIJQa8TWb394CV5CA5dkzRZJwRGhugywrLLRA76NqgxxPLAyaIdmcBHbMuXZ2r4bkSt6
rpecVbB+D+YZeQLfqmFU5aPsM56DE9AlrAQbk3aWW55vAXG8zeCiGkf4rOqGH2lJgZn8UPZJPx7C
d4+bOSnguxUtrSCJufs0lgLhlw4Q1R3ajO8/OsSwfUdCwIxnTSt2n9QelDx4TE7WTNJmp7hSCOkR
mlacgZZNFwVWHnF5bI7YwIiND520R8FATxchAaV9q//2Gqv3SFv3Km4v96H33j/+ZzcgBkrJSJGa
gTX9nBTnTtMXrj1bXmlsMqni45Q0yNTCNeTVzOTKTTXw9icNFlkiYtV/x2gbctoiG2I6AIqzqqiX
3Ry6qJtG9+fl57crHmcl8jYT4VsmhZzu1JQMCoA2Lq8fqftfoDhoUjH1b1FaZpS0/Iiku7xdL2UU
V6mhlK4akVUPAeDF7fmgddYiqzQwLfhTMVY1LDB00kPiYav5Qf9qNKoAJtp0NAi6kuCbdwLuM58v
M0rVJzliYWzRGQBBxiOKNR29QUQ4iVlpidC4SxfoZ6nmN3N3dvAE511jIo+18eQFjtya24DvMP6j
sTbgjG+801LHU570krtnQ38oES8vlIEn7VXgovrLo3hQWTNhZO810cEIWXRCpSmbmw5NKsdtCfdZ
Y2Jpl+XHeXq1URYkGW1//glwJQKB4i8HdtZEEJLF6vOkaIX3ES617HG3eiSTJdNIZz7SF1aFMz9r
e8hC7fWmhY3vxV1yo8hQ4/2EFHpp4n1lAe0RbdMeFJyV+hS69gdYmtxOWvc/76qXS/bSF66Ogk+/
jiQF6AFUAMrfpKc7jeQ19r3SqVg8x8g5yWwlm6XhAoc2s9FG3put+MTniH+zudyTh7uAo/txdHxd
Z+dxPAYQszi0WI9wmaxb77wXgz14m1mKubYTdRYZQhq6VNgOtSizNRoS+MJpMhRX88BXHTHslhaK
FPQYYLYhsMFh2Ckm0L1H1bFIxs4J0ZIQervVfBOWEdfnORMIsiHF/FLKSJ4JY/dWKgsIWAvyjdSm
tcK2+K+puG0QiCH03fdPbN0IM8XIKJk+sv//8gtnyc6I+Vty/I1Z7T8rSPbsHDxEyWMS50ZIfegx
aZwWrwh3AewBF5qdv+So43dH32i8HEHwAFS0ChIhymNqq1rj0EmUmmQHZU+fhY1rNpRNkW6DBb6c
yXnAK/U+F3ffIlEShpt+KXTVrDGGTmy5nuqfEsIZCKMmYCEQlB0fFPUKnWTPwZntWLTJSRKvWlNc
TrimqDcrrSzEumM2UFSPrAUIcHkUFP4EajU8hNCsHwGptaW9+QU/mU186M/xliIzx1GVGwrqm6cP
1IFwA2wqQ7u8MZ3Iua/0nsQsXDC5Lu67NQsWb0Y5vLTPaWa/Bbpsnrzxlr9BvBhaWpDi+Z5YLY1U
gjgZ8cgJ08NF0zBKbLCqyg6UXs5qfIQASMuxTwqHR8r/Fi/PXNkmKIsibIM1bQcJmCFDfXRj3Waj
FYNRxNZgs0laXS3A8HeLIg8SVSvWW8dLfxRqP/0opDstpJsgh2fZl5E5NpxrIsg5RTDLkODlKXjH
aeMk8WxVyR+PrReblieb3kYpLsQAdjIqC6r3MC5l4+WQ2EXqw0WHUVCFRCHohzWBfXMGstjcAd8h
zLO0hBrcdjfeaOByISosWZebfDxaKEAhgBXnggidyIhaKOi5+7rr1wucDvz3aaWKBoLSr6lGRqUJ
eZFAwIMY1iECiEpIK57il9yJCp1i+BhMuhZ8xl7XJqHUMxFThn0oWjKrfO2pg6e/0zhu0GpZ2O2I
AaLrJ39F8Z+wtA3swD0qffh2AsWH9guaByBW5N3vXdXi6Ok4UM1s+VGHXExbxh3aRBD8vkaHtgv+
odKd/ocfwymAoBPvHdbIuPfXrEZfEO8gg3/vrMUEC5bS/wcxocZ6pU0IphgXH14KdeUPxOUHQ4Ag
gxtRI9HZ7uLRk+ZsnZucUeHfWtczIppT/F0yMRbXACgVKo2vbU8pJ7/Z7c7qsklWGaUbDVADeyIm
3T1t2qLIspi6AaJeO2KTSSGQeYZiLD2eW7ZFcpP0F3PhmI8xbnLrCJWj2We12htUAbRv4T+Q4I6K
uUmNXY+Yddz4nVIKof9DzY/0xPkQu1+muJe6QAWZ7I6F+XrcPyOL8EYKfUzqKuDDYo2xlIdeVjfQ
kZYlVRkUpXghI1EzJnEPOcM/LqSAjIHtjEexk9ypm97QnMH6EbszzuuBA5nrP/tn1BO2s92x9pSJ
41eXwPPTKymQTEs4LlcI+Yg9lc9Bd9N7069fWUgJmqIN2VslL1MP/kLpl6pX5hE+MQc06ajoDFK0
lkv6DfDKkiGg2sroD1ZCDFxs/uM2uFLuaJO211WERxh6l35ZUkBius9FxrjM6rD1W6FOwZMTs0n4
JrKx9vFW8VN3wJ1tkzgg4nVH85RLS5EdsGspeO9WFL5JxpdjtkupgY/oCKAXzMovI3Dma+rvj76C
QMF0hombMi6NksiUjHieOutmONtD72oXrhvtrllNlKgXBBY9QWTplXGqxHpudt+bdI7ApBZT4JOw
dR9WEmC81SHB5CinXrlNPilamfrxMehNPxG2PMbIVZvkp/PLUX4VgB/w3sdJA4Ea948jMhw4lh0T
xrf2sI5QoSOX0f9lK0wMJzP8bI2euNEod21wi709HTy48HlGDLvrL1mrqajTq9C8cuEW56CmQBV9
8kspNeRReGPWe7QBFVjrPFTKtgsgkgQ5R+jmIwJcVLaxbiuoTboun7ZLhuSUKS6tbqcxz2FL3gmJ
PI0IMPCmEpGgVQ/SDIyMb3qML6MJsxRTERi4dXdS3jFYXONassySC1hSJIzEiwsY0AY1wvpEn8W8
wPozHqYElw9aAog24W426qq04fGS/84nmqhXGRxKTPCSQPH0KLa3Mz4WDtDqq9QcSZjbctvhHicN
BaqWz9UKOHWG8HG+uifKbvuuKPDfGkjpRdTWZ8ilMvebIaQKJZyo0uRd6XDIVE9Ni1u6j0HUs9N3
Tl0u+bl6ouNAQxBSyMkSuZp2hBdp8vflQk9vEsIwZz2Fnjph5NnYMNVEK+5OK/i5K5ezp0ACJnTn
+A/PLQwt3KVvA6cnsZIjcNkHiHokMsQM9oyPFYSJj47WKbb5lpYnY5iD5LMPGMBEPemRp0OMjD/t
r32XdXwHU1GvFMFl3ZeviEiCzim0Bm2LMD8ZDenlDhFb1APJMCzNUqO9pXRUAGRwrWEFx6Mq2oRc
SIMWpF7jm4aqU+hmObkXs5X3E/Xwiyl7X7Pc7cSP4g0b5DHhwGNB1q8UKGX6TQqZ5LkXus5KP0EL
6UeK7iYSjS8C/bD22F4P2GQR3eUvn1PUmGXQvWhRkDZJCe7xKfalFa7eZTk94bVqLk1iBFIkAyLe
y0JUsImATz0OfCneu5OYqD/DRYKTsjR+ISk05C9WeQkJK3L5nuN/mevA04WF6xWStlEC6ooyQvlS
/5W87rDBPygXLVTFjPt+s/vHx+GtoUi39VLg5rgzTQJ02oEoHzJvDlExG4VaQCEu6jFd7bcSoyAF
OxMnPu0RCDYZpdqUhjqv849e/4jHvCtbcDz6sSn4nkoU0ENML+EjSID8bqk2qAbP3S4DsS80+98D
LCeFbSZiou6vH9IeoGcf9UOH4N0bwjHLOvO7Z3g+RelPEGaKAq2zmSdZzV1rgNvAHLW6djUTwxsH
hsZojl03BwX4mZJp93GxTt687+oKQjkYO1lmS//ooDC0KTN5ScQcuH0wNhV6HIJTwUgIMPnLTqCx
ZnSzmyBDEEhqnqS0WzOOaN5Ii80CmxPZDT1hzL8EDFwRsdBDaidAF5DlGcHHeU5dz33p7u/3AleZ
71PnYQTQpsgZFxc24XtsUQG6TBkw/eRQCeuuBxFay2TkmCShBnZqrlTDi2ijYYi34ypzZErSW6hn
j0UkWee1/8k72dJDDtcxWJHDOQchPqRqSow/gvt5Yh1cV6OjnbRTgHv2zXjMoomtYTmNN6Nl8dJ+
99DbPmblsKV7OJ9D1hV4H2p/6PsDTv5b4L4OkRrC+n7JsnO2GA0T7/AND5h14V43CJIZ/O1cMook
EYgbH90cwVCjnlM0avp93xYlHF9xFDMUT6AXKEY/p4NODv+xsKo8kD0au4CAo+Rn7UBgpz52K9by
+xsiL2fomHHrZ1jfvPk00D6HkBNx6gmtXLF+3Ybq8E1EDS7Qhe+iAlXS6ThMiDES/LNdggHRukWs
jjt3R6aOERUSGmd2SOdWPv7/F7aFMiupzYvdNjUb8iKoMnWzk0BDevP5ElGdnUlbb8JzPOrCCcvp
YCl6qDm9bq31PlNTr6lkTmxjuEUSS5oNtAHr5lfLWzkqWkqyhI6tCxYc8OIWC4HtgcqTKT0qoVnM
cn+y3PvZEd3xxnjrZKz6Zqvbb3HZT5qw0CBymx5MiFUPyHFlv61EJWfpRApJGNLkk1fdJMiE/t52
NKIzp8WUmScB3//gXdWDR1fcAd6kXgOGmnt8DGNkzWk2HTN1NCQC1PUmNdLmHSeFOaBVJPhd2hqY
+Cgl/5LNStiKWpjkV3/rvkqrXvdTwuem07o3RqsaDGoGsSGHvBpMggnR13+yLatvqIC44sFNI06w
hLuwntX0o/wS2MJn7jejDnpnqP9TgsOuZvF2zTTY2CWx1iFWD9fAOkzvjs49lFM8W3INxkYAPH6b
p+HdG0j8I+JE0dz7hRbNmoPkj79GBYWpUk06Q9lYsspl7+EgKDnYqrrNCUdr8DXweIPKbP2Dz1or
rNXTab3oKJhyehWsrlVJ1aa1KLpDu8AXztVVY/ZIpdoazMCq+8RqbJq2Ajas/Xpbz9UCC2FIIUf/
daKT3xZE5f+ox69Squq71GKW53tI5bzkTK2pQK17hXQzW1B1B57mQjNsNPVNtrxkQxc5qFZ5KBEs
WAxbeEsJGF7ff7SqfDIg4R2C/MiL7WpcW2I1VJJ4a4/C0xAs2/AD+LO5AmAjbmUCADpxzUMvSGzo
7KUF++EkGe3NJOFqEk+qnMt1OwTHqWSke7pZmd+Q+l0PCzgoiqu4/S0lFu9fca/We38fK8u91GMI
42HNMBxsy6613L1hiAJUrjx1mghMqbjjObcLbki8G7aGn38YNpsbcjSSIeBaFKnmQMiPXwXL/YCc
JWQtNkz/BkHlC9t1Yb2Qtfp8Y25Y2EFTS5FaaQ1oJBf4KdIuIuyYpsf7k5urjSHo9seD/548MAxE
314cRMTVR8RyHQMcIzLKqiUxhkylycJMApk7Mocj3fqtNJEcdIKGFatfByLvbBB8t2ljkjX1mc9F
3A5ITOr5XNEnnEbMweV81aHlUixiAWRD90FFi2GXDLjp9Ne+hQaVSGznSZ2QwipEuAAhOOmn5wSe
8zfcotOXYteDnXux6PVhTr5yDc/0/pq206dBQGFPyx4nmyagGAzvMesuPNKtlrHcV3zwEPrNsVWM
Uf+qytZA7JIEMPBHRe96oLVrtisIL4mtCxCsryZtXqMg8+QZenrA7aKbOOynAhL/akrpDsCBbmru
DQhSlTFcYOfuN7prXeluX/KJQN+ThUOR4T8vv4nK5cmhCuxePYcQn1W0ZTspJZc0Skb9sxUo4eu1
Fx/XPuorCBmconFqs60vNcNNTcF/j+4MdXQx0IXxkik3VGesDYLYAJLabD1LPayr8tq5KrMp95Gp
aNXaNhR4PQ12nysyC/9zaXSZoYBemvkKd9f52HYeO0qP6tj8HuTC5vvPc74aWGKkv8EdbOHDKvub
jGTnzyTWk04CmxoEj2RLNOuI8/lxsLqbyItkY2XnPy9BUsB06jNXhelkjthgu07Bu44Po9QmLUqY
vObypaOiqWXjCBiiAPu3jBVNmIC97xVwMr2LsNM26qH/162fbD7ucfp4bZrRKJC9pRi9J8W8Dslr
YKFYCvuJVqkMPoEoveKuSKuAXPvdfNfE/W8Oz1EcYjnhYxbtFKVLSJROJJG4aG1rAlxNmKsCyEn3
lv2UEX38WvH73npKAbZNvDlD1zU2u2krcjI+o2z1gNRqJMvrDu76FkZbsJjXQJUH2J/gAAXVtkkz
3E9aVPmzHPjoumaAAVmFX05Ht6qIkkCK7Ke73T5gsLsm0OfXXs8wgPhkLof1kLxAZuCoBPBM8RSk
acpPu4l211a9qf9S7WjlCXX8MgvjXWxlxcDDTOQ6Ll55b3JXGuF8c7VA3xfn4o4MVO9BluEuyj8R
9Lz1UvxUszdG4pHBjDNPaOeM4bjdkkVdPTxSVuLqvGmAClrrWzSRdG1b4VyT+JrjGQV2+OizhHVn
BGJ4dXk3mqjmviUM1dS02rVEklZw1dEH887xi7wLbL3FIaJbkzQyY5Z0I9A0wHosL9mU50Oyihfa
4knoboCFr6N9TbpEhSxNPM8gScSjIjweLsVexXsPeisKWP2q/RaYQ32C4vMfT08KzwonGFqgzigs
8fYUNFXoWOvDpv+JqE9STV32cMomzw10d9VFamIocFLrQoNdSyu3qBFz9Yy4Yt/n9zDqYZp2pu9m
LhqW1YPL8sIU9btcpfF30rU+cePRwHMDGA+XNRr6OOEkpR1pcURVEFPb6OszaTb8/ac4znUchFQw
LGVFwLiIspTnThN3nSW6h+F5Ykax3X4YkpDrgMS7/KIfH4Tmv1wJlVACrzCR/s2CVZsYCvcyl59W
/Qcx18K2s5JEw2/7SDl6c9MYBJAbNns2EaCHhT/hY5zAKSQAtYk/4Os/kZKXc4iQJvdGMxXT0reX
161ycpvy7hszJazecen4sXzUpJMD2RkKZYUYPBUUN0x+gXLiyD1CNkD1Pf0PhKTnCqEyeLpqvG+U
TrgBA3e2qf2Re+yvuKRzUOa0X0AVJ1aOhNjury8Lv/NJ2v68DnYfyoHhSf9b0YP03cn1Y3C4yc8v
TUE7TTvL/DA/DWl314t80O4nRkqP5kEdQc8v0oJw055SQ+GgvLGGy0O3kgomtxZoaMPLob8SQOHE
9G2tzf5/ngaFWWYlI9D/TOqgb+2v1N4dc+wo5Moay3/7Q4t60+kHZt5Rm2VFzGAovWk46uj+PWyX
87PGvQnEcwlyORO4k6RR/UzyfyN4zsXL79nyamJ4Xa9tq1jTmc5VaAoDYQJgL+Knoq1LYZRQ6tH4
Yasm6l+ZtDai+3m0rHtoLP3ly2ml1A7JqO1vB6iNYb61yFQsY4ccCFSj0Q7dfB1p8pURxfS3rTKy
iF1L/LMttCYJpKyz5posuHxwR7rt7CfpHIKjrvVUQFqVN757OFLg+hIKQls116UmQR2angD+Ktu7
eSMK4YwwCfuHmysBDKX2inXme2GWdThRNsGnx9vf6peUUNWrmiKIkl8YaE0Y8d8qOhjcO2hB0rRS
i8y6uvO5L2MDP2H1StFPommrOQjetFRiQgWtDVvg2QNea021un+FrOvmdGU9yczu7MI8bpdMc86x
ct1lCAJkuttfC5INW3Y39EQjfHHng0Z5z4gRm8iqLFVW7hOqs7wotr0S5y/uewhRkPZ+980LrvJm
J+h7Gl/78X5g2WhiVjZIHX/4oDpbn2uv+rXp5luO5K4g4OMKQ8HrbPLZp9xd97f6qximDh60y3Ng
Utpi9T3iFuZkB9KeRdArtTh2EFxGerFr9eA4am1eiJNlCmx53Yxg8n6UnZ82+Xvpf3EEmgVZuEDN
s+Ap9ZPdo9lLV56YR3C+VLL/c2iB8IPt0jegulvyDF21k5zvONy45kFRjvL9/YuCVDVGLo5XzStM
KRDJA4zDwRLIs45tna1Xj6E5dJ190tSMM7HJlsjNsFK28FPLW5+tcdaxpEEE2aKygWMf8NP7ze3Z
6oYDNguSQxIDAy1pzXRTk6TlW2FDL0hE0M3XLbpYaaS3KgNYEnGriP5cZilLxr8SSGtaCKqPehYr
QQaiqW2xOSvTUaVYc8n13Oi105w2pA3aDv9cXqbjBncbm3ylzDw8IRwcSrxsadu8T2PGfO9lhsuN
6VxuiTTPc/mex76aa4jZdO+oRUAtlrUe0fonXFzDgwaewgCJwGqk+vP1pC7daV7ddze7PERhXbF0
sYDAMxlbZH+sKafmPwXbiUvUHd5VqwTZg6tTNUPg79lW2GiCEsM+g8zhWbgNxXNbObLreUlAgq8B
8C8wUapnRQu6ef/O3SBbaOmhe1CffyQaYNbRIGkCNONAVItqWRGN0mMUljIQku5l1YKj/W4S37ZE
C3C7tkSCTgsp4bmfH3XQKD+yGdF+1nuBrglXinRa4nr/A7hEszwgxHgh+Zu+3TM7rAkyIbh3n9PP
Edd4KCx2JEl76Cf2M/PIlnaKJNiH+oFIkk6w+L7AfBo5+IGxA1XM1q4nuaCi2UKjkpXQ6lRXedz7
J4S8E1r8H95dqH7/VUZF18KqD3el0xpHr4pZ9SvNcnwQq87+/Pr2Xk0EnJVt4vEoB/8JNCeqPuZS
moa2s71lwkNk/jjmw3wJXRf8512UddTw9FCQn8s2+a/BDODB4iRcXfTgbC+lYX0BwuKUH1X8HfSC
SeCkrC60h79XXSRYObCQguQI/6IgPs7rNsITaAvpfqlP1RMbv6AooCAWsMnKaK5oDLqN8iI5MKvQ
VZ7QM+ztzGs8C8pAbKfb/dUSwXKAK2hFkOsX0gBnYHwY2GpfOuhp1iwKBm7m3Oyeluw/JDUS64Tt
LTo7mqRVfU4D+nT2w1M+RpQ6JogxsrtoZ+YrywE1hDkkj7b1Fdh/g2uvDXgrA2oZxw9bUjIRzHzo
Sm82gODu6WegX4dmWnAamAk1yfj5GaXovVwJ7cJerRWksPs3dVaAx1jJ/x55rjmqNf6be3oq1yXl
iDeuFnhgSytd7XoXQshYsax73JaVaqyAXAYSxvpNSU/mItDFbfqLbIqKu1aikUsGszS+856tFcT5
PfDGMATwGeUlIxg4qxx5/35QGe/zyo6W3SmtPSAe54CPK/r8qv5Mp9HHcxPuSlqAqhk3EA3jglUO
VXDWBEsEjIREkE0Jwn1v6R3Bc0VgM++SEg2Y+Y7ht7DE4ezuPNnmKd8yIbb7noC9hGfKHbhRlvu/
MNMVOjEud6X3MZN6PCwOT1FT9nU5iCXlvvZoUG4OnrNmCi3hWaiDaMafWCjNDso9G7B+bjxONIit
iH8cJP/2YmgDRCfm2IJChyLaqyxo4PsSXMl98sdJYQCX5CDzoBKhVpLoX/uyXdXrbXb1PjTKaVso
pyi33ixc+znAbLH+i+XJ48Brno9nsjkzGFb/74wIQ3G1jd1dMht+x3OJij41gWDulk2ia819DwPd
Rwuh6v29w3Lr3M//WA7pbG2T8zwLPU1hEVCMR5qNOiusiV6Fo6NHwy9yZjNZ47qBbcAWHajK58Fe
CnvjjCPPoTxCUjeouV84we75dXt52hYCwcBfyGLmyo4jl67HfVVf2pLCKm3WIdDbF5pghKvqaH4H
TodYOXGjgucVbXjY9BZNJC3fdp1Cj5bKaDyU3OLeOeOtKIxheBrKG8zst4jpOl+ARiOFmNSgYSbD
c+uQSnr8qTMPtc6HfVAQ8vzPmTcFctZNMZ4pWUnjq7viMNiXifTGnWi09cOWmmyVtdDhD/PkfSx8
FoTNPD/mVcYcuEiWn4whGIybJUy7CGIqNRqVhhUvhHMyNLz4rQYsjgngU89b/g0mF0rngNgoaZnD
R80bBde7mPxVjjy/2+BmD+gNozjezq0A/xR0dQhXXsS8GZyMLXVc6Ia6dPtjcxflnNm2dVioeQ3T
bhPD6a4rfWqAR7hawQaHkrihdGeokw6Dof2Lqrhmx+RgIGdn2LShHFLaEzlxCdoEh478rHnivIXA
+y5Vo8h7GO1BmtH7p366MON4+sJNRPlOvWiNF/Q9j8b0aUYtWQrtAqGvdmfsxmdAxWrgd84FW2cM
GFUaOEQfwb2J47el90rFVDSv581kMme9ROAL7G1IuPIPsTPtQF+eTOyHnj3p6BGUCLK42eyV1U3V
SUoULi/pkxXqmXYf7j10NmmXwRrvpdNgcQdolcObLy2tiVZEq/okvSLuhx8tJD/1KMGhzULrxtOr
XdMqki2IDBkAMysaW0Po/Tcyw1XV2P1aG1lPhF6m8d5BPCnG7adl3L4mI7xyoLFxslzLn3FhLPpS
WpJ+1Zp2sa1Ne7eVW4sZAKmGQYsT9qvFykynUVk13O3TIb/hyBw9qsEhNXW0Tcgg4bozcGWGMyPM
fkmotSF2buUUiRP2ytsycD6bUitGw0Alurmtwuzuqyl87XBuLfV86JWNSGp+lenm8u1VBKiJtkhj
U01HMBA8Z2ReKBtKGUJkXlkG+2wdbIXK3JvqBGjMX5pL2VtdzTBaLjlfC6muxE+f0ZU8A+fr/kpV
nNmLKFzBQo3jX0oJs8XCixsmlRQP+pS+aggB5HkpLaxfypy3rWc5z312254lDr+vtQgPeQ+22NeJ
cBP8OuCHqmWmE8nxLdsiUV1qVKniZ/QwVGt+Tcuhxjx4YX/pjXfCqdllwdvRvL6j86TIeUIgSBCz
bFsVMhK4vaX6qMIxlQghpVEphliv/IVFfr3oQka6HQ+p96+/VXkztsRSgzoNSYtjCySLIkpx8z1F
scSknLvMhJ31KeXzR1NiD70Gy3Op/PI7ZlPFxWAQlUKFMGcP65BixFfaHcgzzYWwqjuuZIK3htLd
xxISLmSqguWYq8SggZfAFa3MZIojvGfjOvildBPHXsxbaznRRR/jiquwO8ob59PmaHAZd9KWm2Sz
pg5jIL6AkEuKRv9wOXqgzx9klAtNg43oRchGyfFYduIMVHQ5+rnD3vDEzZtDpOeK9nQksdmJflur
xlbFsA8ywEoh6TgpI5cDTp6fm55+DSD3juqiekAk7oFQQsOB/aKHynORS8Y9BmhJXnPFM9jQHTQV
mIOnnkh9Bi4q/73PZMYELBWAKL48cUxkkeuNswApEhPUkTuJhNNNct8bbwJc6usMBGXJsuqnFYM7
hMtvkE28r2ja5WqAe5tzjBbgugIE91FadvWCRoCobYz/ilUHcwO8tAgsLOFLD1PMDHGOzDN8Q/wU
YADWX6zh808wYC/UEbqRkoQbljv2uQEDy2vz2x4YfO8x95sE759uxddrQabQ0qLURew00ODAbFyu
+DxPgktWDG8s609zwWDOYh5uTrt8Zu1+7bt7yz3N+XpDeGFQsPJsNpMaVpkZBDU2He4sKHty45Me
hGp4Baelk2XwEiEF+i7LQg5n+kh8i/KPehFuLuDvtQPOp3Wgm9F6FpVwEn6ov0dsQBlPtOOrpEva
8bTSRa03K0WHjuFWj2acDguixkxKe2ynsOneKz3lbRWO20yZyXqY5KtGlBJjASvcbaLyBVT2A6hO
YEXZjY3C6o6eDs+pzyAE/mSTJ51df5dV9jL/sPn3O5mIeEtw8mTgyoyvfYzCKtR88ob63IDpMk1n
sg2P/Mo0KwDDQSMzVClU6ug86wxn2fQAYOVxgs7nitxIEIikstsMzctL2x+YP66Au+ZHOb5+NJGd
XoiHmf9bEX3f+f/h6Me5hEFTrXJiAJCjFXTI4Y+LATpXpreX3AIziZOJtNoTjCHkPUHN+Zf+jjt3
fUcRf0TsGTiggNdZSTOJaQ6oBlYSklOY2q+HhrmqnM+cCRPDptkHpekFEaC4PivSiZPqX/La3rbc
7Rq3CNCWeTlNuNslrf71PVPmWhNGKL6ab/4EQM44mSkbcxejyeo2H+jccHwfurymOgK6r6i1Y0O5
83whsDx5jigE0iqU/I64GzUqS3qUpxtftkRlBNfyHE1RhR6khsTCyiVfuov6D6CN8f2BH3LY2jnQ
Xuku4c1U87GYFGa1BmDDyFHGKoFftetrB4xFtWNfl9zF9YIRUcGHZ3uNck4Hwq1whU3NhLZO4cV1
2TfBk6WCyhmP5hnfAUdOrizYUpqKBLc4AoAW2f1tSlrrEY9HRzaYQayr7AM9IckgXhJR9QTOPeev
EpVn/bfORvrdqgV6TBMDHxBfoz8Ewf22+SqxDynwWK3nN6YCCHVoky2WPXr9rY5k3jFOB5NbG47K
cpWFKC0wtF82CV09LrGQbBCh4edlTZKBrB1o5ZFUQRv2LweHwJLwuryNcyEB8J+ImtNiiGqQK66L
FPbIn65Aa5S2D9fMKWaXs+/PFDcfkIBYAc+aWXguGoqDb4NDYEajx8B1g2hQ4faIYQTw5UI4uvp2
HczXOe7UzS21uU8DLpOPbgq7afNrm3JQhFdmUVyMdUPf7VGO0rUazUWtbLR8oyopAeIY10FByAGH
BAIKSXwzCaVqQnJVECBqQQJcWAd8WAekXwBompB9sb5CwqyJoyRBzS5hMsbLeLIwcPMyKU8rXTFg
aXVygPyHWf1TJXPjOT4HFrEQXgWoFHXbKGOSiw3xqiTWy/XCFkzQ51cgD/R7EKyFIC3Y0FcDJRB8
wyS6bq9XBq/6G4oSV8DcymB99h+5DQwX8aG3eJY7dAnDNxdv0NRD5pp+VBNv2+E5LrIqGoKklOCQ
0Gqn31n4cyu8MF7EfT/geH0S6fX9Yv8I6sSWukmWIf+oSfBe8LWJINW50fnTm7odKv+4YWrGuAWP
M979T095tsaT6JdM0DRx4dxkCa0LMpSVKNO7854PK80myU8c6YbR6vM3wXl5GSJd+1euRWR4WlVS
Nq8sgxPp45l+aCPwjqoDXGIRbuTTZUPKlO7EeZRZwuXhOvCtL/8j9GQhpSB7gDkn8mwuN71O1uyo
OmAwMEyCTjjFlrD21W7MoMTU6WA6yfhKmxgrRrjnx8AbQDIVEIfTrjpaL79W2jRAOvBbStHQ4OUo
FcQd0XcouszREIRMKYdfbV6dEGMAwJu52yLWLJmpdKEU3cOr8CnygUfAov27/38nRQOCyXRTUnkV
GbmRPRBGvHFnm4jGvtd4924ZtrUgIMqX1IWqmZHATIlV2EKoIZytiQzIZsOBEVIxQZsNNmr7In0+
e1tdBR/HVpXhOcEulUiTTb1HmdBXOAauMDyU7DPqemtRwTG27DDDqbvVzrJf/PBQPt1A5dsEPM42
oDD4tt9HNeCKa/zx5GxvE8tlIO1g3oHR9mvyyMwMVAdBIOtXj5QPW6C2a+/5wh7PHqAc8lFSK+ib
MlpFJjjUDvj+5N2ZqrTho7fwkZUUv2uYpd5Tf/h7p8++dbOqfpy0QyFdK8MRVw9WeX8NesksQw8p
kxe0KjjR+RC4U2ZRS/vhlh44Rds2ELbCzCueKO2kFQHFsmgDbui7mZAoOkbCyYwdqtM60ydvx33h
aYCgnjNmbltXV3B/Rv30QxL0kAv+DtsKPU1jf1iVossP14JTY/o4aymEV3nEQm3MDcxudxF5rXpA
iCrk/JN12t4iTiYiUCdVQ9jBaRKB5ff58UsN6OEbkUOWg7GmhSxpqZEn1NaYr2ZHzBaEh280obQx
35ySr+xvVWfFkkZE9gYxGT1rpzQYZkSRAMuUnx/8MTfbUTUJ8nzOmPiuUuggiiRlwDA+zg/GBGNs
QjaP1aep2Rt5655aKA1uGZQJDrWY2wN736uCqcINbUvTUXaubLl7IwMyahBOh/ZkNGZcy6QwW/Yt
BRLiVK1YZ6bGJCTr+z3P2fkGWT5IV0ZRLP8TE9qbzv8L0PigKEbwIAp6a8DmiOQHQdwDZgKXFpcw
yorgvtHSa936yVatVVWyC0JNrtFJBUIdtLUV197WIf8gKHIko6B+yv7RbNuyNhPeq+UvZ+0xWEYc
ln2Rqsj1vVa0Tg89mtnC8ajESsAMubkeGm/1tLTooDQI6stIOXcRiKdXBCf8/WTtgl6db29aTgIa
AgVR5XOZWmyM0ITXlallU4kSqqob0AINnDhVS+ODIsORUHHsKTSZV5wHTPMoGjITWnS7kww9YckJ
gKZExco8twmY2XmykqQ4UeLiwcOKXMmtHC6gNH4yn3WI8F73R+e3UHb5/3+biiQlrIYK7J6yNpfp
AXFHmnMjHjdj1FWRfcKrWXCTNOGiVyjN8/xmU0LHUP5ugUu9BJxnLxRGTbkDLeYe1Jmzc8pZ+9nj
FQqcwrpefq9PBpIH/gkq9jQyUIuIKJxRqxvASenv+JMhsjhQ5mkX7cg7id2yQOEg5+vUkSOH+e2N
BrBm5dkG+8ioRT4Zblu8/sGss2EJGKCPdHzW4tY162IMyqgdmBwWBurwoNztQTK5+NlLULq/yyLJ
YQotQdGhhkmTA9YflBx8ad161ufuMZ/0Y4LX57ZcG6urItb6cP40/cGynJNGKu6/xg1Ibv6QJDqO
ZiIuYg3gUEzb1RvbxpdEII2PosEPVUu9O/XEJGAL5DbgcG0wbaIEqwr+fYCett46AHbPkWBvmmFC
qoNd+hHOqV56jWnZRcMVaOPR3wwzPEi3bs/ZmzdveqrtuL5uUk5+cpmy4R3ZdxxQSURrD8g/5k8i
f4teDNuGOJN/M0JBn+GTXdxcPkZiGcb3ewe7Ja9zbLPVGLttabLoRMi2rA9NnT06SdBPmAbDXoK9
THcFfBs6r2dzy4o9iIFtqMmuLabjtP3LTZNoChukbkVeitcQEB/x41YhNlhdGEAmx3k9V//DHIM2
dx+x4mQvvdSRfYfnVYRiS9g8Lm3HN2nnTZ+4uVh9QtHUphnxiCiVtzuPWpRNjCC1iBk8u0OD4kRa
HngjZRICFmiCzM5w7HPxwRk/WCa0rTAd22rldIWiVnFSLE8ljG6MYLYzyaNc9o8zyRDgwSjrQZWf
3LHbFnVwV0wfHns+WlQJmvE0g+gF2VW1uC46ZBYYxfNMyXnOKLKat5Rxps2CWfZpCWkK3I/zRAqo
baBnTzm7e5OI9/gc3ay4yB2Fw8jgHcSCCkdcISi6LvLy0jteuGL6zdY4zIesKVkpofOHKiCQfepG
IxqsKlk7jCXlh6Y0PPhLh8z/+4hTjgrdluh3a2/ZfzzA++BpZhj7m6Qw7Ef2Nq4QXR1J8uEi0y3f
stQt3uRiIW3w0mKDDozElMOtRth+b1RHJ13mRUCacbWJomhrnLhnD7jEPkVvkYj+KCQFjBe81bQx
z2onArsLt/nS5otc3lRqfQLGSIkg0TvfVmQRs9EPchYODZgEzCYgCcXSPXjdEuWmwzhb/0MUt6aR
wz8TscZwjP9rTE2T+TWaePupkDOP0AMtVx59TGCDcrwX6heZQe954znRVe8UP1BVGDf0hQhYiD41
w8XWfX5TUCiHlLBMzBmqf49vap5Mawk2snFIZqaLX4Ox8hn4/Oe3wnhLEuovLN/sOFZLHEFcfwsm
yD3SpA2cCLViXxazOKnooQWAu+q9wMC6OefPclBd1IbPTETsKkhE4e9m+wOYMPqb3pYZlAYvEuBa
XeA6sDqs79U0+g5jlWTOjtyRkuVWBLvzi2BQoK2zoY9Wg04u/MthcPryvbO+cq1fnXp8MM8R7OCo
RCoAYq8+k/zCynH90836nEkp7Rz3+5Ul1Haar6EzWHsy4P0jwQM8+Vn/2RDrdL5N26XlvXJwOHzk
LX7Cf0p+fa7PyIjal/AVifb7uokZ0iLz2iTsATKY9OkA9nFE+kBLZsxTuSWxQVDGMODUVpBmFF12
i5jY3JaFGA2FhJZgjDdL9jANPo2XSQxpq7CIcSMZblYBWxuvLScrAQ6WUfbAo7We51U0kfXGyo/z
5c3XqnlMiQ4wAO6lFrLHFV95wpmfD+Ma0a79lLSwilfwtiwT2W8zxdzg596Vxk0ujDOBaxGyiPxF
iXw7NRX3rF3WA42JkXYETxyJYiOgHWDnLDo+aKzMe7LR9OY4TtZG4mJJijQ4kZ6oSFcHKN1ipYjf
SwohFFYHTvxkh/XY5SyH+XDI1NrfSAugZTsP/s9FpRVLKRHgnrCcns4QGvgQ2b22DqTqenzGD/2I
zgCAlqaOXgUQXVNnGscoaa5grV8dTHACiABZm9zOtEccoqzTEQgheak18IzeuaNc4TtFvYJkYks/
Up+X+ufK/qaG9gzMgQizxmBKj/2NrbnyG3zTbsgbAgQw0VVDQgwY8XLtVD6BdkyoFUP6mGIzMbAA
z46MBmYUA4oWApBIqXZqCF8uYE8tQqRTmt5yS84O4k0363XY845VUtsFZf/dbqf9OoznIRI8i6PC
uUY4N54OFn45kHTsqTjDXQYshiZ/0pdumDs3mV6k+2u0zo1aZKq+TcGga5SrKenU5ZQuqC5JjXMj
gbHtKcTgOp+z78wCZX/5z86x9sD5ZCUbgaQftN+i+hN24UPg1fLJxACJU2AQfwCl9aqNtCdUgWCZ
FWOvsekn4X0V/jysCnrmoys0Uv6TFhx411XyBL61czogMVYS9x3NQVwpp9oeeaESJMOMnWQjp7HX
ifK5Ay9t4/RGwYHZ2ZR+H6Xmw5Es0aHQJSPxlva38N22SvvssswlOrTi3NAKLE3T5QpiwJyNRIE8
PtVMigPu7At94RcSMx4kXQbJgofJD4p3FHuG37cXHu6SSaa/yoAranx+8xuNuWrCnJDF0jxaUMjz
WIuKBNEZcvsiPP5D/FyVsA15YobtobcMjxztQLFMMQnrcmvhGNltE0Cn9RebKtWF0SoHns9sqTt0
veao5gaPRYUmLFyBsKEYpiDNzdotegYlbr3ndVV7Q0124QLB36j+soezocCbTAd0XtQhqFleXQXf
PJTxArPP1faJb3V81tzUcG3XOg1s5Ne7zU3VPRq8e921CSeC4tX38L2LFN186e3zmMmMJFMWkX66
o/e+DKP9p2eJa6lJ5LDvquRjgPqqAws4RyAIi4MXakcwVicTZ0gkLOeOG+E2FPkk6vJHFHXiqlUd
ePUM9HhuXO6nE7dja1eDqy7sfshPtjTWZGfadskxe0ncMLJt7/AvFTqBEuxugNef7j/lAx6OUHvi
eCY+BgOS6YbjVMgnAesjvXsAQUEwmDw+YVuswhv1/TncECuVOD10THqMa98SbYx267bzhNvR6toa
i5+AJ5WpksiiRYV1rvA/VHydNUQsA3UGHseYc1w9ITWU1GaJ/Idv6PraGRPSut4SiB/8R6fbQQXO
5IINmNX3BdkJXqek37ZsEG7hEh2FDU6BgrFqqlRr8KmW9CJTb1oAK9CCQySLDxWgtJfja7mjYTxy
cVMFVNvSsOMqp1SZoKd9ivDw4ksGT5zPR+8twI9WPn4LFAkgAay+i9HUsT94rODtgp0+UWrKdwiO
nGiFoBpJFJ4esKQHzExikA/Pc4uurPArNzZEnjbbDTmWClxykKh2ve5owaL2BrqlZN2SVJDjMbKX
2t7FO3lfH1mfvSQbUGRRsEDt+EcoXudokaGWNK0J9nshut9QbDNYC23Ijuy8+VsqW0Dyqpzq7/Bp
LA/J4ICacmnkX13EGnNcS8hXjY2hNoAhQ7GqzbBtfGM5hqZD7RjuK5WrM3HEkVFbS9SYxEisvexe
6ubNRssqEAJ+Ox14ggnQL7crTq1a2j2/x5vsXhyZAZkjj8mpPFgXsRkyxCUJjBSKxuAo3m3KUECR
rdlnsb3tFEi/FD1sQ0Yrh04ZKEHkhRt0cMCVhmzSy4g/Nuj1Q/U7i2gPVRllCCRyqSQkrLeYPSAn
9WH6/9l1ryxPAtHjqqKDug0wogsH8593fdgU0WW554WgX7dPLrl2Ko39GIpXStZxEb+Npug6Qczq
v4fMeBMPTuGcxCZSw/0aeFnOGAmAZQEA5N/PIWltQvUV8Bsrun3Atc3TmLEBFQgWz0SqZ41zT2tC
PdgvTzNdc59es39pbp7e0mC6q4gTE4A0kmqQauqbFA151/HyEl0KOoTMxVxz980W4I6Qr2Lh9Xw+
/LKkDVSgn7yAqEsPDDoVEU86LHCqtOE25qmYJg4v9g5F10m3RHlcG3OlIAyKOvQ3XN11bGmKoHlq
7BQdpiDykwvYP4qvXLuOnEeDkLjo4u1ck+hpp0lA537BhiWO/KY2+ETkRRAGaz/ZizR3hSeFJ9MB
bLeUtXsJPOBf1s1UG9enb6ii8WJ0WG91LYvFcao6nwk0MltegddGahkpWuReK63cCd3q4hDlmjb1
aChfCh/X21mtVGjad/KVwxLpKRUfrZD0CC/nz8rU9uyoyyZd5LQPvJMc4+fIhGeuzWs5UUEVuHfg
QgYFSynUbI9lVHtH9hVH1+EzufvD9bMaER3cwr75yvtQLsR20ZjA0YdjEIEIW/v7kcwV1F+xhKlg
ecoqt9p/c5uWgqjXNZ+yNUXVByciTa6CrEtZ9j6oaNp8BVxarLXt6PD5H9Hl/2EGlF1gxqoGqBrl
7MNXvAQtdoI840rhoXUH/k3UJqUemxoW4yROI0uh7nU5HFVoJPewxs+yI5xSa3eDnc0OUhQjyt0p
rwPuTLxDwdhdEpLBKMjCUEG9qJff81i9FphUBl2BMe0kQSTmRKX3GlHGQxhI716fPrEPsv3uelhr
K5PuMvqOBl+dTEuFjONF6XelyMBakD9VGwBsdsLF2oKQ83lfrCFQAxQxVSO6uTOdUlwGdL4Y6zct
rkFUeg+EeOq7dD3y/b5e0JQGgG2pO3rnDg03ujYN93yVGhqjq4UCj4qtycMmi3vfAtLKBfRGlCO4
ivlhBx9SeMyXYMooPVTFCJoomaZ5yyg9qpHJceFxT8pMMfh5JkKFYmoBcI4LJbkRdavxIx1gFFVp
1nHYpzL4R8LpAF2iTXR+oNqpjIA0LDTTXhUa8wkgdy0jXdnMyoVjbotAN7/jgx9vIfmjc+7JftQQ
EdeOF2BD8U8n5PKaP2l2bwi1tipSMupFb7lOZnazJBwC6V1lxNp7KTknWus88dL5fyQ6O5Z+5uG9
LyCKeaPTPaSs7gXpY0Y/yI5YL8uJXW9v2hL9Mea6+8no30e1MPEHmqCuQOCQS+g5ou8Cps1rJUoq
CMpkdOkb9UTTzBaytsAvizQ+dSFmJbj1Wlu9IkZVNalKhAt/jSwIDJo66YtrZ/yRPa8GQFj22AmR
U7F/3DyFjU1oZYI0AqTPnJLhdyoqUat44kuoge5Au9GIDHSk1AhhqnDC5iQbFYgOWJ5huCH1eQh+
rtuECX9+0Xw0qYa21tooVlPvFzjOXG7/6UfLHicBk8X3C5uaITqgNxQormKGjx0+SYHZO8xSBkaW
rEq9pcYmEIToEvwBneC2ESowE6AucETINA5tdJzsCEZXK5WzfxG7UBY1TV5LWcquN/ktUW9+SlR8
MSBcLNnbDGwKa4bLGnyTzMSWTXRFxph3cYBc3c0NY3XDE4uVdhMWju7znylU5w7k+lAYR76Oud35
rjAMD9t54BFAasA5pt/CrbBbo012TOVbGL+1n+wBhIZdIi1XqF+Po2n4PS/ZltDMArrxNgpEFE6O
zib+HTX+278b6dKqclqdw17ygsbRd/VVAL6j/vyr6DKlyP9Aoq5i5I040RWi95AaSDTv3ixjepwK
fPeCcoxffR9dNz/lZeh7fzIZheBi8vZTH29RmjhUW2g20Wnlkk5Hpa4jRG1Opvc8bbd9dZZ78byp
q6d0nj8A30Ynt3+v7cb2E6ionyYuA++h8vPy8e4k9mtW3lu4oiB1oWjh+m8s05yragSbfLMvywfU
sMtxV5n5DdERbGOLpgiHZJ0+vMNB928jsc0eIsVx1qj2AhnmOuEgHY/j7GNEvluyg6V4UeTusQTw
yuQkjRMNBAxooDQvy86Ny6XMeRJ9zwFWnsz1y04EAHGsMzS05yjrfcNhTVdL1bXWdgR+S2VXc6A6
spPiR0BmwWNmQh4jm0rMQk7Q/vl5fi5/3urjECHGdohzbAsKSrC9QhRvTAQZUUGH8Z00/rp8je+o
Q64NXDL5LMJy5vCyqU2BVIR1nvueBs3wVyR+uojoRusAJiUFRiQd1V+D559CqoSNVpKCGkJfri6r
LRVknzkRuk8Xc5FqF9qZuDgzD6NIojvI/WMWeccoA7LqnI/Q7bkDzajr7GaWirtVF2GMC5xH9amC
mwd/wJcbrV2fmJbpOltnz0jOoxq28rU60sPHY3eVWp4uLlpBgx+MWoxPFrVAkPKowCBrGCv/9Cy2
pOV/oxhUoxyHBuHVEoiggIjYGb6EioTpYAT5z0fwF9FzMIZ4ix8FwK8XQCoe6SfUnlzQG+v+oP6G
s0QyEGTtjoifGPu4UyZBG+lqa1XZ0H2tYHBcno8f+X/MrtcQZb/28500Pmpd/YHVAq3eU75xyM/V
TM3+fMxD94CYpudG+FhIdp2iro8NOm3ulsfhXCCiO/shRPQeC2pcrcZhvikxCCdb8PfOpCa//UU+
9gB/l0HW1kgp8hZBPlrxmqS5RHfM2UimCyPEJWwHqTWKEfZ7kch/bQePZqe8xwhkLXp5Watds3I3
C6WkOndQUbO4Utz/1fm2EHxFuUMNusqw9CV6Q3ORLy2sSaBf4oXHC09hCqHrkKhUwk5I7eVW2K1O
D83Bp+D4LCXPwIpdzGqccVeKK0kQi5pUEMJlyrVI3P59+qjF2LohgC78b1Y/urBCUSTKZgvUxoJF
bvHHcSAJtUOJLMtWvoMkQOA9EKkQm27cWrs5HU4PbQt+jcs+pH7ldF5JfCjWiTllEr3CsCWNbXpe
LU5W0BA4pxMCG7nCkBI5VpCT68TQqkP5U+IVeqhban1NkEB4c/tkE726rPQzN/aLBSC6E1ppKEms
/lsaor26vqLuhBdLdb/w1k9ietyFR9jT0epj1rYrrhlRBTsCczQKekFFeAlbPExSxipcyTlutsLO
z7PJvmUd3Q4nI8IhqMxfF5Qi1wKY1VJ83lPBSp5ZW2J+yj8q9FOwRCsGOc/oUaQYuPVoU63VKOrL
k5Id93T9CKHYl7V2pVK+gWQBvFdm+VeLQsIYVmceHUYWUN8N6TQLitgjgIUA8+JBrRX4WuHNebkr
ni0MoNgLPhq7nkjmt6e3Mrnu0otLNdQsISXofbIPC/MWxuD6IYVpX/OTvsotMjjT9yAvPk32Tibl
AwN7Y+fv+FazsC1eHvLLc3joYyhUu3VwNot5cyHbqaZLXMG2rzSRLgXE+OQNLR6MiMvUPJFwexRm
uC0zIxG6qe2riTfUD45mOYMsZxc9X508V9oS/4+upDlnMEbttrc7Mb7Mfoa/5h0hg4XrZ8AZN/R1
4IkkdDQT63Xc+ma1xf6pqbFWPBxPhYX0CCp2Xv7R7SDhQ7N1TgBGfGcTKT27oFdPjTgeSZ58oo+j
aU9ikTwKFUZxlF2uOk81Er0BsoHZ/7s/uoYXHXn/wQfbYKW0EHPNHO3i/5r5c3JmzmizE1A+dzCV
W2gmjfnlJX+lxrT9c3XJFw99TBYyoJ9fqhQyX70duZ28GrKjo+EiZ2Y896avolv48FltA/7MwZBL
6wf2Q/W0hbHw0jOIF0rYyMHJgV6cWEA8Hwp+6phCzgxyZ43rxfPH/B6jscXxJx3T3ZdJKSeyAkjk
vPNdDIffHj0eJLrkBzcde/zHPw6VGi+alZXtnfde55XGzLAwhg0Afb4Mzi3HCzgo3IMUNqbiN3xV
QfD1e7GBeAMAzhw97wSicLnCgbqLkaaMyd7/vycJK6pQMO5r/zf03Jqpi90kag02mDfPSKbtWCjq
SXyp9cPFKYuNz/kO69QHUYFn9eMMekoD6Yjw02oSA51kwxBeFBqPHJyRuKm4Nak9D/he0XFAwNqi
mHfoj6Dk46vCAvxB49SA10wlTHTbDtcK2N723QqQ9tXiaG3CjXHtYTR0DA0WXDoNYIq2/7FG/gIk
HmEgcxw3XeUQPh0MrRBr1jHDOtNLol8W24S6noOiQbEUGoL2iXasg/DHJbhi4o12/55HU5eOkWv0
X9LYyIeKzx+jxBfK4WcNyW0qZfZt2WreNIuIyyFBiSa/py4HQS4KX+xhmdq131KQC6tlbFrndkKm
P6cbz6FO/NHS1vpG/KwlUNY7auX/qPszA8cM7prskRuJgCZY6YyIDv4m0O+lMheSnl2reuVsSGd1
ELH1gcpjffVUSKjkZmuKJfPSHmJLq8nTI+ro1MvbKNBX7RWjXUG9+Iw6pdLuS/nnh0w23U9CrbAg
z0zF7+eCDx8F6RJhG3OWMNd8zEPvJyZAJnUxtht6hkDgiGjy34qVrJk10eWKrAy4ul2ixe8sKJWw
Ux7/1w221erCjcGX9RcXmt6S7vKaURKWOHg0QjLaxM4DwFl1l9a7phJFY0vB0WdZAtTZWjnhmyFQ
a7LIE9Xf5sS8p+nXU1espQbXjALR2nr8HaP6SsbjkB+xY4MNFBK0YWPJ6h0xul3Wl8r3L0D6Mni0
zImwnLQao88JUbB1/654cYR7cABcmxC6NQAaVJ8pGsNCiSJECYhvVKCVom7crOAb+0K1EJxL1cJI
h2rHsDNWQshyg+OXYv0H8W+Te6wmuneLTWlAI3a7m0dgT2V8XCk1iRjKF9qOcA0B1S6Jxvq6GvWQ
sgngiE+5Bf+BQOVo/BzbLwMN1r0Jqw+EEMfAnK9RgZ7AVc56YqyPDNv1+3iH+zUDeAFM/px6BKxC
+WPbmtJVpw/5DTNJdVp781Y796R0mLypORf1MY6eEH+bIaLqJt2iSbmmAyQgMZxzPOwGqKQ7lX8f
Zx6Z8a0TEG3q5vLgu0pPxxlD6LAQyKuylGqObcKeUOyST+nF6rl8PKGXCyvQ7MR9PpCHOAuPDkVm
zLBJwtEni8AJD5fV6prFoxpIgjw2afbpi8/vyC6i1uazlK2nWHrWG7zm31vUpKRlu4N3skh4IFwm
rjVeIjOUfyqMFXYmlI/U69TNeYEcpHZC5qFv8XVUAdAIE/MaHH/oYy0nX/E26M7GpcnlHbjREo/x
pLJOz9v2/AB6F1J5Xq6zIw7ewVW7atsQsFRK/z3dbt9aOXGsOuYgZH3Pfhx1N2/HzP6stdSa8BFu
PMFWc1DrUdtnvf/feD2dpKQmzaipXBwxPsazdes2Ny4QyVXTk613UeoG81iMcGdWK32RWt5pd1oP
N5JuVKBlOyCwzXDgUTvkdY/WiDaYwfz0kYfxxNA9cQXPXEKYEs4wEG3nYnCNo6uISn5uKJqwdsYh
mE2MMa/idCgqTfsM6WoJwM4lFwYubekX4QUwH1BSgj8nqBePj5t3rnWFsxdd//wKCdBHPl6WD7D9
bXOlJrXDxPnpOOPEwX6tYOTrQD/OFsj56evIJGRCQknfYXB4sXzr1elX6kjYtjladZZ2OD92D/V3
OqOPo6Nmz943YayXB3osVNQUro76UM9U8u9hVWK4l/eL0XuSjcWwpXVCu3IG/Ub8sgr631AcMQ4/
hw2IOxju4ChTfyVZ/LV2YulPOBxebIka3YatPVNWqe/Nc4QB0E/X0IRpKT6CtMsxRltxTR5b6YQG
oTrA73LgBxrG5FMgV4CxRDZgWwQoKpNds0XKn1VXxFqSPv/E3jFW2xJ77BFLJNPS6T2PDHVPJmDr
DOSuLWOfVoR/4Kw4CrXgiveVZiA6F3FGdYW0z1s2SClhfQZzsgpQ4GTr6SZe+0fNvoHur/miyWOY
OK9BwQfKyBZB/2TCtvzgLsjvaORV/mIvIw7aIu+eB12spO1sz3AyMRIWwoOrvlNbMQbRtxJK7wAW
G5QtOdoOdOfWsvQwGGUhTi0hRPST+RqHcPW8cdMGNEmjlhIZlMD8vBmF/AbJcuMI8QwUlAyT6qDt
rhocl/6P+h8mG+F8sjh2Fd3IJEIGVnvv56/llXFSTc6DAJANBgSCxGL11baZX/LO09A8y4Yw2Cf7
vxBjbMmUQCFX88wumnu5P1fBXhew8KC7D+0NHAina8a34rnBal+j/0BtPZQIHyJHd1YjGrHVsh7L
CSMj8c3/A6Ok5/CMTKrHxfYrPhtNXhQqM8gzuBcuLpx6KKGQY2MUrZfLJ7S82LiScPfmGnl1UUKf
gh9YrHvjY4OY6JGvt9unQemMIVNADJwzhWfRCTIc6DVyy/G5aCQv8QO9gDqZAwVWeSdsmfN6JM+o
dd63rp0aYK1U//6EFhNeB8ThggGBnqWubGTNiCWYxY7WUDoTOmohJGW6iD8En+A4bJj0KAuwzsho
klWT6xUMQVLWEHNAzghaVAZ7n/LqSwleXly13M07UKKbBjfIgM1XD/Su0cZBS3LPzvrecCpBbemi
E9fDSiaPy+uDkyXhuy3AVtyFqJ3f1mmOVvbR3HSP1ThPl4WV/Ij25KXxX8XtAB0cBbAo0z30Ebb1
oqIZRr/tyNtHkVtjXo6bt1C+bvNnu+7gk3QATV5NfXOFbgtmpY+rRg4UiwHA+qk3Z9lbjMpqJbBl
AGL8sN09uXE4ugFQROytAbOiycO6gpG4OneGv3RnfCkzP6TmBD5HSSBinPeWesHAL3of3wEK8Na9
SYjWZGjEZnejnOngMQxEQXswcz0jBN+gw78ey7MJe7LemZJPIAT0FUJKF8LIQuBbJxEJBAeKWGYk
N7T5CKkaBumszpj+7Oc9apTHsUlbvCmPLNYfPkV2WPeA2AIBuD2ZJnYeXI8DIK+WHXP4v82A8YfO
j37KLzdTKaNBT3zlHbEwRej/wg7eTKNBblQhPO+EuJ3yIC6zKrLHePhuhaqe/txbqY7ydYhfGFzE
+3o/CzAlTGtsEQFskHApXmPyAUsfiV772rfeKoUWm2ONuFSAO2q3FFhU8HHKls+J+pqwphXnOgBu
25iP/Lkh2r1DKlsbENswpI+OKe58cNiRMK9nNoqd+M6ZDuh+GdW6xlMC5Cxc8dykCI3jU4hwHq5o
7kooAoMpysOEU8s4RsC1QPitJAG0F/AJVY/yTJf556581RjfbSJhqtIBqkJ9s16uOdw6Xx9ZXR5e
pa7rph1UvGmAC0o2Vf3J+JmE9c5aLtTyZC+q74gW/nsLWe5IUicpnEXV67ts2kr1h1tbCCHipHQG
mAJKK+hagmFUnuSaBVYJK89XXTXRCIprOjmjhgdb0pXiMpzN9QAzjBiZDRU5TAzgvU+KGpn8IFYG
/yiLxsGcEjuSGIQ9xEqE0kqTr+1sZ+tpd0JTUvlw2HfEBk4HlQ2C4oP9rpymRwcvCtfucOlLiA3T
eQ6cHVMqg2Jf2CMVnOLjNp7kNYXEmIrqaSnW19VmlCnS29eR+VM6lqCBbwfwvrsjswBsEGHcnBDw
2ovnZrjijyIimTcFkzhddTLA2E061Q4ySUEPKqvkLlf8kP7HxlAWcUv7jZPIYh1+wEAflk0vQD7E
DOOjgvTtr2lSSg+B/q/rj0Vszjs7tgfGblGkfb9ayqBvUqw1+8ty2qB6pc1X2iB+WoML/wqWmaaY
lUvpn241X6sQ4x6c2s0www464iiKzTlFq/NRPGakoOipYLYV3mVudmjX6cNUbrde5b7KCKo09T5B
CuuCIThUCOHb2HM/8P2EwMX2X2die0VEgmNMfXcfTaiO60YtnOHnms65ooP6gSf1Ropb2MATvxQI
xfQJCfSyG74mMG3+ekVVFy6n4PDzs6hGtHmxb0J14XVeEmY4D2MgV80CegV/l10jDB0FsZoyyY5O
+mbce6C6O71Lo39qZFj3h27npHgUJYVrRwf3NWJmmYSlnNaS8TbbqThBMjYbPRp/z7bihokV7HDU
LIZT//FcbZcbnFO8IQMHWSSSFqDdlBr67YqK3Z/CvwkrX5NXYLTw6LTLgEb5KxJDRg3uFWzcQz4C
RI7phxG04Pp0uqpsaqtmrjkcCOv0tmoVCNQ3swYo61HJy//+ZMpGDzPG5uaqAIjY4Hpb17tkhpW6
rcS3/w0BRguAMWfAmwbfauRsKcKkvj1WgkQxMAwPtETxGIk9gDxhK97tigntRPzdrrqPtpu8c03j
y2DyW3LUBVYI7RGVmVXox8Rw9TXvh1Ls39XfRY0c01SZ4tWz8LdzOQgP7hHaS0ECwbpaXK9svpCy
qzIReFrMqsaP2t1hguqtErJfuS+693QJ0+50xb0CnUSpSmGf6hPRqxnji4RBoGb/lpfvlQ9ZeBC2
Pwv3yojHKXQ0OKSf6zfRqqg8XLurazIuPI+8cLK9LgcooWp+lFQT45eXu1YxUfpLpCK0CDk+Q+y6
rslOnUowF6pEvnQk9unutjIZZ2fdzmS6yxVml5FaDrb2K3wyKPJqo4F8nbVrI/23215FeeykA2Dn
nBs7Sq3Nk0tgfIvslQL2CNZWiOQrb9xhQWpA9FHHUcpsMF0EZrHEmV/D0FXopRTPpo/im8XOSfet
UCI32sU8FwZIC7GCqU+l1a0gSGVlUw4SdtTU1G3hJMP7/EW/mdcJunzbKRgM4Qwt/XooXJg56cO+
J/nd/F4HbqOYdI4gWEiQ8NjRbKZ47XvPsjFF3Jx8N6tqtr6XWtTPhdI8rlNpCyZmUeoEwMfEJe06
o5TlqGb7OrI8HgcD0udYK1nUfTafItdn8YioH2n4zRR/W/duZqzAATNyyMtzyz2gamHea9OMp9VZ
CvN1/v+e5aWyvS1l0Szy9fyPGGj+t/EKv9EGNSy4JbAp20QAmx9eUlDXfeULUhlEo+Uxoqe2OQdx
5/EDc7mk5xufo8zPNnZ1VUvcqFt33gnbQbLRZtZuhiuxMzdlXDNZQPECr+n8TOz7deugt7hIV/Y+
T47302xOeqXVOtLlRCl5761PMXpTXeQ05jFoeiZX6FKofVfFKAa1/KN73K3SHwfEcwgMgXCTDs7+
/mnRUrOpvRHwHJXIf8XQ09a4y6XmULenKSGOJDMlegyCG5xIIQ8Vnu+FYeQen2sgSjkvyFOEjJ3H
e+hmKjnipHQLEGiFYX0DtmCx3+CfBnHz8qq76bHHjfG3z+xCLmRty1LSWiDHzyr/tjwAxHp32mr7
wJ6DQFSNtZFON7HRUKtFP9W8/2fW5mHQatrP/O2qwgAX2vD/Kp1OoNxbqd/EoiHq6EeiVGQWmm+V
YWdlGQUaAhSmzIOKhgmLHPKYaatW1MGvWnY0I7E67VoX3IKG/E2d2uh8pkYApcVQ8cwGPIuBLunX
pPTR+y3qMBVLXCVbfvUniX8RQea6SlurDAOUb5kWH5HFY1+x1RKGkeIe8j5HricTwyiaHwjYmTab
i7255wzY5gE/18TD24v7RxCGzofQQinQuv+8BttWe5XL2Or1cXSmX8uFSkix91KiWBe9tSa8gNkw
f0b05u+4mc2yY9BNS0MkLb3gMLE899DcvEonUeGsWB1IBp50SAdEhXTQtUrJxZW1CkX9CjYHmyGY
4YrESUt3UBxRdATD7ZTIxIOjnpUhbDQNUFz4Thniv7CQifSZCBp25UqcN38x/7iCwi5gNXdnghiP
g/AJOvoM7cnT/+Hu5zGXB4hElolnlStPeFRTJpuumQogsXkgXu5dCNTcvAtV/VECZwfdjR2NqSSt
OK0w2Sy6yGxCN3LN/99JxoMb7DVBC8JN+6cqR1v9jIzLlsij5M1SAnVXCoRjHckfENdEvOXXNnJY
woXZ6/gw7tidIHDFRJBX/DQUF6dLz9YeSacpo3J5fmMyZq7tfkoJmYL2exerYEdT+bo8X9g/lnLJ
ziq9Vm1IiW3q24vrIPcqc4HUTMDwxiSq2YAHKnq8B2LgJ4G48BHO9kXzJWt+WKkk3/X6/gOauusO
aCiLxAr5qtggwahDxvabBQF62Pbf2u6DhZNk/DVEUOPWL5kwsvI2xgrewkn9b5eLotwDIKhRlXKp
TqIahzpsvAeKQLGxWQjEqNhHYsfI7DKe8gSAX6uqFI80dbzj9Bwge6HEiENuHKW/ocSfASnpUcTf
kfSUh18PJbsSTqMeqlrPQYZsG5t+W8o15GYXbDf6jr765gc2wM72tKqXe14GpXjlp6tQcjYGkyAX
1nXzrQGYQpmn0vdsljLzD8vUfFEemHSWRBj0bEooV7/t9+RMvCz46aH8yGZE/SUKcos4fpF2jee5
Z+maa4MexehwmtaGE6NBLlzArv0ZcMt6kSF64NMK3FbuX//2hnJcLjfJ9/s+ddWEvmcSHL9Fn4Yi
fQOqWyzjcmA279qDBSZq31qEKNzzAh+m5J62e75Lxm90Euk6GO1Q4ZNlFlJmC3Ews6FtIRgNW9iN
1EphBWfTdfb/LhVmZEIDxl5+J0ZEKg48c3d4sPv11vHPooXMQNVsW6vW5SHdkgyEup9hc2YyicfP
2GmAOss7p/Kiz+4gkY/MBvWppeKaHB0QuvXlV+hKnV7Fo7tyJIC3VsTxMazjhULatAzfUSGWmKNI
TSd06mQ2i17wjj9188oGOvRqiofHem8wPKbHJxshYTymeZsEkXuYVYoJohU2D7KW7HCe2CW86rAg
pGjPP+tzdW0OVzKeM+8DgKCgpmIfPCXAZxq4gFaWXGgjdTBaQPaePbwuK/Qp3cYlwfdwjF9O3ul+
No6Li2Sik8qCX/aYTxsEDboQcKwFaeRo48+GPT2SJqa/MjMiUmtPhU/Lx3OcL1c6nBsJLwKTqsIo
md6ISSj1V12z5ykPc5yWdJRaoH+WS6wtWRHfrEB1d+sDoGRxgsTwcItYfSBAFMetf/EJhjApp39B
FRChSu1NmLKa4eEqqHLQheqx0H00G5E9ITmLxdA2OcgWfAlQxsZNCS6YLa1kTDyC6XS6sb9LKS7V
9A7fS6B+H+yxdgycuIHA27EIfUjOfhGaS5myk1BiSBSZf2BPpK+sFY/DnvlK/XeO/d8QxMWNzMcf
T3JPr75W/wWjpGNZJKMtY1K0YrNaLlrOAcMtUp7ZugxPCYXgaMqVp3zZ0crhzLKYrQNiOv3oT/F/
5sfX03nGxe0aZcSTdayXFeY5cTjtHkfuXLBtaiHsHP7jk2lV0yIYle6o4VMwKNLS2wmBEoOXoaUz
8uiCxTAXwIHbhnC0eBfiD5BhE4Mnrp4atVR3tPKLFxj9psP1GFqPZJ4b1S1ihwZYb9pmMKGWmXxq
NOsG/l9RqlA6l0zNRvIgK2LMXmPGy0/AQCToxSlJtAKefbHGtbuuroj06XQrQoiSNcy6c/Ofncbu
uz8qpIFwpafXSC0yl/lrItwof+oTN3sOT4DwXU7i2z7koAd7Gh54RwhGWrFgTXVSFQ9fxp38F5+T
HEaE+Ab4R53lLJ+Kak7uWg4pfBQXe5+F/LF4m92gemL8BicUNfCJdfbjNjMIC+iExBBZqUNyNVFA
GPX0zf9VgtUEyLvyo89pK5Vf9q8UyttNiCzXn83SozTeaMCzBZ+++7LXzE0IMKq4rG3PsFERdIA4
X5O7zXUCBWhNev8cQIHaOXtl9ICIDwSg5uh1Qtb4POnlxAXrKtanDwZvQRIJg3lewOGy4QklmUlp
x34tM+reNRQW7mxq05KII2AJmPuVavOlMdi/Ab8LCa+zg5XSHfYKSJaLHe7hAP/GAhBIrpiP+gvw
Yyiai34VHQbvfAEk1D4H6rFe1toK9fXla3wyrZqkfJsVBzeByViBk7k+C7OJEZ6BbgGX1iWQFuEA
6gvuxcVuHSELzsmCp+gArzHqc3vO/HQZBja/Lb1cnbK+s4nogHYVUVIojZigFkOqZwN5QnOA4mph
8tBkV6F2ePRmhCmCk6Kao6rMzKd/aCUhaPN7qAwSQmj19jU0SBw0o+jX+bQYOWLvPbE4sHD55q8c
lIyuvJQrD6HEazO0zU4T3MAN5/pG5YW7a0SOJ79Fk1uxqPi+oMNHeYbXywuS5gHxWC+WaV3q4lg9
YVVkFlolPZVc0IM5Q+ybZTvWRQp8gGHDQ70sloG+qBOPySj2ZaRstZV8wXSjtNSkVPgnLtwwnZrt
Itm3j5Z6TEPCYFH1p3aOc/W5XjrfhCeqv2YVspL+xpDB2IAOd+fWnp3Jqkyhm22zEiz7F93mXZ5k
NGR7rs+PszubXd7m2z5L1VJzG40HYktyUnayfU32YzmVlWXuapeRDz1hGkhOT9+gE/kKkQlNn4X3
QUp1s8AiYcLrF8t/ObHVc9DKAxoxPXPSVXeMC55MYE3A8flz/VklqT/0tueRHGtQFw+KHEQVINe3
Anqo3Q6nc3qaMVHSozvBeQmYXI5NAzeEXqRZV5GyhQ8UJBQ57Jn1173qaPDvcWqlt0jRX0mc0dW4
Gdmy/TJSndPHAFVSnGtDdLRg5yoAUXce8YQSAO2DR+ZqyHZDlRswx28+IsD8IOyGqAJxq4ELdi3u
hZJ3Us6I9b1nzT+2mtqlUMu08ujCvjqjk7LtTNPqxH6Y+JsdyKNdPxHyJUiVnjx3lH5+NpYDM3XA
pmzjLlDZzv7PR6AFZy4xtJ/ZSX/nRm9yumIhobRHd5aGPs2M/D1nZbZBfodje80HjoarVDzi1XF8
DBb4dN0urqrNvh+teblq4QHtk7ihuzUYcMos+U9g0IaNz2fzrKlhBJc46uD16E8drqwA+/PkNCd5
ozeVIntXYWqy/6sq+I4PCLDn/NC5Y1iJHx5bfMdsV2YoVxDVYMdp9PSbR6CsN6C6iv/JJG7x2gLY
ud/KK7ApbBTBE6b+u5G5wuieKTqw5jKdamgZNuXGltcAAuSUF989l61qizRW28yxxrsURdY3E3T8
9QTxFfof13aIdvfq1P6ejvzXN3kKjh+f01hGSV+qy0jw9BOoxrQdvTnHEr+f4Q7g9Db1hP7oNuLs
P2st6/NYoyQwwCPYMSA18Htc0rOXP54EOr+/tDQJLb2uYMummAaXllosIQIWuLzL2F4WRHkVgUxs
vVN34H2selwBk/3xTVkOULaqOoaOaUsp/HdMgAffPVUdI+ILMXsuFCIlALa20u3BsxCWOlsCoSZ8
YDJPq/BMlc54m/UoDsnpa1p2oz4GP8pQwCEgQf+wQS3Zx/eGJbHy2hVJc8N7UkYPLmIeXfemSNfe
43wtmdlWU04CJc8kGkCsKFA8D02uBt4IguDIwF/p6YmVLMXdRSbvCTf66IDBIlbvr1hjPYwJRhgN
usO2wN1NJYdLl6xwPKJeesKuXj33xRpIPNI/zdWxCu5VQ8M0ComROgsEha6rRuKaLYs5vdC90gW+
Pi04KGWx8c/+BT7J6HPsWPd7fYk4drwsjnhSseFnbebLHlyzYnl9Zn4IbA/8Tr3dE3CiHZ7f+BVw
tBnltEMERC0d8t/xJlgqeQLM48Aw/RTMeB7ftFIUomzHrGXi/79A91iSbwrir/Vq+xXjza0gMkJY
dRHSSs4/ifnDGW5YtDS/Bsi/M4E+kcwdrkeIUSe0dBZGZ4p6VKc3GypppPIuB9/kqQafZTrgvw+R
uFGTrMAc0wmQNE/ReTOOMPc3qfxBufDodVgBNXsGDYaL5DHeLqoRjD6hBOhjz072ucDT7jqBReGg
XByiKkYa2i54k5LjUaldxw3++MT6AioY+6jHpZq6xA+mxOr7KbWMTRrWIfJA0um3pAIigznhoN/G
z5rfi6S+rZfzF/pb7OPSbZOc8aSOWcoOLGQZxpa4yuDpfeayxlx7Vibk3KZD5/z2a7ns3+744Ftd
GyUmjoet2fRR30OwladE40Z8hZcmRWiFb/5JL8PNCm+WlB33SF5fYa3gddmlcio0HEvlKrZbNLGw
s9MCu66p0/1XWsFsDHoISRXrHAhOeRUqfHRW+wLGb4/n3iMiZeyk2VEIOIiqUc8laRITyyhQ8RhD
Mo6VMt6arYG01V1ADbx5MC6kZnlJgbf2omOx0kq0T5OweSN8XU3NE2zHBNFt0BwI8KIjh07MwDew
7SpRDJiQ7h0ZijY8iFIR/B6rBk4r2yCmhAjTjnT0XcmFBnIc+Bu2ogIQmJJHO+7Qi9LmKXh4rD0j
1Vj4x70+6pUOxsMCgBlmgQ0dtVyjbCRXpcoXflqWMUvdOEN+B6F+XBxarpZkU218+XtG11bmft1M
L6/BnNUJvJ3j9srAAkQcuYGdkyIm2BQ6On/MAK4sVlCnlrKVyZEnpzD1QfNorGpuY5Hn5fRlJEcY
ujXretIxMyMnOgm2G2FlO/HOfV16vaALslK6MS+TL/VJn3cSZKFuFs64vx/MIN/24nBqoglbDWcx
6RsKl7kY7J3yBMoPTFb+FXNXUrRJaiZxw4kWwv/7Gw0g8jl73kugmlf9OeRAQf1IG0ThhrR7fnnY
h2qOxxwnLexHJ89Mb03k4SBZaYWdwEPhfyq22s4yTDiKasUVfZV4E7zRZcaJFKiMPinim8osIBaR
757GMh9cfSTQLfQW/2/KEtBijrAeUTkMgGxaAFU0r48Ax58ooniqhOl2DcImi4elnyk9uvnTh4Il
2pwoSH+gGVzNg0xWuBpL73CP+Sb9BDDTH9IOItS+XYrjAx1BNac60sUkxXNYZUrt56v/zOAgExAZ
GDZ1ix8DWELBeOwDfYxyvJscLs9lJH6f7dQMunIE+OiOQi1A/IZFsPfUtiN3yva59vPSOcklARGS
ilXmulX71q19518R8Uayf3HYVvzvPanWwpqFzkfyFB9Fa7o4uNSTetpGBQEraDr6jf3/5pRf8VBh
gnEENaRzk6xFlaLgdo3UvVHGnhN+4AWDm0J3A4Vf4/YYM4P870nJokHTUhhHlZkU1lN1zTqzUPn4
AdzEnt20PhUUl8sJ5I12DG8DkLuThyTrky7McfIrMeMkr1yve6u9hBrel+toDdVbQMXQETPOsMvC
xvNONsrN9vF7m6HhSNkUUsKoYfrU+qyXwAh0tTkHrpYbiGG/9c2CPUuFzPpbkCjsqGbV8JGEonCx
JOHtUP8jWh6fdbPmprC5cU8y4um6KPpkTHO64V6aJx5E4CaHRraZg7ttWpOfFqu6py+pzKDV18Vx
9GrFQcG9FCUWe+upzi2W2+BMaE/W89aoYcKmUmQpaV0AAgRWih+VKCieZfb2i7LZzQhF0/Vn+YwI
bnVkHUfMu5ckeGh2BW2Nhq/6IvNyu/G4UhNtaEH16GjVzkJNp+dZkgV1tKqAQkuEMj16iB73Kcwf
yV4O4yMeCyLS6bWZlStEWaGTdFdboRUtYPQqhNb5oA+5/tvCU9yf6EiVwtKWRKwAPwojmRlhbgCv
1shqj4iRTKzQjPpbpUgiHs3WvMQRDyPCB6MFgowQulZVcKmzXPYVtgWxRfhwk19+mSQwbXTd9HMv
xlwjX8HczAoHVenKBWMPOsFKYyG+3p8zs3fkBQgzMGotyvCqkrkGdSswqUB70jjrV9mGNjVVuF4J
V4CdasX/mNHvg3Q4aJtDhTYGXDmEQrhgGDl7ne2QbrzD10RfMD+O21F9iEWVboWQK9JbAqMi0fwB
L60IIOjBN+HeZuTXaAA6QmJbgyM1Q+Js3GoEBmAR46eRbzVX4r7lurs81gmQX9n4VFrfENt+R5g9
/28bN1PCOfmGXP6Pm2u8EjELvWsGualRV1ykF/Mf1k8EOh65pyiHFGHy8upTrO5nAbnptL/+Tv32
miEvsRM2JKculFXdKWb9+jHXYf4li4asaKUVkRuMTMDG7mPpgQsmObnBwKJZknSm46lyeYOggwxQ
wZgR86o12o3PRKcJKJNnm3QkooqZ0Gk9GvqF3lBQ8POMa380ohEfRe9oinWxbRjD5xsanXLsePvn
cnqZ3PfR8mgijvf5O2MtffA4L1qgeNp+DRxlUyqQ3cgwouek2fqORW2tpYpQKJ/TMUZsPaG4d50H
Xkeea5LxK42PdR+Vy+qw8jAIMjA4DS0MN2M4gpwlpsrPiBKNKMUEK5x4KXNPHtuNP4i8fQZG+DgT
U/C+oarucUCNHERMKCcp3UAE27YjWYTuH3mFFI9sDbQ/osUp8TykmGtsC6rQlaryb0mfI17RyZf4
WBX02+gY1c2s7cntqAB77ghEi0psXYV4hKsfkP8NXVa5lvDOvQ6F7mNS1Zt4I9ZkWm3E4LCDu0YF
f3PJ/2YVw8RU0iNxXKUtWWu06xXiWCMS9aiAyRPXd7hrZWVJ02bMfC4mCucTvwV1g6ekMnuu6/0g
Te8/cvK3OcOae62joEyqMwgt8qF9Dzdv2rBGn1LxO8ikxptkDah//Jtbk2q8iEhDCprNkDFWllNo
GQ5b5wbF156a235ymg8jxx5b/Hp1AKmsJ4q8I9mChMULO470j7rtFbBGdN8CbtpYZbQmpYQATHf8
ePq6LXNi64OxFZGdmMz5McPBhXxFfLZkC3KlQj1k2xFi960IIxNYqH7JQeZSgIEzyPyqueM9fCj3
V8bjV6znA6e+ZRhOwez3fWey32mvOg3wFCMjrWRcnFeAitP0s1dX13kNagNeP3kBYNbVaolU3Xyk
V15uyfsjJ+riF3xcq1bLtoqMBVS2pAkfcz+1qALJLUqd/buAZrCV0OMTeel69+TorV5u6hM7l1Tb
NyCDMAcXwdj8kp66FMREECEKPBNvPcKsnoOV1srE3LrE0kAvAj0DIXgWTGaN4+lYgtoczOtqF83j
BUUsMSDZ2uLCQEIBbsbuFxYOtiOvyUhB3yL7QO9GCMf0KYoGUPY9dMe3AbptYZ8YHOgRD1loM2w1
GgF205rswGHir0ff0Ci6YKeKwup6bYy6y0/A0Gf8jrW98E+0DeT9joB1lG+CypvTunFf0pIl3oO/
eGfKZ/TY/hv7/RfdBvhu8yxeVevxrbsV0+e6kc9U9Q4lEh/aV8DV67307ZpbOSNIyvJOGvmPg6Br
Y5P0mQRpg9mUkFyssNVVsWhdc5yHWMUSd6P7zItn1Hc2DuXnbrn0hOL9NAJH2fjEOqQTxcARgRq9
jLk+d1d2UqL41Hh7bh4QFxtWo/iEsMzMcP9amC0vAZmDNMA1COaWGfcBYFEpz6oMwh/0mB6kvHXB
SpIBPJjVbPbgmRp3luubgW7UzDWVLHaFhYN4HeDBweTdQCjsBgA7Yhjsyyr1PcEKNfFHsakmaiHR
L45aPBvBzb2TlvkiYH/SoarVwf0Ecsqwx+gXRlDzq4q3EHJj2mBZVaH7wMtiIu1rPr3AZHfT0S4C
KaXtAu8lTDsOwowzjFNiqk5wpE0sIMchUVD6JP7R6KW+5uAHQoKQz/95bDZXVLLsZHn8o86Ct9Qq
RGy5uMVNKp1mGAlqc8HQIvpVo80Dn81TpY2TReSsj42TzdyZDcqNJ+/ZMc1YjwLZ/e/+A1WsW6UZ
4nssWWpMXNnMAJEqEiuJLBudBwhWWT5dDyEYNLsjRMebjOZ55731dzsZmGtJUsQzZkt1Zs7Dvya2
c/h1brOsLCyV9Jkm2bLzOhaVhliTVYILgBDkHBV1zSwmua3mBxXHYfFV5Ql6gCu25Tpk6RS0uDa0
X53deB2/sdxRtcsOfp9xYjVW8RouoZ3QraHmD34Np68wJov4xTdd9+nV/XdpLaJufUkxrlYEqseR
BmGj4N7LSFhZGr9jmU+o+HBCDvfvC2qlkTKCGfWoQwCZB6/Eth1QA9qnG94HjThxcC0Bb9KgmwyO
EpDzygJ2KeIumtQxkdcCctm83H5+7LIi6ebq6mWobpdPWOgKtjpnYquEUkOXS1e+N75g+RZWXwjt
OV8sPE/PAtbKBfuOTdIjRhz42BY6khqrtbFGhunj9hPxM11dDNZ/ifmjOzICMaXqJ7dzwugiDcbB
mIDEZfM6jj/G2L22adK9QG7vfZ73v2ap+HH7flPOLQO4GE3f0PNErS39q7i5JrgJlB3iYxemn5Cp
12znG62+gpcgZQBGbzaIHo7LgVabL83rYU1w+mI/uyZNomVVMm+XrdnsuFCb4Ehk30vMuHB5wxgl
5h5KwRZh8+ojVoAtSJ60Va5gPPXf0ys/uf7RW1GuA9ILmTmcrM/tUC+BNPn7vIFxrTrywx5F9WLa
OfVrsev2m1CG38K32kXg0mzS8p0n5ei+i9KqXQEKUI5GM5YAnVTqxHC2nAjOndktWICZouozO8U/
CCqri/8QaLTUKnE3VkSuOLpYMDav+j3UjtfSFnK8h8k1wmJmr+u37BJKC8RtKySHsilBrTmlqnIF
xpFGzFFhnOqMwm2uaF5nahdBFpSq8zYYzlbgEWpU6+5DKUUM96VkBeyy58oCPevaHG/HZpVsT6o2
cRgQnritB8FjO/cAi/om3FkxboGRHCAvts8Ig3co0Qtf94q4YOIn2mPmCLJ6iVP8/qVvxrQ2hkHc
w0olpvU8j3KEolOEXDT6N6NqoOAkM0KNQQvwXAtcAeK0Y4jcq6dQKGRupvpcYsQ5tzDa7ivkUxEX
qIVlEHxvG9zR7+LhzaEyvc2QNHiFYGCPulBFurhmVgfeD99fWzap+7fEVYTlKga2tu4AHWOvzpyQ
nnvgHy6Bcx+Jlwa2iNHyTbwtf5z+iFXJqzTLbUvhPvnQmRtPEWGTuP4a21S6K2pn5X811xzxaL/g
K9NJVPmPYn6zmwMqMeb5Fd6sLPXRi57lpf0MLeE96BiBUH+k4EFCVGG/pv1rOOE26Gr/C6jKEaaj
xkPDrkhtr4J8jbcV/bb0BBY3s/Lxvy3n2YAw/LKtDbPe5qx6q/KX9fIozgVGt199xPdEPJnyLMh0
wpgS8uvPzvHVBL6Zb6KCmUdElFMBpFnod8VF2X7THI1BZiwqTJRhmLspRpzMGncCgaFG/jaMwXPj
OgEvvrYY+zOhgVobHPXf7PgdzJJzxTb49wQTB1yjjxQE7RTkX/lwmJ00+Y/iRI/VQAZOnA0T9Fs1
dkZMLYpozLCudLzhzFpptIU7eV0ReWcHcpMcV6L6Xl0QwdHld4iRScJ/foMnE7BT6RFOFrD+FDEp
wxDhTV1fW1FonwQiD3J2mZCmckJKtYDNEKapUQRgc99aT8Y4nxrB0rk0NxcNnYXbYDBYI/KcwUA9
lgXTY1b9Z6TFI4pflChr7wmNbuxD9MQxTRvP5Rmoi6VMV45pobjtQHr7K2jEfH9U7HttM0Plr7I+
j87UYQ8iesGvQYbfGH33xB2mbXeHrDjBZOUAXLIaSBNe+wezVn0Wwh9O75rusepzsy+k7uii+Ivn
MQCcB9Y2n9aMrw21UPwhrgecCZ+S8SQ8FP6t977yfroGcewlt0Sh0OM67dk3IYQ0do8Oa7oudkM3
cMT1c1G4CsB6Fj6+EEVtMXwjMhhiw61LM0OakeKKc+jOxgTOx3NI68RxDC8AjvP6idekKwih9a0l
TQUQZqe8MftEkPd2hvWL7ayMaCkHLeOP9u+vm1O0XQm750i157rcuzzXfsFHDR6YeWAAeXY5scDZ
KIEqv/ul51D53jrYU9dqAPWx/dWkhu1mA2Bivg6BX67AlFfwAUuazts4CjqahivKGNd0RX111b61
/+3GwJgvV7mEtEctGpdrlW84lfMJkuwdN+kDE4+YZSUZKR9dxsbVowecTs3m5xmIgK5L8rZTHLJf
Eg7Xmh1r678+7Sd+UjaLu6TTPqwggVD0nFuWyi4l8GyEoE64ZoJPBdfttXMyLC9/MFwg1/j5YujI
70s5TXmy0Co/vU/TR5lmNV7ds8mAh85xOBn/Trz14EObtXe3E9Dj19mGVXVnIKQvwBdEEjUDIVo4
HVvCjqnZPQFDZ6CTe6lyPqaZTp0f6dHlTVPDNIGabvzQlSymaKXLuddvz0GrgbLdT0a2LmjWKjPl
76IcioNCX0lYuB19Dt8R6yTjyWXcWZswEZ/9Yc/XEACMu9tu65OOVFndGnM+7pEisX4RJs7J4MVp
cDyxEd5xu+nM4q5gJVyRU6SRhCgBUAzFP83T415g7x+0hB4ovFCfRDqC9lk5yZ+yQD7W7O7HlhOu
Sxkx4exdYatIR01oaoYcihN1hADWbgLO5S6EYgf3AXJjmwNONZOFJxN5iLm8IZIoDbQz1RHDTNU3
xMagvFQyIyBnHTpJKVUM6GXXAVbwS18nDDBfngYrT5EGV0VOcXRTuxLF7G8LBVfwMqtR5gufAQ3h
ZfzHFmdTvPfow8z0S4yTjxc2FkVKRtnyXeN+exxVOsLlc2QFvteroOENheVw1pVPDyEmhLS+aZ8N
dUgvp9mXb8XbCWCvlpkRnR0Ib6RdR4UKGc9zb5zQm2GaGNPgDwxlbzYvyMiaz2xvTDAl+CpFQrhd
Ogo+PDrsCn+L2qyjIXhABCtybpTouqP+Bsy5D6nYlD00u9SlL0rxHQplDnJpFQCI0VEa4k7Ad0Nd
gEfZ5LAfthvsZQxYzxV8r+Ab+7K4e65MIKBY0p0j12esafEJI13nOtqAfrkG6pK0T60mSSeXmPNq
6JJSA0IDpoRjhga+h7OHg9AUpzSscwzCU9lnuvIePm9Usi3mtc6uEMSEWqWNb1EBxcWZ+sy9oE9o
hbsg8VQ1Oq9LRhCZzbsQH4yf/jTgwktE4iXJ8O7T2tymfHOM9Kh9J7I0UmA3RY2nJPs11KazOWpS
qpP2Fm7GUe+M3GattXQZNB3Q7BQEuYf2cyyVbPI5PWCqRGuJ3GfvQSD/81wa9znzOM4yKUr2iAZa
+9ZfwUKEejcfjHtbnCP+KRNoNgqPyFUXUanUe4LGk/YGQgXl9Y31UlLh04eoutHHvZ1qonaSE7Qv
j+AR/+B6xVVfNo4IE16yqEcaXlFPf7RoenLIaEpyS0zFOx1dByEAcQB77Ji+hXrGJ3hj3i5cDVHA
DU0NRncsAI1y0gaYCItZfPTS8LX078fWYfLv6+XlSMLEv9GwJjpp13/at6jnJja7Nla0CkrDzrCF
o2DZaNmmppPGKOpV4CiymccmQcflmvi/wlKqVxQ6+9tZFFvuwAj6Lt4jTG7LO6hduPRH0p1LmkCw
6O5bwMo3edk8++f9j5alzqiFSwX67lFuUaX0qnF+tIO8s4NMqIMtq13VARcnkzCN08X0gwwMXFaP
nFDaVXRRV3lkF82yOqZllBCR+nNi85ozj7+gyq8WDAG+Og3m9swBa20z9mZEpivuubdLfcy13u27
kMEWyTzQzaRkS8WCAE4QIxMv8vriKmi5612mD53BlQbvBydH9CAG1u+O2XF2B5lqagxT11/qAM5h
KkfoFwfJmKwBu+kv4/h0kfdvhhSg5oXKqM3Xsq/dx+ExoJsiJrcio0wRKrsm2dVs+I5nXypQKnQY
iOP2reqM9hu3GxNZBKVrr24BJnarH/TLQBSN240Ha16t/nrXoJ1YNtc7tnn2HtzlOhkhloqhdRbW
6CqKPnRo5tQW7YdOSdK2yuvpsHCwuGktjUt97Zum+W3k2I1lh1zg0MiE47KdAk8fe+4JAND2VB4R
lUQtRUB+XFGHKgkBdRZ45fps755dD074LIF21uIQ2qjC1P7LsfiNANp2yvv7zMgSVMYUbWebANSr
jaCjE3pAdvces/u2mOdPBYoJHd+zg3FXaVAycS6jLPflT3Euic6IqysGHWF6qbENcMu7dn6zA3f6
pxzD/pDGPb50IHnCFA1NaSm4WEXedk97H5m2oywitPMyOF+9ZM6trzkzjaU2zI8LcENgwW5QmDyX
KN261HMNDijrcFIvNccNG/rYb4RJDN8oZgC/ByNvd3wWzmDxfGxc3j4InW0krF9ybtgjLTMq9JGn
NQyuiCFr3lpjl40cu19Xt9+NC4nCJMB1rEiyeeP9UrTh7hNC0TBXys4VYyGNHj4U/1IAz0owOkV4
vNOLv0AIXLFzoDfWxruw7+YsCE0QGACCaIqmWJSGmGV/lvR4zuz7A/nBA2CLKC7kuP940yCQ8C7J
b3l2YfGb4NkkGsfar4VYPyiXJAT2FkAnAK4RwYF+ZbG+qs9Si8tlerhEWOtXuR3QD+EWrlIv0Jen
ZioRhUOPV4ui28nx8JUvJNJwX3Y9olrlPAPAXuKLbXWQ+jZNBRhtJse4tUSRANAN2XsAGD37X2he
kZqksvR1qwHZbv7Be9X9XkvA3Pv7kp2ZmH3ia33xKtbRPwu5bbvxhXLe19PxibI0nP0NYVseGEWt
zcH5iGMKE0tDZ44yqvYqHsAcqWhlvRQ6PSSKBsxM+vQBF6p1qcIXAe/d+TnH0TkzGqw/HGDBzI8Z
7lgh5WOasePkHjv0iaA+hy4gUwQGTIofa+lePgRbHZqViMeGvShlNYILbOs61HsU2TshPEUgN1kS
gKO4W0H//oyOmW8Y3/xoqDWA0Vtsy26ypLVa7T0n4FtaVOwWAzQwR4YqbnkkfbPmaK+mQwHoB8ea
mtwdYFsJRzt4paVGWSR5Z5uu6igynRGf3NZpWtSwm6j6GX0giwsYc1LvWL//xZJiamTQqguDEVIx
7RLfqS16bnl68GZpgUXYLT2osVoPFrdwxeqLuzvLcmJEeouStwi5g/0NJsUnEMKGvQZLzJb/1eNe
CFNd11RaIttN1nYcJiiJIwKJPOzEuQf7m1EaDNYElum48WrIhTYBq/tpKp3injmjOUeopZpNlC4v
Cqle+vynicxyf7EPMMriWFmkxfYDnKRA9y03aU5KAFl2wVNegZ38pmqatPv6js7FGNoT9jSnVVhl
KebyjzTu6miFtrA7kiWe0YtfW6sBHNmukseDbesv4pmZQPzs33rje54NpRMX1ohFJ46EhqDtRD/a
Aentb0Zr5+eUGMkWjzvdgmLXWaahE+5iX83CAUUBRQt7bjrwrE3GGi6faqSywWJH0piRbAV6FxiD
oJaClpwUGCBTkSooUE7ZALCml7kow4xiYNcDn8H2CEOvCjPTQj75nMi/davt/QR6ompUxC3Mjizh
3cW55zUDM75jC2ZVdd7gLnV8+pwD4sDX9HHPme3MsPlDJaShKhjXw3uB4EMnn4f9W+D7Rbg6Sfih
jgQVm8lWS/htybMWjoJP4PB76LT94zXHYn0GdwMcIcbfRVxQiiPVuG6LcJHqpZ62a0rflcoCUwe0
rrTuplo/AMr3SWeNZQ7fvzPzPxFDwKRXlSK6fGzT87IeXqUMZDS4yXQOPwgrjWQGSD6Xz8W/XtsJ
T1bKHHFetD/0VMum+B+aF2iSFXUwoVZUiHRqRTLZ8BzcQqftwGi8LXGFOB/ssjIw4iiRs2py44sX
M73VmAiegoS2OActmQhMv7tHNA2kTKTXP/CjJar+V7WYC2W+wlcR2h0oTigMEZzsj0gSo09hQZ9k
YTJC5TUKFo8gpTp1uMkkgUSPpIaG4XS9+H1A6m1C0+3QB19n95mPzeHH8uRm+1Ti3TT7jcYouSE4
CiLhyxFMDOiqNa/6jrSwrs057F8vUMK1713lE9/KnlK4kI4F8+QUj5LvZEtDd/BQ3O2giWh10Q6y
pLv+e4XVLdutztjhl3Gnyn9qJPUXhS2y16CWTz/OhJw32GKOaF8uf5sNIC2uPkCvDs6Pd+XrqmXr
R7CB9iDHFg4BKsDUTs+ybTlj6us/RVHpsgZCr05Gc3RE3iqFUR0bOiLKJ6cEUTog4atXD/HYXjx0
WO6lltae4tC9hDDG+uPeyONfaLAGoR8ISvxjMkPrOvdWs4vR4XfSu1tvIptiHal5rW/DRQDgdvWz
/qVGBd1MwdsoCzCJ575PG0rZ50e8XaZy5LD2YGPoTT2a/d8JaL1JUyj5btWwM3xiDGMSTfo7xxap
0MK4PDVF0It5gUNxwjGwXXkZ/Q17XcLmcYijmvuRHBIr4RQfwHdc/GL7MiW0BmXMa+GKuDu/5H6V
ICUr2xzz8H/HX9vV9E1Y3uCtO7HlUMnLzkXgTMYbuHf2XTen1EP9w7tYKEehHjZAxWQhXiPzOsW7
Zk1Vi/K1jHaeFv167yQlIhiy74qAyfg0fOixnz0hEja/enx8bRlOAEu3SRv+dN5u55zJkomRTMKT
V400l22JDf8hUMBuodGLwpY11u+ksmz3P0r6MGNq1qhyvWmoqenX6vVuiNhCu4x/7q/Ce333pDsK
LybxX9PXVtJwkzVltOBVPkvjVBw30WHRif/nB16eKtmLYoQClFPg/YaCa59FtSiooOP3jPQtkgPz
u+Ofpz7Tua1E/nG0H5uaXnbspOUcHeIAnb8Ywt/PqwgyNweQNCUiymFvNOS1zIxTkIJKwxL7YDBf
nHiZnbI7AlXCvb4vO07ji4n5zJLRwvNlCL6+ozWVo1HzusoXO4BreSpvnBAhNbV8MCDZzl66M+K7
fmQn6WH0Y+81fBRHoyU1dYTFB+x9hLzYwB9UG7/1lXuLFgBN+8PguZMzyPtWPAiR4efLgZ/JvCOw
ck8hDEOi3GzHIIMHEgdRt8Q1wYmedATdv4LiwtDkKIWtx3NdfRo+om4aAftTic52iHmRKPVfctJt
QcHyERwPH8t4YOo2MlsigOvJ+VMhfiIZpN48gtNeyfpySEAb84GRMwkOKVboWUYYw1phTeolQcMG
WqQ1XecCUZdT18TKJ9OTwh3mw/CCG42FEq2lkaZDAznyln7qjwHUm/dEx8wTjNUlvPbG5Fp3uiFb
cx8CACtrXmSeOt64Ojkdp/Cf1hMAI+2xXmKZX+5Hs4DHmqD01Tr4qcX+OY1fVLDaCuqaUFWMyIFg
FihMrvGu2JdIUi3RjJjD6iENi4QSIj+oGjJ3G21GsJeF0HGCECDI87uMSKH3jn6MiPcUfVF+AWHD
DszlSFrkKc34GFEwGrVtkqMPYbj+ZjoXV2j/hT0WzTlQ4JX1l1Wk4sIkL9xH3mlBPSrm/lHUN54V
+5CwaGVledrViF7D50Jo9mAH98nFjWgd2x/wcTuQHqNUxxAiNQSiXNFDmDmnI5fQao0xbYnDeIx9
Wb4ZRRfTyOBGxLl2fc3mr20MX81Y5fhBWdGWAxirsDz3fK4a5hrsYCUc/+R2O8gxoXaGzvvURCU1
n3458wt8LmHgBuU8nyFR0jvVQoqBVFMwRIENT1r6mCTNSs5yQ6IpeXnQKRRd1WWFkvHQkUgqz6st
RnixTCFxXSeOaiZYRBgh+nzEf8OrXZJaZiUmTgOGDnBy7o0eamI6AP5p0jF0OY9zotl/WVucDAaj
Xz/RuFVHFKFpO5dpknZ0h9bEvQeo3FmKoCBzdW1mRZfsdaZ3yr7SbRJYdgXgTgPINGkT2h83CMFr
RtJlw4cJ3g1hchWFk3tg/LvSu74N24IaeEkUDmokEwc6TXUsmA6tgLPdV5POI+/rAsg6nYS8LGoa
LQeSS33X99V0jzrljIJFCpNyy7Ex4L1JvR+wsCPbI+060NVzoy3YYiujLH61D8hLm8fK1zElsJGE
wWvArPbOFJac/f3lijD65bZmlXzaV3HyuBRPAnGkvlfiEqyWYkZIr5oRRhME8EQMCJxwckwE/t2M
55yihwsbUz6jKcL+SbB8pjNX2/srggPOuC/m/CkSOT72yga3T2wdzcj4LKXNtZnPc/7k0hOxvOPP
chShs0+4fUkQH7j7H3xSGhpvjagVUk8HtchAPfDJWem3ZWCsCwt2rmz4alcZY5dya744igBabLM0
01g987MULBppi3JZt18zN4m7SNxAiFEymizV+Rmcuj0fQSNiSiRPfevbCAze4BBqHPEwBxrH33dI
Fi7QdKhE4x4fhvsESnhi/xtHDtZ+8hnz0TauIfTNlg3dygPtZOKKt0eK/wkRV4Fs5U+NLn8wRQHh
mYSF7hIp75BRMXoZ5Za0Nt1KHKgHTvvUJnysuExfUMgyddB7MTeClk5yN2NFKGYWDikmcs50XeO4
1EKtO6qgY6+LObND/86Ekmx6CIDmoVQmkc0zL5pmE1MqYsKkZvRL8AF6+3ek5A4yStisRv0QCcBi
FxzmRIt3N+Cdwq7yrpOYGUZOjiMv233Wd7WiG+rhLO+RhvZZh8uCcS6DWu0uF05cLDCKVydWVAqm
4WCO/1ZhNP8QyPR2xyahW6fqeGOVdHxIt/Wl0CGNqZeVzotcXS+Coq8jrlWbe2Hr9r+tnFleZ//g
11CybjWxdY0FA/fX/Z/jKXZlS9BgbIz+2j/iSU1GfX91GKufpcKNnUY+He6f67yx2/uTjILcKF0v
d/gxwNElXinnx13Q+uo8LnitTO/cCAJawULhKyoutIugb4pwrHWkeJjWPp2zvow68I5lRmsEToPD
lRRkSzyr2J4T6SLXgb8N+7EMRPMZ1kV3e36rXGAkJ6Ysk3aX1CESB9X8jOzWLhm816m+IGeGqKce
Z8mEOO7704rdhWeQKrYefOVuVeCUKzTkAUic6t2XF+YdCyuPcXNOPqyyMOjah5mJx5pODzfWQMkT
adfEhw+0jVfwMZRNccNfpxYepJv6SKHKL0+qn9dp3pky6H5H3oG4dHsgkW98hxJcqSu/577AxegH
SNr8sJ6nMvLp/xZEQ8LWKIjdXuCrvX8uYPZCzvQZjiyzoCFPy/WLYxx3R00kaU3w9IFFiIWOzGtY
Srbdu2zRkcy1wf6P5hm7FX3XtR44ceulH90KcdlO+Q0Ej1/i/IaJHp9Qze3YgErwLzv++iIgDfu4
Ua8q3uK/Dxu86MdCpIAMVA6Cr+DTkdClcczzzAZ8DWluyOG3ZAuFt/OcW3qX+R6YtC7mSAUtpHyR
idoegnPFykpQGdEYVgydKnggG9pFGsf0SaOzLxmRKoPf1xfy3tnns2qhBkK97tIIQMMdEtAqxVLE
vT14UNytDexPM6FZ1Q06YaGr+weax/ub1F6WHHEOUndRsxRhYtU3fhF9FkpdZo5NcL5CYcHX4p4f
0N341MbXOlqY7ZJyOSpZKWAPGhhhy/7ssmqrZw+2wkijajQA2wFo/BN9EctzFwNbvDTIsInz/+/G
4VBWKNFHhyMwR+/gfqBMcfUiAgL3pZ9tcmWGF1XOyxnDTTKHb2IKH7W9F4dqx8qPIKhpHbdqSDLF
PgIpK+WBPH9fs/5O3h3yZoeA267oqaBykJ06+P1+ZbvR8k2i2iUc9pCZouLRyPPd+PalkcqHe4j5
NadKx2xPhXIqB5C1QP5xHikadOg3nooVkUFptijya9XKWaIMLnGTkscEmK7bxODW3Sk8zD3YN1BX
aYfcpWjL+eezsO7j4jKdFuSXq+LJE8LawuskKQOSIzXY1fpkA3yle3Vlus1HL3Ous5ERvMymclMr
uPLXVQME1dadJ+065Ce8NpgPe1EWDQdwkbmR/cGJ0hd8AVfv+MHe0iN0Za5xYlGJNILFfzFYJtzG
zvtHP0pQqbC+u2B6QMVfAKtXGy88xafAt2bh5uo3g7qhT6p6aBQjnF/Wx7f21mccUs3Rs/KL3BIb
V3N53tjIH1r/jFoDI2FaMBq1Gy1ICJ8vBDPD7O7PR7KT4IQjBCKcdWjxlnV7GqSTMWO8WC1QYfMl
8QxgwJEjfCDcvlQjvjgWehj6Ni2F5eaFFXkzvM9pvorShRJs6tlmTgvBDlz9KeqNDbB1fbhiWE/2
4O3irwUIgRNdPrcpOctxP+zwf/v2MJKLYrUIMpEA2HCPtDDwbjmzANXVVnpy1pdVgp5QddcLKttO
FRczCeh4ewjpw/wic2geuZvUHqZvh5rL7jQ0ah+bO+EJOkT5bN9kP6PaK0nBC+EBcSww3YdDIQtl
aC/bZ6BQovDOVMPvYP9cAzwNMLhrifVYhqTF1PM0fo60mqaCnJk427DFtB8Ev5WaRjgA1qoIFx2j
xs4I+iHAYDjM3zdC2GZ4v9GsGCFqHXSdUr5IdQEDnFxGpwsLPIwWcLFACCyDtWXpEnDhBtlts85m
JVsZF+3TJdLe+021Sgto0MYYTj55l7+XDdJ7X6+dAZR1npbRhZ5K9YokG3WlH02/oo+4rIBr9o8q
qYQwxn+w6DPhm8CDzZGpKt4LfuwqIfQ7+veBdn0tNLZlW0Xygd69njINV3afIhRUJSDp1TIhul5n
0JuK4gQaRt4RdOBkti/2hRE0MHZ3PS9Uo18RMOD1bk4CI4DJdZF5bwGwAvbnkswTGOjgY0asSxLS
h/FzjkvViwXYDHgGsDkj7193zreJau+bBbIDTakVvxxZJ7NY/I/qAGuOupTqndf6ryU3boMoT1FS
W1W9/yKhw9nJzsfRzVRlUPbI9M23T4BofdZhAu5q/1OnJbSgRTxHRx4jJ09tcNnAoqYc4WyAIiiS
LueuwOfHgWo8sdBiLAK8xWhJ2LFhlSkyKDUDFCkvTr1YU39/TGdFlOaDOkhe6TbuvVfmXbx6FZ0a
yMlmpUgNeX/eCk87csjD2t4YV50WK9+HJY8u1abnvrNRfbu9WviD4k+MP1GHjggGEFrML9qEPnFt
bfMcThsD+REn0ivyWO40rZDa7zeAlsVJUPOd+F5mNWSq39iv7UPJ0KDL4CiW86m1q20GrZCbw0Wr
NNDyLqI8uywmQZ+ScrtLpZe3qY1qq4Y/pxIGx1SW+wh+V2bg/jlsIx2tEkwvTYf+k3Gb4lAEw/bz
L7jsGcg0aA1IQtOQbj3bI1oGcj4DZh87NrQp8LkxXIVOPvtXcYpWE5yKaS9DyfRwriCM7e6owqNB
9CYLPcCm6VG2TQRFAmm5XbLebKMK4Yajl0QefE2z7UXDQ3QCGX6X2vAkHXmw1MDpC1NA0Iq/BIFV
ckNdp+jIrlFqX3lzthmd1tieLW4uxTPZpXDGvG6EbZ3nM8wHRkUXO5NJlRaGTs2ihTWLgHTu4Qwg
gZYs2U+unJAXjy2w8ZyRYs9nyILP7HYCerCBcXCbsZmx2W/X9LwQmvzpEmypB9PbXa9uWKV/WkCW
NmKkm1DsrzfuJcR0FijV8IoFBZoiYRHC4UUolMJrol4U1lzeAcjU1ToWtId8QY6pn3Il1+bxd5ml
w7+W1LS8vwjARdYYtuJhGKIjXN7iLol+Ngon1pQsA0f3gDD3R1Mie2FkdM6z+ZNojNQhCbuX9eoP
VgJzH7yjTKDEmtAD65PEH4xycWXx1qSyogi3V+WuK/HQIBX1jAVOIUPS/4hz0GvC1+nMUNBv8AHt
zJQrBRnT4+3Xk4koy3LWhHW5N1LevqHYZdFOrJahw7bF7CesypIwW0LLmYEYnrMmEK12wy5G0Ntr
/d9DzCieTxlfH5ArcU1DatJg5PKahvdW8rBxwZQWkv/KH+MvHvsSEKqePwMgDOPMu+xgioCnVKTX
7E0SNPCRQDrK/YNGxj2ZvxbKma6S55rrE0dk1R6he1TF68TNgs7tvZBzF/VfebYJxzMWDRkQbWLp
qx9j/IM+w/+d2NsF0fopDsOtiAJaXIg0HZMGNIrthBVZ3hHu7+V0DXu0eQ9rq+YOVQ4qFNCcb8mk
PdSSGI7A+y9XoDeV5kOqEPh+z1yg4y+B+pUjDP3gCJmgjUUqxBXj4YBvikCre/h3AW+ILQ1K3HVO
SNIlIoEFbHU8gr2JDzpqzPtyP30pXkic+razeJ5oPNWy3uwteIpP5Oerj04kqcdwvTn/gSQ23Gbo
uzj57wyQALhLO1mKYR2w8pJBUINrXFvfb49DO9+GRfbxJIQ3rJgpQN06WKYGCBwe9YcQkGObiFlP
sfOPsvlwQIKiTnt51MdAyiRQFqHCv30sLFArgH+2d23hcVgFvgar7Qcgtw6bTgPQgjqqBhWVDT7i
3F/xhzRtwjtVyqqVyihU3dAIQ6eNPlMpKFonP2Ua4FsZBpfglfCXcFqO7HzRJNClV8qYY9Bo2pmO
9TxnpzcnVSatUB4nsOMY+hIHAeVIz6XQouG1U9CttwiEgju+mweGW8U8/eqEaIeSYRyFZ0HJ7qYv
4XBXERBEHJWXSEQowPewE7MtHF9T+QwobteSdyZbWLKbcrJN2le7Q7jg4oit3PTJaP6g1NnMPpD5
ZvCyeJs7v6EPgv4Yhl++lOqkTF6KK+bY/zdUlo/Izx5tIr0D99iF3NnQm89pfRU+9BsZJWo7oj2x
IBpGtSve5C0rVbvGP7DPcpJR9sCZ8G5DfExWjLQVRrpn+RsOXzwB5nM1/KLd/e0TwR6zNt1E2wa0
sdOy7yI4lhmUBSDSga7427mlikYtfd47yuiPnGUfSzQX92zBFZytdepSFeasK+s9sNIlYIPIu/Ps
NqpwAUKwxDDw1cMThK/EWVTfXCIqJei6Pc6jPoyWNE489TgvUoasaohirm6NSd5sDjzSPR9X/uOA
J3V5s68ZnNvf6Ea3xjlCUpDXXYUm56BqfFP5Gx7DkuV4n+z6DadW5kVOo+O5Q9nPC919cC+sAal8
HV3CaCXrPAaxjTUC5wdamxnE850uuZDvLALLdYOeO2j6Gjh274aZc13C4jBdvbFY0N1curBXYLo3
ce6spc5pO1VJBRJbBx9gg5mQIb/ZdmEb7L+N/NoCI4ChDVt96zQ5DCsA+6GchVFGqeKkR/bRvDXA
1X7wS8k9I1grdv8AQbAdxOcOyv2Q5oRnCDa94JBlFsAcdBW0WOJMam0JVmqYCgvTmGzbkwjsEndc
abidwVKAJMz9r8RX8b/FYOWXmKycMQwSYRbTEmhgRdyzWTwImc/8fmM7lTJmUyrGHu0/6wXozLGM
uiKbepG9By7OWBtN/JKJcUlZZ5PYIwkZkFEsrZ2fP1I8hN3O7MHDqPPkTyDXq3qguKwAZ9htNCVD
0eR57SYF0cnA1/NPY1D3L3rrFGAD3b61IgJWj7l+T1/8usMrL6gr2LYFzPtpI/gJBTiwdNAJyDK6
fWjQimNFvmP8CKxcOykJT7j3OJR6LuYX87u0WnI0PEOqFzTJ0QAIdpExoKJZve4h83LTR2eWGVON
uiPySQmzDdJEAQHEnyqb2h9ElCqxsoctSvp0ChzAxeqQD6Ye7PLxRg8ziBC7pUUfQv/yVqUty0+G
0M0Q9M7RM9BdXPKXXU2E5fs8fqGGuJXlIFCbbZcJ+1tpYIpTgNbPl+XH+OhvRVulXdZINOXySpAB
VC3Hs/B9o3LMT3knK3ilyu2S7CY7fwZAFgzdbGzA67BVeKY7o2boKyD45MMOBG0P5KA5KOxJi9Ps
LBPXgviO4p6r8aKsuIZorHffXPLy5Gu2zL2VKsOk7vz7zCuTffTp3I63d5P6F0MLiRU+raCXO8kc
EbnyOoqhbRB4Zft5QTv+I4JR6f7Xyr5/4e+dJz7WrqYP2gAdBp4RpP+zQeLV2BXtzBumSeciKkBA
7uPNSLxr3S/LOOKVuaUYOivq/YJnx4ipya82WNCw1CRV2GMpKCjiIKw0oU1qANVy/tWEevGsbea9
w74U5/cNiVYX/RDz4Cr1uO4fqRHXIrpFC2/CpasHHTGn7wKAdLF9gpx6/+H34ox8saTCpW3vQdVd
mGqivMACpY8TgHfwjQbkOoQpyQmGg47gAxX5ajfJGjCPw6JJlLb/IEaj1ixhOqnjT9engcGTWC9r
kJWnKe+mRW0T+upPS1iFXbhDl1cxA7BFJoaCVTtC9DbWNknYprW2934Y3K7xLDyap70naqmlZSse
EZcjO6+Tnbp/hYe4Pd5UnxMKz1/i5//6lAN0pvGb6JK5dR0oa8zo42FeiBqEdgf8QxzA65O2m2dH
MVfc0K81uS+uA8d6GVLDXEY8FlDivoEqqjuEV5tc1XX0uyUyNN+OrJO87TNchkV0q2xRYBxxVpe8
THV8mwHbp2Z3QyFBpJN5uPfRNEN9ByYEjmKO1wE39cpaHsCF5K+cTEkAvpGShQrK6nmBAZVEUmC/
OtnrDrjPSZUNJZ/yfIs980VesydSLhTG/UhbzzfplOGuXJETT5uJ82xZiAI+Zm9SQNXWQH38NeOe
Wbo+P7RBeoYzFKY0EO1KbCI78+ymRrf72P46g1je2p7ZxsLJt8sRupFyj/09qr+xfzvr+VZtlMFV
BjFxSmaSeOxc3cCBxambL0xhKPkqVuEGJU7z75jIFcyIrlYxudy03gEUNo4P3KnkAhYHTrdL51EM
o5BY0mNXLX/wR/g0uGdAd3KVq9e2HyGr3G9UU6Y7TD43uyBqONWu5GHGEka+Xx+s/Nwk0ljFC6/z
q8CfyOuJdUsRwXHkztZj+/jbi0VLWDTDptoSAEI2GEIxGv/Y28bZER3fIc9Z4cCPQJHbH1MfyTu1
ZzMDmPFHRBWYFEfG1R3dhZSVN9+ih/Pqc10ynKPv+QdB6GT4G372ibKHlST6JdzwMKGDW9HMDjiz
laYn3KEGQi1oA832TioJkkbNUFzYjNDBC5/OqY3KVChlpd4vJtWs04I5Fhne6xSEPLib0uIeRoJ7
RF/hIxD+ps9oQt8EXAxg0UR5U3yyZJVuAANpvFN4Vk7TxEzJfhWAtIFYMYmB0FEhoHB9XAdOtJP2
jbCBLYqq/agf9X6rxEiQf09WnOBTY4JPL/NO/6yrQMopMcmoi76xqi/z7umglzcAE4LJ0ph1L0ea
i+2b0UrEw4mU6Vp5EoC71SHUgsFiVUh/9wpCV7vMZK6xkQivFec0XJjG0OCBkwV5VI1EE8i4gWu1
sYgw0FKF/Q9QYe0mbTm8MJtIJv9921MFnXjiW7lGuBICqVMl68IeIg/eecnYnSmX9YvB6HRz7OYx
QJKeTzENSS297WZCgyFA9ltT8VECiJHmezip/9M0JUJbpyF7G9H4gY0ynn22A9UmNpkFuyFtDNd8
yw13wGvcekv1Yek5zyxlvTOmaKZ52tugZEJF/rEKQH3xrXWeoNc78oyw1psIFajIaTLR9wur8K+D
qCBjOMvBd928JEOsI/4LxEAgUas5sNebnKvvdwytwAxqknNr0epECCOd3kcuT6CikLpWtBpUnWlz
XIeCyQ0o2cDZ1PdOgBFhVYZvM29noC7cxPfALxYN6BBNe4VcF0fDVzjxOYB7DfAOxzbQGiTyysrW
08zeianI6B2IVr8Wk8d2FZSRMB2W9OMFHsokDHS+FB6JCNMkDrTZ7kvHJitXIm2bAoixOUHPbImS
zB1T97AmcbB+G2I4rsWZfAE3ZuV3VBGct2rJM6UBTbcKGsb6WyLRSzB70FH64x6L+T+92h7bvxHx
QO5P/spksT0gl5cKjtzLyiNSOah+tonPcQRV0xKWbtVs23PggePPNGQ6WBSN21GhcmXHLrVPP5ru
4yFD09YSM49E/sOTCCiUozuZxMNJDCNEeeVdUJYSm8Wr9jXLW+V0KsdMXrTVqEd1fyDOb7rJIlje
p1jN+WvrtzlApBwKmbyLaFvpIWlaTgSw/ETKWnW39EUXWvZmMxi0ynBq2bE3t3fB/dlZObTsh6nC
sM9kgMhfiSX6L0hB8hgzTA58T9YyFVRfOGiY99hrd0ynjKRKsfjABrHGaPO/jflioCGSscgAol5/
2YHG04GcvveWN3Z1vba4Dp/62eKLHJVEtSJ5kSVNqf64heYD47iqTCoTp28k+noxOFzbawupIra9
3utMfWJE7dmOV4op6dsa4XodcEmnN1LqajkH0u6Kx/00LLP+i3R8YnRyIi2OtVfyXBXin6IkG1PD
nF5umxaI9oiVUCOTprIngvTrYlhsIxP6nm15k2NiesTwlYVBl10crr1kH6zOHAt9Z14g3ONjnkt8
oCp2znOFA1qGS7AGVMTKBcO8RfSxCs/iFSkKb5JaF9yCPSwQ2LUeukf4AwpuLbNjUGuRDqdAADS8
o1LBn/SO8z76fsm7r6oic3xH0nMGzyLHi7KmKLyVrnmvVUlrI/0RPEmZOmq19mN1UwAKYcGrY98t
D2R2kglm4XeVDFdT8OHhEUz5M9WjDX845i03bbeak4S5QPzXVfTJWFagXXlon1aTT7E7PJOtHZXM
3Xla8W+Qf0h/5RcFmPnPa8ljP00rK+kvECkBjDSlbcrWmFqvNoVQMPDWK5mN8Y/UWTpacOUcqBBE
D5vGs520ysNJBCTILNhKf79Sk/n75TpJaSiST2pRONqhj8QAqe9Heb7HeU1kUZJxW7mz4PDcf9ia
NUwyj/Imu58pcBnXivsjPvp2SIKwtlS+FaO5JO8X84uZuYGGRchDLAUTwun4mkudTFV49s9l9UEa
W6qX7sZ5V47aEwdRcIPBxjpqGJ4Wx1z3Ya2WK0NWbNzGpEOqlg8oEeAByfhd9fowQ/53k/5c8sxg
mMjeF1/beOjqKB135ZdmdwuYdV4Ttb6OQA2/yx0vaLruFOoc+7juB/ftH1spV7fktIQ/T9PYDgqH
FZa4GGuQ6kFaKNN1ga8VckqwZaTQS9hs6DSNXcVqDUmywFrn7bl1RPLwDuCkaku9xndw+f41tTat
hwLN266Pog6pyrXao3fYlNXn1Wb/FG1XZA/urZUe0c0AC3h6+3/U+nhNZ96JsVRv7U9BltGy/tU4
NvmukVkS2j1Z9TAfAC9DEPYn4ijcCsXLnXLBOe2VF5wGOPDaJTBcjW4GIJhoZwttk71mAzAIwdbc
JBv6iX9x0D4D0kdnekojYCsPqDPIp2klY5F57xJ2rsHz0xKiYQJy/b9Rl3+dATPwKun0Fu7RrjkT
qNqjnSTbD54vHbMlkgmE6b8NR5Sf8hTxqEjr/mRvs6Ik78fa5pCj636us5frRboQX1FPo7R0WmR/
2zNL+CixXEn8X+WX+bohFFS5FIMFYLdSDqGonOKK9oncpREhamQTsPDEm2VpxtwtcNbXTva9uZcs
FrydcgK3cHxAKhmzhlncabcE6A/O46e3ufA5lkD1EXg+RSl5c3r3rJqX8rhAdVEP/r7SRsV9SWk0
/zzWc3vvfrg46epUKLkcBFBVUKY8e/TaznZKDG87vWo+rj4GyT5ePpjk46CI/Oq5hEMzLwHdHQyC
DvJWdelo6IjHh/d5MFPXcOcLvAYmkRAKro0DgmMAiuQpJd2zkfmhQtdZHPP7Y+GwsVt1DR++tJYL
nF/tBkWtwJPCuSFk19L0tTVp9OWZnygkk35V2A3YaFhDJkplv27YD3yWuonQZeB5g2xYuLmpDOkP
offbE3NZjkcIPlHAuadFbm8S/ObtFPHx6jnxw6jllSdyFxgI47r2thnLhFfWjhaZXsr56rbregLf
7mtqWiJ0zWQzzkVQMJL9qhWWPrB4bJq3JM5ShlEOx6Ls+6vuLilSFqADxiBjtbCmvwJk8H/Jb1ku
fj5V42aKHKDjPcaLgpSxwU6/Bf+Uw5qtlxA71iT/UqbXRurYfxmjwQk5c9yMOf3I7HE0cJqrpcCv
nahmqKjmGTpMn/s+tYo63OiJ61x3UZKRi4klouOEWMv0sSe/n/M8soSULzJy9X4V9KX9Qk9uGrR8
j+QsS7hc7MwlPAZvTsAq9OPkrD3qKzS8wsQXvzApCjq+4bIRY/jL7xjx7uGzkPXHDHuVua7Rilfz
Lh9v16scFzhy/54igaduQLYYAuSuDw7qFTD32pnpov0bLS/S4PFTpmeBnOhYoMzujTPPQKQ16jhD
AfHSbs9cHkbewZdXOuyoSawd11Xxe7bBtRWql1UtwV2Oz28YxQrwbPzpU/3qbf9hqC6dN1Hn2hzb
4p6oV/etVuZEhMZDDDgbVem2TlFAdGI7IZxRPSYO7qIYvR8Q7YaTymTShE0XHojNV/0rnGXwloEy
9CFIUDfWVqPQYl3FLwajSS6CzsYxb1vA9SRN1ZxhhWns8J9sFiPWcyd53vFdpmWkWFwOvlA1C2p8
QkKs5LBxiC2QMxQKfPBvrnKSrmhMdYd+G8YB2cv05+vMnklAK9LkvnFd3bUrruax/UW4RQS3/anB
eFjoXUgKoj96uSOC634ZRtxfnBQzBmfm39rjCv/vnPRrq++Qq3M+7smq9CyUXnlgO/RX3O8IDgHm
xft446Tr7rtwbGLaawLiP+Ossfwknebsl1Qt1fZGi9rCDrO48y/jeIlzCq94RViHZpaoI1v159eY
pj15g7EQccEm/PomoKb4pZd6AEMFCXbrEpwCVlzd2kBlng8497WZZhVFwUO1vj2K+Nfo4Hang+Ou
3vM1W5fs4UaUbItEoRCIQaMizc8ycLS/6SNqhxfMGC6HLCijSfGpjtvNHMWzvk+LYHZ35Q1q2PGU
bD1jYsBsOAEYBcJha4NAkFlkuK30g1k92cPAEA+4G7jNPKhh1ZKbUvUHCahrna1L+WI2Ip1uZIBZ
IVMx5xfNaZ8xzBbxAk6KYpDDbMLXRlLHhSe7uWj/yHU2AOF5e3Eph2Fp8eL2eLrF1wqZfFLRZp1Z
tY2N+UEIczhxWskGPCxGkPj0aRVAlQhcXYsc4r6jncLyQwKeArTjSOrDNyzRKFd51Lf82RHRPZXL
ZrMAf+neRxkp3xHMinH+C0YVNJZrTR/7UhOH4Uu1QIAGYaD/cQAoCQFzFsIggFS9aPqF0IMs74rV
21clWQh+DPt2+NhYUdUfsB4lDaUdULdZxO+xhewZoUsUeQ18YFvz6OkVXjtqWBwx6FACmaIktzbQ
5ZAKP8aveCKjHUfg0AJwAOELQxLtgblY0iZe5AQZW4Zsrl8dqJOwEGpASQaIRu2A19KLMuLsh7Wk
yL/p7ZuPAOgjm0XviNql5K9/FS/UcKefBJNouSXpETqSQgCfJEkSRfEhFAQuHnTnT85lmbqXX/vR
TrI8Gf1wuiRXiTCgJXt3vdUzUdcqjdYIY+7c/Kp6r0qCYheZQ0gwAj7ct6wIl+E5HHARXlHMMYxg
grmOlT0eodDOt5an3ySZHlioTgyP/5zXP3PxBr/QlUUIB/JxaWw/tl3Rlpp1JjLAG08BsK3TFe0u
4x4YKHoVyQHsqwmlJwsroLpke3Ngzswcqnbpf8wc6TDIpjRmprJcq4vbY7uAXARk2ILjDmpqLf89
0jR3snYPo8JrCjCAwJuQJBCfe2bYK7bJRJg88Q4uIiCUaV0sFamqFSrH4RSuvMhKKlle4R8xgEgf
tujXPJ+6AXM7MHIfuM7QCPQ5WfF0uc0R6kObfsGLg7VMfQnlJLTJSEGRdiQTomaLZjSO8D0tQt70
r3ZqOcS8C8oAsW0uXQaTR1y2TlL4BJ4ozd2MCdVesDEzDJZTIwhfso8KJPY7rFRUhJ5962PydaOL
uINiam8yg7V2bYWqY0Z5q7qNEQ8/ufGDOhazeJ5Uw62M6Q74GkOAgAzlaF2JLR6LnPuZ/j8YiL4j
G8mrMFki+2TZm/LIsC3TaEzSNSdMJ4RKS7zhRNfkOPchMA7PkvqXW6dOdrvQePdJBmXkQ4UqOBxN
Claoouf8dD1Rsh4PWxQMvlV4G8ivxtNEbi7UId/wsLMFNoDu0qQrhaWMVQgh+4rhy7/lYShH5pMy
gZEYfyVihn/nOqRRme322OLpUfeWFFjh2pwuxsrKCetSeSsJKQS8KLP5uMxsxP1r2ws96PYNmJMc
9QXsG5gmzYzSXv6aDRa3jSJq3+otGy3iztIMjCoi6c+OXoUAD5IvHnB59sYFTQjtzIKUE0kzUCWE
e1y4Xv5T00LypE3QCIycSx2PHdjq0UZgS+Ehh457pPARZQQDozCAc+DWL+gJgS2b6jWIOBCkySnD
slAvTbDfYe7HWCn19da2N/KYdNbfYQgmPdithrE78MRKHYOmNfOpyKL/YN0BoBy97YP+/Ul11cE3
c3hd/LssfuvPY3sCuVpK9gLxYfibgLRxxfdDEcVTxMLHWnaSfYVFDKGp1OKu+96Cu4+ngz0KFv4j
NPaE55MpcbcojtC8XWG08zubeVkMBJUrAgcvz6dSBQmrKK1wYwsu7kSNbiC//sBuTUpowcZe65xM
IYFPjKtF7Ve1MPtTFgG9R6sOg2cMZUj5V8YpMRfjwL5aB4cxKjPuSDF8YGQsRbDfAlH3Btcqk8lU
pKDFUxjhiAPkgoKt4tOzd13y28b4wANXjWVPbHKc2tLf/ChdX7scBKa1Adj3ivD7VDj8Sqo4Fvpo
YQE08OcjYCNI6UBJ3mpnbHx24pPp2vM8DRfBQiiRI2b4LAgsR5fqOwsylRs7hpOD2VHjh64qd4Xv
HpzmJk7UJTItYt3T1Ze/7TWW3cfi+RFUpa9RKc0RbVraGMNcx7p6PO96Cbk04FqNvp72EWoypR7e
5jWsrpi/HyzCo3xb9g0QfSspu6A37nmsf2t5blerf4Da3SihhKwkv9bFyOAcygvThJ2eZgHkroXF
106lChwSGuL9CPxYEo4bV+e4PbAo15lSviHopqqOxvulr6AQ1IkXc+eGhfun8U/Z9ic2lYuNPArz
il4aOgcFZC+zf5rGbS2aIKVrefS+H07U6eFbAU/aT2VezMjymSKZbpkPiw0chnIdghJ9cQEORo7r
vRx230uX7guuCrH6oHwdRmIZYmVmkcxljcnNDN9bJqk3/6XWh75/03kn/4zkJ3i3Q1fD4AYsQgar
8bwEAQzzfsLrUbLu0djLt/tuhV1PuoiUs75GyGLy4/eMMQ6d1dw0W+xO42LgwD0GaFIiiywuD6VF
jauihQPNbWifmkzvlMSJ5pDIgLHIRHue0crAyB304RC9j2aOhT+V2SRR4WQEx1pPA10If6VjZDjv
lEyYNQb8HwYOTIpNPQNBgSDjmEAsiv3iNBxl8PxGZ/quu9esR/YRYuLKnXSv0wkY6JyxNXOGrbMC
aK21YlZjTXcewbb7PfcrBXQ54mxwQGwlnFAEhK1zqlHe0t+bYBVhGY3p2Kk8iLKrp6xuqRoPxT+k
dkpl5aF2+S0Ee0AvcQTztiPB+E36IBBzZ+TNGgo6bAWj553SJA3eAYYsXpH23P4BN6KKAjTSXce1
XwuiCJqnAg/f1acs2sKX6cyCEaH9CtjlFYkvHw31IOX2fV7j/tZXvtj2XGA4c+A+u8qEK8ZRJ91I
GoMpJwoEkL7CF4K0Erm4s0vrYfIvlz6//3NCuCeBw+tkYE6SwFYO1LyfOTuZHXE0BvoPcQQ4prME
DCYNDARIxahVnctp5CEmOykzG01J5izdpzjjL24S5+5GE44lZGaxazL+qFmZ5ZFxN5IFEuqgXZaK
k5dAkS2vHTmM9KoVXkqzZs83GnOt75jMvn+m/slBtHyiekpi0CWN3TYGoqlkMmspi6vGxlMRISAN
WAW7A/THWRPtla9rDKb0JVfx7rs3zF1n2+2ZXYdo0GUj07LU9fNwrABVSnwEeGXA1vFrerG60YnA
oAnYullKrWSZCBbt0CyEKu8i5+sdVi3W3iVvmEizldZ0EHQRmZF5Q1O15uRm8clrvqQGZfS+5hQh
OelBRGyjqtx3pDkO7KY4wlYOPCMaTleuFTMjXfvp8ziU46oZiLMsDHsR/MnKefA3SksYM3cRr6lC
StfRJ6dw0dOKKjxlMtAz88s3GPqzwy4oMMFUYqB8ZcjLP41bzxMWzdOqW5GVXW+YHs6cgBpAWJo5
X0oFwog0XES9BdUIAMIpP3TY15H+MLqgSLpRmSRB4NpDirAlP1MmsK1poQlC3s0Pl1l4PZYfdeBH
1klVkAmykQcq7gLQ6DMyJdjTr/FCDzWL+q/DAjFYXCMlAvgbAJzbxOiWuyNgPqbYeqmbVUDAOH+o
DWPoX3m9EIqczi6LYLlvR2cVd+Hxd6243z84U03ZXb6l8vX7tLDTr2qWs1sga2GhS2bkJSLq0iUS
NcmltXQ7gPMeneB42ktZniGqYqhQMV1TO4k41S9QhoYpRlngKIlZM06/65dWZwH/KsiF15GLdMrF
i+QvI1LQNt/FfNl84OwQfFGQb8HyrIBf1mMGI4qu0/M/sqh2h4OLQ3Cpyu2zwp3f8rjVAXWYMaNg
8qxJCI27nrujvjo3UTb11/yhXb8cwj8FwqOvpO9tzqXOiGoOFAxsag4jFtCDebRpohuF+whKYhm6
QxMQDBSVkvSBg5xPMfsRXXMGAAqSWBBSeOwmhw0hnluEu80rj/hCZrcH8P1YZqmqoXf3objFxRr4
gevDo6aSutPMbgW500bmZMtI2kzSzZ5qlZnFE+M+Cth831tDoAM4K2To0e50W0UuMPO2wDbpKVXz
OYVoVNpUv8wn85yrbC907hV0X4dUEB7I+5mx0IknFUMwpbTZ2PBmpQtxQ4foW6RgDlDH4/86g4XF
j4djeBblDv8Dwfl5uYlQsOI3Zg/t2DwIlQ/PxbnE70muYXS1M7Nl3Pyn0yxbWINZmL+kxjmdtA2r
F7rmZxJZhEBwpqDdZmP/Sy47K7pqdwKuCUpWluNNPMZx+9fkJPr8MAG/pKI68bKkpHCwjg7PKqE3
PHch6evHe2dTRLhpUW0y9Fj+qdN3O4Ao5MqZx43U63WBEvYGARPXJ/n9UTs8cxWt45LEqzEu/bLc
fVSPMAHs87XkSy/Qz1MdTVUFhBzCiEZ5gexq+COMXY0x8ZeUYuZpY+NJdMKKjAu1avgOQatyGO0y
b7GCWq3Yx3yHcf0Q3UPGuDx4o+wxhlhTjsBzR3T7OssUSVL8GANRH859Ac22ta+9BIpjUMTrhODs
wMuyL+EazuJTCNX2wbH0MmRx2Fp1SSP6PBhrSbWA8wQQWrIuJpOkqaF/MFNUlvXhUmmuOaXbc35C
wm6ju+pZwKG7HdvRdlREgo5tu/+uiibGaYBrePbbVweEtbVNHlF4onFaf4lbwlnShWirgA3KY/rT
jlk+/3qx4XR0kAvZlN/YpTiHhVbW6WuUkKsD7RNwMeFsAS+1Qt0IeClJl8CRJVC0xbpHpoOPVia/
GJg+xgmYNz1AzP6p61w4lqaN1BAMm3Hco9g2eZWH3ddlij+2pcy6cTff8+gvDj7Vwdc9FBwHMVIC
nKsyXqV/hxzCvL1KkevTfiMoHcCkBlM2ui/MDsCRjCDMqkHj+fM9vKzUUMANYFqQV/YcCXNEe85m
HFMdmltJA+kpmXPw1gWW57ZcuNMjxnDT5a4vI0Wy2GQqAEONhTZpLGGMx4blY74FKkvMeex49wSi
wKPChSJi9tU/KNLMkIZiUXmwGUoMqwDkwWDzCine+NGY4nwVJLF7+hup2Lwua3Qfm3C5h/+wLVUy
I8lVlOkOQnxl5NKPKl4B+uEdOSEuxqqBVqxP44JAvwA623AVQGXRWzHBoyipIJxyO0W/JgjJbAeF
k3nhZbxMmwd4rtMFBvyXbdUOQeFIdX9M0GgTWcBKMqEc0rDCto435gZ9y2QaX71oBfImFAEAWfDB
jFI7GvSuMJnpiW7S1eJN8rcCVGPSNPTxbJ8rl3oSS7JG0Srni73Bk9/hH9OUqLycIYU2isrKr/20
J7oVbenW4lAObVNJ5ZjZ6DhJUgXMZesXcLEXAo/gwTdzuYOIIrUUiI3kMuBUMXaqyEyn0e1KQI9G
cPDqUHjf5WPCNosQ5z7TwD/8ipGpc39hFofQve56ln9TrABzRR6ziUzrP3ew6CEUDCM6QdDayJ+W
QC36yzPAR/xPz+0LO0IpoEjBc3/RkaAhtIdC0D10RGIUK17VKXGJ+u2DSrcsTI5OdB1S5hVVgeOL
YnNGhV8ceQRlQNbLHAOgBgtnUbMdOE26fLthPiw95ybuf4O0f0rhwkF5Wu61XVavFz8OiFj4EJvO
NM0Wv0nSju9rUxEyG3OuBgfyNt30FJOBztjD7N1Qj3irQbvrYUv26hZcw2WT4VFymvNoEdOht5rO
5lgZppV1irlWdelZIijGO5twALOsCvgSYHoDb1qQuTUnP3zzcj8pxC/Hj3Hi5ZiVzRFJoNDOrqDh
Clhwc7yYhIaCJ1uel0XYnqI6ZuFzAmXelNjC9B7v1U03AZzSjyBmjWKgfCw85N+YCyMB5wR4Gjwr
690UCtaIRIszC7uiamEi023bpHjwmkjlk4TajfFSh8vGa41pYwBKpdWrc657gJQ/RyzEAHa6gy0Z
neAM3ejeHl7BGDUGD/vZh0oZrwW3NzLTrMoGIf41ILcW7sUMu/4GZ1BnJjQ4nSCdMbrGpOY4N5lU
XLSIY+mYoI0OZInO5w77LEgwnII5g1wIx/u0BbjvRmQaXxprABeTfq6ScF/lkQYC8EGhIAGA7TPv
w6VPlM/3UyoQSKQltOmpATRXK19ldAYlNGM3pYeTWWIzIYE0yPCSq10nLb6a3hjq0z8Z480J8jb1
JaboD4eunccdPbtreJ5rE/RMvy2mzkkFnLfgSTRRlz8n2xzJqvawT48Qh6LffUnS5NZMo1KPh1Rp
06iHcJ7bBlW32CbiOIqouVX8Q+82grICL/MIukOqUdgRW06o5At6GtehbpELKojxnu1Lf8B+8XiA
KfjR1zv2z5Kct7nTMsZI4boWvLJd4Za/Ou7wfv0ChavnhnsoXT7IjOHwbYn8I6dePsNGKPsZhhqa
V70oOC07kKa8ceEivi74mIkRhu32x0tAZGR+Q5NliVarjHmMbeD0jKsEvtEStujc36el4Q/81JXh
8uuxXNZ+0iYMfzZ3+7i72vwuIAT7+Y35TfAwZGmwu6MIYgwLEm18+o0id0Gd6aRJvj2Fi945CVIc
kefs8uExRSeUBBtE0xYjovj+XOr1zpAJLIFcafi2MzPsQZW1U6RWoUVtznV2HDTgVSLOY88002CG
qFovZbR5OeMQPFgeNEGms0DNFadE/h0Rvz4gE75UfOs+hHlVB7mtXsVXBEHZrx41zWxKdBa++R0i
7pcxWyADkQEBz8pzYaeCif104gC6vUWFUe2UWREr1c7J5vWRawVjC1BggNnymv3yzVVdxOCVKaLM
ynH1xXd7DJZislktgK0v7yZf3CJxGLvsbtQRShaohs7VWjjXgSDD9Y/IOhx2d9Qqc2mz2FC+SS7G
157+lP96L113BSZFbdPwR3K92kLPV6mHzPPuFuW0sLldCuOxxQ3Y1KQVgTDurtyIT6z22WwSdDnI
DSfPTtFBdORmg6aicCgDjGpsMy8rmR7ADfHyjpURiwb5Est6M/qyv7PBNoziJEXDjPBoJAMlg558
d7VvaQNzIQdmOhiu3/XIkRkeiboCNfXBBKIW3nQHgId6YwkxvlarQrScR2AO/uTSpzqD2Zv1ZleS
frf7nqZxASiDUBoDu23WoN1ClGylFcnPEQ8cLlWM4i1GWrBzv+xthWqG1jg/DA4omFY0JEywDXVT
smE0ufYOXOn7zLhj6R8Kx1DenWU+dD/S1oK2r+TImF3wH5+SFlRuEVIA6scQjxyR8TINyM09ftNy
HEUuKWuIE/ioZjtI+lNa6AmHrj+ni5ax9f5FAtxNjoQJWgGml5IPcwBnJPPKv3seY/r9L9v3fk5R
I5s+jR8v3dWhNnawAVCEEy5SelZ1ScP0BA0jcl3CB4a1tpVzGHNN0TEpu5ltER0jNi9MvHHxWuUv
7JixxkOPrNo7dGb34tAQQIWtiNs+dMV9M1QRb6xi6kD37N0IwbtUfFkvazjCEHx+xMbEuTHcD6if
G2SM1IM2LDzvscqhEZOuiBoWH/KFFkgiuFglXi+YByfC006z6w54pZNG/Wa2jG2bnE3xNZMey94s
66xBQ9/g1a1cngUM+N1Jtrwa7e+6m2MUksl+JdmD8qmaJnnnwdHYrb2XPlK7B/vGfGF6Pg00qWir
lUGIGxRjRtC270dcQvumtXP+y/cml1v6qrmEDn5xGpzVT+8O8deqUP2JSnUl5bFMkhU06+BFgCsL
9NRWOey7rtk7msyXZpOXtYUHxYE/45R+rG70vIHi1PX1dnWVufmpeyYI22R/L1qvTTHHcdSCCM+0
wcRHFVp3hh7LkhiqkyXZ4TYJedUbNdsT9kg4TrQI+OkdHEcj19n1aCyORlPdVCl8KIXtJ3nu4QOu
BRQ5oUVIVDkL6epr9RGrYHywgkUpK6tDlHyRSMGAVf1C7+JgPX3klcFRZw+uFfkdqmNW8LWr7A1h
x5priTq08HbhlV5FSS3DmAUwcCmXUib4oMtVhXu0a8yYEfUOfsba5/6dWrjxgvkWKEWyPvAFr270
qAR/Joc1sfTzPtzd67fXp+34nXy/6ZC7kpgLXvNWladsDg/WptBcRwZKPyLa0feDgOq2mFYdEDsd
fGPWydQ0ClpmkevcvAqDAbcndS7IBrvUSQlDXOa8VSZO41iRsmydBcKlX/4l0VBfG42JuldErI5k
DoEZZ1U1q0Wu9qqb+Q9Hfz4cPcU7TMQ1ZXR7Bjv6i0400cbz9V+9fEWaNWR0YGY6DWO5eJJYk/TB
doR9UnRzfoeGK6MRRyclzcJrCIjVNGHHobb9wggu1wtHVaPtKMjK3uGuFrJfcZqs4n4CPvZnXL94
QQ/san17yDWsnFjnqAzi/xdwDIJc1nIzT0XxyMldny6sIvE20tVjONIzGd4YcEhlOm5sSF18pCWs
VoeBv8OvcgqiUwvCGL6yDOcGzsIiT/QVHR9WVmkL2mCr7RVwz1pJOWwCOVFzlMiTh+QLL5CAwCF5
IZVJVmeu6Qd+UkS9lpSWFLvwlze3+U7RkO3boz8oGfvwJdcyb4m43R8z5RXddXiiuldKoJObyfGR
fdafSPGDd+UW8VtXps0Dag5Oda0l77ONRHvBPczPEisQp8NdiD+3oTVynZWVcOaYc4ndudzQKjjK
N/4td5hpSj+zS7fn/K9qxoqBktMj9aZ+JzCF3VfHGiUs7X54LI7LbuXcZS40LuDXWXTQqTaxoDsI
o/jKb3pEA4te6DaQoPTa9eH9vp8qFy4sF3ktHWAMYZ+zKl1yLbE01MLblmyxYbe5l2SA708/yb4F
4F3sz4IoLyy2ZPVLdjKodXOEkyBC/3jghj1mJiJtwoX3wJZFPmHCwIYp4YF8c1+PKdb4TBI+gdKp
HRSFAQcCWI9UmtGtoghISg4Fg39ifX9WKjgFe1Q9MtBuVEcpFwfwO2ik4m+LG3Exs7XdBFCLstr7
NmDqgLXdaKvTZSk4Bkfbg4QY7fTt6MbQyK4yjOBo/GySfENhLjU4bl8qPc/SFbqzdtq9FcP/5C1i
RM11E7u8BxfA76citJwU2wKQfnJn8VMo2lRpfwR7AljZacqrLMANh1jHJhhVf4Jd7e0VSFNQfIaJ
O0ngZTLRmN14EAbCo1ZFr4NgXqF0PVhBemSLsRqQtxXHIDxJoZu9AJesyAhIT4UobRu4284UmFpk
KvKW2oogUz9hwO7CL3yj+SRkOj3mvE+qtzp6u0DjxXcR+aQ8vq89aBqkzU04gvZmnKrGVzrKR7kG
7FFus5unaQPFOf9tOGC2v2EXbM6SKvKzgyYuQaiOrb0DiaRucYYxKEFXAeMDRtnClJNw9avGFmOO
B+Ru4QJMzE7GD0tIbrwLVDCF5lgTJXyc3JeiS6UL/P+F63YYeUT1f2Ca2jvEqnebwkqhuL3S9zg7
EIgYAouUiB7RYLflDW/uOQoWyoZXrkSIUNmBw7ffbpIVnj4lOPAeCjLFFccUVqCvOksojw16vz1o
2LOzJvIX1iDtpabhiYOkZvreGyF1d+TPj++zMswLfZcNL/xpHOll97bk3JNXKxykrhu5dZ6n70vT
nNnTyJlqfdBhcLsRQjqJpYw0tC7zrvm+ao7B1Y8s4mGNcxs34qOcxuE2qMzqhlR00u2gIXHU8v41
oon2GKfwMDi/GMQR/+u3lKFbiifWBjrYJN66WaQ4r0vWcLgyUbxj2XIcja27iLsXOw5gTi8Z3GpX
YQgJY8KnwqMBwg5NmdAWLVyoWMCkQIPWcBWo5mVe1twcSok+/aX+7dNiu08PSNuGiQmgyg2MP0wV
kcE5eHrcd1a3WFtg4xBUtUVEIt3yYogFijNX9uY8+Q1QlioGmgMcVp+WjyHwOxTE8AWdcePu13aX
b8h0+8/m9qVCLsnSFHtTsFxFptqUWEcId4geENtVcO/NnUsX15VWUURlNIPgPCz5c0c6UJcyYmj0
MIUd6IMGgRhB5B/RVS8GzXY5Ea0VMtMu3OjUxWeFSZ73yRv38bF/BZajrLH7iEB7MCtX3uBfIHPW
GqDa5sj6xGJ4cgiHdgChRK6pOHQ12IDduhEdDI71tVEvFqQJnr66/M717QN69WcE9w19o/zI8z1i
zYX1+ysEwJjtCyFRC0gpio2PfOa65ZzLSj403t7Kj4lmxipVVc8G+oS0PXPwzYbnW7aeXlkydgGB
xZ/592u6cCikOonflQHZKI23PQnYxXgJZOUKZI/VXlyCCU3iO9VedzIlYynmONA4vrOhoGV/6gG3
9mMJNrIVfajKknkawfFYobrB5qNUium9YTx2apcL/z7yUVHDaW4GuTa0NGDZnxKYznZOw2LjBvML
sH+WbgA55sOZmSBgg0bavxmTxKMvLsf4BbgEow8cAzE4IXdFOupAOHl8C9hUl7ylHoNzcoI5gw/h
xoeEJ/L3kwstSrteV+yTc5/hUfBoed1t146HCO8NNh+9IpC9vIr/4Moj1/6+2oxNZTnMAR/0FVJB
BGu9SucqMoRuqaeNp9CqV2FQ1k/Z59xfUIjDAGZSKTlcfRjTN1hNORrVvKz5IsaEnxpGNDAHTgNq
blrQI6dLDOeZPThImyPaG8O9ipKKmmB3NmMfZXN7M0PSeSVIsxcS2z7QVhXcTbA6lJv2dL8LbMge
9jaNWGcM83JVEf/dvO1txyLTnkC+gNFto/psXdZB1wG1Y9m4yNffi0h0N+WbOUgQaM3md/XRQyqb
WlYpywFHkqgZFtyvnhdpOcz0BDAuF7dbSwu4ZmYa5Jdu5ILoZRtzSVna4vWvf+HVu361vblW2q+4
JurVFG4FB3Fgc5UB4+obObtX+6sa8GF+fr9kpoylDnRhU1T8z6wJLF9adBweFlXSJshWpbYtPNgJ
ptOyDhVMOObnRsu67AClXzE9OL2owwPDywe+A2rrl6E8zwNgd9/SalpBq4X5+3xXAG9qNqQtOp+C
+e5/FXUmoC4yF6rExDO9iQbDmcl+4LPxLbOPkEidhEGp89MND8xwZuDrf7WCURxQaB69wyeb7Xpi
yK0O4W0FhbcTNxqaQnJooh6z3MSEkaJbcUGn5COmR+tBkkJu+hwPEvM1JzSAPXCbzuD1/ZkTe7TC
KviEXraoSbXdg5ByOyx70YKBC0cRV9rP046Se9fV5TV5PPwTesfReQJ6Xtok9YgogELT/5cetz1o
K2cWHUHAuw42MVkqalHgP4XiYbqQI69dtQ2f1dro3zu0M74iXSD4rFP8ZJPlIKk5vS8NnTcSxu/j
vYmZNFQiTkApNhirv9p3TJwHqA1J/BvbczXYh5Cad5UKYVOM+T1Fuwjk9HugOyv6miOjRvtvB5NQ
P/7rg6394cMvuPe5yWBRBmss/Owfzg7zHeSoBGllie4Rpfzza96WFgzzd6BOIJoYTa2UKV6jDbTg
xlof/7blm9oFcrsn78vAK14y8ydrCiPX8GMnnHwERXi+hgTfnHAuKOHU90HF2m3HWg2Ekd/j9Qe3
96YjlDiQl39inUrPwmQBNJgjgpCFuYyGYLCp+ET5U+EuieFIR+nVKQjrdZo2TuuXn8qGcP+0yNSU
6/qlfbrffr7w/xVz7kf/+ykHI/q7Nvatacoz3P01N55xrVXW5vwVDeo1tFb+Jq/iDPomfRyGROZU
GTj1EV1KkgaM/glHB1dWn/gDVq8sg7GyuApCdJgfuxGN679zQc9qlFIMscG1+jHeQTBdyBxiBcZw
HkAc4HImlgAMbPr5X6wUC8ivg8tNPnh1SbPhaA3zZwC3HAWh+5r7pTma+bK/Hifh7TAPPFEziJBv
CWnLn8xM0iulfUSrZQnVahJDYS61KDNZBIQ0/DMbxfMXKXIqb1z0O9d6PWlux4rWkXZkB86gL/bd
wpdh17PPaxLLOhJP4TEHav/Ht/6KZzPwujitxjyxUcC9Zfe3havdhydOM/8xfYO10I7a1uL8GADn
K+nNl59j6L03t+cqFTQ51mZtP1AU5OMRq+6FDTZ6IisVj4a/G7cYwmJM1d0dwfbyeuwaq9gCBxWt
u+qnc3EzHcYWwYfEQ1f7g9zNA4kJzUuF4JR2vilvcu9CNjLhOG5JKSDwNFOGXmK/xq9meFtpEIZ2
ed4xNCgK3bZXiIqwZJl8owr0QU1cuPDjGNx4UzxO+CWMm1dlRfTFDuuRtjNMp399J/j9knLXpuFR
LECz8Yt7MFPY8Y9P8ExwQ2GQPcQ84ZnLhLC4knZHiI9PwjdofiK3LSHQIEBNHkN7A/OMPGXD7XQp
o5VK5mbXP84rtIvcxoDDbbbZO9g7Edf1fSFTc1/RJzhpDRaf17fbIi9IhAGqi5hUbW9xCxpcsoQm
GhCkARUOIVAO5Ny7SxMlexkptr+SL2gm14rmcdiEf4zSYXvwla1NYR1rhiW8iSYfYKM8hPlaL23n
DWYOUsnxzBAqugq6/xUVt5nBXJSTnRPD8Ep0aWIByZWeUSBISea8CsY//LnrtALfi/zTkO3F/haZ
PO3duHCQi+8Qy05QS2XZCjemlCaix2ntD8gG9YvjN04yRo8mdrNAgf5wbEyQ46YLc8fvrLXNWfW3
UnnYglcbLJYPbAtOUc9uXtcDP+qWGQ/G5OlnkpMk07/mFehxeAIJRS4M+CXPqKvVPp+8UF9psz1m
tokFLoJFh8WSdMVoQgi1AaJ+/1vHWNnZbgk84ULKRLARECAgwxBHxlN8EeI4YW43Xx1QvZaEFwKb
A4d2AidGTOk7iLjXZg7Y83xTt10F0bTxRZAC4PKBmRoNwyWo3o50Mot1jSuZA+we/EmwZGOTBzfz
yC8fLe0Va1A9plJUOSQc5HXCUYlvpb5j65ne8/aGAYB+wqyOxxllQ/NK2xHCvUZ5uvuM3OaSJRHs
j3og3LtU8gW9PSvUGcMjYiXKpHk+c7v0UOz/M4QdHcaOUgstRinwxH2+mTU9jw+4abhvdllb9p2L
sOI41B/4KpRjmEaK1hgCesFxa0//NvTcf6dcNuyHvc2DAd0ScKEdjk+EN+q0W2Rip2IpeT4VE67k
5R6WXyMy2mI+wHmFEroZlIvS5dpj8HospFuwZkyw+aWsYLGUxT81vQZYHJ55D/KH+exAaIxAR69h
T0HYe3Q+PcVM2KBxb6y40ptTne7HWOt7vlM3hzFBk8z9pZX1CvrXfF0Op4zUHI8yIhB8xfM4BKJt
aCZQcBAFxJlM6MFx58069MuvsgWA+/BENPLuSLihzHkfqksRzp5byITSsissjpmLYMbGl+wflur/
dpmPsq9PQHLR+/V8nuT3tLyY00F0hmFDSE4uUxkM1oXqX0Z5U8HpjCX6X3u2PooFJH9oJYzUFQ+6
QBlIq8SDSiBIqwQtZ8sF5MQK6BgS8yADP+QOCVv7cGbn1zDp9Xu30YCbSIvm88E2A5zbY4bIaXq5
LmaZMDwau47l3AOgc7u+/BsLPIb8L8m3CZB8wX3cTlFSEt7sax1A1s0OIQI/Bnjrn2+Ib7qLKxct
80lnpYEwWRDgMPO5qyP4p0A4pqgB9piAWgjMmq9oZQTLB3+iFrKTLZhb0CXzZnfOm66PSYhN65A3
8i7PwGQB+Vh9YRfnyvx1FIApGbIm4hVvxVPKzEo6aq3/zlpOsKQrFTpDOPkQMJ+Zsx6fGZvuW9OM
tSJngSwHdiEOTtJmzwMrfi1PEo3xoDR92rNQpNa4F4vKG+FyHQdIZ8g4beu4vK5gGuF8Y+92VcC5
TU6xxiEmS4rg82SFR+S/owsoj6HoeuLBvrMGzqwtX3rXHiinM8lsRsDNY15YVi2LzdBevLk4EJUv
KMeSZQzv7J/QrSvivaUDOOUqo7cQMm1XXYMRUY6eF1G1Ekbx3OBkxVPzCQtDZPhLjP/vEUMyUJud
Pg/mKOxnERLWkY+Ff8WymHuJJP2bBffT25RyTCCECLkrsG6RdrWxgItYnrju7OYTzqaELV+zfmX9
mfgDonfhuso/au/0UmA+g/fMUkbOgTq7LX0CTCdWTN2eJ3ocySxp0aU55ATb4KSXcB+9lIKiH01b
SXutKsGotHnUK22EtchstUcQ8mxpCrK4sluOXdj9n8+4EbSsbIIycECxg1OeKnlZJUPtjz+ucg3O
9kf9K/Kv50Yz4y4+g7Bo4xo0zhJwSDFasK9Y4q6tb6MfGAAZxVcNyzR82GNnVLY2rGy6nsk8+etu
NrYi8qpgv6RJJpdhspTEd++brcIUJnY2AoxiCk9qV6VjA3XRFMwWpJzJu0zy4HtTVjAulUp98tLk
fsSeFPfsrmbpXwrEWQKsp74VMd2y0V39DsIUmJ5UntnYK4sd8NzbK3Hkv8wpwaQJD8wMHSeqZkjc
8WWtwEpdi13eebNqTbRbrrzHqP7nzq5MBw+opoYaNqdjBgGHpl92Ky02/BCc6fk5RM9oqeEb8A0x
Zisx42qJEzRqMRh1ppVNvGh9edpXC9TS7Py66oZmKkGqd2JMzbgSbuF3eonfnqi3vLj9Vyrfb0p2
1qTcxrmYBUAQtDk0fQZU+fSpZ+fLFrIDkpBgHAOOklWktVKAQHvVIOUsseEWpvlt6NIGnQEQIXil
ZKmCz+ogFeVZK0fbOtVAQs3B3qB+44arSRohpH6RmF6rLFqXFzpNE9ctGsvkN+KwGmfzQrIiaEJQ
In9I4JKo9J4saDVvlKCDKI9Qiuj0W5lu0zAkwjx0ebEgUUfRHiW4RQHiH+8c1D8sQf0pxpX9jTPE
V5VT9qp88n1I66mMiUwtR1gc6h8CQmniiN9dnIYIm8A6lWiQRhW8+gR+v10cjajUDShwTNuVl1r0
+wmfdNsbHW9aJCv5J2/P5sWatYd9ymJ9MoAlWoGz47shvOjpkPOxTVzTDrrdaWPS8pLRm4o9cz4m
bJtLFobj9VyRQsZfyWJPkZgQreJtXE8OqXSB90w5LH0m3rSgZJ/7OsrKQ4f4FlJsCzUxv4Xyj6Ko
m0WS/ND7K7kk7DckUkjoWfXzGAEi+oAZR8bwLDqFtOaRc1tc8557XQS80kk268t/NqIkn9b4gv8e
SxL/G9pfeTQs7aFs3rIRa7/vfzDcBnGo139MkW5PKzENuHt4IXHYXl1MWagZ9wL/AaCLKMVXIzh/
YHZKDulVnpA9xWUYZMHmPgwghzVfhRLgvPLg/Lzx8IzJSgQZZOblix4mYlDG2TffOc+5VM7JaQgU
hbBwNgxk8x4eMdNQrO7cR06s1h1DbpbDQ2rI8lTdd4A8MBmz58wHSQuHtO1O71VQo+9FW30J6T6m
mOeSocCOzy5H+JGxkpBrEH8oHLdF2a0HttpCUiDM+WDYGz9Fobk02o1ihYXRpe0poOLrjWx9Lp6f
IbblZBjEhTeIc1IR/sF7EAVxA5rnUYMhgOfq59aqnCAPs4dXHABLmQpDL17Ha3uNyDmCE7k7Eg8b
XtVN0jGYKY1gbAsQxPbnZPgcTw2VL4WIBTxutv78OB4q57r7QgOX29z2/DQ2kKcmOW1UC78L9hmy
Vn77cvtrUyJhpvjIENrUjszdy2AoqBzn9NwdM/cdR1l80ujRmIzczdgx38rIFEe8ovVBRc4Hu2ik
qXw3b4wfKQXfbS4lSLUp2hgJJLRG073lgB/bW5iECXSlAl0q+Yne0d5mKKk20OpEiR3ssqE/jY3r
HkAZwE3NI1BLgXK5IGc/+7f6cDMRvqTpfjwNwoBWuykhzGpZYRfUU+mHqWMpkacGie/Cnuaab2WB
wl/xQkFVClBdYEyDB8XpF0OT91VL/6jq5jQ2ZHBICPgO1DKisPdMgLK2bOkwMCTFCWnLXFXVjnh8
sBzfoNa6MhxPNdKh/ZwOnk2bLcat+En7tRmnv6pRm0q2Yso7ps0YrVWh1WJPMYq1LqafhZcWOdbb
j1soX0qCTxxowmxS9AmykF2/QCutwsU/b6rRzxDdHWqC5q7b7v2gXCn+/WYIiXV0kSwN0WzUeTtZ
MzcD73wXB4i83OWVNhjZdFBlAYmEeIXugigUEBA7QHwYuaHWEjUWuQKHqXw54cz6zztGwpoARB07
K+h0Zf/q203L+mAivFV9ItfaCOQhUSl39Vx7g6PSGhtyWymBF1F5rMmDe2CsH6Vi1P8imN0Tlnr2
TcdTB2VXVOHCk0VliW1L81rw/MCwj+c0yAUC6AqXH/dERimHucvb3ss6bzYbXUK0vrJ7M7DkCdLf
bTBAyXfjcJdNX467zqZwH4XfRWEalAWQ3HxjLR1CNYUlwsjtP7RLpE6rFHag1gB+pM9ORJl80rg7
v4DnXzPX3evhJfgwSn/FIRpxv5oaSQiD5YLRv20RY35joWPxedyiYRuEgp7RQsfN5bAes9paii0c
HNWzJs+n8xezO8p5dgwXfx6XNiFT3/abhhzPejD3YSDWzTJPlr1lCmdbA0bHpbQCE/YFw1I12XPX
sGQuPGaiRHoMqRyjxnRxcFH3tiIc87WmRo6dd99aTCW0sNLlliKy70C10rU8f/X+mycsveoONsRB
a2wNM++/2EsG4OV7xXpCts7sjUBTZgsDPoMuMCwhwaROCwdluXpolL0mVfsocP6CnXlWOey6of9S
lIh0322OWnXiiGj0TkE7lETP1sISjUpFfQ71e9WWSDoT1835JSnF0cdRb4H6G417FzNJlCFBKCbU
/gkxg+tbsrqCBG9RMIcF8iZWD+x9G+U3RsyJHPOqAiIXOLlYKXMtMRb3efeRlACJFjX4x/c5XBYB
52HdUlh6SAIS2KfrjTfmSyPx+9VUY4rrwyTyCaM2CfBsNuU+uSg5TG+vJP77QoWW4PY3oEYvtqA1
MUd/r2cSXGGCiaQKDNY1Wrt25gBUjdTFi37xpvuXoqGBubSwg87zQsosZX7vBln8/xJ4qKU88Jzl
wtjopysr2CUjgGPEyMHPN5S8YE6GwZDANuEZN4Efo2SXuYnzNAAkqEgLAVe/MuNICMj1ihnGb3kN
HAYVWRYBUVJ194ltj3l+AyhxStc0LSRITQo5BzOqCzf6vF6EdQU6Y6qm0eGxK3aqOdmlUb2Jjidk
0kvEJNn7IwryXPyRWjdupvtNlX5TpoiGSupXF57jYK+sSIqgF2BjnU1bZ7h0TH0QRdrjG7BSgI7v
yR9Qa8ZsH7RrDJO4Z5YkHi6oVjk/kmF9YmV6ReSZbnpjWatXKztD0kYtSKzX8GeiylRSJs7PZCi4
MBp7B9wQ6mhukhBSBqjX7DOz6XCn1JIYTJbo6euh9BCA7RLE4R94F47D1TQOcs7aYPuhX4Wz0t5F
8SHtQPx/Twr42ltIdwY8gfpO25fP2qx3AjbwA2rTBaFUW4XMQAT9tmUr3cWfbpcan6lVh41ZekCY
DGtCjUUpSmg5WWw2S4aru1bv7M+FceqK9TTwZhZgtl2AdzNX1++TB+me4st9wgpDH0fqYS9B14QK
ACVdATjE1agdBULeyzLhv0LEWuKyxN5Hf9qaNgtnZhlEpTiZMp8jpwJTZczD3VKBKAhOlwwXFrDd
xsnnNuoRBONhrkqpcIaN8iCzZgQ6gGn2usJCkw6VHZbUw3TomPXSiz3gv0RxZ3qkdkWYwsSei5Wg
u+7jgRK9R4FgZjo3qwlw16OGbU52N//e/8QmH1H0MCjtkhqdG3u5oICC2Ybg1pXNXUjq8/CrV61x
SyFb7F3e83rlA03r76RItJu9I8BfZg2EdwL2tay09cEGgAvXAJ9LyUSTFIRMXhJ62G4p/E7Wyp0P
U8WCC0etcS2B+K9YhcwhtAmKU3lhs9sKdWVqj1r6Bt55wkgrhYw5rG9hTUTO7kKbjcfIyFNIzBoI
ArgqsYS645mg979mDf14EHr3jCOnAAORCfuDgKQ8ic6/z7t+IZsGloUaQLM04NuylFPldkgaNlFm
kHr9Be7vrXOckMuJEZhCvxI9mHrrKEdHKQbtHYt9nEo/fUr6MMP7YMoA7e87XSDkoJwClJtom6rH
4FBR6+FITsOv4PzFPfML4MiFt1zx9ljZ6F1wuJnUM9pN+qbY8MCtNvGnyg4/tzh4eYbkEDC8nmHM
6ubNwJSw86d8INq0HXsOcvGJI3qoLhtvUKWAfhx/r/HrBi9z+6w9HSSi3+uknYasYr+vSzY0RcY8
nsGUvqP30x8vc3kmWqPE+oeNxsjzr+/14X3erDkl4pqHHupf6pCwvyfke0QtNLbuTR6LOyOUqs7f
gcsrzlCkdZTr2aPEfEYiYBD+5JiX3iQ9vIVAvKWMNyKgb77GgUpj7sLLkf+E8hM3y9IO4nEGh7nc
4Z/lAqdbqPg3X942bcAb8uWXgAgn1Qtl4I793RFXT/23XYZkNk6kXFkIaXtb7FXGhw/GccbsFq3R
DCDXv9nOOt5ZwI6Nwsro4Ixjgx7G5rbzjWuUUw5Zdiy03xa4J3dvF4D0KiRxcbAMCrzSv8+FsOom
TBbeeHIeUMsq8ndAX6yH12C75yaGqwylv7IfYlBR5yYSQ5P+prL6PWfmapZnSad94v0pPmFFRLCs
xXrZjTBCJnPljTLEMfnTwbqmAjsMois/q1pfDiHhYqDG/568VRkEHwvtT9j+kzcb2fO6fIxlpUFj
CifUQ4ua6TKJB3zkgBQNdS983vsM5EB6MIGG1dUVQGOQkztPpWau4qbaVx0soCi8uPCrm6x3YwzV
Y3dEy6JKhUAWbUL/sZrkwTBRTbCZKN0VscFPTeOYtbiHajydwCZK1fSpEL28iqkOppDm7ZylL6l1
Tx/T9ztpiwX198khuwB5mo45gaI4tg6CAtHNeG+1N9fpVzDCV/yKS4gH77l2HyqSEQwRlpY/S4ez
NydRyHX/M8gPUyZ5VWkR40FLZvtMgBtOs+P72DM52I6NnozMrFl43tlfECSkvrwU7WPlL5hop+Qr
OCBOEbsOscaXyra2Od+azQBv/PQodAq2FdbTQSYH2NWoD+FT+30S+V9vjc31slea1spf/oZmoYlH
nrow3/VRGboOn3R1goDaYcJ6FLkMJZUonpMb1+4Azg1k1HUn2ijzPtID+WLmaAMqiNAbkJkAB3Y9
tbkrRJb3q3ClswXAzKsckNHq62/1xZwCFxJgW3I1UnZrOv+tWHZ6LLE3oMb1RuJqII0MPRKJq48p
CTEPEPpp6qhzvHj0f8wuJmThOCDO+aC2dzq8Kffz0YG2M/LUv1BrZ+cYIE/8i7GnRhm9Qgd9O0LA
CEB22NbVMz3YBPTqt2bokssjqgNPy8dhnLSm2xZFULJ31g7ZT39oO7/ADPZXvX2asV1AAJeWj6Ck
KCu2k+oi66KUeRgM7Dj62ByoUCilAX0a/1SXRTyCAlTl35C5vwlRYjTyBMQxkctfoegkZMvJpOJY
Q9P9XyKTzyFZJfbI1LojZuwXF9yZjZ8XlxqhzaBrUNLI2atxzC5gBW5ecthx4eupc9KqNgPr9Fxd
AyQUhSQIr3VEB3iAwol08NFo6+DId3fR9GnIxDQ3UhV0FaMcnQypgqG6MxbyCrf15xC0ihktWunN
yk+4F1jsvpC6HTPeLoLXDLu/gUp1WKcLa3xgYfJip/iJhyH+l5qp/hkfwTxAp89LwHQxof4xvoCh
AmZKdcctepwKuQXwbO9IvC5/cjE6a4MgadTvBnEGE44Ifg2yUoVoKZ9GMI4pSFuuI2wtnWHNHyqn
5LVl8RK8TQ2nwgDyI9o2RFXx4laU93Pk2nbQQw0X4hp2qSbhMKSS59pfkfEJh7E0Q3GHaebxMEqa
jetuk91mCPGbfjxBXvZ2VNTJwG0xxpQjZ766k+oviulV0XAnLOzAM78lm1IUJiWetvOFbPMj1UBn
y675hpcjCCoPKExukcfsbN5KVeCfmmd3AU8bp9sLPBiGxgqpv8PR13jb2XB048slmPTBliqm39vM
dk1dfQntuVSrWSGsLC4IH9LOZQNV2XDqi6cY1zVyZGv+UwEF0sBSEUeTaMbGPwshweBVSZoX3Pai
je/sgZynr7aUElDxh4jngbpioUcbIPwNNdsuzfcrf/m3Bdo5fKSHYl6WcEpGcK23sxgRpYuKejn4
NmtC+GG1BAplxda8AnJW8ABu+1a8/QQ6opxB+jbKW9fw3QzE4IPZDFJb4zRvhT/yZrq5ri0BlVJJ
34ba8KZn89+b+3xi7eGSkWSng/JtCKSBm0542el12JjOnngt8Xrj6kNAZsHJiMdDXzoCzH6VwpNi
J3Udv/RFokNNc+eg2xIS6/ed6Jd1o9Djn+A0uq1/JSO9+B4iAwocOjVUjbwzrAgJkBZrgFgvMLCs
7LJsD+XxLVzrQNJSwEPN6tovcNOkYo33QVwwdsV7rO15kwXpZ2fDhfUYONs++IEVybQNlBlquH6q
WF/klE/yHtl80M38h4XvKNC8LsZ6yQuTnJSDNCrT5ef/0JFhL+htwocqto/FacB6mIWcQH0a2qKz
zQtKRtlq5I5D/NVXJ2T8hj9ZCftKlrqlIkIVq08sxMxiyaOj066OV0G4MIzgQmquKC2nDXthor67
FsHE4REWNnxq2RSAIlg3fMsqf9pL94CubUPXECZ571tgn0F6+OjBsC0qTdkYjSACDM+b40D/9DLZ
59d0oCeJbolYfzKOXth9TUFfH0tJ6SYmRIYvFyts1V147hFp/FxECo1Yw71SWwMRTq2HRGUB2wlQ
PVWoZRLCbiikMefL/EUboVoTObPJUQZrBPsppFkx5ihUZL9OEMjoO99rABZScz49L6WC00vN6QDp
MdE9SjEfAzOrX7NIpBF/ljaPymu9pvTYAZPmwczaBpc7d104hY/aNkoBn1ejAlgRWI+OCLPKOBTm
G5WBNO5lJLuueg8LNo+EolcBfGBbghFOXhTURe52nfq+d9DMbq1Jv8eBr7OIkwU4pFeIThekeso/
HyU52vPWZtKdeSET3dCNyrcI/3lOkd247adkq79xVXSe/ti5gQDsQLlojxqt4t81pl5WW1escKn3
6ZsxtYEteMzcFsxTJq3Arbzs6zXp1ehBWuf+YNXERsSV9xPZgE9itctFQJgvw9IKH23cS437DyEC
R9YG7mP6DgY43690q/Kz/ct6nPME9tlmQ4QhyvPaVxb87mrQ5MtTMIMVLDCX2RzVa+hkznRY8KY5
JIPfjIVdwqu0b8gK+p2c1QmwGiv4GXi2NJFY/WnULgDq0MPcBo4Qbr/rSsHAhU6AujcTj/NpY0+z
fZnZBkglj900U/af8ceXOawFcuvV9Ofid2KBV636AbAhZfgziQTPLHCPtSFXUQ/xXTbx8yoXvLri
LBCAMgy9fJt9U/pudos5t8W/MDjdjASCOe6nOwkdn1vcww6QkBYycsovu8ZRT8Rfj7FTs3mE8Q6I
AALr2U57X6e/Q5LB2vv06yOLsZZjTgpczSXRtNs9+7BBx3IXImX55U1WUyWlNQa89Yi2GKBk1yai
drlCStKzcwIeXbLWUzxN0SQ6gvqZNYaN6r3C2DeEEvwe/g298eDdlR3gbF0eemSzjQ9qFDLcvgzr
P6qssM+EW6+fUKyGfOMZ+RSoA4gg5u0A9rf+jLvBAAjnBKAJ4hhJL8bwLfFaH803jB6RSRlKBwPx
82V4isfzRzXE46WOUj4hLX3o5MuUJZKe81ixaoe4C9O4PMnkYAxA6uHibRwZejkkQi8fwH4FaWu3
AcyyhVvhOEZQksufFQjfKQpFgTzND8xa6HPbuNRY4ObN7b9l86uKzgVLYHv+QEUgiL0q0ugk7sYe
JngpoHoQWkXo2oP07A2qloU+XDTvQFJydfQH1/XA/QeAsfZ3MoDukNTmssqIe7NnS6asQcRjcIfg
lucnLarVHY9K+6of62RUDHg+7CPFLybg6NspQ3X6H2B+R1yJxamaUtviVMsBl5g4ZScdWHEnCMju
G/PgkC4yxmXRQI+9FjneDAM0Wu3DK3SgWaJMBcxK458z9zdM0PvZQGmGWMrOxhpx4dbmvRVxUzKb
2CpNG8jxndEEL9X4Oa9swSPn8jAb6SN2DWI4w2Gr/1ajwsOvcsLYAJ8qqVQktHCYNp2nkmgmt9mC
eyFzRr2wm/NHpTiE44bhyQxA+ZqY2WnvOlYnuWoBemB0/bF9bARDYrYVgO8sKFK2d2+fD2TV6tml
JKAUkDrW/dUtKqim7OCycYCVnD8MAUcVG8mvXef6rDVYPkoVjNk5wVpkGHwokZXoiz8ZdvtaaQ71
DKZqEDsP2Vs0Z0yFNLlRYjEGuJ/O85VNQPj8dgONekkByWruR5TaW5P4/SmNLOJqFfZna0VBZZjg
glwHmXExiGzCqnj1sbcKTbQCCvMal+13/7aXTL+63dszhXw7gSUh3N1Pt8OBAIDLbAyzu7jNnJm8
svhJ2jWpPXKqs8A5QInjsA4OvA1yhJ+kmSiy/m2685BgrKjN8GjW2mMKAzD4PoQDfIR5uPSza7yx
gLH0R8Pp1OzkHOk44oVPmOp7v9li7s/nAaWC/3aCIEe1xe2OaBS7FAJcrs7EwB1jYpwaFBWVmJT7
YCb2ZcCADdzBd2NEOnljk7drfLclDJl0Nw19ssus1c0Yp1dq9U07O/X7xuaslLe0YAdKvOhnFFHN
Okd9aP2u5+ixKKiXnTj8+bdOsOdLcZShRODY6AoncTWTs6nUFYD/hJSf0x23gQO78NFydQjnct3T
6YoOP/6etMnePK2gg51aDhS1biuLn1A5I5EL1CedE9wJnoSe0IBoLds/U7H3JyvBaLW+qVLGHxGG
EakSh2kFcuU8IkwCEHBrM5j9CfucCmqgRdEok4FLNI1wQ+ZyTEu/P2JKDEbwgO81xWqdKwe8Z7+G
43XdmfA5ZzVT6R/1iF8bEaNoCRD1G+7IO+6XhxXvH3393BiYf6XGOL605W6ypn2ChM+qL+M+sG0p
lGtURnKaUYqcoQS7xlptSsP2Vn9BkLowM+61e2IVjq+KOj+qIvQ8Q1EfgevW59hiQks5htlZB6BU
RQIwWlou6BBzlrkfbSgFI7BTXn8ALByc2CEd1V5vqX+Ou/u23/kJs7lB0Kk8v4ood3gcLu8neZAK
rtYuqJopuS2zFQSDo0ByQK2ZCjJ0jPQkwBAO+TbianJQW5IqSWlddONGAzyyFdtGljPbrCKeaNUy
B+uonYkMdNVTjyOUh1cTLxhlC+9vd2lHavCYruakSFDoPvkmzgR0H/oc+gkBFaUFznbHzQ5dwqRP
UlUMIT2gFgEAb/3ALT10T/fqIHRMhrddCyw6iagjHoWJ4iLz4w6RjY5azbtbQPRi6Zbj9hgFUNk9
Yt3E82/4pasFJ6EOJPbv0oILlxzezNaeGIkOXT0HkQRXxgjRPQ4DAwMDXYbslk0dFcHF+dRTKEda
2kFKDuw6iNOY3w7En1d4iOpWBg9TK1xBcq40uwVI1czhHfe6w/pJ6XMIJh6AWX2lZHUFh+MR27Vi
Q66Jvhp1IQQLzmTjK8rFzdNPrjs4+cxn5J7Gwo2Zps7MBDs/pRJfcfCPUsoZPNlipA4wa7m8z/Hj
hpdSBWfwrik4djsk9WvPH00Ono1GPCuMqo+XicgBOIjKHS8yytBjWpSo3BkVCmyIBnncRP786WAK
DH4/QO4D2lXvnwrv4DJRZxA2y8VUYRnO+r7ksXi3KT9NLnQ8vfyoJ+yd8IuhKJXKiKAx0MosDhAE
GXk5dqxqe4K0qizVuhW4hZlHCnk9pCWw45VFhYpKxkonr3fleozgV0exscoBohjpnC6KoSp5aNRi
Zdk7lWpCwPD4/PVbVGr9bnpz+ZkJh98t+97hATyb7qgnoUepjUUIfieW0owj9/b/VqRe2ZUhYklx
O+sU/KpOzHcOzepZB6E4vbtm1xhfyPBCve080YnH03IriFS1mZC3A9Z+unfYThNsPJBq2anQ2TIB
8nijqArEitF+pFYU4cSegadHvrB1iQzodhXfdslBnuMfDRtLefYXr3omNPkaURIp76vhKeO4oJa8
VIJTwqKM3wa66CsZ0126bmEVDipZDt1uTHQdr17ZCSN7OGJUrS708WfpiJdKLNfDe8EV0JaQ8XFl
3xo0tss95dJR0Y9gj+e1jdUeS0W+nMnif85f42s0U2N5eOZ6nBcWnVlxdXrcvcSsB0X10ZcXbOTq
dEymQreY+2u2aqgXoZD152PiekZ0oYF52EGImeOY0TVuvfiw1irFwrbd4SoKVWZZt2hgFYeh6jIB
smnRpQ5o5AJvKaVIyUfwlzEs8d+Kqu1VJ+/Q0gOjUI3sn16+AaFOiB/h8lEb54v6bGIU1DBpNy7j
YjWn/pAN4UkmvM4acUoce6gwHm55PSB7oi9NZmqUyNavpwDKMWGSO230aVqMxBDb554cjvobUYPw
VF6H9kZ6iSCBvO9CaRweBs3Ol3xSp7ejQcBx7QbcpvWmuYAeZwDZDk+bkLPioAKjgorVMnXHBD9P
tbaj7BgYjHW7Uqm+uOiGSXx9+YpYBPQamyU4PKJsAydXjE7iMYdsWnNJJwuyxvTQlxXXGfyw6f/M
QG3AmapFN8fSS0pRZe3qYmg4bITlBVr1PK8GBGf95OCv5AKwKnW+YVAuOUWW3zXNRPtrb5/jY+85
Saa/7dIGy1OCWfejWt/MVCNumNz7Wm8py2PCe9FQtJkMETb4H+eIAlH98ezxYUJq1v6N/YSEkBRn
5tOS+ntraDtZVqKS5u524Aq4tyn3MRhIUO5hiMNGaLfhCVdK0XQxr1KGYcVtl/c5/kQV2/9tVoxc
czVv0qBPk+H4qfbIRgOb0oD2WS3SHrpOZoCDnSbNI2RTP4Ghp3YoohIW22/cPhiPdB+kpH+ZPCA6
ogQmBMrPY0VtNhztoCns3LNa2k0KzAw3bKNW/WZMfAsHmzChh5EDpnrh5YWVUn5ZDkV6LXqeP/f2
G/jhZ3rOD8uvLC5YNmsfKhebL20qExeV7s3fPBwmWRQLiy67OxJCX7D5N6p0J+SAoA0/RPSXx7H6
w0SDUOAZjGgndFoz6+/pusS0o8XLasq46z9O3aVH2YnxQwAaWiqC4qxz3OC4wz/UcsJ7Os3kM9od
FcnfkS/MRLbmyqpoxc6LITlhC3oqS6A09ymcgXtrSdSdLwx/9ZwCtOSBH+c6Rr+qh03ZujJPs5jz
JS1Ql/X1ziBakJndymNrcTsxvBIUSWc4+/Iq2nD97CHXfWqU6A9P1Z4ExCPIlw8+BCTDsHF6DhBY
bZTXaEVk2AcksT/Pf6wQxkLF5TLRE0CRAUrX7VC0MPa3GxuoQ786LpRROsoY0RtiV/uDuNXNDH6T
NtuXkdnyKTjGEtwozYkNIJOU7w18Yg5jjJYap5cOCOrREFwVBXFQBSfPREbpBt61nsYI42T1eDju
c0RRU6rtND9Obb7eVSnMXNLS5s3gbwQHZj82Q77Uosf3v5LDAsOXTSZfG1cTfaKCYJ05H9RBHQpk
zrsgTpXjbxHQv2YXyhQm9/BVt33KNYnASCCn86UumfDezFIC4o0+Mw6I9saPa0c1rwFWprwtSQnv
ai9CZpbaT+1202inaCN++fnG/cORNOA4FIzyqM/n2kIcJBMUFFw9LSeq3GDprvxMS7zXnvBFhtf7
ZAjeMaKL+xaxk+UQq58GLg9xI4ZKgAvBOIbzkG6mvhl3oncFGwweB0rnDoNVNgMxcJbzSEwT0Ly6
hddu3lPiW+6jIRYyKeNe2+rmaBtL7XwkbtI4TXQG+kfJ/xOjIgR+U7uzyPJHXAS9uQi0fdY03tgf
IOSFhsYBvQyLUgd0ynzEyj9/EotWVBgK45ALzVlsYbOjZ3rGEzmkcFXd81M5ICg1oIOTFM5ltVK9
Sn5ORAxR7DLehb+nG05y+C9mpFyniJ46JIZntSqCuCiy+ITopHJ1we8Z5pDro5AkgR+o+Za76dE9
Rr2jv36I3Es1IKiQisTa2+RA3sYI75n8cAvdJ9hpxg5MPzuFrfAslDh+5Yd1P1E4+9XpmLFb0YPq
KD686GXrigM6cUdmKsd/Nc8XBaw6WfCFGkJEbX+10PKvX5V9e7bCtK9ce3m17kITgoIuOv9+29Tr
3SawHcsVwYOEBkxP+vyQ52WgRmhzHWukVOF1zY/jXTunQnAB8sOxozaJYnNDhjks6lkHa7e7mnsc
ndliYpvdXjGeyPTqYuSo8P0W3KME0JIYa9m8J+JkJiQYCXuViEc/PeR3vkGnJyn7ui8G2DkX/Ue0
ttgClNuuZfLWjTTqy0xG+bmJc5SOQ4c/D5K2ucdpLuZnavGtPqzJK7wXa96u5DH40Xung0lj35bP
UWr3Eg7pjow10mZMyfD6p5sB9oQ0Df242L8NALeX8Nx/HQUZCly8eyroEFlY1vtF3xjopQ68Lzu6
AoP0UKTVS0x9/x7eecAbs01I+8YECLkW6bbsPYWf04sri4X3b7+rXXblu4aglL2y4ojoiFHiRzBq
98Bqr3KMa6oKzIa29b1LZbg+CkJnrmu082PNYbO9Bo7a+a1KlF6Ebxmwx7MblhPGUENEWV8iAakd
mLMyrFm4FsnVeS6g52Q7kM8eIuB1rBm5HeaYu0kNxBEFsJA5/8Vz0gnu+RblyBLwYhBXiM/UhgAS
vQKkipwuNnm8X//DuR21UKsb42dk1Gx37ATR0MDOHyhMJbxWnnUr7f7gq65dNessVbLRgnLA3AcB
F4Ol1ywivvqtpsm5Kvp6cmPPtcT4Wcuo8BKJ1peI4QQbNAukac/J6Rx33Yo5B8s7+FRGdbu7JYGZ
XS5t0LsfErdo3L4nl248NGOVLQZrIQXvZocJwhud8XO0rMtCPYPUmWzM3pHWpG/iKL5fpWZN2fIc
h8gYwtfZ4eqr968yXhvOavfQbHSO7ZeAzhNIOO/JyDB6EXMwY7TDcMxXwk2N+EDiYdP0qrJa3VLp
3S9SsThrWYQOi2z1yHFSW1yfsSoN3iCSRBaJntvHJVLE40i+A5wK9A5XdSAbcc0Clqdx5iilek/u
2+zuIFWbs2s5mpapCvPJgDIaS+V8eehrUTClewYlGSEglZ971zqgmtT2pJ3s5hwXw3PM49nD7eb6
Fh+1pvjagD5B44D3Qb4kvdj1D7ECqHoRHk1lPMjAiMwvNa5QcpDNX2AFCnN7101h6rAytsLp77Fa
OkfLiFuOVBkgJwBlwccrxMQHagxFs8jSKAMZuW+4O2k8AjOJKI4epxKMSGpWHThX8VbU5kKBaGNn
fqjaw5JT645u5bAFMiZyQyna/mcd+49D4q3WJQpu8E03WAsAPGwLY0ZjaIJwZFVJS5fmlEk7cJxW
bzhIU8oZg3u8eoQqFtP6YrbrL+tGS9v9jyASnLwXAHNWCsofOY18ukEWWP744CcbaMOYasS8nMuO
Uat6hiUxxdTKZsPYio4hI9GKJ8EnDTsmG273KxLYzGlfZaA9gKas6hem6oWdNqDBzMoswhNggweF
iU7I8IjpFYXfY8MfBtrh/jtPA8eEmSf4surbYFpKp3MEY2FtTQgPuhBUHcVQTb6T7HP6/gtcrMC+
BGsQFUKDEn95gg2VmG5RVPrDQXph+y7VG/kzqfAi0OOrdA4EZikcLY1jhGFnke7rqBv5ijnH9h8S
U2DB2w2DXSNORttCgJKLxsUZtN19tRWPzYM2n3ck4N7yUH5s1lUsemM6QICA6zrCpgBKd+JtxQYW
XBxxbvrndlD8K7mjjObm5eZp06zV6UTntJuEa6BCKblxEeTL2iC339dix1x/UJ5cI6qaqDKKGeCR
2kqhIfYhn++MRhM68xkxfjbm+7WtBbAQZe2NwJs/5mFO5hWwn4AMml2fjGBTcuBWmcdyJ8Eeta1R
OVw1Yb5gUK3TrjB8Ug4dfnVoeLms5QyAyRFAM0ui5DbezfjfCowxexFcPFZhjJpOA5o5wreiOYqM
0C95k/WhrfiBjK8kk2sHGPWVjegbZFP7K/TNnoQyTnEbaZ17BfKt0Outm/N9PsfOkyyNcP58xf/w
S9CYjW9t5Mj6mnSUc2/AvB2Qk8UKxFtP9o5d/9wmWwLm5f7JrxLr7wbY/rqka25ch/ftVfvnvhBX
DlPT0aCHqvXjQPJFRlknEXBx4k/cmhMQ/V2RbtsSX+1dFpPVuQ1HgRLREwy7EApmVnoHn5D+CjdF
5rI7WgShFXxZMReCzNxfxG8TjOJLNv8NqAD/aKr33nQ16rFAls5OB/FRZjTLdHERWs2/dKxxKPVP
bvv0JQeFSVZ8lTYB0Jx53vmRjPdYIeQO5pjzwNBN1T63l5azS21uBYr2bBGkFkaCrtEtLaNBzOXw
8juedDKVnfrNVvytMkFf4bmFVawgrTnxOjgF3ZtJU7WvJf21vkgQJEPaa28OhQlgDBmWqkJyYr8y
xakWOCku+3CyEOay8bFXUg/P4ZlrL24KzYglu/pugB8XJA3P8M0YqrvzeiaSwFN4GeIB5knmXuZg
V+vjZUeoTslUGEdENfQP7g6gmFnXuhpNFlCR5lWGz74zZZMgZOMYX3qMvm/k2vwoX8qPtbfJcfK5
VdKFpQ9Vw2jP0plHZPbOURpVD2lI8px+uIvTNIl+kxPZJqEkziKB4uBDsuVCr5RigpobBqsdFn3B
4KK6RPfh+1hNirs07uBjQloBrdwoHBG6KTzncGs/2MLvptvQABT03bSpqwMYffapPpyu0k+HPABD
JvIDnErXY3TOcvttG5c4591hLgHeNgITP8b0qPlt1LusTNuoZP3z3tKZ86wXxtg/WRpyFOyGBHH8
XfribIB46YvW7+8HBiNFHL8IFFXutu6VdXGbKANENc1uDQdcUe9J970qZrie0o3viOO8oKxA0T0x
A9Z8FkTyhxJaMoOlAAWvl7nJmay3KktNBEwZVDVaLruoN3rGjT1oznAjmhkW8v+i548O87wif9DH
ov08zVZ9a+4Y+kc3JgWT1v57vlBEUDZUWIVEGhMOk7enxqVyN90MpHAN1Jfg/2vNHXm9XkpbdKyj
hDKldqkB0evnkkgNu/5AuAo1n9el8RAhI4fWdCcvAdbc1uf+3QIqhIW4sRrGeb2zLtS2hpUgGSxG
8Vn/SqrawSBmuTTfHOMRNHceuaz7f8iBW4hrK5/TGHPC7METRDo8Tz2LfoZN91u7jn0FRwyLm/Eg
8px52+hPUcSGmzQPcwPY62WjkUFQPiYMI7YweKSLhXQk3klP7AcMz4dyPA0RXSfgfhU2d+5t/5Ah
G5D8KdK/Y6TzLXdB/8RUlcKTYP1zL6L9tkwFYKqNo28bx+mxvRCn9RFVAFiNid7efHWn2+5owIAT
BnrVCW2soS3z7LL+EhMB7j6bQecYyzGf3OP0NJLfLzqNA6I4GXBNqP8RB3RjwUdrNm3oOk4tLJ47
pwUc2MMRl3yh246n4niUNS7nDMQ0eNtKktwpM6svEaDKFXbLvpEU9mYchugU0P/4ZBydYOhefgt1
E/hsGEelqi1l00CU6zD92T4Epj7Xr8/Yu4lUIpyu7LTvKDfmP3KW1DWOkVncPvikrN5k0sHTSJYu
9y4H1iV9slOtp2opAwVwSAyXkly4aFLVsYGjC8zBkA9+CoPg40ysrc4aIDplOXHhJhCyknu/TZ3B
tLJ1q7dsLSSDQR1RdGF5lQCiql0bFEB7p1r1bdRZvw/CAV2BWekKJ4sZAEbr1LCCaGzjO/ax/lvQ
wjgI6EX61oXW4+ivCiz2J1tNLp2CsGpPCGkbymilY/11DOPisBRqintIRz7PxC0983PTC8cjlJHJ
POh27b0utpIEQRBO6cgF4Y+h+1QnkBFOz2EDlFgTjG1LRHQjpZMyC4zrRLxI5CwQ/pfDTT1MnKtY
+E6Mv2Pw4TfpqW2nhK5XTqhwlaclCAk6vVwy7Z8lcwqf2ysCFRzATUd+QANSmJFro4vDcFgWhX1C
lcUcoGLZsXFg/uQQFIR+XUv2kdGVzbAIafhJns4yYtqnklk4K7sIoUdbyr0mzi6p9OijnMQBulOf
A6t/B/is+sh5V2v+Hn53fNmVP39JUBO30kmFoS/Ox6ShgeX6M6SZ/VNj6Vyy83y3O1dLBoV7V7GK
9CxYwtCudE2S2Nn5iLYEVZVjEwwm8gqan99OKqam2ASwoGs/cOtdJYnKeFgzMlJgTbJdHTPC7qOY
G6ACiJNRvU3XiwoEdMGG7QxJWDo1YV8Ul5fCeBjMmBPrP/inzMRR6v90hcas8zRsjIEQYyyjME+i
TXqkVL9BjZgO8GD5mpxGM96MAj7JWXvLJz6o/aPumY/Drxb/iG8/MxtIPIe3CrTIGSZI5g0GOTYR
ivpm0RwOWF8PSXTKJlszz541pqdXllfXwwV5s4vD3A93OBOPORp+A4XrFPgf0YyfVOFL3SQYooKD
7FhKmmTpnx8AqY0LNO/RQlOTrZKGnzliBhuvSS6JdVibgVnINmHb7TbjttKZr1n0t0px7ikSDrYp
YaCgF2apmd+OySqSAraY2c0o9BSJv858Pb/St8NiFhLbLkeBr80HXQNfuHs+znbU1p9psoHPRGjg
kcbIdpNlV/LpZ6BZo6q4rg/+rigKb+yeHnsGfEbxrA3Nsa4ple2BHsgvXMOoKcKlHST5ND5wkaUc
HdAswE+o1U7lKUlypJRdvnT/hFf0NjGAM1fETuocV0DO+aFUv0P+qAl8X3Ix6g8xpa/kHXCz3lGM
EpGwl/ocYQgmNhuW16WBj+wv7aztme+0cevxUhlcutSvj/lEjpLkeOSrsQCGL1IQqN2F+TCerzNf
oIf4LrAfIT3Ju8OgoeOMSjZRP6arH/QIgUxZys3hb1f0YdOdplzZxStumdg2/V6l5Z36mmDIGvWl
8OO05FD7ZU+naiAdI0Hk5tuJj2mlAgSVJnB/l0ZSiWKsVg06P3kEmaQ0AqcqwfjuvY/3ZKORrv3D
uFcMei3yu4i5XWTs9ciaydF6zBH/4L0rvzpDxWQQ74+GxTDbhsKoNBD9CVntu+4ZsJ9/gm5N/nTS
+7ouv99WzOmwALy+S39CW8CYR+2J9ccaHiShbVAZYMUL0HPkiexRaD9JfJgs6JYC708hnKMFru8F
4pR/66lIRy5+/j18/CAreq9FsUOxho9yy4hj3jzZAhBhF0SdHXNlVEILcxLfXp0PbLwDFBHr5B6z
86DYnmbFCTzmK4B94CQtZXmYIkx16Gy6qkCl7/3o8gvSwJ4/GokZlPv/xX047trDnCnBrJS48+Iq
sk6Tt2qR6kqbJWDX6yWvunf5feD8AWMv2ydPkOja4SfNarjxrISCk2gkV7kP8wjmuqYIPLVxg95k
C03VPaCdSkBzo0BpL1vzuC1MMSDiU08kG2URJbhWsrA9/CC0vqNcqFe46VD1sJeY8d4UUj5QYhJb
GKlhEZ5YRclXQszs2F2HVHeHZgfsaefxZ1r002d5lbs1K3crKtnWIIcqHsiIAdtFZPDf8bOoCOAo
FV9/6dhe9xT2xmCq1fmY9KfgDlj0SQPfurkCosgmXBk0f0ZM1RiMGXvEJEtlNPRBJemeT7SELbjK
hCIKVCBtLK/aV8ZKQbS/0RtGpk/HBmWrx3v94+UL8MAcMhaX3MWa6dEakvnpa7JvhUFsWVuNQxCP
Tsklwxr9B5n5v5Q6rIHgcaDRpoM7EmRToZJXQ/m4S72CocGJ1Um3rQtIYZdoSujEs7gNtqKLz1ln
/2ccszljUAHdBbWgMANOePeCcLv//0RqRPNcov+FHQ7+gO45mgZz1z+sZBze41mg8umU5uiy60mS
PL0wFPbrwY5lccIx0fupOTgAphYmHyQPWGM5laU49x8n7n4XgXWrmgRrktaC9DTjoXhEolFhnXBp
JVy8v5bSxczhgtWzvPrKgVXQd9QUUAIZSrRvFmHNP7gkprh4tKScotq6+ZCqC30aHMko0pkhG3Xa
M4fmEUFeAmNR61ePU5Pvxk8iSuQIr1oMT7GbQFiPD1V+Rfdf/iU9qrR0mtbYuiE3K8CtXOmOYBpS
bR0YSXXIb1zLcNV0wzBuYUuf7Ruw+zMf7rYQfAP1/x/Uqp13ZT2wiNTMNiV5SHKLXovsVNvTboYZ
fbfPKZdIcyzDUv33yulyjz4BTLI6pDnm7/pGmr9+LSbZwyIRGapGh1+qFedR3m8Xlaatir/DHFu8
5ofUUYvKZjEyo1cm0NiH2Hq0e34+5DOWVg/M+o6jscPP0EY6GPH2s2iHjgmyuO8bJj3kSnAXVTrb
PXuq0uuLnOZAeen7reHLh9j8mQeSsCs3zHkJ8f1zI5KGCJFFWKcqu/25Tdfn9jbyPd8kOvffbLwt
vspJWeQUcID9iQBSxeBX1QdTgKb782zaIakK7tCmeuqBYySotwC84U+nGP9/7aQqPwedGMUYxDrP
hsnIf2Bui0Bju+5URI5NbDWPaND5Uc2SNhN1mHANpkLEuWXF0iy+20NgtrNA/S4AipSYH+FSVyR/
m4XahSJnF3P4C4SwRV6D0g5lJJitdB1mXStO9kV2hZ+QOgELynsY0dfL0FZ3Wz3LpnU7Yq1QJjrW
izO9pV3EcblFOU0K0k8Qrc9WvxcjI9jS83+XEsZJEkhw4e5v/ILtp6yobQ5xvcXHTZgPp4tMr2LQ
+VgAecOAbyd/gIWLOp+RE66YM7RHk9K3UBDcV+6iTD8W6HlbWdB+ij/3k0MOnvSnzADuVdP8RXyH
/lUvcpoGnHF82+zAdC/dgywnqYHtHM5eje4Y1tpJUw16Z+0+JgBVUiq+ZJPQT4JaIrrTglYz320D
wf/K4x2n2tnsZy16oZd7AXPrchuMIYULRF74fudrytNPJY/7LinUf4OzDf+Q3hXicj604d4VG5gu
ECqyzaPkQoKWFmltD6Zm96b4/digYFCwcK3KVE3Fw2WvuSMpPdJm+jY4WbxHcBEa7RP9PF7UY7DI
ePx7/nnoiV0WEopYvI/91HjgsL7CHXK/oVNyVOQwurCIK8rA5sIeZ32buVNgZG6ztad2JBAG4E6d
v64fGfhDWfC75NogOvJF2F/LfqgFQzCAJzwzeODqsg4GQek34Sor7XWHW3BN/98voDsNHKKT70dv
A75728WFO44JS+7jti6qQyaTfQLovqUQ1+vFawXhOmdQNiijCtEDP/UMdv1hcIS/vZszR73S1Duh
78PaZGBUYEhLxgXbmz/RNdwg9ORdXIexvcQj5yOrh87lqgEmh1cjmMMQ3r/53pd9fsgg8RSoDKFM
pEuNfvysegDKGQftW9uoP5v85Et4YxNqGHHRa+XMSWsN6yyZa8yaMS3M5Q24YvzLAe2DJPt1BQ0A
hQNB26iCIxSWM4SYxAPhvnhhyLFLUYVluXc7X7NGZzpEZfimKLn7U42MTOenZWSJ03vhBTSeBZIt
dhWRxSeNFKzFD6VN/BWW2DXQ2fYqOGfTcJOLl918h5bK6p9TQrzdHODYHF2Qdp38RXP6d3rNyg6O
sXW2XfTL03AZeyRrih9cyz5RwVLYxvT31ogO20zyjF2DrqT5xkr7w0KHsMoTRAYThEIUkNul0k0S
X48KCSVDyU3wqFHfzOW2VQCq67J6b3kt9vulz4WKpJNeprG0dJQxJFXhQzlqCINIMfSuGXu8/tlA
QSyKah1V5/RbGdLBw/ESPmvw8lyeXqjU3fLVMz7hBAllwYjExCTA7P2Nxr6ueUNvlLO80kbTxjVi
QR6OCZuXJOULxYMJ1ww7fh/ocGHWzY9FP3Z8hi0jLWGZ1fg+cE242rSSzvDiz7a5P3St5ie8wmh4
yoChRnAtn0VjN9bk8+X3+UNbcLumY9eR6nzSZxWvg5KTDoWJN8+Bvr5tJx8x0EUHv7JnBZQpZixk
LOzKVO1WhOvf1768NKKqquiM9HAr4pjdULrk90RDX0Kd+50imzlzJ9hVV3Ybz9MQC8gVD9QVnawd
yoekji4wocMCOaMkX/9LrV5ba6kH66mA1gZb1JjdsHrRboOMWflQfxjsbjlh3ebAdzDPAeX2pdIX
AYO0RfKyjtEohsT0YXCCdweqx3avEI6f1TSnFF54YC1N7yMmmAn5/+Vz5ih6LSOpnWNvrFCAHq2M
4aSSlvgJwxlwtJzYpZus4pQ2e4yYOoGd8Ev3oLf64g7XoF2SuEK0g/H6WpP1jo+BQzxJAakgyBR6
guHRZOuVKU50xp5ApUxSgOfeWjHBH/eVZDnzuzh7COCOpWBViDjZ714bBGeojRksVcfdXFVI2lh2
k/iAry+Z3XgjruuvTyI5Lo/Akst1iQTKnPmw3IBzzRZ9vHrLXOE/F5JJvzRdBcaBD9+LsYRhA3RY
TWt/bqQxsaMy1YX3a5A7UpNEW//ClWaT0hJC9OyMrMvVo/pqZeO3OeFXK2iy3UDKQhEGhwsYF1MW
75T5Q0hQhhtZ2zyHn6i4qR9KWUOoKwBVYLG1UEdo6emrW+5rc+uzX/uaAa9NY89E4hCVfibDdSQk
QHxFaImt/kRGyzrVfflI4HA+dP+6eswgCLdoqfZ91DSloI9PAqj9OfD7/Lj7uUNv2/lijtdyadTo
WMQ1KF6lYsVu/lCoQKlViNnmTqnOA/zzo/Cu0V2ZU0MBdUPgHJp/zuyDbzuQl6g7FvHVyl5RV8w8
HBRsChFHYi3oz2eHEVB4OGY5Jk4V1k+xKxEx+0D7fh2j9EPLAM5DqUey5WJ762htlRFpdO+oIcpk
b2bRGbcuR+P867oYxnUKczn0+TMmvB7cUuG8ViyRPVbiXFG8pf9tXlAgS2EdockjTLsZyYR/2nl/
jdJH/EbogefJ9/9dpEX5Fa+DMLe5EPXyc87G8IQBxgw8jA+CvHAmPsPSAssY+2mDlf+5rp7owsTb
jTNJ1OkYyAUasnjD4vZCIr+vuz6Fkbrf4e6ihaDq8/Q3z13pji0XPNPHiirGkXEJeo2TR38GWQUl
7zaKQj6sBDG+CXVIbH5oTXv8OBORWG1o2B514f1E8loJBnbANvSehz06dcOFwZWQ9CvuoYsd4m1Z
tJyLm9Ij4vFkFHbWjemTgVPdEGo3XNfO5XGbVJLV+aHVEusjJwfTA8ethpYuISbTDKmx8siYTA6c
6X6dbGD1MzQjSDt1BLgnZhvfo9M9DjwkSgDDfaJM4++yIidfdHww/bwCQhaLreDPhWHyDGfBS8o7
qFX81cfD3tXikMq5AR76jiyBA6oNdauWqNKBkTZ0kBCC2aCqIAO6B2Y3MW5+gXUGiiWCc6S4tMxd
TZZUr8dKjPCE0Ljn26yYjPsZpuUdR7Z2FOBlkVIbz0PRiIX+NTVi2he9g46G1eY8aUm8bez770RS
tAg1y9rHE4YUf7zvUvoNGzgH8/HUTtIEtSrc5ghw0yVQ3IAe1DRW39rsjKzJNO+339DxwouoIfXu
4FLewk1gFa0QwQWmk5a0g0JJDZEhy0AhLhUdVicum8pCzho4HG3Mhqu9BVIyyrI1cYKBiwu7fZOu
w/cTwybD40F1VksbgbfChq2IIqVNuhtTeRLGXoHArTpXBS2npC7YwLJe8K2FDg4h7MgAG+LfWX99
lIvICozHzrPPfC/Bw/MVncawWZfkvcQ1lmmorPzbVQikSdVqv04U+TSZZlGw6DoyZ0Wp0lkH2Nua
1bZF6nHPvZWYsbQJy2Bv34NJIop2+FvjjFt6gUZZz1gfak9HESRjW3LnkyJTVsOQq9zkfUR0ZvDd
+fChD/OJz/OXJJDjuPE19xEYgRawmu2ms7jo51y3VOnqJP2eb2XRhYsBouVpUgKcbY2S39seVYuR
ZVQMuI8aawfjnV/hiZGp4zQzK1mBk4NWRsidPcixlAD5Tpo7gAYB/HbKhrVNrlsGHmMPI18XgFBj
W3Xvj8RurAkSfv+tabLKaRYK1NDNXIlXvODToa2IAMRLf1XIRnqtYIEiXU1heVkj2yG/dav9meAj
VG3Zva/v7LEgGH3umOUDNNdEdpW8R9WQZKCcN86Oti7s7IU5bXBlxeWRe1z0lZfLjX3VIY4e8C34
rT1XKYX9BJ4Zj/gwiqH0YtbeUFe8YmeHhg8KxsN9jCT6mJf2q0t+Yrq3zKj9W3hxBdSrXey9Gvk6
uSs8rEKwOAooJao51krspMmUg8YQdiy0e6Xa+L3hdAdosYllTGtLdsOjkwpPiidFJM9nc/Mu+LnD
ZI9o0BheuQajPeT6l/TULWphGMY6/3oXfTsoqixKKFrADfXUYOXPfIy6ACwJG4BAeYEh4A1ICgkk
e02EnEIszFIgANeYBplCxp4eaxmCgYhnwg4v9toiVjVPSYqrNm85pxBx9TE16kPo6m3PFvtD01V1
kYmDgmcxuiJSDCXL8aObhRLtzg/pIM4e18XYHuJPTH2QWSc7rS8c1yKzJspPbtljWhRzRnPyZTZk
9+bpi/t0RGw3yhDwaPdw68HbXkEPg4LeDMIG/hyeMoagYJmh6ADoxsmpnKgqsvzCaWtjYYkOGw8U
WzBpW00cnJQ1Xg7mDllxdkDp2QH1tUhD4TxVa7MNS2KEn8Ip/dsLEJzPdYAIfT7WejRb964WUZD4
Y19h6r9HS1rGK1Ehs599HOu5/OXQPBQMf1GWdhttm2n2P0y+E7Zrtqlb6E0hpxWR1pl07eNI8LT0
4cO3gClwLkEW8nq1DS77UTX5mMkiPAWdUF/DUtl5Fxib7HwL0PGgJRGozDaOOTmlIAGj54AJePlI
VKqkpo546r+Y+oAzcZMDGZGFDLBzo7udY5Es9SWZ/gEq7PVb7b6Q5hph50lSXJ8TijgI+1ITKbHC
+K2JFCtoobWzbK0QMCSzf0Y4XCf19RazrEmb+S2IO3hqN9g1+Anq9UigYaXhOL5YT5FQedGq6VKW
RAjtONnGwevbUp7UO60UyIjuPtyamWyt54zFd3iNDzKOZsx6qvo/CaQBcmdjsmViyiQEr3T68u02
z7YzNlJ+EwFexrJRvTij+gA/9d7V5+QiveaBUv3YkKbIZn7lNrWpburD0O9X7GAkKYQasAmsEHKO
9TAHektJ+ArX6uHpglUMAyiWSS/CIHBPf6HRBm04cvEa6SgLtyx2I5tu4oPgffHwxOwthjiRqSeo
xSaTaKMzG4YdsMBZ/f4Pd5NhuG551dZOwCFYkHAWLLzfehoadecpP2WGPEnmzyl1QJc8eqDigXhY
D+tIcAhSB1/blRh9xb1nnQBt3tkViTGLh+aIICWTuDPCpLHVsfKK1+lsd2fBt2vKZKCUs1Vvr03V
Q+t+sKGkUKFeebjawV7PkWJPAtXUN1UxZ0RhvyrGN6Q9RZOv2ow85n54RWkDjKItUAcaN7/SHU/Z
RMEGcpPK4/Kw3onKmDFHRVwbg2ruhc6YnT70cg/p/TvEF5XGjezO4dq1SZyfxIuHRTW3Tt8x2zX3
wGwgOBAs0zFiLVX++rKXeVMln5LIRQLWZ6ywwRJ/ohBUJIS2k5slvjB+7WwIksTpDsvo/Ptxmojs
IgttfkQXoxNaHQ8Tmuu0HZkfGpojxQlpg/u6f0/Kn46rqUCHHVkprsRxLvpmyJ6vauplnJN6CT53
eMWzeKizwI0tWo7+IyNfyHZvognmdn0js4uIppsAed++5IFz62jAaHEP9D5h0hMbGUc4zvuPS2wU
JhETcKZ7+O/g6bJ1UjBIo7tMZsYMcTere+x0ZFLEtlaJpN7OdvcY5XgCFv8q18FsKdmxrH8M+ALj
CzIodRI3/n0Lpcl0jE2beWTJS+8G9ZUiJpxLLXjmT28djYdGJia3FaNr4YRUXsOjbhRjkOXRcY6W
IB0GzbMEGA2Qml+IDLA+OiuwtY3qdf8LJ+EY5LBZ8do0iPbCSw4UFPlnzachoAdrgpBHX0TC0vo4
1Yo8AIYONLFJZ9PS0XFfP727rIs7dQsKnnvMMmqFj49iUbSXuxqcLklbFx3yi7wtaHwum56Pg6E8
uTYM1nfp/BPuFxcl88/ZQF+JRHhf+GFOApncrk/c2TYwdC1f0hAa1Mw95FH34dOhobDX4w5gy+bW
Fc27B65twZ8+UA1iR/mkHyK0LY3Wm2tJsJvJZ76wrSv9G8vRZ7hu/QNbnxp46rKR+UYNKwADRDLa
ltOlTjjPEMfQFnxa8AtW3XYbW/T/TFl8oBmDfpKXBEIUGDWPumQR/IDSUsc2Ysj8hiAH+iPL2tqI
pdikyoRBKl0YRDoqtop0uhmCigFlfIXqlSBggytSnd72n09h4zC30XiWRMl/hTwGSl3TFewlgmD3
N9wSJ+AJPaQ8kup7c5axFnK/0XADICXIRNnF6EA/UzMz2KU3VxT2wdIhyjT6yTUdZbZ+Mse0mkyn
8XZEZ4OSiWJMmDuZvzpzdH/FEhoKCG1XiMJ/ToNNHPVK8ftoQICYV0sdpJzsrk3gLV0Wo7lMUzYh
m3ADClCvJ1hw1JJeWNHV8keyL3CODGByXsEA/9fA2YtK8xioI2N2XXJuOecAqQ1ucZs/01DKoH1s
Jhp50n1u6cHG/WY8lJSrd6aHJEkby0JKifBFFEzKu54H5kotzm10/4nh4ZwbM6kP04JiNoyTP+7d
+aOqbpDcDeKHZdyTrzRqaQeWguN3LvJKVi84LERbC4NSHoVsmUPS47O0ddWpwRU8RCxwKIP19KWx
CbGnHkzMJEvs1y/WZ3Di4StB5m7G/RkCS+y/enaZMcBjVvfY7fOWXqm+34QwQepzfRdwCGDD3VGJ
6u8JgSk+oykshEk7Aw+ytMymiWV9f1I/EtMwY2LijkfB4GvHAX0RHSxk8teLpOMr8mzSGupR6V1U
4q0Ih7yMY6rBpULJYi7QcsXnj4XrcVdFC9EDtzaBo7Z1lZvcJPQwghiosM4mES0ihiMenM4irq/a
a9En1Vw+ig+FCxaf0grfuAzzGLQ54r0v1J4xyqV7pMCup6cG1xRxHVYXfLDbq6wLGYEPAe6kFHRD
UTfysWipo3KEqmNSC/BuEmbLoBzKcZUj+6MLmtVzgqMDGnSX5WW1iglZhZv0zDyUgb5iRu7Uaj/0
atQmBckglsQDpgldFKlG5titZ+mKGm8Ksd9Ct/LGrMvYXYgruuxn7SBfWKq8idc6Db0lUaLFVaLY
GlEA1bk3aXl6xcovKkKP+phRzzc6vl1iygWU/thQ/PV1xv/ju8WFPn0D6H8FmqMfTgtpLFyd1DLS
MeMUtcBM+d+FJlJuDryJ7sk7o6/e7IQD5Y/VLuOit5cRIPWWR+k3GEMzVWI7PWd+MdNPfamIRFZq
1qSpzIB0FrNQqcdcLShuTL+ZvAXQy0nBvCYUj3dXXhC2CsKRVwaZJ4DeTHp/NVAlsm2T6m9/HCSk
CqLwJgF4cPd16dRWhRoBcuCMRDq4shgNlr6sZsjMZmjkTTG1WgeP7eTKa4dos/CulYqSG8jCwwNW
aB8lAyVi8gSn+UFVtp4xSp52Gzk4SwWcRv/JhytDqFtzfTSCFI1ukATUanqaE5MxWdVJzXv3bRiq
M9gYz2o/ui6P7O+T3brhRqWewMzzS03+26uJrjBQe9fAW8lNn9F+KNk7INS/V2tpeT9Qa2vYoOSs
LAltWrzkJoTHb3MsGtpoN3/Tvz2TPU39DslDI9TJ2mKyAQJ3qmMlyHVogrhL8pJ+HICvMUl7M51y
a76eia0poIL3a/kUhIP3YM4Jb5XUpnm/VeHMe53fFd61Zg0l4mj1NrQfi8IThQU3OYBgEPTjJ+Io
V7P/T+d/qdAQQ4HGvoo4MkmPdDuEqGgRX6xgTULiMYDnsMmaIlf5bUOY/krG4VSWmZovqWubijXy
cdAT6ZwOKP679M0UCnyx8VTBZxIVsox4jhvldSejP4mPYCmSDc5AsChpcd9LLY7ThXHnnJ+axyEx
Oozb7MUQAZCdUS9Gx2Sv4oZ1lNpBTUqICfS1a3oL8EDNaovz9BuHP2+2J1dYj0a4Nw+uMzzY5ap4
enJsXBAWgeHFC+AwRDI/V3P0ktDOSoKIKtTngTct7NyoAvSzihjx6FSQIpqzKa32lej5P0IHxSyo
GNe1mU8GbIu+mmDRagrJY8XNncDaCvckO+1gaDrRVjYTkrYMhM+LEwiXeWl1hciXnCCHyAUdGrqH
+KmJqNyU68HtaL3BnWFab5aoY/OsifllsuAzegYVS5+IFuR17DHGbq/sK5CVA0pUIiru9wiuDh6a
vezxXY1HKl9YfuyzUazQXS5btJvLYEJ4YQqJWY9UhXh2t4dLI0QjMt5B/IfV61Wv3gwf4PZSOUT4
UX1pdz+MRYWI4ZsFlc6ecxNbO75jF/B3ATkd4L4MmJGu4Ky15S4uPWg77CY0EJ8TuChB7f9lOlO2
E4rCFcryFoMY+7Y13WJ3FldUNbRznyultdgSe63X+Biye61X8TOmF8TeWjMHhOoTjDG6kDKcJswf
3jUZ7Rbigh/ekoNavoKtePlAVVo6D/aFLMjdSIoTwdDGg5FeAgPN87QcMKA1ccczpFNmSr9dFKMC
DQ/RX7lKBOodeB8MiSKLLfNxle/zJq1XSxqpR59lwI2wI4u+kPczaYeRjlPMYZbZvFjoGRKewY1L
qpGew57/qU26tdV4Wj+Yc3SldnrHwIZ6sg3MInN5XmU9UWGoC97S5Yu0LmGZa6hsazCHOlMufNaB
XpO6fGKGcGZKmbqDUgARe3Nvro1D3PLUIMtCdyC2SIvEb0Iz3898t5RhQtmZgxDGrhnERVOi7E0S
Lr4y8vSNDgRGcYWfvkksECR3uEnrnia5xbyaDJ/L9R6VrprSwW5twaN3yqoBh5MkGvnyRGOIvOUJ
RziCj2jNIfetLPqkM0uUUGd0xSXvnXvxXl0tPGDenWKkC83Vfpv8oovQOLFtk79Mr6eAYQnF8V+R
qw5n3q0vtOj3OzZW7mQACopMnVDmctRb2cKqooAZMTD9bcyuUblGOkOiW4HeBNF5WO8u3EUPf3ES
2gUBc/m60aqneklTPIR7BGfcCoIlTjXvwmHmY9pyqT7phhu2TVrk+CEBGiDlKTCwNLltr9wlogQ4
rzWAHT3WmkjwiCdsqijcwZMypPa5OZEpJfwKgqa+0OzK68RwyA/06jQRkiYMeO4LhN9Gzlehzjhp
Ai7bY6juve+6mDkbSjdxblEIEVtkUHA5pN+Vtq9yZWdC2lQ/NAYzenfOirf8vrD2rbk0iBbqsyoh
+54sCago26qoDWeDneemXn385IxJY49e83/bnmW98muqHaaJ3hY8u+OQbkwfu8X5wgH54xk8pqIN
y01gqzZnne7GxJ5DSI4j10uV2mUF7hcpfs1oPjGbjRVbbcEABiHXRYA1xYRVVRTpFW4m2eO5UBsl
Xo1ElZjMDB5cFPVVn9OS5YqjbM1nKb2fUSKI0FY0411qwSPP0ODrsBhr5XWVpCKkrlTBU0vljGJp
CrBCDMhkW9BaJOG/0DgAz4p8gJ50hw4hiGd9hRPUXSKrhMboiPc3E5WHoF/cDEKsZgST8zcFRoan
3G0eVXVbchjPGYLwjzFQjDcDSu+4BiDwfWO4/hTolfivurjH75XdtZBYX6J62eIVF0dg84P/SCcr
ggUizPgsgoYdjaibrJcCP+WBTjlHtOsGuodIHZboSxBGPPcjIJBV8FKCYWWd79XZtNI9vzJndb9I
FkWwPrbQzjVo5Atp8V4GbMlZMAIxMaqYG8MpOmCVniO8fRliUxcBtYrcAkdNZfi+Dh5w1gOG4v4H
v1zl/PRRS/2K6szFnZr281Ljma2qMh39bJKzZ57TpvueR558wxv/4yrKFl/zig/Dj7fTHLd2ntok
oQz/8Mar2Ynwuw74/Cu7gYLHRTCePp5Ift9n61jEbRFVyEE6p/tb2AICnohoYenRHC3gB1dS/xnn
Pm2Sm0RXn374dvMSCZfHy0tqmkwba6Y5XuE+PEDiCSUyVtQwiGyhuDg4smDpAR1Hk9fzvBNNQzhA
Q7mJej+EJGLx/5oXFCbb3Zc+hhDwSRFRtnlaSH78drFqD2wXJNY1PX2wyLr9GotclJthzzhQTxaB
32hY7H8yqNr5vxGG14sjQ2rQYL2nG86IWnDwinRK8M1Wqga+PFUEKRWfidyC3MiTiPN2K5/zcnF/
mrP7dKxLtshmK4Ch752+eFyhnSA3D48Pu85xsR0fr8e54Qy56N71kysUN+TO7RY+NVcekKkjKhim
D0TBnikbVR/sKy3UI9pQI6GqTVHnL6SOZ2xvKkVKkb3BMzVNybkp7DfJ5rNqhQet02ptkCxlfU1J
Yn41T7xXU/rexnMCXl76PxS5Zl5VEk5pwZIToZX63Y3/tsgn6u01YKMfecGglqZ+JNbt4FXcfG9D
jSkEUR40tWoGMYSA89vT+36y9s9nvNds5z8RM5FZhbUWvzoiAdb8PPHg8vU8cFnx7WXOGRSerAy7
6ofdINZRXOEA7i/4OOExrCfvB6dI1tDVPLiDnnicR8kL6/nFl19lmma6OuFSgRTiIkcNsR4eEafc
OBfxm/OxOyPMUZnQ5EKEV29sV66zDTYH57hDJl3c9WNtHcpMk6tFiUcO1oYShw++cHIRZIftTDS5
CpcIrQgnuJeT9f70z1uXhF/Ntm8iRuFqXStkZFIi7ORFsz45Hxvlqn5kUFvUn7aEZAliol0mkqXf
7T9LbWCfQIo3qy1vAvT6AI07t6OVHVrDunmo+uPpOxG80xG5Ms1hEN3Zh3m08/rftqP8+ZfljvDj
1q0KITCi3WosSeCmlAC9z7BcSsgn00N+YKrWe9JtBS0oGozBQJJPHUqQk37SbyTuG0ZUZzfA5J1k
Et2ozg1qkOHjKYPqvDIAU6DZQNwuEuoQ8q2fSbcKL9DVkixPVqe0o9AYd0i8izo1ijImipSO2C4+
RAqRChNPzhkMnXzg1VkxhDQLyzH+esQhLecLeN8IFOb8uI68WIJddvwQfhqtybYcFNU08/UqRQbu
UFiRSRuEJozO6y226AswMoWhRGgakZb1w4V17YmW1OuxTn7pfeHNGxhEL+sRYMQqjgJKd98gJ+d0
qKuPvuGzOSQnKfuNKm9o/2D3p5YeF5nFDxmj2fC9V794OW1zF7LtNoeGtnFJ+Qa9aCAnzPqFF+Xy
4QfJionZY8mqqoUNrD+G9sUGGmHKaoVOtU/Pxb7jHP75wrtdTn/fYt3f9QtADMJkmpNz2PxMGAEc
lDrYKbaY7Rkk7OPSD6vnW4yHItFugStRqlswA7KrXYZp5W89nNZdBj6rIhl3Vgn3qIt3CdsIL7Oi
VkcLsg/yqrAZ/bbU6pbp3Fou+dgQUPn6DertZ52cvNB6TcI9TwlkDrFOIzEZ3cKLXeHlUTf6WKen
mmMNuLDdIXj7DnMKCXA6QyNMZzbDb6klnNwwRddChf6auYpP44T7aFu+vatxv318NHVWaKpsjGDb
tYZyVO1PJkiRFkLLypKzQN1A3jS1nwACPkuG3D8NMTOR+IGkJjarN/Yg8oaEIhtMJSsYDosI2qRC
EnYjkMk3FmSQQOsAeYi3C0J6ZvdjBOuOY80S2g9y86wnvbLScJnHzd3zV6fGRKgW92dcY5aq4J+1
gLsHEjAIXgvbDX3iToSmjlBoqxIbxXXVly0mw11IbIPXmqxE0p48n9LJ0/9FSmMZzs8cP5/2wxL5
9OW5h+l+LNyH2kTMGklqTafnKtsH0uJJ6MFAE2/874+VDG3xnkD+yUC6w0A00gT7To5WGkzdnb9N
BFg8XN5E01asEbW4PAecajbFVum9V116X63246amK77Y5e8nF8RY7OuezTstiXLDAWDHo18Oej+u
Uwal0P2cKf004rZXt/TsdfeQlHhpHitWut44TH5FnjMuiJzhX3RpIy2gWlAyrwJzPWVGonObMQTe
6577S7UqoNXwGLy+ZDQ2Sjo1VEePkYW05S30hzzaKc9vQyb5VnR2n4208NM51mz0dVGLcPL/6O9M
yJrXA6BDbyhbbwR2i0HPMn9P8hWWHc3dN7BzxIMBcJxwVtmcUV7Sso/vVGfznvmKE2iVF6G5RMCI
UZd26DsjraYo4O4US/GG/CiYTP7Bi7795rzPwLbxlr01zcsGViRz49I/udd0T1CTp1R5h1qTTgqd
SXhfoYbzBKgfS7yCE9J/sPl8KdJfs39nUzdaWanAvpRvb+Cv3OXg8Rq4hZWO0s0YoylGfD3Y97kZ
JMiY8FxOFPhU334qdE/Rem/1/3zxykCRseeD4jHjLfdrPJlYs9Wv1+hBZO3ta2AC5ybxT9nugwFi
nFbavjuGlXysQJ1dbLNvm9aPJGoQxJbaXnYZvqme8ZYkhwjPAAGL+3HLqn9+tPpw1xk9MSIBmrun
s7UorOU6zRIJHn+BXJelNAAQVt8cwUrJkV67k9XbDh4IoQMxPrSUQxVWdz7z/YxgmMi19TrASRjf
/NplZBXmZqpIMN4ShZkaDIIsaU3n/ZdPo+PX1O3P9F1ejLfADS5+WPvsv4UJAZHlKyOWdKP5/9nZ
juKRYaWbxneXwHGsuu8i10na9/Boju/DOyQdzLVM7nkjf4bWhZIDcXGh0Sigpngt/3W3k443fWfO
9rq80O3Nmu+l4EEvsL/REK49XT8nT3P/uOvlmIq9QOytSio7rDMbhWQEBEzdVEB44CWk/+TmCWXZ
w6CaczqV3Qd7jkOnSgoN7Tg8olBJ+ak977fVbOdVheMQAtDzJAQnuz+3f8wCUXMzcTYHSISds/QP
XUfFqmw0dZOPtRD0WRciQii3SMesWrlXGbLqL8ouqiKnPgqk8ei7rbZ/plAjiijhQF+V3lROddP7
Jwa+XKpV0cLHrRfxTY9Fs5FkZQpxxznXEjlseNsJyP7RNKHhUKs05caxVuoeP0ZVqZl8DAwt49QL
bOt92dRhSKJyfb0A5aIwxdaRFa/suF+8oa5e8YPJIp0aSQQ3qm6oLINX7aw8e/uRLSExZEjN+wp7
pl132C1A/eXZS+S6HPrqwIPZWrPlVakkrp81Q5T4ya/yFjyFgSUxdbKzGTsvBtz6+BXqbiKSOzeT
ZA9QbSu9BNv08Rg+/6V0C3C685SNbJvGHyf81/5LmY6wbjlorvtCiJV4x8ANe0UZZtMsTiTYuhtL
gg1qMj0Ltw8w7b7AGwZwILyNfgoJID+ycd8rp/h2wyiiwBCSDQT88vu4mwdAKR1UOYRkpng8GH2B
AYD1n56YuMmUDfavvX45xGEiixGU7Z44zMh67IQ/WedfUmjflc9y9kBM206X+JhPnAT3k/iAl4O/
CQttAlh2bdujLbvtGT5fVvMsdUtEjMS9aVsMJI3bUIEuRUywVSTkjkzuMb8oySykOjD5wv6nrJW4
muJtA0CGkp7ik7iNoHivbLYJGRYjVoTuGXQYty/Hcx7AdQjGzZxi9DCYhy+R83OB1d60dH756zfO
h0qlnmpcH0MNxyzL+DpSGTmFCX08B3U568rDV88FMBReKI7T41rEBrxcQohrwHYw0me7ngn1h3iE
9NyIT9VTyF5suREOW8C7OJDKAYs/GMUkJorkno4Ll9K4i31Cd20MZHiQ8J0cBF4/AsEGBSA2XQF4
5ZoTQJsOv5R1eSpe93Hrv6a2Jy7FB8IB13BE6nmTjn7xlW0bWnBr7eIsmZ8FHf3XKtJatxgrLwu1
3QqvKtdYqHHYN+0sY081rbPCH/jV9a9TgLilNWBKvwzx7c6s3Fg4fi10CaA/Oxt2dXCIKoqSdsmX
KqM4HMdeAxpwdhDneG7qBd2VuEKbueJ7733NX9IDPQFbK6ddvkQkfaXa4FPC3GCIbOHNmwUIg329
QNjJzmLS1kC+oy3p4P47uGrhsb2FHRqD5/GE3B5/t8m4MtRokdCmY2SUM5Qij4rSKZH9wAqlzgpP
PL1HkpViJIIExID94ootI1vf+KGjiH1tqn09bd2669YlETz0y8vKFvyQ2ZI5KspkwEKaKfMtFK4X
tgrPq0HdP99OQWQqdA+3o7ZnLTedMplc6Jq87xGA6RZrF/YaTqMqI8tmEKPHA61OGzwXNU3i8FKI
SNB/TZJwjJsRvPmQavkWR3a33G2lx7i5aZeRxYRLHJwwaTcUDXAm5DLT2QxtN1OFv/p9BysPf0pR
WDwssKOFQZBxWnLPifxArQYm9yQIioneu/qItpppsj6B3qwhNi3Fp+xl7fMvnI2caGqTW5gQSZLk
IfZswQWCaJnYyFP2Rm9i9w4pYhAcJP1/CF0YFw1lANVvbns+5sbYBEOD/PExUDMs7H9jefHZK8j+
MxKqFTOaaOtrIq84YQwnwTaQOA5upMTA0gvUIAJjDTv/e2qGKm7GQj49FnXJ70s86+kIBOdhsEL5
sAkPkQgFUVjQr/jRTpaWN9f3j/o5Uct53upYcJ1NwXCBZMsKoZDFskjwzLcYeZenW2c25g2FnLPl
yYn9L6JWC8WN7MBO32PmHuecFEgmPZGRVERnS9rwkCyyh1Yg1jnEeaICjmdFa3qqvLSBpito7jRV
EfE9oGB3IzshiBTuo5s1kdZhIsyiLmHFw53LOBQpCbZ+mkWTGJfjy6gcsLSKsEYQ+gtluTmBJTOn
Y5CG3TvH5gFe0ehcC7mwtj66F/heMOJr5sF7D5soEuQhsmZZTWZJBns+PBIArxqZctrRogRGgBVn
Oae2VtPjjJ/iSnsRX4zANZ9FUnMhCQvGOSKDS23C2XLogDb18VqIfowhWZyChIlTkxvZE3l/ZoFH
F7lGBi1KhpSRGpuVjVoucmYbj8d32wLXwRn3btSCBeiFeJY8zEvsFaSFJ1Qxnsqhcm3RI2hFHr3B
/BQe7Cv1yFUvStMKlkzXXfVMVIREFp0i2vaINziWTOQqTlM/cln2tVkKWksYpejjrMHe/faQQUpi
FZ/1tUrkVjfyb2SDeAAwt0ATE3y5jlDs3MrAHeoKyvt5u8exKTxFC1gDCV0VfxlvDQMB4V9MfRK7
5NwhIcmF4c4tauHIMc8bOISxBfmueDdeG8nkfamKmdu/ASrDQra9PySJudwWGGiAB0UDx+j1uaVf
pWcmTYCOVxZwZd94KZ56H9mM9HLvWr1mxAsR0JnNpCHhSpnW7BapGmI7ff1K+Ppr0P3frNWaXM7W
mU3PZSZMFINtjoHfHE8YnhOJoe+Acmp8AvmevD9NSJdMOzqRFwRYOZzlpvCQt2xwWrO+AniYXsKv
aHHmfGAE9JA7CSnoyxmlH7K280wDDPWty3vZLcZQZ2UdFOF72AmZM0zQV2p641vnGD2fEPwc5pML
ADMHMlly/9OLGg2kV6q8j0yeXBMaNqYKvKr+7YyvbyMU5d6CXZMJcWArB20I4kkSMleB/9gDoXta
kLYdLqHNE3NKs29mKsKXk1lVeav4kP45xyEgF+rvrDjKGi1AJ1MrTiDfRUJqSiy9Pujr6OqNoh4+
NftJFdTsuV/Fmr9J1JRdKfs7zbgxf0BhVEfhqebH3rdrGUrtLMaA5XrESWSaAzE3xngrjDF0ASAY
faPMulUhXRY5KsOv7wsxsyKfcBblAdegiBCgr03dO3M1IMbu2dQ3vX7+W5QP2lDzG9ydcG736FDA
MToJjECBa+Jt9XeVi6R5DIsYQOwiyI8o1WpR369XPk2dh2yh3MjnG0X6FgIDuMZN5TKv9JjfIgza
9xsYBJA5hWJbvl7lau88qIrSv1P2CfjnUEw0PFZUpA+p+dnbNqVNqGbrTQNzJIAEdgGf6dSbLWZv
kQ6KHFAXbXVx3dAyOWF2GZt4OAuGUV0WRKQdiPo90zWpzalB21ZVmCT5sOJ2K0n0VJg2Ksxtckme
/g11Zxo4Ra/jRJUQa3prw7NjxE7DQJCMAka5i867k1fnldqwC0XtvcbT7mf8QEU7mVRRUyTpTGOg
BFPm3d/iWZlADBwzn4lwRxx1iPAKQrl7FSy7PDTYKBmZ9qOZu//SarPFDlbdzLGMEaVB5MSijslM
dDfhy0CbfCHjrvwjMFznkdh3LLldfr+x5462vIf+Mr1VNnHCMLwdjiCxFhMdztV/2NbRM4ZGXZOS
yMVULNS8weR7gMg3U9lHzQBkm+EV3KGvxflRkJ8cGtx9uGE01IVmiIC0lbsLdLiKG5XV62ICBb34
B9pHZxpmtL0VWgBek6gRlrArjvvXe3rd780fcACArEIAoBreq8KCezgs4wp18g4DQxYTXd9KW8O9
QVqwTPqf7czX9EbF2SFoKjEOpjHbjzrFFUIKzHnGw1J0tw7P6n7eUW35B1FbHNTiGEAa1SJX/Rj+
SX7iBqUuZ+HqGJPWkI/uoy0Gsxf/QKyLVwtPbZqU/e+QfpumcQvGh/uDqvEbIJ7KUUgkBDVL5wv4
Yi+BCuFIh1h030+QxZD/rw3QLzOl9CmyQuITCdCym8xfF3TCMc2EbIvdwP7NiJ/GVqjKWZ1ckuEr
d9NGsm1JbLIY01V/0F56LbojcvG274Iuv7k3/hjd7jKMEm8nWNg8do83bWoaCZZKplJtwoATrIDL
EOH2LkdDkFw6in0fS89B4QbX5m+BzfjAXR1rMuQC/V1bDGdHa8as9eGPdgqq+QcbBQ7WBnKFpYzI
8Z2Hmx7H7FmBYUjPz5zt5SyxpLUqEiU/JqFwHxKcjWtN3ySHNAZAaBEUShiBo+yIgOlnW4ZKqsxL
lYB28frgesj9bRuC03TwIgRz7jIosvGk47kgQ3kYm8JtUu+C6tRii5bpC7GE8y+T7uG+F7H6GLIL
DeL10ApuX39esSYHBxLnU4/NiyC3DHpdqbZDlBC2wUGVrqqlsW40FMERdSIxC2sn967rTSCN9XDj
1YV9tPsXkej+/vYPKpHN7aRHNNzS+RlrvqWZdXXwF+kktEWSOb76/1lG9FdgNlITYxwRgW37JPzv
r4YP5FUHWzZcHYjJNjBinARVltGSinXhfE6HK6G6Q6SJl+MLuhjaRhLe8VN1m/8heN8g3YCgEmws
V+eZfW8eTkGSxgnbx/G+MNkKULH+e4nmeZ9zzr/V1Jc/CutNArsEZAEItULRKTkearOncXtoQxnT
E4Qke9fSClf0sGmI6OEU4ZQKrq740lI/2k3/lqnFr3w7TczZAEZvS3SgIUs9NlXOW+LeAnfNrhAH
NlYRXLQyH8voo1uCe/VFFtjKN1WWRL38zpdWG4Yx1G99VQBEGbqYKGGA7Pbu61s6V+1JBnnLE8yR
moYAXzgznGo21nAseMQuGCLI5uJzKdLFazl5avVPpiQeRrKKa6hZYPrxjwtiMgxado9QsaEIwQrI
eBGork4sSuKBrE4OY5ndbkOAK8mBo3QW6tYDjG3i3MhNFSyXMUUcslJpXdnbsZe2Y6SBsJlhtg+7
CKpr2w21jcnjvRMS4OgUOiXkpzEuUy3wrS3UQDIb2TE9oigDboEPlRCoJI84OH2xnJv1PESzUcuZ
FYHaeAI0kvh8xZ30qrELgLvD1CuNbK2gXbDiAWOHmSjJQj+2o5XZUE4/aidXgn/rjHzvARp2XAb6
lc37RUsHdp7Y7X5g0tw0y0Pz4GSO7gmlbOMoLpdnI5elzYcwZOsBY1T7dBmWaU+hhnmiDPSQDKTU
Hz2UKs+6eqRvmmDC5ski5vF/hRvGDq9oYcxCNYl90XKkql+v80ugtp8h0lxxxO9pM9QrbxyzW1xm
1WX6quHSHdf+hEr8Y/sATpYvxK9RojIL+joZ0ouoWtWZllh8wKhKpHqveRnl0BQTgxDkyX9QviMG
42ZUOUXoaQnOGQ3Ahr2/1uwLzJdiOnq3DnmoHWczkLHFDQ49YOx1C4YIsSVq0P8Qg5M776lbF/BB
WJssPYni8bNMwn3dK766X1luaopghyex0uJfVBqXlqwsaxbcHIZtvCvxOq7dWHIoE7qQuVngWElo
/BC6Sst4VoUhCpFJyh6fjXkN4RZ9/pKFjc6mINLg6ZPM5DfeNHtLPjf/jUSf3og2K+ZORPSELwdb
liGI8hQ4LUbZGkeWT1tC7PueKEdbMOuNx0ktWqXgnSnHzC9xNg/RZOl7ezfH2ZzDp5fn1DTX3O8U
0zEmm108pvQZXw8/ZPTrfyyxZ3KEE0MPvdJMblzZW/EkSxvFyWMqDpVjRqNPYJtG2ceZI9mZtole
2vMVBPa3Q8eH4p1p4vGeLa28jMCpHp4SoDfnuIcoC+8FudDDn8rjtwyVIv1DyQumaB3PM/DmlG6y
u6apmJ9gP9MrX3bI92mVfMJ0VPhyXxS7uQg/mEvXkkKl/Wt0jby87bCyIg5W6Ftn776P2xrrU0j4
zZKs0XXf0efjxFdylwMbqLxuyrAXon6vqT/5Hpf9gaYSlVH1hPJsi1lzMfGszI2UUbcvHFkHP6gK
1ZgfNfqmPKkWnMn7nXZ1neS+E6vwsVKPCPVDy/u9hCUsodlAYhpBzNidhzEiuk72fsOtf1OI11cJ
Uu1cr2duVXUIO12xWumvx6KysT3h/4+3HOu7TUU6XfXLVJm1jBNH7hWzl4uQ0wFvkizF31vkU+46
zneR5o44GHiEnxnNQ8eupoN51O9uE1RSXStyJ5k4daTXLCg4Q//qVyd34Ojyq6a7V22cEh+NWgz6
KwLfItjzcPVu09o/6Mfv/W0V90PH5MLBhFvuitu3nqKvVXI09zA2iZ/gk/jSNu3siNW0DGmyPu5e
frW0N8DATLTmtz+8PlYkJRwZ7onK0x9McyUCvMPzhoBnYH+82RbjQoQ1raKuJ7pZbr6DVp+i1VpD
GIBGhtzRPFssE+bS+hDg66WiWJCMC8SfbkoFTVex20lmECA8lX1LxVDIZMLI4wnDNL655GVWE9kk
1tTjQ2bk6Zd93gU/eWpVM48hgV5yTjE9C9xub24E2iZDkT21G6VPLPrwxo6AyX/dLJKYvci4VTAd
SKsaiQf7tlOnkplU+sITzuxcO6VlmBwQEv11Xr0R+KO8KzIIjWTS46mVeZIoePaSrVnaWWMmqJ03
sNyzW32DtaU2mS4lSGNVhQh57VmXDXEw9KQ1GQuQuPV83WnL6z8TOeCAooLeUzArr/Dddr5UlQbT
p94EK2WDzYw/TYjQBeRMFLxDlv/z3mhb1CzEJ1TyeQdE5oHzoNVB2ac4VnuaemXTiOXu1jhokyrS
TufFDCwFBSw2s5JA4M49sKiwyNNSJfYE1fuOBs2fYwHGadIDxp2I15FhYhewpqIfNUvYf2z1kuD6
/sOcUZEr6Aos6tNAlvpN+WrUiEkRu4CG4zHUbJ+oOaschFxf7vQOP3zcAlaROknX3JWzAJIPUHY3
pODI6Zqd7+5PkWfg3xmPg9Dh4kpQgYH44c624eMdOPnm9+DiSmX9UxrifL35RuwkaRgEjOBhtGa4
plPk0opCiFk28wstugK64gTj50ytBtWqPNe+olVkBdT98ScIEeUdQoniqm+OWEewhoisDgaKcJun
vf5uQUSjVYCxcrrXvbnlSXKjBS5QzcI2H7nX2eD32pXtVXmoZQ259Y8jMnKBEKo4aPkZEbob/lMF
OVU9+jVARjFhl+3Q71E4FxRy5h+Q1RL231Ift9ClwL7PKisuE61SIw38ly8Z7en8le0lIIt8NIst
Nr++dKSuyOzoQyw3qg3NQPQnq07uNPBPbeNeGOGHvg0CeaEBgWJTibWwBBre59uDSIHjhjgxQCSG
lLEKFwBQL+XbA3QY2scAq1IKOv8g7kDVaJpBQ/v/1aLgBrVohl6GdfsZxL3/MuAsyE9qlN/cD/sI
xN79R9PIXsNmtkX1RzIkdEMcb0M104MPeQY2kVCaGRJttfO88A6fUw3dx/y+fXQCxII47y9EC2ig
Me1ECmCjuNc6PWUchEwH28hdNU98yU+M5vskEgY0QyolQYYPTvJZgNIcv/31lVxmKqodGWi2yHFD
wSy8OvFViUrxKMreLDbAqa94CsB4U2yaHLcgFjmrQVxxhAOE9S6IrMHPezH303PgpBe3mCHhjzoE
gdTB8C6Fu2Us4RtyJnqvXQWjqrDzKE1+LKT8QNR5PfoySq3qVdRcIwZV6W4IKD3cDKMnsl7jXIzO
F7it1ZrYoIo45igjRDmB/8OStxPYUvkye29yBxzPLOtD0aZKxPyE6fgffc9H9H7P/XBcypkNT19j
VatxF54zjhr23GK/NbdtF7BpPliAUBmpQQ1RyBfFHC/Cp8ZZO5ZhsNGIjfkrUkhVec8iX+jwYV/B
tUbdhb47Fxiy2acGhk1vPUa9vDg36/0UWxcrSr3SvnTgRtB2jPGhNjk2p2V8loeFOFJ91QnWHhLg
QWunQCtzUO2obsF1R/NOtWW8nXp6CAykLBy0JVBO5XONL6jXZh+7OjtmN8BnWuzDjTsOB3K6WsSZ
Gqrb4C51HSxihYHOk+A+Fm1nlPZWb/UIxLfqzDkuePsfH1wpNFpBFdIAZtvdtF0r9YXyMCl2P/Lk
eJ9SLnyq2NAtwSqPfObJSz2TBS+6Z3W4QRks9syscy3sakePZv2Vjm1jJP+CmJmOp8afyrh1VgPt
t2OqcCwMLdgWn5KAXjSF4fiUhr0CWZijtvRUhoB0yS/a4gakybL2mgR8KP7ezJw2nQE6Z5Zbkrd2
0zL8d/jytkUPTS+g0E4Oy1BtU6cG5jIqIL4OFQ8AlByFcAxcAGe8BUJejxYGp9Hgt5YWST/GsK1I
SYCsdFX0KeY1AYvWtUPzG05Ar28TAhHCJqB4vILyoHblqQ9A03e8k6Ju5NekYS7B8v/ij9k4tCH5
ipv+C17or5oSDXsBYE8wiJTI4alOceb3eo0RMG+HHaqGa4HWtwAbuUvhyT3pV7IFO++xKiLueI3h
t69iP5EInGXinK4WEfUoyqXSV8lgZwu2HLYnJG4wlohIuPebOtqCJpc9i4PcLBzT9z1RP+h6FblH
qWBd5Sfax5JHqJ2fIh0JTw9WKj2+m4qr3RsjvQF8MbwqfAkFbehsZsMArhmCRMm0KwDhwRCZUFxx
7xnqQ/GtQ1PYTkJaiza8vo47KL1aO6GRC2IuapHaRpQaNj5TWxc/08GvhKq2XtD2PyzVZoGCtBit
0IIoKTGXquEtolZYuIkIXFcrxuzb+mb6WSCNCVoYJuG+WUf2OIXG0j+FDDoLevTkh4tVKApyZE+J
12mWbLHDJXZFpPzMqDqTvuN3WwNI6BHjGApRpkHGJwVIyzSMiIACcJVWXx/fVqJlCacRF4A+F3or
QEvU6fa6Ju6sXgBYVKXwOEBrVU9e1xquVXRh70TCIPyVAGCbbNn60TmxkZqD+cyN8JRko3qIjPRb
c8gz/QhAAXOZBT8Tb/pJU1Nn/DdAZQmgwJoMNhY50n6/tbjQnrmbp/Bxu77upDS+HmstkAdLJXKr
lcGxh61qB2HK3RcG1P4DmuvkbUjmYp89aTHNsiOAaC5XOSbSbRCQOrW2shzI56Q+ROZmWlzwoBkm
InLos+3PxNf9TEJXxIGFJ3SY0dnFL8/z9pIbRi2fV9RbE79XB2gUvQwD+6tyhz8PznhN0SMgbETV
MCQCEo3mon9IiYv/FCiiCyYnGBBPdDxcTS1uFSb4jUYMpU6tLc2Tb32XQOwPUf1FvHt/2YKCK8Qv
W7L4jd4lsOcuq8ZdkPasCXH8cYB7D14d9G92YzFLZhxaTPsR4zmAA7z9k59p4iR8sFXT6jWp9a6m
6k6LiYM7urrnOG6Q5TZRNiwKEip2gM96BbCxmOZkK7mIJS5/Z2X3xT4jKSPfAaLFFha57gZ5493g
ACqKovx3itxC+b2TFNOC5fH5bris7DoIyP8+RKyVV+9j81B97VnT2WonMJM2VJt9E7iOlsd74XZW
i+hAM2ON2wKFil8JWfDwWQAit0SKyXETywhMzGDXHFQq1StNNj8xUgPIIh5o13r77skN+QYtNkg4
xK13OHsF1sWCSoiAAWhUWnFGTLOusShmhsycUUovupwuf+ZY+bWrDkoB+VzoYT9Q8+ucv0SmV0Fa
YEOUt/6YAezUqDZAceFLa3z+P2pTgXdFmfT4bSOZ30fkyW9J4tbTA8P3GUsIDPcRr0ty9e388AvV
gBEFiwzUsDZvTnMMVd9XDAXclBIpvW5zdCDLrJ6O8vre8pHu38bzt4Ywwa748LDEmFxyAtR23757
6rtuDnFNFe54hNL4N0Y/vVfcRWqsQpPnIutpxPACS8HtP8K8dDnI675OYH8JQQpefPQSJ7yqunrh
jYwUwNmbXNPIrYSRhtE9G2SgBDbkdGosyRO5oZJdpn1zFLMZp4W9k5gG+/NXfKRYuvgf+IeTJeEG
VyQ79XwkGOs0ZddikrL7u5Nb5Q6WxNFss8VCs9VNSEw50DJdpDL0K9kGMQlqZmsYG5E5TAtrkzsR
TDef5tceFHAr6wD3SEfd97DtOfz0OzCo5RNr29joNrcAiG3ly6mvZu9Hp4ZlIKxLsY2EyJakIHZa
P2cjczLTMQ5Mn5IdR9WhsWUE6ExAxLYY6fCjcbhAlEz6ZlUk3RmYI5ZaSaAcu2roawdl+FMldgtr
ZRPp2YByfNZtObG9j0Lf7dKNJq1iDoMKcALTS8KFOhEJgMbrlU8XwWxMVgJtWLySG7cZ9XnZAkrp
SK3rQsLsgUTTO5eSDwY4tWjykkAZo6p6SxpX1RmuIsJSNyYYYJDe9lk6QYOexG4hIVw+jp4F3p46
/SQdHwAalMq/2Tt1ojimqjOukcz8dC8wgPYtM/olO5rjfnUwR1/chpqlVbx1vPETyaoMk+xmk4Gd
ChzljmmFpEj8IPp7YqDccPMjy7zlvl/RIHjK6FRc9rkww9KSci01NxJ1r4GPmynVR9LQJ5rSSTEH
KAtJoVUStxLJVW6nx5cWtI2d5GwGrV1goy/9WMUZ52bp+z3jAigW1dNqdXlg9tFZKBSxbJQ4/IeE
TOBnYsSWTQBfwt+1z+F1FTw1qkTKtk960G7JcJGOOb+I+NJUgNpqxdJNt6atpHrrXFOYTLKLQpWz
frjV2tumhLlO2F+b+E/z8/92Jlq4i4LQrUHvS/Opblz/b+8tgn/QSsYnURoPmTGkLyjS1I+yiFKv
QLR922a2u1T5bd21yF1g+T7NhWNFCYfAaOgSZbHpmJYv4WJiXyDgbAwoRBuAZK7btfDfkE0eoapf
hSgNPPJu7H1BSfKZ7LUZV5GmChI24LHVINSBevJu5in2lzRpRTNWGbRDK4zh9swHrZwHY7PFfNuL
m9qMjopzlqx3uh5QaCgx31ubFhPjGvkTKwtsbX7ztpxlStKtSnf97ePPV1EwVA+GeTJ6ywKXgYkV
sjryZIIjQ6L3qb1zYWsCym5OXzYIJE180+DsjCTyKdncTXpGabmuru1dk7qUkL0GrBHWDu8+7pCY
SGrImM0cW6mvxqJSQ2mxOJwVF6/klz0L5S325FmaEcLalPcEFcudFnPZnVSsdkPeckzp5GVVelV2
rNiFLYP1B6Dx09/UG7rO3gRcAJjOw3dcv79JWC0UHL3A2EDUhIC+fi+s+S9gR/kHZDZghbkU2FU7
5PbCPx3yYEUtp03EfU/NncIJ2gehrh0/6IxJWDdtpEhu621Xj7sSkZt2pcEDbdYKyIv/fSbYc1eT
dao9/bZ2GGgJJrDRFdSBVteW+7Ye/1fkYlZWFnkg3qDmxJdutWuXjsYf12sL2mket08JVRsgoIgH
BVQYCUCbjgfSLvmLKNZoOIOG/BjjfmkhCeW0v1D73AqeOHBG/Swm+V5LKl+0cqRxBiYIWjrIddFt
kW3Kz5A0VN7+8mPByWsOhnBkMdqpv0sgSod3bFH9KNCdTuHKmsITKhVw99Xjgl47F7yBBPyEuYND
mcOv8bqFIz021NpOoCPiFT8OLlR1/fo9Q3VpUA5XbY0upsJBeOhc1NrGVyDK1uDcYUE4vYT7IAR1
uxF3jAWLErB34MWrVvwm39jXgomdYAEOwpuBIBDVXsNBAA3YnP/BOuN0ZYM2/POLquvh26Txrh0t
9TSqkvOWodwVxGy6zM7vJyLlfvgOw8wMex+xoGI4HT2S3damt6ZHcMNQGO19AfJtYbmUeJKSPDoD
wVsKoJTJ5ZHOaJ6i5Y5MOJCF7Y5TwGwOxle33p1sLnWZEYRau9X0+TrNHtu3lr0hlQPDtPa5Vsl6
E9XDQ+0BgkI+3cGhje6Edpt/aiREwVsVsQJYzkhIUtRCnenveC3aaTDpzoesQNGBEOMvHbBgv10o
oOWUZXOd0/14qza2TRx4UOi57egqV7JytlgkwcRulvjPNAPEE1JQr9OhaFToon4tW39ABzvo7c0J
1P8l8ugKy331prNhbyP2ihsFJkF3BujJcuxmUWDbBYC2LtQfPmItrhAF/78zr6YnioUO6FH9To2L
kAPzRJjytzPITmVuINtxBb2pjtM9SDPiOS5pa4aCEo635uuyNujhZQSXao/uOo8tqslhpIXG37Bx
Or35ol53YCAkBiBxZ0YhKbZ2o7dad8fgFgutcYiZJjkr3866REF19H/ZmrWkFXPma4YAJkwjjS6B
RADSam8JRPHuOoxYUdC3eKstYDvl3fwiC4ccHFkUIild8smFFQ6zlXtk0hQ77Sd1GaW2UyiXprcl
QeJnPAXY/M2282pVP3WHVeDvQyoefMMbcClQEEDpn9AFheRBhP+DGQittbL04PGaLIydZrj7KR7q
vvs8PIszSj/LDKrFnvwWbbTA1YPnwy6VZM7Xzz/bIlYhWkSN2otdXfneTwGuh7+qPYA+mbLpTrZG
LfGNu0Gq5t1uNt8kFNQJgB5J+JYB6/yvZEc9FT3DXgtFOKBxhZbP0DXDGU/2blO1rWXA0w3YZHEJ
0AX8IapQ6BfioWFr77y3AOQkqjkcr/DiHFO7nr/xLX8cqlHQ8xcSTa1zGcSkjYwjPrQx4vu42KVm
VclQoQGGYR9w67FbbbfnU0xfHQ1u6vFKZ1zWSO6mDCpGbxidv0C84B16ARkty/T6zrvaZcvVgym/
s5WzyBZzDbXgmaGs4qyv/6EMEAZWBsbeN6aeYhPRBv5MY//tT/e4rCEQE3HOzwjaY22IXbdqOT2t
Bzia+S4HadbLK20L1Orm8o+OlsS0K+6fx7Aab+mua0QYn6929wDdNKNksU9/e2FUA/GVHODgRrdl
CWbVeRnnf4dpKdj1D2QGUyosRw9QuCuCpq3arj/do564a99F5Ck2gf7d0xkyzhz4FGfEVNZYzZ2u
L5av3n5lEWrlmeBDro1/WJsMzzuvF/ImUWYz3Cv6OxNOsiPmduzbZ/NjoxHm+vrhctMtDhv4eZaY
LZmGPNg4NE0J8/YUq8YxUyc8GgLLjAycWF0pujYnpWAdD2xsODAIVHtCFLc1aHcCa37H+OzQemTr
68fsXJp6WcSS+xiRyFFh+u31M6sLik2wwXjfAqXvjZnyw3OBaoTPkPJqXqxIOtUc8DdtNNhyjd6T
9pfahYFnQl9KSA4Nl3bGD5Jh0VSnjUXlI4mmPD9Hhrj1bbtwukGVtNEb0BqYYpXH22Ea4SkSxi6l
7KpsD0NQRhZ3Pr1u5cnj4tE0o0UMBkn/T3LiNVK+m4evPUE7KvUO95vXXdL6owrFqkH4LW41l0n7
ZaZOg38PnfcFyuWwukT4KZ+YfZd9f+rUB7b6O3GN1ld+ksa2CZpSdpEYZwtBI/+wEik5DJR+vMbT
F+Kg6NZZddEo/xuTVvZoDPuUY0RWM7gmtYVeIuzfLaFnIxWQBWnhKltk+fY9BAcqyy17AcI98YSG
ftvLJYftN6OSQp5ixTmH6NmcybK6vZMq7AywC0zMv5DfJYLyNYVmaS44wY8o/TPO19XJXrD8abWg
bkMeJqAPMqv2HXP0hz8QGNTsP8G4xrhaCSQbMaiXcT8ZhM3ZtpAh327q4VkHa6TTdaQ2Fg2F0CLG
0kE09v8519S0qTIPnqpeCMVR/3gMGgvyARm6kUMNj/CTGSqi+l6+8JSj5W4rZ6NLiDYtBD8/ca4l
9kDcgKGGPcgnV/Cz/JT393INc6V/kQlo/A5trttezw/RJ2Vj7bIvJKYTzEYElhGFgs6i1E4A5m+/
A+X7pSf56LXQk+NvRKOsv5t7xBewgOZhr25PQt6saHLxvgU7fefqH2WpqSlN42JMcsx1GWfRdrN2
Xlp5bNfEtuukHlNQutDrKfrFJ3oEUX0GP64ANSTJ3zqNMm2kHCydOgYTf70azUhcoeTdIijRyAAc
sATwydlizMO2p1KJ0+ozMXnrU9GJozXVMZUc8t6M2sdli4iKr1OYO5CmtyamDEuUHbMc8crVXjSK
nPn1i+3J3+ZkZnbxTTUJZk9sf/XIdfOSP70VdTv41iDKEe9Od9mUYx2nZC26kQ/8V9tmPMhfCsFZ
2Rsb59/3xwUEmUYs9xVSOpgC2xNfGopAl04t2jrnKO2mzIV5x4X0vWf5n2L71HllicepDpyXwhwF
1HFJZI/403pKj2fxqvIyJjnR57H3FLIRgCT3daMZbH7TcrWo3Rsx0/jI6lGvft2yhXAXzX77bA4O
p8Fd7B1fRPZNnXlA56YY7ziwxnT6ed61rmnW/GK0GDEnuCvuervHv1TC+zEY2Nt+YFIi4zi7UrHt
I7pXxAvhymB8nXE1JGJWcaWI7FgKQTFdh6Ih4iczvsBzNLOZcoVziioYyApHb+TlzYzbcQicFgX8
sUu9LRRw5OFsvy6vR+24XMjNXvuPnSkbdDGV7O9aYcEBahH7Uzj4C2Kng2VEeCa2XDWXjAsaQICF
piT2uYowX02p16rJg/CnHbMa7qjVF/U0Qjpl1nv70cPlO7eF73oDk8kInVYu0xxqHa42RBilyUfS
VC6d/BLDWy/mWZXCPH5Dx8ET0CmtFpYtw8wF+/LS1wGo3Q3pd5aMOPxm4SpZia4At1KpExZtVHSR
X/oTLpcDcDpgbYWXLyss7KgnL4mOc+sgpl+Vj39r31T+qHMSAkFRVzZ5jt3tJMJRJ5lgPKt2mgH9
YA6et+azClbFZVhc1vpjGqQ+6w4yFRCr3EtDoR6qqa3LJCHkglI8fTNdq5mbAA8rmBudOvZUOpZH
nJbdb4hHqmvOUU/Kw1444j6bDIiT+tAj+Fvnk8vKNyWumbAoPelG/WvtJ0W2QEgjwI6f+sqVpql9
ZMXG1xLYLpXBnjhabbakCMeStmc7M5mpYjh5m4o4NpeBqXwR04nYxDHW6WRETYhZ9aAiqk48b0To
TSaCQjo8UEH9PkItr2cWnq0OBbGs+cKuwfP4IfiIGcNgYNoHrzhA+WK+gMvDCPf1I2W30p7yielZ
5fdJIa3IDyBQfncx7ML+8aHMXd3g17Bafx+v8/J1akP4LeA4JsqbGUsjeKEgnfeHbFde2G3/Lqeu
wf8vEQ2X6aBKLFl2R80RZkrY0l0cKLNWAcpUqRdg67XAWdOMehM07mqEwyOkj/bT7aa+slSuMZ1z
tR/I7CgQvHXcZRvai6Ch7R25DJO/WilgkDpOSOCeGzqNH/mA+3ARnDLEbnZW55opBC8Vput/tRo3
EqICeRjnYEi5zhIWSWJtAPECohKuJ8aWl9jT4K/ewNGR5WUOXmlgX1/+CDBhGoY1gRGtb3Q6yY/k
MVCnRQg/siwH5UbmcAS3eONyqGbtw8NZ1Cjm6rnZggmK1LVfBQ5a1LxXKm+S/a/lW+Hy3cfdGDfX
FaArJlUT2V9HRo0ScMyQziRnlxcmC6i9zIOe1nF8ofp2ibM0PXcDRHY15LRBws2Pdz6F7PXnXJcc
8vYmGyfFeqIwFgOtGOWHGnseKSZ1WHnjsUQCX+V57ePUn5nDchCplhwEWDE8fLD/Nmo6b4DBWAoW
tANwi01MX0PmILJH/njhYrFLJXZ/EulzVDpIjMaV2pF3NbHq7VDVMMOIqGA5MRsJqLiaDpM++4EH
Ym1jvI76UYuyYFlrRJo1JcJ65GYsygl3TK9oJ+ReafoTON1WXiHB8ezgo5tu8rRoy9PaeDPcf+/8
BJfrm85cxv0kHy/71VSAswOl18KubbHOd06dZeq7su9JRrSuIKffhgsF64CiKihUfndh0ZtLs/P8
pXlFpXaEymhgA/cE0+l0MYZ6/mD6amHpCkbXCly0eaWLp7/d1qzwqYvVJEIaizUUdJ56jfEXU/tG
6JU6s5cNgD4lac0MLVzjO7NFKAs3Py7bDEc39aeagcHt9zk0F1zQYspVOMeEOWXVrTHxj9ux7kup
dZ6YP9MeQ8HS7j2XLimQjEKnFruDQyCKXP7NjRZQmVID+M0+0pnNpEGLQZdesBZoc4F9QX+C8s9q
YYBv0oVRYoY0AacL3qtLh2JSnLuoq+T4WboHSrTpbEOEGVdumq4rFlUG2JxaFjONg7nYzKOTNuWx
oQC9XQfgD4MDnHJXTMvFrM3gJhkKYuf/ykZnvXswPZAaipNqzM6Zsc8CbmWfkDXuwq0pQCv5Rx6L
b/uB8rRUQ6Pyo4rLyKAg8qpwIfPGlvPG89x858hGmbNwgks3NDIchnrtm1TdaVIpVxECM4jAQGgl
CHPCcCqlN+msYLlZa0yn4LdCHAMXKakYg26fQEbBBX6wOGlJqRe8XtOONh3Pj1nRfqMD5vdXn6sa
Y8tghMzCRB0TWLQuo8TFCvMl8Z7lBRkDII5Rl5jDVVeFWgM9VnPio0eggXkHMdCUjCEpRqarkemu
mBpGzV6FtlJ+hVJjTxupnOHQRk+YB1uz9/OFtY4nrBvWW0D/MANrUVFpsgL50CFHKAbBhHNSx67f
A4tLaaMIToQB9dJ2ifv21AG6i9ElIfA8KDoIdpUR0Vkdr7O1DXXUjGtpLxYtrGdArHX97WcKLqI+
mTpkVoIKeHNJH9ktH7lFlXEZFnZWbUZ8XJdu3HVU5Wo7leNYlRhcK9nFR5h6MxAxR4mrIqxl0BbO
aG5MQpX8X045a7quCwE6h0sSolZ8nvxHmz4wON8C06v2nVNHGrz1GJEpxTmQLy1B0WTp/q1C/D7m
B849u7P+LVSMKB2RZoyWxjAU+LIiJYbg2Rj8Bc4mo60Pjgk6K38DUdUYrNxCov6OmEeJlpRc8yjE
FaU4VeIgmPTjyfwBMcKjHAni2bm91xWR6LlhV1SIWf2W8UF9uOvmkyHma4VQYFFYKs8MWItYRCxY
Qg7MxdY8HmNMZ70HTvGlINcb8FTD1M2AcNt3JIPhTno0Bzoy/tb2GSYMWaYgq8qGWIoknx8Ld6Xv
7hIsAcb/CNJoJvamuYU3JyO0ilRz6HEVpJPHhfLgK3ygZEv3EXFCg5uod/lND8cFNkgiF2aQ6GxD
oCa9jUSi5rRlMCoUVb1ieqkss/SDW0PcHdFsgfLwC1BX7MhxYB1SH1AhVykWo3kgih2peCb/jXCk
aNjGJAyPOKWEhsNTPLDabQrSsL0gjdd4H8QKUQSDS1WhE9qIP9jb1GRfWLhOOUo6MeN712vz/W4O
Ze4Bfuwt0iT24rr2QPsGlRrNYawbZz3KaGzr6guY/iIncIA/h7xFoHUsG2UszIWlfJ5SXYK+vyEd
S2zz2DxYL2444SqUT4R1+gOpiAq4u+KKvsCXjwYu3Yvj5Iit3hLeP94cSRjZNcZp/xTupcfJhTgg
9lYqFjuP3nsX8utMZtszgtS5u9OcWHdPgAZshVxcyQyREaANx4HhQ+MXDBu26Cv+bZXOv4IO4MtL
vvHlZjIh9QutbnFsNzIGlsfiyTQft3UEUYFTyJJvbGjT/M07ssLeXyZ3tUWgE4WoHCFQw6CPIWj9
+Z8AkLWntANmQs/fJyImvMnB3iwxRx/fOZKOxwSvFwZRWDNn+qHCrdhisYqvWDSdILFva65rxbRV
P4X9yvMOkQsncRRm/EBa/KFLptUKiraS5cOWcnpGqreLCRSQvM4CU2N/5BoMK5UZSAlf1dMhMgLM
qVngrvGhmVh66L0J7bzOFfMDC8G+MfzXX8D39XZhUWuWNErKKBO+wqvpxFZ4DweZPH07Ho0GAQ1B
ENjK7lIUTWpaxflx8lK9i4rUwCwEpYixAsKDq/zjyA02qYuuMfJI4fg5JwpeB7ZaNfTRXHS91I7a
iWM63V/lNVfNsuIQNLquv2xZ2EgEyzRGt+9LEb7QvBiZHf5zTLxZqZw9wBM/GNyRaMg5f9WQWDJh
Ub5P9SB8rV4KIZ1jdYB0XZsS/ixNo2kT2xB7iqyI6u8GB5LHdZlrNzeM6NhEd8Fqxfu08qMqdJb0
aIsuoVIaXJXMLZMyI1qQiUPjJX6epeM5gJfW/LtDVevf1fj5uWyYjUHwjbirDBAaaPWhbr4I0Haa
UqiCpdnhmws4jIN+We1ziEZN2+3LJ6snLWSs5obE4xUaGiqntvG6DdfmsbpcUlrGD9EG8OLT17B+
buv4hWxp2xl+F2S0s1vh7NC3+XYqltAlQvucGycb4ISiSLdt4kcmsgcWBasd2d9DlRdsQ5lUkJ0t
DbesPzkOVRjkF46wXjeGYF8omBXze5pcvY75dd2UZoddBFT1OxfnUvepL5HvunB/jljcuNMVfZqQ
z4EkAuJJwZWexDzNzqzBjD49/yUi9AwOSGX6lAsIsqi8lMQ8avSD315/CH2da56PIN3i0pZuHhVy
pQiaCOUjKinF1HCoaTrE2UIE2V4JXxmgg4RCdwLjGau1gzVA+ym+hURebiQGOsri1gpZvJ74Sy/t
XzGlr/niOOwmLI9N2VIMequXM///4NdBhzLFzoCvVi4is1SQNjphjmfb4xCt5FUf81+HFbFIQBPg
VztUvZfhIfwqAveCdniEiBfxdVH2Qqn5BF7dj5t4umQPvlkc0lX1CyrZZ5a35t2Kf9dS+cruvWqg
tjPuVUfqkHvAtifOPMUQrzm9lKBd7vyLZewCvS45EI94XzxX/CvbE0cs6ZgIN92ndtDnSS4WqBah
cHTwNjGqppVEc5ATzHvsDChmb+uG7JIPKhOe7v4vXteYEXSc8JIb2BmmB9XbM8koUe13o/V/5RIu
Ab2Rrd2T0SX0USb5HLUf0M2dCne7BO/vEvCF+C0XnSqegsrGiby2p2ve5sJGczOO0G9oG3J0UCDK
YJpE1mPK+nRCUANpIf9sLUgOV1XQfnm1Dsq+8VTJOKM9Wweb96A/zWoGS8SCY90cKqAq2+TMQSoA
RD00SDEBNrzkR+HbFkDRt7htmmArfX0GLxwdfO6Wqfd51AadkIc9XVrI078o9hd1+gAuSm2PNw8W
fRtlZEJHmQ9FXSq+6aqNQSSrEA2YaPI187bj0AkznmgcmYNXEs98ySvekLhlegQQ8tScvunPKWS6
Len5ElJbS448eES4PV77MiCMkRWbLVot0i7U/tGA47GR6U7Kpr6WBj1/pkQ9b6JuMC9N21LMGJTL
REoK6OpIgf2KUXp0a6CcpFaDsZIEbYNk5iu8nSrOL9m9O0kAv/lFrj1fO/8wJYQWGc+Piv7mk31R
AGffkZqqj+hOivLLjnUPDgMBjbDh4iUNIcz1l1Cep4TR6IA/Ed7KIu3UmafbmAdHjQhJbXTRczgp
u4oeu1cucneeW6Js7zvgPHqjZJjtJQ0fXWEHg23vePVWW8AiNl/CkNZ5Xhch6tOfhVg8KiSd+GZu
iqx4cdld8cnNHmiQeaWN7vDknXb9OvMfGbZBE6BLYN1tOJ5mdysgxSGp4C4ZfDtFChQo3GmO2uV6
HkoIGw2aeLYX4w8n7O6PzdvV8pyqmUIdtuEi98hZGTC6Wq4Jda2zIMZEdkBDd5PrCk5Cr7n/thoA
jDzAHkQrpVP4cJixV6qBxSAS/tiNYMJscj5oOSQabRXttW/T6kBLBRrukuYy6Cnuq0OW8a4fTyF7
W0qwPXZjlUO4bG9+MSJF3CcxECfHbsZ2H9heMsce6Lu0i5j3SWyroO/CAFORxZuoVwDvYrtOlxmk
FHNMqaIzsYCD7iKx/KerstZB7NU1TQKqLhfJa/RayAW7MA5aBkF3FNdnhngYfGhR2AJUzwmqyBqx
ykxQoNcFjhBh6ve6htLie4k4yFGSis+G9Jybp+oBWkwhtNSP/6V503klP3n0JIz2eWofTseF+0mB
Mp/EVZo8obwlfdFf633WslO6QwkpBpqIv/B3dCUTHUNOX+DLM/Juc1TeGt+Pd5G8hfVCpdfp832p
kqYWMohlHyATSYC11N6A/rt5UEc9ouwU7pm9qavrPExUUlzmr2ElMkfK5Y61pO43B8RfwdPvWHX5
1JXUfPtfjTVYqx/ndAs/9zUxe+heEwvmvRwwBPzcYMoE4nIB7jqyiRGtuZo0zumodGLM0LQv6pwT
g868MfV0x0r9DtlWcOItr2e6bCB/fNkd9HPpTBKe3gSZphR94hf8GrsWUHg7oPbV5WQ3ovdRioqO
GtjqEw1dEruD6OdbBG1JfOX2+qocUQDWX8WmJnw3xnU/HzmrHeExEPbwuvZcXp41tQsTvGs+ThLy
y98gkpx/D6as9F+axL2gg0lUrsIQF45In1g6EkTJ0ECFQ4yiyMz1B9mh9JBOZps5pfocHvTRmits
tmoCGt049yLU3voXI5AJhfpRHy+ki/2u+/39m8s8ouY+ESCI2521sYhEZOfNCl6ZVg0qK4F27d4/
1kCyiX+VOPW4mvwcliRa4Vok9zr9MVnuaNeJSJZfrrISePAO/R9t3rn0thXfNVaFZSh6/2c5M93o
CdAJcudkP4hNjG1+QiOc7/NWbOPyAG6/1zZU8W88BC9Igy6n94+phxwJ7gs627Ykqw1RVGCc3Yvj
SavmfG+v8ocOF1IJfUUzqRcHzLmoWNH5BQaZ+ws5RZ+x8BVZ1yzWAprUTDSe+yQ76VzukVVdRKTy
rSM2vt9ARCxcP7P4MPdbMMPLA+pmF0wYQ1BNrPmsA3+KHOk2YJhNGhcPC56HZ2shnIWPxdDOzQRh
JaDlfQgGsPxteJoByX9WGH4ci7eYBafksDC1qLAh5y3QVCfssEkFtyJLuZfZYiId2f9JeGqZQQa7
5A/4fydn3ST/7nRraFJIvnYsv5rQ8RpRQEVP9yFWxZMMfd22cnEZab3vQwiqPLumw02jDnfskX1U
5LWAPxvp18N296lkwFxP6cp+0+MxPhkMwGsWMDpFmlm4JG+AHvHkBQCCZ4Tjc/3+95LAYbyYjQAB
CkcwNF3wv1Gp0tapgqjjtbnWbcP0ck7eBFG4Bq+bG0uh3bWucAPH6U7SlCKt55FIgF9qp0xbasfV
in9L4bUSSqURgw/oVBi01R11OEGfxOOSyTruVaCYK7M9/CczFaWOZ6Nh1Vwy5D6oOpCM9B2CcKte
JoC6D0apKa/vTPrTm+R/Tc5tOlrE9MxqTiV0bctGqCW5h7lsLoibp1hruWKCVLjUGc1yPe9aTNgY
lnmeON+XPbTnS69ahw8fCif6lLMwmOWXqHGp0wAeDyjS72Lg2HS85kU6KDFGY+pI5AgjE8jBnCO2
v8CyM5HAWpjOGiU6yITOS93OPbfWG3guHUFZmEx6sP0FGaiao13jbwmRAMTwPtqtm7pKgU2cpsgJ
R7hsMD7jD7bhVtvbt+0GQ8G8aGVvS46yILnujA3sWnEQGQ+s08ryphsPxQjrZkCgHwXF87fbUBRm
Qas4d597AZsOL9aRBpAAnGW1rtVyAPqNPzmvIznXvF/rAIjqU3CSYJHyyoNATgb5Gly2+TOODlDx
SYzuwhkzUAa8QjR6SG1eBjiUP+H84dx9i1+3XOUjruw/r2QTVYildwtUWV4Ev/qM4MjlkPhKulXE
8GD7fRasV/MpCy6r425nAnJrgOMZl3/IfJ4SKByRTTxWCi/cx4V/g8Bfp0pxGax1xYCiOvgV2iom
0x+UYRHgqprSxUk4tU79Ouk4axHw8yb687YDNCpc0llVLD+gKgGZjuPknFMkf3BY2oXvyRr3jnPb
J4yx5Q4EiHmZJN/lUZViBDKdNyVZ5A3C5Ue8VasnZgihxPv1S5DAMzALjvSGZG2OlIVLenkmERbO
oJdxRVNBO1/YkvPRS9PAgwiaPle4yVC/SPrnwR2pLUjJpLQv+KWW3BfGd49VEzH0OTDpWtaBVibv
0+kCBTIf1Dc/z9wrEIAMr1S8cLkp3yb9F7YFSzVgVv8S2kYhgOcVOuAnWsXNKSu1Q+DXv1YyU5y0
gtNy97iSa0zC+M7+kXRm5Jx+YB8OMyAoiFqJ0li8VXxu+V3qoz0YcdGiw2kVtsVymk1o4nBa2AtT
FNRlHGVS6x1bgwzzZDG0+Mm7hgWGlBu5vj6UnO0uGqGHopgpapv1nBch0TF0CRggewQ4UPJUqTKB
z4N+8KZfIz2R77QaIAMO4KAbFNrp4NSMG+KHm14pbTOYWW5MTLicyaQIhu2lWddSehri8N8Il3NS
NAb3/HsSlkfFTntR5000Y1uZO4GI8Lyh5ze1lBK8TWgXSpfr4rKTWpXSincW8Yf2wpUNBXGK2IdX
HJ/SubAtbvnWLHEenckyPNMGpbomlz0hSuVi59jf4xrUTYuPyLJlszXKGAh4dkfiBW/iTMp91kRn
1SqVgSfssLKPUACE6EVtynQExfaVLUT8FDtZtFOlDYablqP/8wkXmIpIVPlqRdW8z5mtZZ0W9GBU
Ax3hBrP5lww7xJacdXPvfa3eSb/UUiQMtoNLRZV3a8LXfA0rHQMHSUKZjET1YMbvQ1eSMe8oZfGs
WHuz66ifm7dGezigMi04ZKQT3ZCAi670Gds8Nu6TJE40iQcEBbDDLCXC309aiDyMhuqG3Dc6msqh
m6JTnJlE4XBKVKGLv46+jbeYybweW1m+Hjywczn7OnS/0VfzvCYdOfuFzR07jXR/iifNut5TASjA
QuypKEfVp6FktRGTK/3JZh6Mi/UFU6ogoY43+WXfbZGIb3MOPhWOo9IlmXF2FqNGwcqUQwubQ1Ub
JruV82AFRsGLdapnT0pr3LpELDDylwGA0MLJQ9WN1LVmWaOrTT4xl3VHkh8O3wrrwgedi5lH85Ul
Sg6COYc7Z/gG9wOaBlJIEy8z+cEgscJCK2ZOs4lySl6vwhzXMxhwaoSfiBrnYpAeTWrdyGStyL0h
4DDle+MzoF20Tu7BqrmzKoFHA7LftZglbHgJwAONhxT8+9Z4HMHAqwhE8CJormdJCxcFrgnK8QE/
5PdctUgmMSUpqhOSwthfjhIdedt0XHas5fth3C6iYn4ABMg4Fa+GiZNacCB1ubvdvA44lTDIQ7EK
V7Laws5YP+GOJ/wzzcvYIZpbWJtA6X2+Z0IJ/NaxrPeRwPmEO5OQMIwaP3cqZ7JuAKamE47T8vhH
susbzClFsTOsXy9jUwF/VhMyI624NNYah7Ywos2m36vl14fznC7L4q4JCM0t/XYDKMeKjI17zRfr
kfN2aMgkZma5JnbcsB7PmSM1FLSueMa6Wd/XplfgeDNxbqjADyJFZpOa4Rz7EcnnB1YEqLYNphJu
Tz09z8TUZ4YoFNfJK8756LdEwKV0iaYGXTMjPv7NPJTtI2UKG6ax1VYT8uszkyBoWfHCvSv9spap
U6HC3vzxwBi57Noe+k7bRSDI+tD5tjMqmkCHgZzgJ7FVFWQwRHDoG1/yS6GdC67B7cVNGKESUvFk
beBc5UtyuxC/oX2kI68ylXq/a2QzvV4QhyL2j2G5jrzF/7BLqXJGt1J36b+i2/YcNlH/5bmeQ3QH
TDOSMWQ3/EP+DIKJBYvmdReddO3yEx+EdD37Od7J1NPWGk4wRi31nSKqGCXSQdu3IgYNtqjzv/X8
gaE/ntsxk02ifXrjTUSJie1L7FPIdAxsBx+hwHpARjpgfSIpYw/ZL+Ay3NBym28M3fPD+c5AJV+f
Q2pfuaTs/iVspZCrYl7jsyfx1yf7CYMOTd8tyGmcnnm/sANQWHcZVAkbPorlFZbCxp+Sa0fhjFnR
kdc1h+N9FYVJdDVJTWZyGucn5Zta0P9VhjQxbvPaAdYAjhb8pSktw5AQcduIjfpqPsLwhzSsTmdZ
PaTIu5BKRq9ZllnMW3zh1UIi2Unx8/m2hMbLMCXBJqWwFJWWV95RM5LROwdGXD2UOYZbr8zlGiYC
ZRF6g5ZBArBbw6W1I6VLuteC4ZpRW+je/dgWZw97vZvrILTkvE3NQ3QjEPUwA9gKtlAm44izrkA7
SFMI6E6GbEPKj5UeknJLD1RenT6BWKosBcCwhjuSKjUPdmaxc5ZHVq/EflbJoUpHYwCpazrybF7t
btZ6YSMEzcU+r0G2+ZuTm4kQ1MazjizZDHlgwkzu4juPAWKpkl4dwJrojrLpKU6EhcdC8nPIBVTg
qoRFTA1j0to8dcS8azPP95y3+LTBzZJzs+XLJNE1EcXSgU5H9Q13niAtaZ4zJwwzGfW0vxZWljHp
9NBjjU/YgXcL4IdyZnCJXQwUA+v6rjBw/ApdJMoDWkGoeSdMNc49U9vc69PkBW7I6hWiHevn5K1v
JzYsnnw9o/YvWwlk7VnyFUfPktJZrmDUENDEl20kuLkwHjC2Vq3Y47o6wMs+Nf4YjtkPo6sJsooS
HaF/D51B3nVE7LvpalNywN3HYoQ2pn30POI5XJFiJYbRX1dMu5fMwWR9uPIJIbolhB7BUZPQZMho
2sJbPK4Wa4s/4VfqOXSa3DdFakVp2BK1XpFewYMq6owclGsAjNUqSMq4HD7YqlanDABbFOMP9LOp
BnwR614LHdClQpSABwLLhuT8lF7QMPslf6OD/8aYLcNmQ4NqFgwYhqbUd8V22lBm1z8gDuTfVTjD
wpjIvYDEzCGhQjO4XACsDUy4Ttpq9h2qscFluf79fkK4xo+gpqvPxf+AyP1OA0LXpz3o1mDNEvYe
LEPloVru3XakMLl9hisCbH83jUX19w+aN8CtFlN04OSgluC3S5uSm3XMcna48FaP+9STyEyNZN1Q
mtX/Hzj1J7MYFsajLuDi9Ig+6UC5Omt5ZajZW5Gh3etLD7iCdJfPozvWeK7lXN/SGPotpQy+uW7U
hprwPJbckKsG6KzQK3nDzP4D9O4fOK12HGrqdYUqVc0Z+a2lYr1/UGNkGUPQ60+ESKbmEpBoUhYt
TU7ckKMy1mZ0XrqQpELvJ8h/cSdAKykCP8vfj3aALcRfJftaPHIxlxGSdI6A0y/yhmTarejZXbfd
b0PyW+8SzZOvl9KI+uguDy2gdWNWvTicytspFDdN4hk2J7J5Yf89YnspxtNT7RMgs6Hua3rbLcpz
bqCwn+NN6KD61bIf3ca5jpsMHoj2znOtUSyHdIKZVuVLRRx+XauVQ0YZctiCOfgrzEk87Tjoov+V
V/ik9ZOUCB8z6l1gL8WaqdYOgSZ2868C8qr4M9FYlQV1LrNP3W6LYtwZMjqis9oKljpq8SaltLl1
xBFWXHQBsQ2eTwvJ6C55Qvi7CRuMDISPG5qeM88AvyH4LQPYav1480Ak3RRNfo9oJDll45LWDVjL
vKkzC7YWesIhSeReyV0g0xRap+fCl9+W1g+mJl0M5ULj2JsLzRGynXBwTdr19g7blaRSxcd0ayPG
DSwpVaiyVl3rnfJH+vrVOvrum+Cs/HV2N4u+7xg8BS0JoyEFIJ03JVd2Pe4tOLvUCu5V11+CHcJd
YmopLYmqUR0XxRcvW9flIUDuQvglVZkpwyew9Z7QVF8dPprTac+1mf2gZVXhrpnogmZXAUaxO8io
1LtTGt+Oiqkg4FCET5zRllJKwiOcJ2UWuBBuEvOftqheCMjd+3e50Zxp9CVDo+waQ8yI+hF/x9Iq
qSU0qZH4YdmUOj3hIJPw1Rp9TAkOYu8eoAhDAV6z9mHJ1mAT6GtUfwKvj+VCvZITP3/FEcI58ish
S3eMBSatFmkrBwL7GiMOsNM+l3TXhoTCddgwOSMGHeXDiaQ1Lv7Y1at5jZVV/uETfQZaISDLNfZc
V6mBll2P80xsWpgnu3xSDtUb76XfgE1dOG00Bhe7WGEUDVQG1zDhhsNZonp2wkJxSjaGzgdQqlOJ
uzmiDMUZe1pAjwqlrbBTOhHdUaBnjkV22c0xmwXOuehQDYE4TOXglScCNN3ZdapVhZLAAqxXd6vF
BCg8tIkmk0GK55rSM/BA8t/ktxeZAhUoOdVwcJS/UXo2x7OoFMpL90S3YCRYjep+HHMk7Qxdzz9I
enizPS5+N+yO1xpnzxyZohk66PSabTPNdCCPtYICYTVPKKQ/5t3Kg8/WUo8rYB+Iswd8XEoXMaMD
36X0BzJzLc3xkXU8nTsrbMw+qHyDBE8ayVnlrCxlcK6GO1NONlWxw7kOirFRsQdvXjkMwta/5o5C
pCIFW6yO7f3e6RNzyemxD0EJpVFUdAgy5L0QcUl3hmdz0pbxGLqTbpeRuMeJqsktSHHIuRLremB8
zYwqOxZz7PPRYkwrvW6/dJkde9+DtLRE1sfYmvYlbzTux5HzMx7IN0E0/LjsxdUw8/sj/xCMtLxD
0/tNMcSGM0S4qu5IGpCWuSCYULcD7YeifFI1Cvt/bqmt9aN0+l9m8tO7DA5rUP26lvodqvezIK7+
pFSripP/kbqsRGZDzJB4zbP2p4PaZqT+yehfuwdss0nzGeors84jQ0g1IHhUpwmjaOo+fo+b7j1y
ZvUTAK5vWCcLmkoPcgB4eZznfGEAMsFMfNv6OYVZhTJ6rsrpJKxtbpjd56XoeAi3vSx4pDoy9vKi
z8mr4yEo+iwtic9rmNN7ukB4eAcyrBQSbXnk7StuYqZ0sfl02+ypIaIJY2a0H+29+uzECoQVPN6U
hmG0Ll96FuphyaEpus3pEqo4LDIQc25XBKTaAHo1450o72uJpuC0zRC91ijs5Lv5s1sfi2MFInTb
0AEoNq92Vw6hWRVEnkBl4K8agVMLo8wRMQ3xpsgF4WTtYBvtHL5bysqdC4xOrykyFyEXVxH0jgbK
JNkU2EyzYNPpze+acO+aFN6lZTpKEUddZhtlXwgxZOr+CroS5MPN9kDS4pgeDThsdaCsuOq3vyEd
CFfQqJ5Vuj2MO2l9gc85qEprKHwAuAZo0+RhDtj3cc0YvSEnGOoYxh2NyXUk5JhSuCqEP8sqXyAX
t/RntdtYuGe7vI6D35GBcIrVN/cr82UD4F4ncRaNPtK61BHfGxMgkRMzvFCKY46HhZTeJgZFN9Kh
QVFIKEX3Zx0MalU6LAvTibXt4cixxgAT1ic2p/P4m7ExF+ERhGTC127h7/jIaCVgfqpiNFc4JcvX
pInoZW0aYQKaM9cwqHfgle1Rvd3QDsdVqcEWYiCHzHcFjrhOl89K/EKsYjcTgRKwG6/18OZn05e3
uVHtuWJInnGyhIXHd9i+cG/8KtJao0zu92ADST+fsI0B3T/sDbFScpJLZKTeju05zC9AbWRFFaMl
HrXJSPFH16HKGb7Nyvj5KbCvhE7gdjI3/3qf9HR0YYG8H08Pxcf3MgUUfwiNOayu5RV/3wOdZO1/
jeqv7SU2AbrmoXfVeGk3wRgpl3ITq8Wo4pbNltNz+Jj5sD7v+/YHyfxaqxEQ72U2VNDptn2WXMz+
CJh7taXQcSU7xfd9uGy8cOnk4cFlmkjdDxGq+Dc3anaAaQTACiuHMCUbzqAv1ZxxoLqfmv/bblgP
frYey/QFYK3QEdqWelrdpKWa3MghF1wsXyHWPLpyvhILfRwxpHWixTn38XMqIqtf1OcpxFp4NcPl
Ggga/TfTdOLihzrqujq71fZcyjULPW5+iwmWALqm8FScRc2XRfh+FPSq9WdxxRf/1wKoy2Si++C5
zV0Vu6+FMqZXkYjj5O6er1kI7p94gHNviq444dENYTgiIWO+mlD1NB05az+9oTXu5QE+tjC79tAz
wkRk1kBvVPONkMr27UtjAl6VhCvJf3wSWGFceJFRlA40Ofi/rn9d3fZU4N9gwrKqNRyCwlA27u1i
CRy5/M+GEdg+63A4vM+3W5+kAZA5dy0Hp3pa3PqnWWyK1enV9gS81pcPFPFsFNNgY3JbddN0ri8O
Mn0dB15cnWrUXXCwQ6V5GpgPvhSgDU7BuG2RzyMoVBtCHedDTdB3bVPl4+LyPBG2BDoyiSp0EsfR
IVvy1OGBOP8MlARCXhDnbi55xolNrk7n6rY0D/VzE4ms4OdwPEcrJmglUMu4L/RteFrdmD609MZm
+RbEWmzD1TLadz09cBX9IcGHvMROoLqjy1xBHbLlbFuSmJnoTpANTUD9u+PiM6sBT/bY12uTP+zv
BxOjRHpQLgpK2rEPtE2cYItNZZW9K4QMKZUPpfzJE2YMoaxa0pMPLtnIYmeJJhG4/W/h/HTz6TgD
2mVF6kuz4U2yP5XCNf8A+8oUnxq2XGfPv6GfwmBDebz9YGL6yEuPFnwSUftGaRd7xB6L6iqqWq3a
CB0j66P80lXfc5Je0ZWBpt3EXAn5GII8kZ/NeVgfHWLFze+se9P8/OTBELCT5BPDK9WEuIqwUuc0
nnSt6G6k1tq0WDOBEyr+HVQxL1k1HQNfdcZk2/YhZVA27cIZ8QiG5S0D2p2jqB6GzRQfsAStgC4g
gB9S5uhqeD6pWEFx7tvA3b95TspslLC6Q4CfcEkNshZM6ZBvw/AAEWL3NCeI2oqCYvG+2TZdSoRc
jlkpYZBo4aXPhedve1sd27BtBv6r0eBE5RojYNW/hPkVv2wjucDu2yVlCF1A0qwogsqeQV5XhBMF
86a9ASKIw/BzUiKTN2pHAtPBPwmfBpn8FOnBEqcb43aElm4Q68F18xOVQ5MGLwB7CblxNyDzf0Ur
ic6h7jbsE1LcTd8GMNmPcKrxJtpcNXXNLz8xVFDmUngcpkh9B2qhZC+lNS0upQ+BGjo0+tDuVW/b
Dderygzd19Z/Z8M2aA2tI3uUOYTp2ASktcRiq9/lsa9FlstVsvsJYk6pot3FirEQt9bO9G0rZpu7
U+E4vQHOQrTmZ7BZP4zL0pZrurXwml1DO/xDaeXXEzwk0cH3w5JSN1YYlHiOuPHAt4zUUa4Tkqnp
6LiL4UYmplSPoWL/wHm1/MCGsAlNWAkvn5fMVbWor8gyahr3UNSOAK9OF/w96z+WDMIp6YM/R/gJ
UIMbMPfvNlB1akP8akbcdWZ+yksj3ZmYcWNcbzHzu1bIqnAMjEzYiST4rNiVdgKD9Rwqn1UUxQwt
dcieahtTfuaDPgwMqM133J9Pz88W0AzDziR5dWWmOY5/fQc41TdIS0Zr3Z3jlEVsAuXnP5MHRv+g
OYrlRCe3Efo+2Ggexk1lbZzQZCt7akHKxUAQQrqvAuNRCgYdXN2hco9PYxhI2of3sFHZ31+yZOm/
hs4F2fR460Q6ZanP/Ge3BgH9jdbg/+wI4HaV+lbTQetJxz8biZp0MDVGSYlfPpGZKtmLi+9HPlPW
RPNHHf9Z2BbL/mhHH1ep2nEFI2K8AmfnaONmkf+TkvxxZKOM3S3C1bCU7AE5WbngItQQO2x5zOqL
21E1iFcJOAWiJcAE5dmydFdl2+GAnrWR6DdR46DSwtoxOe3tFKkCiIbTQAgn6+6e8If7pDHE37u7
N896TCzSI4PtSds2Veg6kxWvnFp97l5veHiFVsfir3zliqCCxycLDrC8BYX7hKEkf2rgU5YWJk25
nd67uYFqJiZw6vIVMgKQSWg4tiEe7CgNaLpLcUWH1jWs45WqDA//RIsGL3PWDtImZlSXS6Wn/o20
hh/OAAyfMZQKLkPQxmcKud7OKXfIOSi3gMv8EiUX8YIXZkuYxG3n8BwlcRYGgZBIbYW/WDGnZVoB
uBnCgMrmMKlqg3U3WFkhKo8r8BRkfBUBX0Ym7PO8e1Ktmzx8TCrQIi9dDb8pKL+z/H7Hg4YAa7hw
QGJILiqcXcbDg3Ji9gYMCwfJodXORYtETBmpPyFFBpFxL6Gs2PwTph9ZWXAr/lYw1LREKh8CpDLS
PK+vP0qeZQHXywBHn/9Y7nnS1zDmcvQMbLvB98PlKH+MtyMtAa2dF3cOPM6tgH52AyXvEIgKcmZy
haM/Ubs4B5T4F78CI4mxa1R5x4KMIwfY1G9XJ5xO36GgCWk4kDJzSnmxZmVuX5ZTFg2NBFjx4bZ2
MFolyz3MuvGlGTy3norDPCtmbYYmO9uqwqpAHObD/SOFKhcAa0AQO+B/DJFMotIysRKxeYhRZW9X
nq3Fb/eTlZ3BAZzO2pCZIzW+dTx+p+9ez44heR7eZFr+EJVh/RXIRq2hbKHRxvVmJHveGYsUwCAs
CQhiBU2SvKJ0qg/3acXtDeYyFtW9QvEtLf+y1HUPDkeSVvVu81/RfTmC+P16sVgRrk4/e4v6e4fe
/2Bga2ltRajemAEoq6ZgHnJ9QIc5gF2Y4S0MPomxYMUpOOIdLWWMHPdCC6Q4S1MXdLcpI7rTE62l
0jM+kf3xUfArLX1PDBnsYD4QhubEunEj68tACR6ian4JhTbAyhcG8XHYS3HGEwrMZDp/lyiSv5gk
uCWQkjnR/TLXkTBnsPGhcFXtN/DdThrP9AYuNC1Zr+gMsZV8o2rHDRFqay09BA7fX5zmgjpe8GLN
HByYhIvxVmtzwvycrQ3VptbZ+DetwznZPCxQuPSSY2UZ+dnqFpbi1YsqCEQ45f7gCb1ML1Y+pZaG
zdJRuEgFlXbV7qHvkO9wk6VQNYlMPEQ7IeQG1ArpS7/M83pl0H+QAo2XI63ksjcDp/x479Lqk2vy
V2eeY1ZQOgwfE1sAefQofuQqZJ7fAi/suV2FWaBOaLUkmnX1hnn8ziz1fSV55+sFolNsByxpmu8o
tdmrHHA2939OQau92aJd81XEmgOQxfjGoYa3U5CQ+sgrDOcEap4jdn2WhTQEltbFLGUYYE/VUUjM
QoYHq9lgoXhCpaBeXJj3bjMEYDwRpK3UeNfwvh0ouXAgB2d2kHnqHKd+73bxgQOH0a0MRErr19v7
5UW6gV7ORsbR9mLbyInFv0kaTkFeyH1ibhMawVACu9ueJsKqtAJmNKRHDQtuo7v+j+yDJVYQZf57
DP8cqUXBzJ4Oa5dQQVhbtIGJmVxb9KL+vHO0sU3xd+FkI5ymIsPDqo7d77HrclVGGi52ErMJcG9j
JqQHwJDbgk/B7lU3zv9DRS8S4J38aukhPj+GIIDePzhQeA6eBCp+pZpKoN1yHkmFgOnG+3PyV7sH
JQKFJMyk6WgdNL110X0RkhBBocQLh+JQkedL1Y2vXbbprHNB7/0kmdLQWBCQITFOQvJy9NCPsqbW
3cIQ+t0HUnMSaILL7UwwIG8NLw4MV52YLuftu+4PJTQRre6mQ/m0Dms0un9vPxpAxlFNvShxl5CZ
stNcOM+L/RTRPJ3oChKmiK8Y6OO0jmVg2eh28eqbeD7tXWUkmDfOQSDVCKC9zreLanhA8TvZroXF
LbUK3kt8JhsYEh7knzolKuu8Cbm2zJUXCdoUpKmQPwMU2Yftui726JCmtGzQ0kwdvclwiGNk402D
hdmt/6R2J9ZqVv1cIuFMFbfZLS7z6rglCFIOK6rg82baXxhglIo3A9k6RMIBCe5jRRS5abHpfgHn
o/ILoxHe9yAocDBGmsIf2q4JrgtjML/NjvH6eLEnBKwBY1mETMwxMfVFOoX0RjOWv91NKc22/9yK
pIcaKwDcMl4+uqd5Yd83Y3Kwr+JtO4BkiclCeM1ZyI0xgbMqz9EY3FV12BflgzalhWdUrEGHOwYo
trDJmtgQHD9nc2MuDsg1S/gVhZVQqlDmqEKPnADEQdkVNRaqW18kxvELvQWXDZiQAYzPaFt/MYUy
qZP0ylD9Yghr618naERN6sZsVkLh4H3wcGWfhLK4tTePSQQNC9OptKHGvnf6rYSa8Qhf0RcD4shW
R57Bu4AR0HeYo2nloaW7XCQrbcSIZKoHBakTJKwtxqG2Eh19tTzM38PN53MaZsmQUeoFkxVUX0GD
thXBqx/bCkNKyKPEB8fcGWihk2G08g7ib2BB3RnAXc5k12Io+RzKXv+8I/mJTryJd+KZ8/kJJMi2
3MdOxH0M3nKR968OhAjA4TJ5l0NlgdJGd659j9YOOBPNZlXWzfGKI/QGPj6AV176YZbe/9zggRr1
KndJdc3R5BovSEA6WGnA+Q+DNlX1ABcEX3jPXpQwcHE5FxgYojE891tO/YUS1mjmn7yq1a6n5mtT
Bw3M8tWOdpiTQXH5/5RVVgxBvyNp8of+jjmg9HmesaCLC4ZHN7eTQRv3z7ltnWtpFH3+udhEtlL+
yQcUa/jVMwKnIWPDuSFElW4ZNzoODhTeOb2wZVdI9rjIcagIJiExmQz9vHJUf2Fe94ybBMAwVed2
7u30muh5HMaIsNOxFNeXo962brGciEusoDRUPZLw8B5Jyw6fJDZymo41VBo0g2zTrzFTJdqtbH13
ij3FfcWBEP9uYr48QQUMxWbzpVei3m8qMk6mfxjn296228G0K2m5HNnu4CMiTcRqtkcGV1qXBU2s
ahw5QgGFTr+UPvalSaUozaSIehxOM90GaNAUqh9HdgG5i5qZCQKlpCeqI3JtwS5bLGC/BtKOHYRT
SFQIQDYT7WUPITbQIn8OWD++unqtzZgAnfhR6TifMCP05t4drFbTRNxBxBePjLQpYUziARbHGFTg
gOMzYxLziqImVW50uU8LswvfbACS/L7BJyNIYhHxQ94GqInqJ+ZESjeE9gIjZah6NWQu/xknepBF
SIPViOeskkgSa+TxxsIS2UzY+1Aj5g+yu4q3WWlKvqwrmMtKxar/n7bcLWlxT5ryDQ0poPIDrgy8
LaYxeaW8NmFUYDm24McmfMRU292ZfqLwn9c/YFMdl31BJZRE201RyFLjBqpWhWeozw3XipAxIiWW
6x0mwm7wudjb1DjyctpqYSEtAmp4+J/t7wpP8eZ9rWwFrLrN8B4RjfhoKtfJ2P5x6wmBxGLzfd7F
CbNXbMYyeZL93T9+y6bSdZOzTC/tSav6KFGEvpPFEfPUwX1FLm2aMX8dufOVMimAxZq2t53tgg77
EogVYZzYHdrmAHLuYFmbSChuVOLYa/km10y+0Fwfs3OnRkDbTH5+rIoi4e28L7J5z0tMtBL6kxh/
KFUDl22f6vo8WE5MBYKR4j43oEZ7LxmCaHRFn+IT8klj/XxJwdL5r3QZ3NqtJSiRZJdSNRSJCwVw
+FR+c/nmnNUSTqdxD9Q5ZG9aw+vWnsLLheHWQE0ENkAqXdX9SzAlzB9755uUZ256G7ZZ0szCM1oj
tFGmtqARAYZYBGLwlw010EUq6a9UpPq3vbqFUUbMEDEJrioIZNq0S1QyefvIf8Pk4EKYmHxUUGci
IHF7yfJ5fMFArzFT0u3MxCCKWmYSOQ9Xx0sXk6yJKuiVok90nbN1Prr4ED4nTSTGsY6JKOa5nFWO
7ARtLTsjxFfhNrcw2aBQ7rWXoQWk2u+pnD0d1U0APpvk/gYWqUPE/zkxJq8LXrUeC5tEu8PxkRis
SRHzpf+MX31zUn88lQeVc0Azb9hu1oDrog7HbfcUQrpbN1JDf1HLWOeDZtSNTm3OkfCx86x9ay2N
aHspZ2/kyHn5JmwRwFrMFtNqM5NN2fiIWLPgws7Sd+LwdcVePfStjp86TTF0OPw4J1qFpXkk7gVC
Pf5zd49c8PmXD4CHhPHbYzzeTg1aox0d5/yPkk5I2K7stDjE0MApz5+o4JdiCQaYuLBlZxCZ6Vu/
LH3q8F6kq+45SUHZG83Lo9c9BUVh5xG/KTpRWs9FfZHKGL+YcCYn1ncD3gvsoXSK+WBeNo3NK4X8
gqeE47vyNAqWuKLpL9YBzfYEIE9W4sHWGrOMiP9i53Ez6cxiAkpPDJptlWcJfIc/0oKajGXyCUPu
C1CR39cQI54ikjrD3IWIemmstwlYvYPwC9R5VN0H0Jp6MP6KVYZ3Ee7Hjy3GCwn1hTL8D/Bw91oW
m/b8TeAqV8ELfPB6ESrJGQIaSS/A2LMg0rv8JE0GvvH7YzYlUPF6Q09hAWoBqx5964aAvP6O0eAL
KPKna3bzs1GsSuXjMbSFWPm9gNvBLIiNkffku0/xYLHgkVmGM8qnTmuY0mGIkq56TIfv7rn1k1SO
68tK7pKTbw634tBEtv1ZFTSiK3dAqkCPrBTlqiU1C29/SkOIkrD5LIfUB5EhoBcHmYkCN2NB5aUv
V+obRgO5woqTg4QuCqrktHORWuwF1ibI/RUtLOPo9qwr37XnkM7Xu+ue71v7R4FZ9sjpetfGvApL
o/jEX9JCOhCi7ZKpReOL5XrtLJ0Yi4Geqb/YnXAjH1PyiIWyvVwqpPnWrRNLloUxmvE0a6n5/U0h
OR176HRlt15Rfpk7+pplOGebJyqrnN6nVf44FrFk9d9rnUZ0aMDboqapriNGS/u4GvzkI6YUER6C
GOl/2hOgy2r/l2UE2pm6WiuQ5RVIn1l53M2K4ypui57/UUQQtzDBKOXDdvUdE/ARNyitdLEH7sK5
SlZ9GPXhf/YamIkUJ8O/IliPoyqX8QR6tQB9FKdFS6Bwt3kUQt6Rk+tuhrkyQbscB38wMKtYlE+D
5VBsElxh2G+5H2WI7JXM5SOBITDrQiqZwfwCrciMKPsk44/iZmgSa8pgSPBityL0IRUerK9+/an9
HwHa+naMUdmKMYrlkqj2HeAMCVZAZ7gxQRbCoRDOZFa4IGhCf1sng227XhAZX0NdpCz6K1I/YOZ6
U+9fRvs9RM/98dSZQ0FrQmxBQeDR6XcJNm6MjBa13kHAbpu3lhW3vVH7Bjg6U95PFXTVKeYt9wlb
aOuIjtOhPasjjnXA0kObW4/FOXwJgf+fddXz4LjxN2irhOabmzawsmjYJKz9iS5LA3TlntLPGew2
IahgVkhjAa386J+jjE/w6DF57I7byKN56A+PTpzWMg7hNECVyZv0WQfdC6OnHXVZP/xmEZO39zZo
COfai+MJdcpPvLzlCpgziUlt8qPOUgSnVG6Nf8QA3mU+FhquJkAgxB7uF1kTf98CqqKJwrIwk6sK
YRj8/Ve2SsS+37518m5pveDsvMzVufeKzoHjS6jEp/9pCNWEf1ppyunK9yAG3efBEzkQ9SyxqV27
g9aIgHFsoaAsr5o5H+j2iwQqnKx1MYFmsFcYdN+fdzJBZC4NTJqp3/YFY3bu7MBqDhgy1EaVX/vC
9PFpmFiqGbisc0DirpJ1/L0YdV+E7Ynsh5z1sd7mFlJTYRWYF3b4UY1p+5165+vVxg+G9drwT+C0
5gj7N2YFvIWIwN3q7MIpoE8qDjVpS5hCN1aacp8s9WadQD7KHvkBI54YwXwCakSi28mMvthVjI+Q
iAOSWWgkWXegRYSe8hVL1X8V10VXWULCUi5sBh6mWUQ2JjrjQb/0VXC0M93wMznmxYFU2P2RYvzO
R1oJSUBZpRU8K9FC6OGJd73SjeJzLkkuBFKhq//zM6aWv/bbztpPvryMTpFriopwI2hFvNFQsJ79
bMzOy3nM3awNO6hofjxB0qwy86LEw8TW/OxUXr+olxT0ACmuBd5Uv3o87ILyN4JeQ9UZjnIJPmXf
SWvjGfE834sATxSYhM9XTMJ87FWyBOnLMEiJcU/q4SuIKtU2uHsD9pD3kRl0jr4MpK0Ytq33hxej
lHoCia6+5HBY+vlZnfaVK9K3hzUK8WAW5vJw9eZGGOvgfIxrEDmzObP0Tyef4zrvNWyERezCX3lE
xmsnG0qzjaCB/VEcbIFhXP2Q1ZiaTq9rVB0v9Vx9uy1C5+tVe24xVpMtN0peaFzp/4BU5HzlxIii
QZ+AIqctKcOe99Fuk78Nfl8itOoFjzb4KrS0pLIzC3DQcdc2P+IO0HvI48OiffsBsrZd7sYsILh3
aqV62wsDJ5/txpHjod+yyMB3MJ++cMamtPw3Q//IwyOKvjg9Ew6NFC6JpWojYsOKGa3MKh3h2kEm
WTBMNOnfRLv0k3IJwxHj+ySFbIh0tavcE72Agp+CO1sGR++juj2nMPdTCHSSBSQ3WfUjrejxiNqm
ke8vvcii/9fMtMq9WQDO9GWJoNKjGSE7oL052XaxZZcSPgsepPtzZTxWtO2C1Ap/UOn7hUFprpGW
40aGCJv3/tZxx/5KO9DnGxkPTjtnSJSi9F+evhR93swlWH8T5rezB1BQyRJ0QjnYWDwvH9YJl5ef
/nTLgrLGda7g78aL/DA3/2C4X0NFRgEAXg58TCDatfR6z3iSP3loKXDHNaM761V0+9LA+/frS1E4
WTuS3am5+z/R46a9MH/MSPz+sx/CaVaJMOcpE0xkgMNgPWq1FSXI+hWV9Yj1BhZ/XIVXKzr0ym5f
eWd9mYxvlLKrqd+nmRPY1MRuCT8kDzrELc6dibC/xErZpqHCXYlFqrQcetYkueE50f4kDBP1Gzv2
qgkqkKM8h/wh2ZVLE5qTODjw6GC8E7AIzjxuYOoOpSotG9tR8hcAvq6EeZ/go6VnDWivNoVjvfyL
hLQF6MUbfU1f5DHfnvmSbxwAW2R0avNSTqy3gwVNbAFIf30IfrL5yxcCGHwG/DUIAC4Fj6z5s+lZ
OzZXCH9RN6A0MMGcqUR+t8kcvultmKlMzyEYJMHrIkdjHjwt8+RAF+waz7hX2MCWYT10oZIkHqS+
atXhchKYaIJ/hpsdSepvp0Dp5SZyS2wqF5tf3n/M7H1P0IZjpBRi+L6i3XAiYejNDoiYLOqDpjj7
I42i+tsuaVkT8pACOP4xwuP1Oyf2dooY/C6hfu6dnoQIrknOP8cCIKJQdMyLCYV0bKWCusC0+gnJ
x/8FnidMpA0FFVQWIfBPO4CTAlxwdDH/EUEGzKfhCB/SmXu6bGUqHCvnYXGAMcOQ0E7xjHg+n8lX
6mdf8MNaGRBl9LPuPKPa+W3sJMsR+K2QEfhzJG+P4B6a2zJw3FyLxkTV5YNEYzcHVAeeDJOkz6Ch
YRAOehDgORSzDekzK/0dgAAUqFaSEKs65awB6KfNjlcxlCU/pjekcK2phhqGrmWMswbdYulVzybW
HFLvBN0KQwM74Jw86IDPCnDxDpqzsisM0aNLDWNL2d2cM3xCJx2yuQTeLY7QawBnP73yZfAYh1vq
hF2zXDZLoaGjNGf83ltLtt0s4Hbkgejlr7xuoCb4MvEnw247VhTgPISFIbLlekrceLBwTeljA6Xz
mJcc6gxI88wUlTnPtVDVf6zy3jAfqHLmaSynNRGws0LdoFFok+sRHZkWCd2hhKcYI09gfnqL8ILa
1rMaMd73uIO8eJ+FFxoyKsVMG9J1FH5Zstz9n0HSktTPZa4BqENilhlAnMU37BJtOgg9i6wrg5hQ
mCrW4u0dcNmo18cJaNZ8sIQTSXQ8t8BvWdwDb9WG6eafJuakrvlO+5tkS6X9s0zpCAkd00PxIzqM
Jgt3ucEDe3JdCgGrc0KsFN2E9zKcxJRrIiOe91u7+gaWGduOc+q0cJqHuaHj9f0UVAHFermxFlgs
jZHVlY0+XAH+RAc5oa9CXac3ZRENgXSosv6LCTUIQuX3ldAZRB1LtxiP8bmuotVpQ99nbkVW0tdd
5Bc6+FGHGtneZBjkdn4HlpS0/q51HRHVfHlnR/qItmPRnqZNYO2IIaHbY8Cd5k7v8+oJ+L5nANv/
EGwzHFzuSypxVCRNrflm/NFHV2DdoZdxDglSipZe9GJPKH1WvYZ4NAY+W0AWg0Y2cpOHuVKqDo0S
Im+Ix3617q93IJZYMMPHppSskeis6PXUoqQLofWitf9zvYIMOPE5vI+L5vNTunv//uRHbCoRRiIJ
TrfqBGVl3BU0ro0d0v6LfJ4t46KkEOgqE8wvANqZ7MCmvj9Nbm7Vw2Q4BTkRkTWL+V2v1TVz3yhQ
tZcXVW7rE6CvIl+vqnq2D1NpNjmtWvnOKEcQUzOPbUynKtpZhzSQ4tW/M3y4Xuv78TUIn+rO9ysr
d6clZQbFFM/gy8FqFGER99l3qINfPuF+eptqH2qBE9OJ1+rUkmu86+LcXSPp2seq9P0bvRyHAmZk
47h5GQBYuxX5mloZ74sH8hsdQ4h9khMy1yFrCo39BOc2RM0jQzJcMwrwnlL7enbMorcEiIHQ1m0b
/10y+3w0CjLRxl+aUEXG9zYJ9Gz9IuV1sh5u9nKoaccgd/7CDk6z4bLQf4V8YP11Gzw6mdQm+6N+
aFktEPmcr+Mp8igqER0SOoplYMtEf2GZGAlsY/B88P+UYz4K8fAkzTAM3Cd2XUCBcoQU0+Hs9jbW
dZTlbyv0WiS/b0CXN8fiNTEmSL2CDbLAH02Fnn/nfGXO4MomykJDamDk5DEogpWmg9IYJpFpV7Xw
u9yEKq6dCp9PsLhIwvVbQMWcK36CXDUscYisYPuSelwrbZ0mHQ+fXaF3CLHx9kFuIXFFpS3NFj59
9XVHZvavk7iETXnky797PeDf1waAg0nImZsH3FMi3NffUrljzT761nTspTU8LxnTleDCsCJj3ztv
ax1fhFV/berxqNJydgY/LAOS6EblfHkFshJrpubr36SKbY4a6UptEHMIX8wtS4omIVVM67UZBvtz
YPGXbfRDruVS+iqCE/Gg7xG6AW8tQ9bkdCIt0X1NTzJL9CGMuhNtu6Ooow4Oci9ZhI8DvWpaHZ4a
NtJyljzvPWixVkWxYil1BA5zachKqBl8LOnp5BrpblpeoUUTWiewUeVwSEKOX06t97uZ6ght3Q09
S0hBkHayJM8zzz3x9ZSC9hcaizdZLjIYf752G0N4n7wgSHqAX7RHkqStf+opBa5ktPxBejLI/0zN
kz6ThAZtP8xlAUpr891ziW6RCOy1/SD1x3LeoBU9CVXc+Ijs+0kAJv49w8fMaQS8JtE9uv9anywS
fic098YStXLOryDXDlkAcYe273A7RVoz1x7LenFCUD3mTbRUOu7phT5apfM6j2kXQ2nHIj3DOGow
WIBKuEQfIywEziyjF0oSPJPFRjln0OlxRa6aiI4LE0TI60mprxGMY8Vqlo31hKQcoXziJzbG1dEs
K8/z0r27yDU+sCvnGUud8uP/FZp16DnvaHnrASsAmx/apgwVp+Qc2q9NpP1WCWu6Nq01eYGDTX4s
2QBqCKcBQir8gpDYOhPS7Zw/dcMO7AmEJB7qd/A19OZoGHsVOvIyJTFvPgGONbUviTX033V0cxAo
+Pp2iimx+vTj4VIpl+ubD8cWHEJmNBSY/lXWq9h+oI0e9LMPhYDPtNK6qqxcHYiwmmeKMzBd0zSM
i9HDSEdL9nPg+sNhEhTQAcXsYAz4yazZcP9mDZZ/YDMVmUJYHs69mzFEhlmBZhPn5pq/ruskxYu4
Y0nWN6vEolHqrJQfVWnHY1F9k7qtJGOti6+pqR2myM2MHIlvKjTCDqnt7UxIwf/ch+eKfqR1r8Dj
wIcTsCIC9rJJJgRKNTQFLeAvbt6clLoyvxkfBmntiEgFkmTcYgKGkfDlv8aNwdVFWzdemKcLKKce
TCdNuCI7INr33ewbm4yLTm+XvS+72Qru8YLpkHys7YwI5AmXjYgWEcJ4j6GLJ2p41109vHUMSTOG
iHyYXvBBwwlqrt0BAqE7cGQSp6b3Vjvs4/lP28d+9yZFh6tWn49DYI5fEJzPPzWTVsuNiBrpNl0Z
OsvLblibX009qGLlTtIgumB3oeNmqSmkMuI9i3VYe5alIQ17JqLxMpjXLAprgMXDL6Ltjp4F+Vk6
qRXLoVD1PQ5+ko9To9KblxVfDz2jHCTxl3UNgS2TdvZ0DeRU5rOolWRNri3Yu9sX4xrlXVxCuD1T
sC3BK0K4OBGgnOpEYj0EUEtsG9UIbCeVs7KS3IyhMLcIFTvpXlZReXqzfcEw4k/Qd1ySKEzqIHiJ
YLd8f443BXxpielnEyk987U9PgtPUh2h6ddHojJy7xuGGT62GIdInvf2rS4arCQW78ZIttnz0zKh
7BNXCcv+pgVMhwchdxvxDVVsZflNzwciftkQLaf0l+YE8oKAUXUnAGS7v6lVdyfjbzi+V5YNHLBi
KLjQSw5ZRL6vvTiBvkKhppn9+qwN3UGtFY6Nc0/RiAtuTVlwRJU02zumg8ANXPLPsml6s2IH1eE2
0rcI860NHTiWWtuuG/0Q9hQkWTN+yu8d/hkQSZE39HcD7jNvm5Xfr/+2SLuzGk1FrhGxl2Lt/Qmw
Gt5LVzHVtN1H48EEMLm+zOk+/k2iXxe0st+5DXpIbjSVm4j1+NYw3pPNxUgHdG9qFfYC9Q5Hraep
9WVcUQXVJvbH52T2/UU76hfLLPKil5IDgNQVnJjEfBoThyAz5ypnO+yEwhp7yBU/2gHyqLZxkZcP
I/XNJIr4kRznhMHvyMlhiLVQvP4tXK5YZxfeHc2nuBh2uDSO2RQqFLdFwD259cfBcit4KvonCTqr
kBZlaCoITgk0BqUy8hylbq2tEMeuaKWedQJ9TNwiNcLt2CIhEwL9iaDRmh0W52Y4AjNqKGe3q+GO
ULO+1sAkN1v7ZWLeYoEtUuPiaugDx/F5dNKYkc3c8cYze6RGzN5jhUnbNDN+d8IcueBKSA1tdIy3
buom2ACIPPvZn8M9upld4D81Yzc+YqzCtDO07dxV7IMoaRATw1JqrngnhIpKwPcocxoeEDs3JzNR
DLiPczOx9muOT2RKnsH5RklpbLgu7EY2P4NcO0Qhcu9EbHig0MjLxgiOztkPmlB9JN00CztSWxYA
hsZLS7EOdJJlaT//i9a553kUYZ+FCcjMrxvQHRjE7nZNuixnj2qXRc3k4lWWFil9ySJ69bhQ8/xn
2wN7wGMge9998hIUSi3EOBUzl180H9uC4xccLfdDLHQpJ1RPW0lIAOGKYYTputTMHgHy6ITbwavk
FUGnZSLn1bfH/9m1/dyzCOeDaMUhETlfGZvN0iiC1pS17cC7i2tP+eTtHbQSGvvegO9jQbayFO2+
Q1zF9x04HfF6/2fWW+8p3upT24qaaYuXKAE3bsKKktR8hCFXaYKxwou0HXYuUlrdmqSQkOlBGHhZ
LA2VpA7lIgmzVN2qXB9PiJ26SthvEgG3DuWW9rsd4ffnfNd2dg2TSOR8d9mwEPiI6fGEud2WavtC
LL/L3I8WtL2TD/MG/A03DpA3IzzjmmFl1lMTU6lWTStcyNZaWAHIbnUZw8U6m9jzYElWFfWN3DcO
pD5CqPdK4MqLIMj3X226guUPeo7wMp9iXh68zYPnrm40BnVe38KvKbuV65h6+6AypZ3ORvn2cIWi
j8mOx8s5gSw5nY07dcuVdqA7GuSSprSPOqmZabbrSx2/2ZeWK2v0ETi5rzDzJuiuElQfC/rAMNqZ
RUZsY67cHRBNJtOYRjJvnFopexXL39Q4a9pIaqzf9MFmH9ieRWuajkMXu+w0ci/JL/35QaBDgtHv
XaH6OsfOCY19NwI9wLHhvU29CiWq7dC4+UAHeiJhTlpF7zpFD9XFXe3cbQGZMV93Xrp85zvbB6fF
35WSJFMlwIyJfVqZONbggXFkyf0hlAfA7wa0ONf7/Z020VfsomrppxTuNuhWAdNO4URJL/47dqUc
AAgRiaXO0J2DAGo/WgnfTS5SFTtJTdc8ldY85iJbYvZRMdPmpyiljMPfxoBx24fOTSAX0hTX17eg
y1mNnUkj1npu3JiK6DW3jKt4XZPWZajHTh3I1PfTYUU/wNx/YrulITb1yZjqWBdeSMobIhEbGjA5
ccctAGquMStbRkoLwajEyBcYq+XcluvsImxDMGz+/ciJdHCN3gW+6UligE4ggyxyFdkZecYmpxnq
9+dXZY+TSv9B3xu7hoKubsGgVNd/iX+Fwb3BE6uwiFSAQYXa7tVkHt9EXmIbeOTmhgZq1e/eYay3
umtQim69srL45Rdhuti7MqZ9o+0FHoBfPHfj1yF5xOK8T/0KuhQH+KedfPHBQCakzZM8khRnN2AY
egdBapXwe2V9T4OM4VAlc3pwMqMJt2rgBhIxpkha8N71y2cCVa8egbHAcHWFrAbheK1zPhsjxvLG
7ucdJLKGcrlUjm/j3tjNok7q5TE9nj1IrgBV7YvGfk+afFnEknu6ZUpnXuWipm31C/hxu1HLWGCN
62xQwdle+MJlw5+cjFa0PQtS/KlDB0A1in9ZteIpmiuqtEqe0KUoft/Ua+zYJ/lyt2yHZQXCiG05
FOZHlM+R6zgxxB7XFwKIBW215mC0j1X9OhzofTDjNhUIVyheg5N+ddUfIbzfflYt0i8RnK7eQsiF
p7R6kHpjnV1/HPl7OqPo9kPvudGiV4AOCNk7F3s5KZ2ZY55oSK5eKvWBVjAydf2iymWg63XVJJ2x
G8bfEqvXbjg0qAGr9SWn4+CAbs9JpGZVdhczg6tiLaBuAEdxIWkZaro5f/Gt8K2raRQ5Jw1iSQei
Cw35cAW9nzS62c5mlJ8Y5XUV+iH4PkiJ7BoemkgnEktXDe/pzu1YdbGyo97kh3flsgGAtZWNaSxG
R96B9E0kkle5WJ2vYpLW3jqBFfSkltuzfvLcBnlFQ2k2ImInT6WIjl+D0530/qg4Ot1RPV+7E+Mi
xVGbUlQtT+icRUWHuStmz78XVIWhZJ0yDGPVsQOiYmFnw3/FeaOkKi0tLJx5o6KBLPsETjtTXtKl
i0uFJQFbZH2lwD1nxtOqAUT+z6be/OAvPygnP9rCXJRqyb0r52BRSPiKQA2Q/g2k+iFnt35C/26f
Ml+E35gHrzMZwxoVVN2HAXWVCTqiQQzdCDFRAZR+eTmEdjv98A9D8uHPTtdGJMz2xzbQrwuRjFIH
dPwLAhMDMdCA6wkhfnQe0kLK7/NvzX/lIpKcaMWa1NuuZFLR8iKuhQGchPsmjiD/qgsxwlTdSG//
UygiZ7I4HcAyAhcO5d1jAt2ODELr6iX45zf4JyiNOhzC9wfeW0drS7N0C+6W0AD9FCu9SW4OGF8n
+F1HGtEfaRYB1NDSU6tBR27crLiQaivEWliiA0QTsdcT4k3vZr74xIUj/WuM5e3psw/lTp49pwv7
+VI9IsjsblzKSErotqBCeZRowLq4q5RvutAohTwJo+51C3uG9MwV4sC7vzsCYN6y7Lz7FM8+teOD
PtwMXElLK2FB1rJQKypCi4+A+DPqcZhxIj+m3qiKmY5dKRwPWzIjI/9uXnV3KtSSKD4CQVRdj2kl
QGJ4aZPzCzfYBx6SbOJ20zVhLww0pFdCxlWkK4t7eGPp4gZH6LEiiPdMYuepevF93DxOIJKMV7xv
ewowIes5am6ws2zfsQ/o4YXTUMDgrlMFMlsiG483Kl34LupsnidsUfq2xgQgRBz1Fzf5563c78kL
/q0usIqn4+vyCeL8CSTopG/UohMDb2YUmIPjtirO7zUVvb5rtSthaCCams58O5ayjDB0hu74z2O7
3EvEqrcspVlEY4wpc2rXrVwhdZIYALv+eZtV9GoIDAA4FmFRLfDK3dxqijfi0G6IqW082O74T6jp
b22HZ1MeNLfeMoYNoZVN0eiC3HrIi/x8oMAPVN1uDEEQtNsEytTqKDbVTjvIoOmbkQPAqYIUoad0
fOnI7fqreMUmKTWvsGRaiKTNCw4nOb723zMPwEj2QOtSYGvjhupJ7dye01pOYSjldMCWUuj2b1Cc
KlMvSJBk596QkwE1TzkdUtpiCbLQoctf4II1g5H5Qlq5ME4NOO3+iQf5cA9CXYkkdjpVSOyz8ja7
wmvQrFY3Q/EZDCRhOepYFTaQ4iwuB/+ftvRJNU00exP/QoXsSKp6KxgedWC8dUe7QdmpP1cJCrtu
FEPK+2IxzIkvoxsPWv6hv/YWKT6Umy3aOYFP35MQqsbws/Sz8STBvbh0/UZM7rEVaMggAcY02b/J
bQBtSZh6gN+k5rmdvK4P3pgPMq1O9Y8UkKqC8nFbYQztVERJYFCYglbbQCSOo7GywbyYSA/bJvSC
zjgbgYWCYlSaRZJgf6UxbR3FgED4uphYuJ16kAijXxYsHiRSRQnaVeTlyxhLDMoIEHdPXkc8uX1v
hTOssf1yN9x7Bd+2takxIisPf60Aw1rDEMkFnqon0aB1xpFYRtqXRv/+mXg8m0ayMPD6S9kOve07
quz1qJch+4nd6i0MAis/L2VdHXEHwmyHCN0GnQDrj+c62Cr9+kdHAdiVOVDgVA3nNE6YbDruhYyc
VMx/Y42+ERAd32TnEzTxYQpMmh0aNIUsYKZjsyzedlXPi/+V4LUISsQSQiiFSvZ61A2ls8PgZMna
9bx8yN6Dnq2i2O7KZ7rN9pIWa7ngsWSlUCXeOaULZbJWBEXPgsH3BKQHUbGQz+7GSsw3/iDaN6ad
K/qrRna64FD74Mnys4YxGg1Kf1NlCvrjNYR3CTgUjpG86xJKSiYoIybCd/GjjS+Zt5zpg6Ayn7eq
qtUbICJT64Z50TfUCq0irgUFejUePvO4rBeaGUORO7GKxzlaqQcrbQzWP6b4Hm9pu8YgUoS/z0B5
RpUeJOMgH4EhlGVvM8q+XpN67LQF1inYfkft0KgTKHqi4wG7RRlMHU+eDdEwkgRkIXSOJSVo1CRU
fHJFYuwc3NIxjKXIzl6IkjYxKjjF9WO7vkMYeHpEl3hCzPkLBG58R7T2ETS5Xl/iPHBAWOH2mir6
QYFZFI8ohTjD6+p3zg2ibu+7evEbuspbIxlkbL43+edXGrNKLa1yRHF9w4Lb8w+50fyVdSN4SLJ8
IsVQEOcP9cRIBt6NWNUruVyTY3PGFVlhOoDPAOIngHK7FfxQ7ID8P9xKxisNXfDgjMli+PTpVkcR
D4Mew8B79cJqM72OVjvR6yYsmJAQaWFGoeOSNaOAEYbPxpM45ECocA69hG9jRUWWgEccIIiQt+pV
pu7o/KRYha6CZiDEdC1ivcq0vH2XOqdlDvyh6BjokHVyUuDrtO9YAsLsS0FUvftAJXIHDGFG0Uor
ScHK3JS62adtIjS6NMwYYyqZWKDghJr8XrYae8HM1GJS1/44mfkCneNCVhgmp92rL6W4xs8aotI7
3uzN6WMR53hyhH73ZOpxdS2Rkym4GFkO1D3+6hjPnQVyloSZ+aiSlyILcz6//AaNvqAk/8sgQ+Cx
5Gnge/2b1ICvlnO924mOu4VGM5guahZfns1ARs1XcEfZ6nhhS6IdCCEoN8VIoHT+1E9XB0M2Pzza
9tkdMwA/I5JsfIrQguklDwpk6TSPZ0QykWNLyYY/6rIj6DpgCMTFN1bzeAtYLs4zQBmUA1gRwTzU
Zw8Zwr8V2gSsxWfCem4x2DJxlnSQUS/R6rTfe7Uzc2kFTdDq5oPQ89F5ecHd1k/aGS/91FEZxmFA
chIlyWjgqaRkuzV6yWMo2i2DbwevgrrAdKFTJ1bp+qwLGoGYY5rS3mRvhBaECzMRXKmCyn4/8WDs
1XiV4AX4KQj0m2ysY2WSWI/lOGSO4DcTa3DWX9e/JHrXdKVF8rUcJsCNWhAolOdoBJ0adfgqktq1
WkvVdTUflHfqehRkiqmG++zKxHi4RICpWBjMKvgYiJLjTC2G59J1iHA6Q5XIg3IlWOfyZ2kc+Fe8
I7u99+ahbInKn0/15IU6FgVaxoSsxMZEGd/fIG334acGi8SzkSX2XS2HUGlPzwbgCAIjBNtXh2MA
tGpjEJbqoaldBdJemlxajhliFVoSVjAawfXJOoVi97+Ovm4FGa/o6qlr+tpY/ooCAmpigwNzrCLM
af3diZAUTo+QKh3oPfkcpilOfsZJ2X+nN9P8QVnaiIhn0O4lUfJk4DrPWnJsCqNbCY1XhuuHtuDP
xM3xzR3SMrZOPqxHOGNrk8Cr5uzMAyh/2zxyNi0rcINB63n6Vs4HiRMfPvadKPhYf+7XqQFHV8dM
6B3inikbRhVpZSiXgsCGuYNgqAyMUJWeztRqzEBuhd0rweT6E1O4HudmZDxdQWRiuCxOy821K/rt
sJ6LGDPih5xPqYEeoh8FNUnk39HH1zOuyc3ZUxJncly9V2EsBdOvjSGmbqs44uG9/Ou1tOJMtaol
+rc6DgWKtEs9/X4ItSEJhpgQNdoFe+bafOxH229atbHzkE/UqE7fhizlVw/SgyaNS6Y0YBBnC4gJ
HC4QIjvRshhOTvb8A3X38ToVz9D3+cH5k7P8kC84thXsjpWqQBaOXkEaPQifcRQIHszdwXAupZhb
tG2EH0TP4O5nK7P+xVmqXoyE4LBT5WN3T380vmkYoowy2LYNt+EV3n+ec+TM5UgLUODmxb+pr9aa
ao6baM4DFArtF8YuWbZXJXPPB3a0nxTxlfjWX4oJhqTp4pSvlUIMTpvHIqiGSLIkKy0dudq1Me2C
L4XebZ/w4tZSNHxDx2W22kM5LSAAvX+SrRGggIuqBHSCF6RuXporGU4CIhhs/QBARPNx3hZMMt+z
2x/oi5qQi3AN4MwEl7DQcmEoeyah03X0AMGB60kxYwQu0E9l6MM1XjRFmJ1y8spugpB+fOAoJ3xA
E28zGWuYeGwst8DJ3UvZR7QpaFAW3y6C4eHz0kCVNRSsgQYYsM9GoDO+xDgHESvNAVdFip92y25M
576WnB9vn7XbUBkIHNxKbN4QZ83WbO1H4tgGdHxdnXjZPw7M3xi8lBR7P5xKxE7kaFkemG9WsHOh
iEN5kA3Y/BZ8j7+s7bfxbNwtfbGb4P+mZyLiSlkuANe6HtaB+CAwNm3R25j4vg+rTvfSbRBK3fne
jGDl/2/PEAjyqwsCLnE+fiam9ByejQoA2LAX7tUQNnOoY7YfegjVNla/XB+tF9sFe03mQIDAGDLN
VQDkkjttUov8zED6m1hQghelF/JzQT0N3mOe2pwpvu35+2AqAsnMyqvNUVpZdhou1ZWUEoss/wTO
fpLFgu2WyuwLpTEYxOnSnKMX44r0EzMDoh8q82Nyxr0kxK04vhsXb22Kq3D6iEcYZabXH8fHqZko
wjSoY8IHR4lA80TD5vJFTvP2HwfdizuqKv4KdlWN1YnshZrzo89yiIQJn3JqH1nUg77xWjZf0gJD
quyj+9Vhfxp1ErPdy+Vgb17i4rkuaZ6Hiaf6+XoJKcjWLRqWunM2/9wKUh635X1ZXoUi4yq/wtp5
Ixwe2Sh8mqY/wvCTqTxPe+za1ztocR7i3bQvZhLIxXbutPVALOrdTdhJlBghrZOWeECIkVJncbBF
LM8OY8VMIr9WP3QQUvbyFxwk+nAwSELQqg4VOdpd7dKwd4zlOPIC4R4mIirCkQJEb4ntEcSP5e4w
3geuljhORun1BZtpYmwIRq982cBt+s9NQAEZN9MJL15kRNxNS4ECrVf50oM27fJjIDMhawenfoac
KJpCQhHV9RVkSO6cu0eyhwoekJvyGIC+jY9+FOuImJG0Hw4PjLzooDZm3i4sxdVe1dZXXxRcXmJP
hdF4H2eUtv9Ltteo+W0kc45YNR1AJXMQjCcailTkiDoJ182RDzN0MCNOshnZTsorL6V8xLzJBDQz
vyFnFPkuUNKteFfdzlhn8cRy0M62pde7XjXhGqlwmXQuFBPm/2XZlCt46opDU5INVe8x6OToORxk
LLa5ZRmq5o6TODZnXj2n3cZfe9iTAk7/eEtQP7iMvuGu35ZJo/B/Ig3wVwnLILCRRpOrrT/boBE2
4q3mBrTw6m4+O1aM85SwYQtdGKNsEWbPRlbZ6vqIN2sgOBnbFsgsFahcEqynjJzNhpJSGU/nIcgy
wsqCmw9ERl9gdhl7zaiAKbrdU5zsEadKsbDxOsXA9UXw9Krc+sKEUgDCQI8kJ79q7aGNsaVHR8yU
x5ec0edow/esurWv7YJmRz57Xl+UrtK1fi6aF1QjgzsnAKN18QboErAW5vIRZtJLK9tEC0E2l7zk
YrfeqAIcP5E1hbYH4UCH6ZTIhI/7fBQLnmE+TwRobvKk0A4sT8Wenf7rtojPvE4yr7DGbg2DQ/xx
CBvQvhDYu8SWhOa4lj84N8GJxe256xLzEQ1w5/orW893qYO7s9FLjRImt4epR17AUa53foTj/9oo
3uIaje7Od3c0zbuSdsdhQoYy6Hnl2H34bRcrWiL7LEVik0cSPYcrLIM/uMl0RaWtT8Y732mc6VQz
ayJdgNM4nddFkjkR2OGp40dJvwZp7mbbMHd1SFjY9I8riAiEUblymT7CgZb4H1YG6EII21qI50B9
2KO6OiNBeGXCw4BUm4pt8Wn5m6XdlNwy2T2QmhsEZJit9EFk5eZd34fFySZdoAnmJ/VT+z0fHJYC
mfTQZKqR27324YRy0U6NChu3neaRkWxs59vERo3OBaIOtDtl8e+MnYAPqwYIMcmV/2rhYBKSpxTw
rrlUB7WaAfYnbE9OfmtF+s6CeHGGzeAwHuruLaZBy7hdwaLLYtHpxdLC3XvDUu2MLqkKYiDQp4/r
t/TKBLtry6FqLiQnHDN3CL7y2asCEyzLs8s1XADU6/1k1Os6D7cYc/7GOWqvOTSYvP9yZcNOFlyJ
cPWfcYZadao+ITbw4tvWDMabCL2oxbTu+uHyrJRjzg6WXInh2PIxmqxfOaAtHpCUVe7RevWrKevy
YydLq0muQHuFMjLCobUqbdYh+4lyFMKooGrJ4nwcGm3FhzHgYBmTefB2PBCIMbmAmXdtpbVOWqC7
9vFJW4iks2vElGK1rxUVuWTCdSoSbPS6FdtoTxIl0kFCZeOGFu7F/gA7PJ5OUrtEqZhLtMj8Q+tI
5bnHhVwlwUQevOudpvWPY2wnvId5eqWNZA+T4jf8X38p+6xACA46knGRkbO+dSeIwGn/EQ/vcoDQ
MWI33gcszf4wnq8CQewPv3RPlvcJ4EW+WXlbT43Kr1m5qmhRX2TuN+NbOx/TaTK3k/AyK+uRTtii
o8Gd2SzYSMMlmqfDd6FhHkSlWZ1WZJFxsRHEP/CeQ3pC245qRUQYwcxRnopJlAmjvpMyqgKwSuKn
yJRA6bq9U3p1ZpHXe2LD2VEtO/M63PdggFijLrXdBPzxpvAVDJ2Ev1ABz0ubdEh9QfS67OqjJDwG
xNlW3+7Hm5m1fI0gc65JoUNRVHC/4u3byxMa1LMz4ysbXV+1GoXibBRY8Yb7zgowwQE4FjwJNp4W
N+ShboRc5cVyrp6sG0Zl+aEqBIY+xNFXuUYuYtpOhNBe7aaur3Jo/5ImeGjf1GuS6a3H7gcfdv7/
fR7I4SZlIup6/w0unD0v1Nb95wo/tFP230ubRfSzIBlPvrkgu7cyrHiW+rQWgcHf+XYGM7CwjZbN
nqfQPwfGbjmqQjZ9WgT/sZj/vCeDI8/8F/sbM5hC4qiOERRyOo2/UROGJfEb4OW1himqzk8pHDeS
kSWC7J0btTDgdOdO5rEkdAXHAchCBcqr83IxYiEBypjM3lL/0Fr+0cGKd5cnFi/YSlhjycufdscR
A9RW+i+MjLPPeTwAoluDNtr2Ey5xJY2tJ3vvbolMDUur4FVsLD86a0txdMgkTSqDgBNhEaTg1spz
yZJCwp+voKMz1fIIcog0Y217nVk3dXt3yk5SnDd3ka02XnwzWVjH5wJ5pm71zavVcC3ApNHC+j1G
59rqF4XCLZYb784UksP24SsB4sHPgEl8S08wNBYls60tGVGb6tLkUUnSrtdk9FyFN+N86xFz/vIX
pcihqaQAUKj1EFyYcsW5mnDDr9n+EEGRm9e1ZzCKr6mvFaYxFdgbXuEBzouOMT9POiC1mfyw5udC
6gWYn74KLnpqDD6WRW6piIB4+Xthzra2z4YGfgkX6ovBsj6O+wTVqbm/rLtFQD54/EpaHWNe4Rm4
yi7mbHi+EKvtvAoHLlrZjm8MYBb9XGkUVEgCKSUBYCNKKVTKvOIAS1xpg811FG2ouS5YQpg9djRz
p2Jup3N6+IBi7iV9fnUlTqdKjiOQOuCfxtNdGF1pgA79CLyP501QxhkaU7FyqQ1B6LcI+QHzFBYV
nqijElkepVcigZWIvL7Cl2/mPmNVOGIY6CSmNtq3kJUTp+GFqQNan0AgDB8JNIt68RLPXckY6sL0
GXTqevGzzJtD4CVuzdNdmeGncxh8n+fJ6iTPZz+PU/MvB0P+inpopXAYjVlIR4u6K8h0MobpVnb6
9G7OvtG0uL3Zkb1nqGht055I3boXH1fsXNP4KjYK/oIeMkZQfqPteIwnBsaKCYANiCBzY6itN0/2
CbS1nc1kCIzeLYnlTLDFP7d1W646RB3WWWpeR6yfV7vmEF0tS++ujCmbjpia96hBVGjLdXWRlZ4T
CNsNegztbMyBsN3wqVdapo0spUnae3scwDRZjT/yo9+L3h5jRPeY28lpFj5vLH79e1jH+3Elh99N
7kcUKVJlDIw7/uuIptxhacx3Iuao2ImFXtxecYTsS2tpwgKIACF9ZahgGCI7SSbif33M+iZZme7z
LQj2r9CHEnt1E0Qa8XRQ3JBB3gm5VLZzDg0Pt9gy4iMzzts36OaxITTGjUqWdijmaEtzGA/qZ1qc
+Uwiy/9isZd+i0Z9+tREW3AWcUEM/OHuLOfCyVXBlqFKiMsQ70e1DV9oH1A1Rnw4J+GfUYyQPGBG
6rvNsC6csygFX6O1WF99tjpYJTyiCnSfMsfYtFmCQz6b9xF99qt2dzTnmnN07hpPo4tlq/V8TKug
FOiA+2GEA6VDr0Xl6VisOFjGLKNXmuAR6fonXMjcDTN7ynrrWYUKuVqd/UJ1aN9u0R0h9EfhMxJo
l+Lo4sc7NHlaz2P5RHhYaE8OmaZJS9AFt327uyWQocE9ukKBNmcS9TBxebfQg75IjMWe6mcp2XrH
PCYHJp2slf/lnPeM6tPtJr7mZ4IvlE9mUcWiURhSNTkK7M4Sczwwp2ghP9fH83fmGzG128JB8HxE
J4T9OMtgjbHXvDDmFCuMCLGqpkjZaqkcyylYIhGgqtDqVtsRlYpuvW1oUKcNZyzlrgC/0SIh1S+6
HrYNhx/g4DZdNwhDOJ7N3j+BbNatdfJkOKTINCh0Z98Ls3RhXAvyPq72e1yJvyU7XhbUuLYqXOv0
WW/gwnAyyurFBnR/07j5zIABiwB2Rq5ZJj2m9Y+odWcGrbxwV3Q1iU+XNxtRVg+ijTC66PN13TUK
llbV5DjfZPrcKWC2OJrXmdvja2VDAAKB8K3FF4evtw8YDr9ZFOxmbA0Rk2x5RL08ZWg2HzVDa0dR
SdxWoUJA+E1ooUz+v94svkTPKMniKulR44u1kJR4K11Ahxx7QmWlktk4LlKU7Ci+MfbBu2bBTvOE
uW4qAKjzTI+zcBydF0c/1C6ccEppfCuB8mAXPG936DQS6Ofhc2WDHu1urKzJ3ltc6j5jpa+w5M6v
IV1TQpgBlMlnRXoqBb0v0KxoVx91fTftQK32IZoKPH/9/e2FkHLrzJwr3/WVfg9d86zAddSuMisP
On8cC02Cv3g5AmJ7967I/Ugx6kXPEDQ8iM9TBfKq00KyaUGKj5eod7gE601Nj0wpt5GAUlcvmGKM
vNiD2AgOb5AhhvZfr2xh6I+G5BQ5jfZSxZa/ZxvyhlRZWUFC1o3NKOQgi9z54uI6x7IDt3zTzXV2
NbnQAi7ZOo/p1UUHbxttVASA0t/miRF7Z75NzFGCb+PQ+bsWxWHZnURhLOcsmi+huZcDCOSbBSfO
LUFwfVbhd9ok2gPho7d4u3a56erRINt7zebU0KAvbG6qO6D0CC32yZhU+ch+v6lhEckZnfNK7IAA
+ezF9Lr8Nyp7xALzKkIGizXyrd+QAAiABVo6ZTt3JhH74Y6YrzLEHkSfV213SQvgkc7IzkNziGXQ
u3Y0hBpZBPm+qc35IEMVZLKM2RJ3P58e9fcS69V/Ursn2AcTC0TaMOCtWyDVhNJtmnRj5mF5Y+5g
hVZCXt75C6EI4akVX2LzHDeNyBwdfdBDtf/eknw5yd7NghJc2OtdKwW0oev8epfQW5vl+XFC5eqJ
ZYmADDni9961uyaCoaw89BIWf22eMRFZ8feJxyTUcFBpwYdsoIlE7+SfAqgBOdd5aIXVZGg7NXbg
wPbMqMjycTa0z8x56nrdqBWMeQXOh7mX5HPNOighsva5EPloT1C6391VmvTXguSkLWDZJF1ipt5e
4queoq+/x3ubEu/6TnYcfe8Aw4DNodP1sXCDnnKu7xudGuaKkbk5SHZ1w8oVbGXd9/HVEd2oZHJ+
VTHwG1uwnUq89R1p5GIGeU/LgPRLC/fE1n+w52FjykqP89xW/GEE5A0Dn9wu63u/BwgU74zMFEmm
HIn0nvQO58rDAlVXtiX9MoIUvhzz+ecW3v/Qmv9kYaA+fWPFYF0aB7x/v3R2qcyt4RK2OILdoErO
PQbMOmJ/IjmmLCJmtml7LUQHUy8B4TFvFHk2ei9JEqqjygzLdscObPwj1xuDXVZPPQjZvlCm8T9M
46CxbaPVdTd8aK+G3zas/8Pwwl/6vyGKU54QciPvE675OIs3V+a6wUzwVNtd9Z/BNLC7fOd0lepA
npcDmemLzPZc2W1Ps7bDX9oHBLZ50CYPgk2sZYwXwSwrLr9WAUZ9D5joleN+TdeAXR5szCaeUwC1
F0+ImQGLALSTDV6MKRRus+jg9uu/uKIodBXKbL44u0xqKbG4ciC2L+kylbOdI+ENJASiZcMFR3DV
i766K6yehIiYa4USTgjXA0Kej5AHRHA4nbAJv4tPpVDaS0AD36SIQZvL6Lfop0vy9ZIf6O2sX7+Y
cxl1JlrpAYDVUgXwYQQIlhu8cB6NDQ9r0IwCem0FHbD5z10bVEaGO25b9mhonk8OYehA8yABfxpg
mjm3pBv7ct7guCCv4yjR81hHGw1ht+fqtZCpJ7IfaDZQG2qRVNXjiT2vSSfaG+wc7A2dOn9NuFOW
qQBK5ZJQkPVPm3DcXUQF9gprLF7hGSO0i7sJcAP9w4HZCa3Q0DdT7UedSsuLNC3rDbNAsRRiu+HC
6oKod3YMctadJCC6zsmyY98NNTsXzxL3pE1xSvp/4RxFmdU7FuMNABYwxpgk7AbynPGAJoV2oDjh
kAZOGziok2H0+eeO7K+xY/+peDfV1lDS79KiYWzaH276k6W+g7alD4A9Y2Xm04IHPp0OhJjCkrgN
G+KgDSA9gVxW0CxlWKTbibGJYDidBBeCasyTZTAoyBF/kU8TtSmNgknPZE2BDrnZuMtNAv0Z9QYv
do6m2GhYwc/2wYFpAVPlg7xUSrBOk6XdkkNTY9ALJrsn9jvph/JQwm8rlwNWdUycZNLqnOUMMMND
k4cYYqqOBDpJPj3eiv8VQ+BwE0RLBjs9FScPdOXxrICrJTuD8pnV0IPoS50xs6H+dSrTeEMs3usB
BUBWwKKZT5Dc3CVGnmUeFbuqN216o8qaYtleDcISe0TeGxXmcd5y7eK0vb/2lxIgVE+ilYpvWcAt
NRyW5jZkgr4/Ws61ZA6zhpbAD3kTLHHHVOl5Hlk5Qtr3RrTGdKvXqNN0RRRgdaYu/uha0BNPYoy6
f62dfsrHzkFvMFjwel+4o2g7Rl5XJTuuy20G9uBLjZ/jlVZw6Otsu2lR8M2F9V2PV5uAbxbLb+Zd
C9fD7pxjlm8947GsDkTnnIbPF7xTbum7Tr2JXf1MTnYOEJzuPfDX5UUkFRZrwHKPNCOP+qq1feNZ
VbQ7k/VR/PyOj/1y/9PlHauFTtrPlLF4nCqr7X0hmgl8Kagn/21Rp0AJUKtPkp/2oa6XBepOskHx
91KXyx5laXuawtIkCrntkOg2fszQO1utEPOcG4XgaxBys6Z/7oB+ZxGTy3k8IXl2qCdSLYOavJuj
4hkRcUajBoCXGHnCQnaGu04y4QLTLf9OXDsU/VVExwA//71vY866s8j25Gruwpid8lhNEqy8i4nQ
jk1jMdaqYXMcNcPZAeI6CS58/wn4x/nyDzJ5LKlm6THQMRyrBa35XzVxIZRsh6IzCmPw+Dcp4H5Z
ahoIRDyOpVQ28qas/PT29RPfrMNL9puzsmrCpevgyrcutoRXS+EaqXj31Iep1of2PFKpx8tQYCS6
35eoeAATu/lCWM+KdFRxOsJkQTY9Vd3wJarenOogChYsa1S4rA7Rufb+ADOa6awZfHbteCjk4f3K
EMVXc0HLnVpiB4MQcx4CMdhUXtda+z0OHw0Wyjp5OwgaFWtnO0gP27D0VysiBrrJU8Y85Kn+rBz7
Uzm7JS+gS+cL87BhZ7568rFUNIwc+OI3ksX0P0JCGtLo9Ih84ptHGkR7sXfirSUnW0bkV0qR4tS2
k+aXbHmV3qZ8maS4BjbZc3Rkdrh8lAzB2UbKSr9aye6bOy2Qzr8X1kA6S9jCaRMvTsldnL82ZJ+e
9yAGCmZYRvgxZ2DLUWgUkC6E0sZOAdKzn1tLIfQnU3Sho4g9MScKOg97/B5MyA1kPfxbilB6pBjj
f/KaKRpspXjxdshTZOYeoLKuhx3isQcxr/XL05HflurBHlGYYYGygcPip1UOVaMIvmCzY1aRDCu9
P0Bp0yc2MyCmwqZ8CnL60IEKwAwHkRdnNM83CHahMBLRQ3bqIKBXSvHa6vRGIoNPBqoWCD6cFWQ8
92b/PfpvmuY72iFJPEQrkmXkrnzM5+GtkaM0GTh4oOhe3mZPlu7SwBEZHiv1UbU79p2W5016H7Wp
EV/mqsZiUKN2WQrsA1f0BCUJTKYUpYMLJ8j6eBh/xGgXBLtTR5qepHadhjzeE+Pl3YxO4uPZNAcT
WbAwfM4m9mqJM3F8pnic0ubD9SZp3PwJKRIjy0IquYYdEqgh7+Jq/5y62cfR8V8QraUoDFT5PXiD
1KO+WKSL3esNwW0Ekf/nzNEqOrg0qUYUAyCC11KWYDJ6R91xVpE1NXX/B4dtHugqQDmv5Mz9xBSd
P6aAZTXxjuV9YPC2OTFIuPYP26CWUvdEBQQWlM866X6yH/2ZaRPpvZUS960xiPzKvqbOp9MEpljx
AKyoVx/XvJNtm2pEPL1+fsyAxe8U+EaLyozpugiQOtL98SNl2eewJ0fsP0jUQpwlUwOnv0LINNCO
SvIyQDnT2mWVyU3ZDSweFmQiQhzzEWn5J8Z9nztBVFnMZEB7X+dCugp5DfDgjjcnhyCBL5YRgNPI
beVdmUaH8p5QX5S0Sjf/7pKRcIEryvGcOP8EYUEncUyxoQOdjwm9GfwNLvy7zeQng8jN65748THV
NnW4UQU0L8/Jvk7Ri2W5Cni7J6aIuus05ueUgmU1V4+/CF4XR662Qnih01rovACzXDwM4rhA4l9j
x/AqBqhqtFbjENlMICpR3HoObSDCnhqhE3r/UeoWG51R5dwZ2KEuTWXpJE41ffjkk1kJErO23tJx
aPPn6oCilbZF5gw68dOZobW2tNUggAoLHlhIAo3FM9uAD0Q2COXMpE7lcA7pYl2vT8eOEuT5GhLw
BPjcplWBp9iJahNtC+Yx9aXchVvlY28tMQiPr23YI1IyK2zyNKirsZv8IHYd1ee4GX14M3GRT2B6
K83qbZJBmLAkUVWR3xakIk9VX6IY7spjOoa0cN2nkWJJ2h9Q9DfbDgeUXY1kPwnmf/I+NKxLUMn6
LxW5UY++EvlWqMLkB4WXMCFziCRDWWjzbZ1IIdtMZy8U4biXpELTS3TQSgIjCIj5oV/jqF1kSJkC
U0vS0pdXv9Z83UzWMszYWvWdOznV+uWqXhsaygKBuBf7gE+1PNZ1p3i8ypnoBIt8iy0Xaf6ZR5Xn
bY+CpH2Qu6KCrGIBxGtw5C9DJwUqqiT3WDj953DskDstBfLCAvbrHxk1tT281uWzxB9gfYUl+GDV
dtEUHO3dwZZPXU+1yI97hgI5FYK+YWKt3A7ajg4btLCA3nYRoFieCHlQzokuJKRWS9pTfASWlmvz
VTJpuOWPE8pggighxBI+xSeTepDcYCf5GXDpWso4/vzcr+e9RvxazdUWmIIRHZ/PYW4mX1DKXglm
8cuBQ96HVIbCiQWpFs1FWWUnwa+v5BXQvZqOfqpAuHF9RYIyhe+6U39fvfI0l/lUkIt5/7PwQl3s
Cwse4EH+jOXMmgmlOwKNCj8P4IhdCGK9mchwGN+/BLpRZDIk1/NqFTwd60i/cBHrfTox0Dj/HQ0m
KaKDAT5skzE2S+PIxJ121zokrB2A4fR9fRaOJWMkeNGH2aXtPsyxoEDdWEUd7aBUi247f9bVqw/D
fDgUP8cEw8w1VleI9jEmULq/JOZNU7j6AxYqexzm3w2EVZpfGsGuc+kpGh1XyEnlplyMZkn5SfK2
iygB3tg5UQqOgWNmd+oKjhV1eTCG5Q//v4G2Uv9PcEWZlqxO88xR4lQcxvcvROdZJTsm421xq1BJ
MLb1agJIWm8vVgUD09xY5Dg+GQM11jkHqMKaqKpAz6a77VsOzIPFYMsgisBtBtJRhfEKU1OkokW+
Kk1VsGaS+y2l3Z3eKzNU9wUs8cZkuVfzFFQMbkCAgarUZvlz2Tne0fV71kPfMkQ55v5/hwMUey/m
EAaUINahmQHhktjDU2PZVP22ujbtQXqLE+VLLJcWT+TMAnNt82+tjktLTvk21EQDvrsbvFRhX+3A
AMmTRDf+ZqIc1mjHxLhoqlMa90erIN8puLjZIkVj8+YTie8fkTZ2eB/pKn/T9TWbBhtKKBjAI6sJ
xgJQlsQRh3Z1TP5XRB1X5Mz9VzrGl04lTOu76SrxVd3ti+JJrc3e2v/wA+DW2C07Wf8z0RagPcb9
vazTVP2OgHlJnw9mAq4oxGvokuUpsqAE60FUft8WyJncd9SpxqzbkMk13mXaIqDy8HPJ07XMMk/Y
5BZCeYhXPlnmPRYwU33/SK510DkrtJDwD/c+pEsxutnSHTcmGDjccsASA4E0ro9AcCHnnyctpa8G
pwbg4yziseY2r3FboZ0BrV7wclmzjYbY6BMcQCzp9mLujwVjGDKYCZm60AyteOS1S8QPUuujfGRo
8DWCZh7a14svMCKhS9HvbCtHqliyNU4AFlJA1QA1yCe5XTLUxQmhfdVPo8lAa4703fNBuBk5Lxag
UP1gLJlMQDx50L7iqUesL49o+jmf+GSEL17Hhz8uvz2Pj4sOQjY2zYPvR9CCaVaVMNuGwf6f7t9r
tNptVcLy/lZcNJ1kJvY9Z15OGDKqlR69kc8VoqxrCfplyB2URxDHlNaKPmzL9aRatatVmnkl5TIt
DvH6r/6fB9r3Zo65JZCgmgHtpF4ngu9Q9I/EKfjdfiltg/fhGxttdDcRWjG81H+QIqRknoDSPQ6f
weEIbExAjastw/4Z4HgO8vhXvQW3ZtWcT6xFX0S3Onoby89ujE1S3rzpoEV7QisbIPC6wfPjxj0M
q/P3sj+hJw4qZKQ68y6nR7M0Rm1EQy7PGjMAhRhHXqU5iSAhQVhWMtdWs3mXm50jcR3ULiTyXOWF
MdosD84I7Cc5KCJO0fbDbxVLSf/Cnsn4BmDTO/3Z9gKdXqg8NFDEKAY1RuvC6ynrd61EA66OR8KR
tdUEqhyrhyCa0hRjsoGbNl2Nlfe7DIJhHHRgoIh8544Yn2UmxDApHdNxI9Gbx6hL9rAaAK2NSEPK
m+8sBjK6Ae5T+ivJs9Qd3mIOHix04Nf1v4SsZzw3t9sBDFdTUhbG8oEo1zimPrvkKFTwiAy29oYP
N9SGJDhi3VwLwEw6136ah/UPARBxTohz9/lMzKZbCqoqmQUPH7SS5LY/Vqg9sX6/efjd+NVRGB2G
47lWGBG3+BIKiXbCepbohhlaC2EYNvyrMazj0m8IJbrbuKEoXVXtivs+pj8BXBheW8ML6LUDpxKs
8GzUtRe9g3cs5z3gUmduP6uNukKsQg92CahUOWiggKLvMDFS2ARn47YKutkk3IHlV4dih1eKQxyy
tY8ZHYso/Qy7wKbhzIiFSRE02c5H6lppXEmtyusSWnYRDarjJvnQM+t3bgmKrSFPqXEgaP16AZEQ
0SFDVNfHgWtYCnRUASHWFRnuj05AxLZQpLNyZwKOgBd/hja5p9BtyOkVYwb1KvtPH7JNFAdi/7OO
JxQ0GFfBdo/k7BOoWX/G6zvm6OcokZ/oUJWDGcF8vmIEZtTjDp7g0uc5qSS6FQiFl16PCIUfkM7E
MY2ngyG1jMlqfMA5cWJ0JnJFfPmw/mkw11rnXZ8tam2FPsZl9nj/qUGhJ49x7+xXo4ixNCh3oJDU
eBAZg+Kp2pIwjhp6sc0eETQnf9W3OF3yG7tT8qHJswTi4Mr6YbZA9P7m4rGp2tuswU/YVgsFaFD1
F6uMfvZaIplRsy4zfW/BlTX1o9sIzAbtVZxso+zDzVfJqpT4dnbtss4Ony70vNueDDeSdzUFgoWj
/O9SLWYGoymukKo/EW6k1ozPxmEJLBOljNkBLitMW+Ir2T1L788zGvYCRM3/toM7iz0jHGy7kE17
g7Pf2mpF4SmSrkk0u0iX+WgWN6hP7zi0lmMcPOlDoj29+GgAK7DdDCBpyRZhF6yfUxZA0LsJaGFw
vM1IE/zH86sd1wFFPUBrxcXsJptsSJXvAWDVfj5hKGzOAGmPEWDsaSmGaZ6IBJLyn+piPPWnsSCE
J4ba1W9gR60VQrw4SiN7rTqoBfc9AO9bLAsRAYbmhvSnmRLGOsrGOydrcuifskWBFNaoOb6SvbXp
OPxdPeehlAW58WywGkSkLBBPELk6nuUIXE/AFX1br4cWypAvW4nsm/76+8mJwKFHNYax1rosDgdM
Td+0sDjoBPQfq3nZWNlOgdPC93kJ/a34N1VWA/yb35FL/l1dISRZWtStPh5u9DvBRlcOM06KA5Wh
tXessELxxj0bxE5ggIWH1Sn1W0l4hEy4pigmwnTxB/jS7otKXKjJSbdd0PiROTUGY7qoxovh8ZAN
EaS5fZDZ6hcZovJxYk5omlwjWEaZVRo1Fmtcr356WmFJOsxxaDi1rK6+d71+hMedauYa2s8kzEua
dQ6ermhpjf1ek5AWbbbzMh65OucYmE3Lf6c/z02lUzJU5kkl0M3Xkfm+x2e616/kpx6byz9IDQ+O
sSMb4dJT+W5wKD3t9R8f4tKt3n7v329pBRmQZrD5nJrkHyTMOxwxKPyz2qhY9Gj5591zwqYwHRUk
hLsP5xXm/mdx7ekFdAiXfE/gLKLZpgbCmwp0pdLPPtvai0pQGy44VTbjiQYbUHRbGJ67MfN5kTFr
/MasElgEKMejvliT6jXzF963sGOrz+e+musKdIs0kLgTknJkDC7jYsviP6WeMENhbALGKxfvcZOb
EvaKVb5Y+M2hxNLD04a2FhJ00SsBUhnP410dSMSRXgcR4ID89qHVv1PaHL+fVrRtzzePiO1h9CEL
q5KWQLGFwgQ925dV1k+qfb5ufhaF5RpBZU0RE1vhp+2HB26CELNJzOxN44qzO7cLRNttHSRmeJd9
X4lfy7HBEI49gb0H8DNvQaSmU7++ZzApFYTjGt8fu/z64EZJsB5fwimbIV+v/nt/OBquW6+HdbYE
EjKJE7ymhRDPz6YaOw2R7e6vR8Q4oq++ptyQ34G62z711TTseoBX5jEOvGy2k8RwgkT+axx+8gdO
Gig9PYHYxyd0guIHbCdegQ/IPcXOEENKS39SZ0iw1uTJ/btp9nmmFt4kGdy+rY6YRit77KKul6J7
zITPgkEYIt7Lz2KAGczKBWCowQ8wBxHDJMICuw5oFmm6x5KUhABvLcL5C+SLx7RDlcihSXs0QxO6
ZWAweivM5g/0yj26bgs1jXVd5+LHlbI/yUGNdbGjX03O8fAwtyytehIy9NCbkSJw4lv4mINukzKo
0SxqMNFkBicLIC/scjaTDnPEH8WgggtpnWfCqWgNRSc+ESSSO4EkSZ49txgRPgtcgaaVF8Aa8TRF
F7s9BbDrWtBIB9ssKEagGV1YL7NTM6b+dANTGPZ04yX4k2pOVqJWOD1HfUF/OHcO/mGLfKuu22Ay
sJK2nBCnOZn5uN9QjSMmcA6uqESahWqFgtwZLmWgkVolWxZ3FUZq1ip09Kiv2o2lY8vHJwx8j9Nn
k2gwctr2IdJQjjmcNxSP3o41UwK4D7WnNVyzbEVIVgJmIDAiSE8TU/3caA+posqnKQbqtspTf1xV
CTfAgv3VIVFb63MxF53vLDNQS1SSJrV1AGNwtsSKrnYQbUtgeLncBMdC+nDF8X9eYrBlQibrS28F
1JGC9uQwYvMh9piXhetiLctn5KlqncjlxevKUc17e9urz+ZILf2VwHx3qHd2Y6rc41cOi+Lq8SJh
nWup+GWdKiN+pGyuI7i/PmL6n0hLMF4HAJECpk65Pka20EWVfmmQrO5yTehDx66hwopamIfV9AFF
2/fTvlhQsuhKfP3loooKMr/Dbl0jAMcLJJg2PVsNH460s0majJRDjP37VnKnGvLdflIQ/RMRQnVK
SfYqZwTFyFF4+HcF2g/7gkBEJ7Oer8rcoe4NFoc83d28JCSmD8C3DIojdqBku0p8D0xjWxUi5Lkd
SmWKYXb5iIgxkdxsUR4sMvpfPUw5QoWyGCrmlDgPo8cbiBuYKClwKWtgqQrZQIvohO8vfhj7Ab0W
DHfuF2Q2YhkqouYSl2SjtKVEfRw51ELSbrIoTpDapGTvVaPlPSvi9o51tqobMmE1y1uqQioXNrLm
JFafmFdZVeomsm0r1JxfgzTlcXmw1ypqj6SHJV8GVpFx52X6z/ITj0wmuifgP9H9+H1AEhz0PRK0
CLCEYubA2q7mI+zw/bCm4Zs9rCFWQmvbMEqeCuKmBUuyDn1fwef/U/8/yOwfDhQ7hvfAf88L8Ocd
xn2unJ7nfcXgnWnFzNZDbVA/S0EbKjJlx6rszOamxHdgkkjNb0NjKW9tEhPwya9Wfmb4C9dqpDNa
qBk8CU2N6LQV6MyaVxOVgF06NMeESlKb++0+0Sch5Jyvs4p1GKLTzV3FtIyp41lJr/T0i9MVR1W3
467OjaZphX8yYiBVCOdVWOjXTCqc2NoWAlWSPj9ot6U4gTMmNtQxIKl6as9YGl3rv/nIBasiKCzL
PG5HjVFJls7INf2Zkp4Hfj6bBkSd5intYqY5aF181kur4xM8qFsdgQOh4YM0i4SjodGN/i/ONuYL
O/pl+eMo+efK3A6ORzlQKe12np+ucS7cOjmQfcITvzhJrFXdja5eI1cgUVRwpLY1jFOvPq7dENX2
CdtEYZ3Qvj41x5Xwzg+r+qjUgMjDD+5GuH3GasRTeIfcMHWFnmh8Nd8lmXPVIi5jVTxBXucWTVmD
9mEYwjUK9Xi24Eqz/+/uRWevuRNRIhRCP6410Oj5DsDsjaRK/BJlsw9XgW3DjQgu8XJsvr0xMN5z
S8WWgn3EIbqjlpeVYd9myHsmkSLIKxzYy474pEo9B7FDuTuqXiEUJ1qiA6rGRcRNJNSJoHZZRi4r
1nngP3mFK7YOqcgoNQHxfNJDoissBKTpfI2JxgAmCAvf/KqdCiJH3iVPcLRFT64LAMqZg0VnI6ot
gZc8zK23bhppkVnBlSyCC4CVgHX/0W9ex48R0Lb4NNpt0VeRsTsyZTn7vDwfwj7GFjiHD52BMP2s
LSLZifM54L3sj3BmYLgCplBISThZ/WRTtiK/q2zaKR+bdO0LA1ruUqPJBKsl8hJ1voymlYV4SRC+
KQT09+b4BCHPL5E9B/7BNIRgSQBMEg/4jH3HGENiE7DVT5RQ2c8mC0tJM23dStYWVtxuATNwQ+pB
MgjGcJ0AH2VMjUWXK3JlLMrcWn/0YwL9b7EpmWfYmvXsZgy1HgQsW7/4Qq2OG77wiGrqqzlvJtpF
36rSXEfcCFPynJ+VT/FzM6UAEmp5Dn3lNoqPwdNysI7v6LetAkRzWQnSH6bL0ra/gGyYivSCqhzY
ux/os3KyPJMogkrqD72qFx34wmHw3Ghr7K7mtaNIePfOeeQ8s/i2KfAeuyr3PgyGnn5Kp50i7Lu2
JNDlgkqaPnHsmi8WaIWa94HTlmsLYReB40dIZbEfQ5PtVaSAHlFYtPzXWOJUwI3kgpCfYWCn4Ujy
CQcMxZpIhRRc2zJLtDPjQNsSmbOaUBh8vYHv9kk+eXjNAa+2/FzyPa6e/InCdLjRcPqP1uphFwpD
nY4BFWEjwKs2agLTnLHdUjeLw7LX+kmrvyYpbPcKTlWSt3I+hXCou7A52a/2ORYSQuIagI591lXz
hl1N5bGxK/bLokrq9HnPhWZMxEPFGvS4I4O9wpAx3Vq1sC3xHZQeEZWphaGNjhnqw3wl1NVy+Wd2
MVG66QYlm3Vbq3SC31J2lXWpMl88mXLz0hmRYMbnJhlsxqqbEipNTXf6wdT4q9Q5L71/a0lLyR1f
h/hm173+/qfzytRNT7meTtc7HAfqNxQ2WwFdJnoo85Q3LgoYMHjsDGABZ5BBBveMxev1VWkKdNAC
pmFJQATwpI1yyAH/27YlRkhFZw5j78gBqzUnrv2EB9Va8PzAjzIT9ylihgVneKes1QKsd7RNebeP
VC9eddcbnIAU6Zvej7TBlMPtZVsmw9F5W9OiRQyh4IJnoANR/HYB49hEYLG7D66k6akTlO51g1il
13dIdE9CWPnqZvz+twTE+qRM5MELk0UwypCk+zpiY13oIdejw7uUg6Gk0UfsFh8OwGhKU+80aHwf
arh0+VZCcUcmD6gHIfSQMRmkGSJV6nfcCfyrijmggNY2gpJ6H4fqLAwH1KpASW4UjA6DOkMz2N3m
/731iAH+L7O6zYlYSsqZiR02FgHALW3H/LEDG0K3PBc1wlKIvhR0Ucl5H54Kmn3h+Ks8ey33ijgM
lNdIPoB5emHt3rt2/7yauWnY2+ETqk5tgRQEZ+7RVIR8EdP06XHXpgz5Ho34IFQXj7azi+DdIZVP
T81if0RcxkiDpltavuMJqCnlYKRC9AwsmoE2HXMp0ThGB95Zf16P/VrTpD8CRT89uFRfj3mWuC/g
QKBuzuYO/s9bmKiistTW/Nxb4S5ITvPwp4LyWIw9CaQpLpsIJCv6c2mB9PRgMFS0SZj+VsDvwQXG
72c+RcSbDefK03UnhrgfnAhLFNFGnXQT9RAOaB3XgoCsItDMBAs+Xg/4hS+8W7sKHZQKByvMlyJY
axyIu6rtc3TZA2gf58dOO7qyU9Lz5kDTeybic7cJGbboYGNrA0nchfMScY6kwhPPePaYun890w35
KZBdDEBrXkMbLsA0ijkv/b8+J7OiYSXSsVQNa2BXgt5cD7lWZstmT0rZVzWLuOKTCCd23FiuUoCc
8Ha665TAKkGcsmmPBXgWTRKhFqYI4rtUrFHWO/cYJOf04+3RPIhJBhDCMOMyq/D9qiN1vLALK/HR
R20hoBatw7sCWFmOlbnTePfKJW7ZS304Q+XyobUzvehPlejy9JCjM1A42R2yuJAiWQdh1PD/7l47
jEHsb5UUAX7ppIjHRp68NtaXOtXCH5l5A3eqVFqghfIlEAcwsVDlqjhi73vxgKXFM+XSFY+T2JeF
WfNQQXpscjh0kpgDOxd9WADTs+FCpnqBMBqM65vlLovvVtz9r9zWUqyRfPrw6am1W3yeil0yU45D
m40Hhh+PVNnXAZqwAkRaHOz63jtta3r+NtA8hvbvWwvRcZL22a9bkSyBmFFjnYpakGrzSeuCrnez
g7wZpzMLoNMAfKaYWfdtkRobYUNBZ6loV+W1O+Wr5MJcuGME/2Yz3gyDqfjRVugMFaX5/9HDHmxV
gfC3jxk40o2PqZaIekQxvmYf3P670naTEOogACCMFzqnVM57k2PXpzP6eEpvkxlBGC3Y+Hu1AScL
xyfskugnlrf+LGCUmBIuwJbnHWP8Y/qRXrU6FgC02Hn8GTf1HYy+3vq86w7zjn432NzMW4tE5ixC
FeTXtDiusz5MEwk8/D9IoSfdKc1nDMcvZbyrGMwm6Shc0EBDgEOFVLzfij5D7oaymuPNW/SMWWqT
DQRwIj0JLTDzzhuEjPELww7cr3y2tLptmgPiSzYCylecNIxDjTeHo1SBU2oe+DsNHdFpILRH3ZXJ
XZ6XyHYNPog0fy3E2n8QmvOavEhjNn8Rw6lchU320fS4QB8YTkIdWcmz3aSIxAxgWgnYTSZ3d+nQ
IEVoCdgf8FwJSC+VwD02FyFirAnMotXkM5GrgBJh8lglgie1jLzzZFoTFPE7WFEY1y7yZfejGrSE
mY3OKxwfC8yF5K7iy/9FqXzTZidJk+uRdNjGFA4g0KMJlqbtR+9jtNQZSUfSLgvtQllIVMmqZf3f
P/rxk4Zkf7ODivXpymhH36t4/wcylqiWSOGiRakEolTVG5bj/fTi+AntfJE4FIXb3++KGTKM75wY
pbGkWoeMMiFwXH8Wd6ME+0iBP8+n1r53xCCgQ4B5GOlffoPSglKIfhAaPt00HXegi+ulOnbDudbn
woOu0mtS1VuyU++3cYskQo/6Ri4QskJenWG18fdLWEFjh9sQmxXOStE4FlexvsFqlaKKMuDZUckf
800QUbzgzAwC1dxrpWbVT4ZhKwC/c63Z1r4FBLbn3zMkkziseeKcH5UIazHez+8EVqj+r7AYdXrS
H59ZEYe+bOYZLbGGpAkuuueraUkx8LrgXHbpUfgtmiD0c3IFFeYesj8JCMj/If2s1LHlyyXDcJVC
fJeuqy0O0w2T0IJ5wBhgYye/KebSqYt54mBwZurHyFdLMXnXfZRadOc5C5ah72TJPlgC8K/oNhzc
cWI4SUsjW2ZcycP6eC6C2teL5QAtuc9Mc5EnviSax0oeN6OC6t0ZQy1PaIlNb0VtjH8Jj0anxIPO
KRV9P7trq48LNWylViPXLBOJ0nz0qr4EQvW0MdZg7p3kx/GU4Cyz5ZswhBHZ6MWBl+yuXH+p3aot
QJPliWORtePtAgqbR2hCINPPyiPCWMJ4+TZVxRzC3XhCOsKbNj9ioC0hu9qUg5RHSsmA2H5nmmTS
Dczjgfabxl7OB1sboM/V/mQXBrDp6nwb0hvO6C0pEDDUaX8tWCuDwhMTkKqvRyXLC+Wiub+J9ISG
GKYVrRioPi6QCgbLFcQr7aTQFct8RjR8e3pAe89JtnlkldDrV1bC3dkESYGdRsqjwW6rhE/nr7VF
JwlzIcyObnEEkWL++fF7COnpT14tapyr+5cCcapWuc6ZO7IO+kZtWZpuu1cRy5GYRFUZW22cFL0l
ocliAU+fZnfJL5aX7u6j/a03jGHCc17/8xzIFq682r1iQhXK29OjJeWuN0I08os5ULU1n9IRDANA
cvaKMnu7zB/eZCswrZ5Ln0pXWkU7odkfXsz8lHny04xTbd1kWzXadlxApVUFnI6iioQSzuSlUj5y
GV0muy9TMllYe/ooT+1rSrThwrHsazJlwRC/38bArhdyHYrYdEF2rC4guMkDlG8aVf9BgqjGIwHJ
QCB0S78WD9mOzYaSqkcl95JzEY8emU84/71L4hhXvY/2D5amXYUEOzwP0wqsldJ7r1AjnihBYm5j
VXEGj3vsHMfWIAIYv6kp6xCAdsdfNmOrUXpzlal5vPHdOkeVy6lVjzlFCzfzT5uxQDnTwOkaujEQ
dw7KQQjNZEzBZifdX/L6XE5eWF2aFnn7ezBR64kL2xwDkLFIqdy8twxBkqOxibIqUhhjoEc3r3+v
R6gtSm/+IYFqypSc0bJBb/OSBJ6zPHOhr+dl+mlLiqPZX78PZLB3BXeJ6S/rSxPcmx4lyRFYlyRO
VY+cXnvNXgQilkAq8/+VU62lMJzKeScn8LQ6WI4zQqyiOlj4OKTHPKd3e0LbP7fEJJhSyCN9TcMJ
jq2sAP+P2j5Y/4VJPNgjD2a6avOc1UZmu0v8lzYkF+dBTSdMjkxCtK30am3WmlTH8SrtMdFRL2Ve
oFxDdPbUeXWs0XK9WJEGRhza7aK9CyIyQUpNHgF9sLlF5KYrSIOOiIrJ1fm4liu2ofnRN6y884bV
OW846cbPxmws8quISoEJ3VvZbFMIoQumgAvLw/BVcFyE8OD7/qBFDP5ayWxAWMMZpbWw+rLNRRUO
GFyFIVhu1K8sEBoyD0SdE5hAq+Y+v44gtT8YugPAa6ofKBx/IOc0cr5vwVf1UR9+3zmYxCb94tEz
JkpR4YDDJ8z6YITyvD8J9v3tLcM2CmBS6ohKny27FgrcE+KgINZiZA64GlM3nePJAeiUK7LGugFd
Lvtscyzat8nK15Cd5NHZjm7n/VZEMFKfe7OAoYIPhYNr9PFnwnS6d8GW0ovWHLdO35ircia5Z3Lc
6GPNDdF4TP8c0vjGu0W2Zr0p9Z4+AaXzKvC/fjFwc/4vy+DUs+NjSb7yuXZcNT3RVwBCP3jWrYtp
4rvIP1uZzBKpsA3fGU9IDGkiRCXN3ef+V/y0PSNHdoV6TutB4YEnpIdCKikjrr4oKi5kFxytyjTA
byidtcLt2G0ujU3ByTweVoSdC0YgoHkKpVClmWcXt8UmuBn9dOYCSM+nOJdC92GHRvwqX7Hg10UX
iaFs2FLJTwm4XdVZEg7q+sxpeCkNwdkjhHT92cG0mXTDMtl/CARDsbjg/rZYP+L07dKJsUGOAMa3
Kw+LpulOYCeCfVL9KnDLQHgYpbZfv+l1UgEeSLnf5HoK6kdTxqVQ4HfDXUtBZVRFGgACr7J6ffeI
k3ZD6d/ULBXvonavFEH8LdWPgciJQUkLdc8a99R/SwWlcyy6BrazdukFNeyq85zsCu3PthkZUg3A
qsDoYT3DgwNCIC1AvscXvGTGVSZGxzotRbXjUuB98kF6wdJHRhqignw7W/fc2mib+t9y883vI8Kj
Df91fgfmL53Rxz9Zy3kif3XUySdBZcqjJ5pwHS2AsEi8DxtqAU75VuV0x2nz8rSvvGI2TpvCAP5H
VEZA/lNaGOIp281QbglrlLmQXCIqZmq3ZcnUQNOXsc4j9nbKLntxxQ/G4vOgpKzx0noklfMOQTcM
p4Jie9VpqXzNF6EsRJuX30dEiY6Elr7QKB3NaSyvssahWILAXmASU5oMac3DGrHdklg4FqFMrgv8
llix6Xo+KlERx75yApUSZuoXz5K1EWaEmWkerQ8P2V+J5/VMY3bnyMRY9ngMVDZVQ2qOq8+lg62j
oduzgeDuo+R9p+TTIneKR2Vw1i08EDt0sx6fkyFbSJaArGBM8NDYIDPWsHPY/tcfmHI2vXIhsuHh
bfD9CDZAOGxwkySK7n0qwhYxJy9EBpyUuVFRO/9BAfjRO0FqukCxq6gZg0ZDKI3mfWou087q+vgF
xt4TfXBfHofho+rZcDQgSFpCN+COcwohAv3qDH+YRcisq4y37H+EjXMZATRsz2L0Cq4fXh0+kf/c
kAl2GtupZasBFuN1VV2IVe7FciaS5vBQkwqXmy4D2LvBk3LfTdRKaCqpMpNeK/fNNbEnQ6PXPu02
DdAQmCDipLrsPOgS1k0xz7VjSXDMEFM7wFe1DIqzy0ANERfhYM/o+OQX4KsqXlY2nTscA14wRQMT
eCXqt7brZDIA99j4djb3laqXV73Xeoebd1NwCQLMj7MxdARAGndENSnXtITrn60QqDwlzknSfz6x
F6arv8n7Ejmn1IE+cNt0ldPz/5DW+VWzd8l/65V0aPxXalymlso5gb5b/pI7ccxqAIIl88MK1of3
IjOyZNvhER5PCHn9arSWc76B9vLvhQWfcj/CSAOedGzP0c4y2Ah7TTZ+f4H/F357ZQ2jCpK8+NnY
gJUe88T3JVb2XB6p1magDfjAtxQUb8DaLsYlN5L6ITe+Od+BwJp9b4ebh4Tzv6vhCz1nXgeEfdHm
puauKxKBbTh09l4Ep8/hqaCAcrw5+G39BJzvcKmmA2TaWNWF/YiY9na9bf7hWkwq9mkevH0PBsLZ
r0nFNdADXrYw0geKWPW9A2IhkwJLjhq2vn3MnFB6sS04yH6jQsF+Gb2KAgYsKnyvirgF/YE9mKc/
2cuFg6GaVMLMuUtiOaupbz8hSv6WTP8ED0T8WfCGutZx+Cu1rYDbHXKBSGvc+C+96cEY3AS02H46
anPcH3dkRUFW+LsHmllBsstJKihMoAmPfDK6khHccbZJgl14gdjPa3NrvyxMS4/m+rcK1+CfBMe7
SXX2lM/0H+V7MDT6KgJU3w3i98ajsO3IzuMS88c+Y33+P2sniqjO7Jk47BRLwC69vAf0Ss/jPdo3
Y7u5OhORIbqdm3Q3Uje4ybm+albD4R6dlLaia7/PO3+mi8Dlgs0iP/RfrKOHElElVVXesN1sHOP5
69UKvc/mBkCPenlKIMo06Df+yD/+NCppMxTdg/ZZJokV6RIht3//LwGJd/nGJXOtqJFZUL/Xjd7c
OWKA6Bo30MbcNr9IP7z7lJbF4KcN7QTuF315/dzIQOAoK6RajWNryzJZSop9XISJ1yWVsfDC1YUd
zQcuQeVFTTC3Vfrr+slaSyLgTC0/g+Lf9SEZak+9kw5PdUaJptOLM746uuQ32HXw2TiG8BnAki0K
urCmEijLTZyHsjFJ91afh3dpit43qDLm+CP15UyY9cD57HY4mvOJN9Z3VL00T6CXvu9Hlz/1goD9
MkQgSSZ4dn+flbamO/KsbfQnvWB41KLclhw/MT9i1g9DYigmfmfGKxMn0w1ZxUt/NW+8KYRiWFRP
up9gTFClAa0alpVKzl6LLME3GF412JFFbqGu+5Sg+sx7mN0/SQwJxrbq+Z+/Z0pBnsKkwBspECy1
IlmLLUXLTfXtRXbEFry9+VKYqlu+jQr15ZTZDYGhsAF10DOjQ9Bi6bOOFCzmrXurR5YJYIYrshGi
bU/Z5CmJCVN6Ypi8G0jvOmyd+JG/kQ6l1v2hHd8aZzOlbRHWql0U0Eafce7nXec8JJlRpTDuBrEb
wxPQzg7VQICpHIGndwuS6mTIaUWesZDOF0c6oJirpvMXIUjg08SiEftxJ27ZMP16QT0OGaVFc7cJ
x8c3AzLwqhxHCLy+vSKBdYtuWrppAvBDgEvD4Yw3+FFU4+QRiGGtpqncFvD5F65e1seAmpaKFqjm
OzivJgRjl9VcFFIeWTDrTREcz8sAEuyeXB5ovWajevxfd68R9doEqYtWFDlr5O4ncXUGvBW69Sbi
ANipmxn3ma0MBkPAx3YgI4b1axWlsC2e+LzN3OtZTbnW29iM1+wJqRfEWHbWduW19FOp8aFQ/LoR
DQwG6otDNiFbNd3W9B/O1vurQZ9pZqDLALUQTogWjaC7tjd9evwsqrQo3AHU9StRMgEfQ9mZUKH9
QbESLCSoOnHw18uiqH2Mm+wtOclTV6ICeHP757xO7PKh8PlUbngxZxjw5XmXLJIT8fKECzNW5X04
2PYSqdecKrZvsjacOdfZMeETBTDUm0qI1SROHY2lwHeScf60xh+RgvXwzsZmssjZY8K+5hAosGzP
uYpuJ/F9c95OeUE1kD/kugYO2Dk/YKGBKW21F05gsbcOjMfiWNejrmSzQMMYt854yRLPG42dTy4H
n7v74z1A+fu5sTlWbenTZfuylFiDPzaAcTcN+gVuAYCjtlT/0gTbjVXj/9sq5saWv9yYhyiEUlxD
vaFKpe9zuEfHtFUKNcBNMQDb5OmiF+7NqA4a0Eo2J7Qgbu0WcTfzQoOsU57GM6Y+is+HxwgLNNPC
iURPOCl7ZjMVYW3+EDA4g+YdlJtH0EnRSrSNqegVEecnUszK0Ww9/en+GKn0XcUDdwtULIlOTtsK
jIbF2nK3s2knueCEcV93Y4slu1nz8lcMXzDFWTeV8v49Du4z/DtykiTG532ecD6KkTGOLNx89t79
lW/DNIq6XK3Nz6WbmGNogmOhFCDPGdcPe5swh9rFDHYIvR44opcRzAUN0MXrnuViaaiDfYXZkxtK
/5jIsHIk/Ms+J04hHRvfKzPYfkG3godCMZ2d/z9uariRyJUYXZJ+IDHtQXFdGLbXzwmJS8V6Chyr
ha2c4p6mj+AaYUXgOJ2VatI3aX5Rzq94g7R9td+lkjcDaGZBCLLgFhaWMK6HZgpgWT/P+JzEcuPS
XeSglm9yD/2uALkdG3iao69TRQkYBlgLZhmvUuyqHCo43+BtILIGSJzqKmRBlx11/rcKyaPuhFUu
hrfH+/6n5lwGM4qXiWtHyzfAAkOGLZyyYqqMbwjmRBpAOejFAO/x97ze9vgNk/vajNtbUXtaWkW+
8RxDXPyZZr2M0C2SWxSHu6zQo6aF8R1qkasOfKJ/5PbSVdCg8d2wc8/TaaZKWILPhpgNojFhQD9K
SIDurODKICDYXTywuPwWbONzv/7Fg06eJG5xB1py8FirvRqSzOPgwk93BG2E1i01hwNwtZTFjCu3
aqPavDLe+KQ9WEq6TZEw+P3CWc+ymi7ISSNxGg05XQV3igYE/craIKRrVf6vVb3KBy3LatCSCwix
4uCOngNzeyEW74efW1Adl+NKhFMi//1D2WEsDBbBAwdWrQoCnmXkX12Tui3Qr7ak8jv6lR5leivC
vmwimmVKVB+HCmiC762+ycZBBnZFuz1PudYKubfkYJEN+NCbhWek8ba5G0/oNa0SzUgGnPdtSLzt
lLkatjVpjC6c8uS3HQamglqdXXwY2Ot+GKp759QxUMOrEW+mwDCcgTWsbN8mFV/+aiXiFU8gRxzT
YD9M8J4msjnnWUddxuRmWk9VdETRS8L5wtEPH7gC0Shj87jGW2r1PSay6gA5qM1I87imnDazSqpb
i7Qlz2h8qW+ksysJ4bYK04ZBAIPsjsF9dxbOZmhaY3WRo5zyzEhPY+3spCIapCl2ENf6VGP8hxuL
MDg5n5Q1ih+C0QaPPPS29iM42UexnzvgVLqP4GC5xkFwPychjVvNL69BIj3MMbQluIOUDx3IMUhW
X58grJg7FjeYyJabcqjWOZnJd2opJf2ZpKly66mw9BZn4fzqRElpR00z71pXI9vyFT+uhc5kG0e9
mKcRdTzXCjA6T7odk09sWKWZMJumtl7Fqp2GsrW76ztIo2KZttmfwLgcsPl1RJmFGn1DxfkbbkZD
Q3ImiYhUjomdhPvOctxdHpoMQYVKc0Ppx1/KMvLNqlQAM2MGDnLINb3OYl1kgcLkiGw+i6R34IPm
zdXmOz88DIou6p6dBmewmjlJcsweJKDT4k0HWxQHBsWnMZL65Yv5bWzOa64hTWvKYIK6HwJKyexp
piZkRgKDQgca3/8nv0NF79GBXjujMdAnwAGD2hjZIUCD3st+/b8oJ4PRw0yJ5ptq51V7b9NUPbxZ
BP2FdVlquWhR3OOLhR8cOgQUpLF0Ip/rKYGFdHPCFoooBMHUU5haX0hyZkIOr099b3UtO1yq7EIW
TzMxBaD6yDJKO9UZK8yN2zkgLH98oj9LD4FdqEA/ZS46DWQNMpv9/509RH15D+pP71+QR0vW09b7
F3/qTuprAB3o+K/RmA5Tlr2hGv8SSiRyIy6yALwiI2fF3ZbSSer0ExwCfeQ8RE9Da8y78xfGL1gw
Yfdz7loA2WYBhbpltCMF46+BNB9tdl1vwGaIunzKCrqO2HC6tVJQfdkx9SKlELyVyoZsfwkNR5zl
sBajnQ60JI4zkmv8nckTjqzueg2nGj1hvFooJ3fJMvDFWA4ZlCmPVVt2M8CFXsmyqSqWhhTmybVU
2jkZ6wRLnrdzNty6/VPEandMMKjCGIwqrawaYCdDMvWLFDhNxQCw5R9nfPBc/yrIlLTUlr/wLkrH
MmsthCGuYKmQEdPPzB4HDtSbkoX0yKTTZZWHBE89ejCD98irRTSgUROACyzE6VZj3jCtN5DqT5oU
GwDrCLmK3TMPWjKIFFCXTQJh6/ukkh3kGXFFKI73peb34u8oScdOvx/lrcXoekNHuLWOi7ZSivxU
fjv/VRK/CQInTwtHvAm+GTDANmyQVn4NN0Hhihdzp6azrTfV05hpaGpstRwvimRGbjf8KIXs3qUc
aPExktSlR5W9kwktcGaV2m6eThWyTrbCf8L04MmYqxPxm4zLOPwPawNr336/fH6RIhbljoFBDAY+
9es8D8cNEKMQYWrwjdOsoqh4WSm17KRy+KlpMDi1Q9Gh20+lgfKYg3yqzQak/ZmGXBiOkD03KUUx
YN78wkJLgha2IAKHrHgUBFtE9hVuJwuk3Hks4AYIHiWirTzdHoMOJUmHPunfzJZHcVmJLRRRmHOE
BDXI4lpAH43QSjQyk+8bmsLyw2SehYthk0yPkYVus1qSJgYm2d7XBhX5AKac5MZChTRSBSUPYAk3
cT8dFyCNqFeheF5fz+GbeozclS/+ddcByENDtxw+1JIrPgawg4IoxhKJv/sNjMzQHk3bmTehR/5w
YfwbpdMhai0m5bx2RuObyrrMrjcV9xEshgsk3jBuDA3pfRwLYnP+lQ/nZEWl8UuU7Ue6kx7m2xJE
szo4+2oWEzh+ZFqWuo3h3nF5CpsW7hN4FxHkRns9YEuFfGbtH45I5R/P1G7XMAqFg21BZHkyqzeE
94SKpyAKqU7E1MZdvfOQBsoyCcZHWfUYdiesHQJRww/rIW4rS6CX7wn0JeeTNU7Vy0WA6zyTAeq4
L4Nn4BU1DI+XMIUUwKJ2ddkFstxfZPAiK7LvmgVCha5z6ljcrqDjICU9Ml6IN0upiaUV7Q79NJ55
syYJ6K0pje9Rxfo593PFO/ldfKulg+ZXDXk1dMKzRLfLcMlakPZjLQYRdLiBDdkoD3iAB4ClqSZv
WjBKhAhIFvglIRBZ4q4tC8gLV1pT8cK3hr0wv2bbOsWvZmCJM65QxfGLJB/Ak2W85OEgl5n7REXl
i5LfyYSPfNe1MA9gSdTX+N3ELpVfbbsTGDDk1eer1cuRBMRvjxg/aYfxuDwQPZiK6ZIHbe+BBpeB
uc8pa3u4BFW9z9esK72/ADQ9gvHQ2JbPFKyMHnXWq/AaaUFMd7p9BNyc4SWy8vfrD14py8v4Uc9W
Li8LT/wk8qy7SdlG+/VCXowSRKzqDjuf3TuwY/8Txm5/tHYjUbx0cYlZ4FNLbSD3QK2T04+lm8xB
slOGAuRLG3ubuTmj8EdbafknIAn3AB3Pa1rHyztsaEGJGYeu3EiQFdgyHlc3z6SK+wuDJQRXcd+b
L7RRSKoJ9GwSYue9u78oLuRBlQ12nkpr5Wg6LPDP55gA/ygyXZHAkDTaXLkAIDncjGiZ+MUhTZuA
USH09Be3P0aIbsxffXY81AogN6nhc897iog+G2Gcp+CVbo2ChlQfJjkbU8khP5YPFPT/0xRyOESz
om8pAIOvUzdzTKt2zbgsSyjC3qQ/TAV6riqYnHoJplC0obu5rNVhB/cli3fOuUFrymWhKl2jvZ+t
bTspV0gX4iYXs69NjyB3sTQA/QoTfk5AIm92WnAJNcwoh8wmjmrS5nN6VSkN8c3+tYVgVimtD4Ka
UmIUBww2Q7ZsXdNFR6pjGnqQox9wuD6oXyvRWidmRELVruR6672BojMusWoXiak59wA8gdjo+yIW
NHAAOzbod1WnQmJAr6kHG0ibSABD7eSzX+M8mP3bI34kkRD/DvOpnOjBT0G67b/C6w5omXq1mdo/
jn6bS+GF7Zw4lHO0SAR628KMqBAED6q7Xtv7omw/yta5XtoQPKS0fiYeRj7kIX9fpeLc+ZqdLdnb
zl8Aec1B23LTlz/occdGLdMQalWdqUz1yIblYmCkwgP5oJmDUl+uV2JDkOt6AhI/n9+uVA4AwzPH
cZAo6fD11/Fg9bJpi1i0NL1j0D1e6g28cJHGFHqLPkOCMGbgH4sT8pkMRNCTuidab2Cr9/VsJLJ+
ZxpgsHQKFY/eCKtCMtLhfGF929J6m0XC3Et5AiIltXsfnyZGo2OUwf7H3zUCQ/0Ne1sprP4ACMff
ffjMBt7SFGuvl3wncFJQmniM/a93kOvO5+md0y9V2CpEIcuKzIKPJ8W88VVLF0Ak7wjDid0Id5xw
VkM78iI3Ornrk6kyGltH0ZJtRwNUxuB+GsnP7D/3IQaZh4G+1xZ/wijV2QkDCiQ7OhxgLI/Vsir2
/Nzxt0tdAftxlpyt03U7mtPdZc2+ytA+/y/bphxNpDU54VlM8cMxSD2k5ai8bONbvX/SRuXr4n4z
dJi2T+b3t4CVx/raVeZbAwk7Yy9Ix7KfAgKYPL8KVhuiLriIU553WKdUGuhWAX02uVvEyf9qm/gu
IBGxEOkafR3BmPZdjHmnYltkgOBUxUiCB8P28FyREoOlqxtMSpzP71oGYiCO2RmRBZTbBDzEBreH
CETb9OtZ0LCKVx6aO8H1XZBcOencaHj8shGD97B0amFUvIrN0/d8fnFQq9ULDOHbXvmGMuCG5QQ+
pxLxOagTcBtkNyybfj7cKLtOFJ3q1MywB6FBt1BP2f4BHwzF6g6Z/RHWrzTc68KQB6ZpHBRy2FLD
jQ+YRRK5CAdD+cTj7VGCm1gqxj9dIvvoctk0p44k8n0pIZsMT9ja65On+ygk/ooyNRR4KZCuTpG1
mG+N39n4jdTq8jPVbsrM5UhmfyDEUzCjgnb2BQ9Sc1O/VNimOlGPNByQ37qNQFH0s+JvG7qsKA53
d36SXKabZmoXv4zNmTzWnCKO47xFzpgYLPebuBuUD026AHeRLmji241cWXlM4uUb4N3wW8SZR7s4
DXF3yFtca28kr4jxMS16s7WC2BekQS8PvKaryFr9Jahb/QAXR4wVx6ZC+ROib3VpwzYu8AowGWcW
8ggFT10swo/MuJQ9dlFf5656cc5I0L3mOpqySeD1vL0+vI+Yz5FyHMIIR/DQABKbFGrZQBKEg//b
vo7CnryRqjJiuSh0CK26Wq7XPZxG2+8wKGqghrplGYOHy9p+8muf+pX4heqnzq+UilsDXoeLsg9p
58QH6Srts+RcrUyOJsI+01GYs8Rl/mtXxaLnCyS0skLol1sm2furVNmfhb8u3pjpcyG4j4xK3ubN
yDk/1Crp1y+duCBh2AOKxqO0ZJzGsLfZjXV2cAhAYfW63wOVHSLfhSoYpwxCPeeeocSlZVSqTMnJ
WYpjC99qF8K/TYvn9Tfu+wKGyMXPotFtGjg+lP7MeUASgb5FwSSDSGXVI3Ug+3bkkd077dc6KKKU
a3hk8RUnT4XCQNRvMRvqA19YoaK50b2n/oun9M9z70jU+Ax7ccUG7otf0u+qepFMdyyFnP2hROeV
7lkQ0PGh7NIKKD3bX1nXM4f5q7EQfTSnAoSq8TiBkNyNd03nTWmnhKR8Uvr+GGGEGzzXUxL4Eswf
CtedRD8sqvPX/I0ixIO0ABAi+3MrMxq0ctuoSpKlphgF4+QcpUf6XeK9vh/b8boRx0oxnH9rDuue
NK1iO8Lmfsb0tVS9//NX8Xxf4skcyZt/0oJHAq7468W6Qhx6DMa2cE5n9KYJl7UPditfGwv9A0Oh
8PEiNjKvY3cL6CnspnnFAghf3WRKJT6rRoKHlKDY5mYp/sTXIl7n7dPNI4vLXjZIuzn42Q1IhEto
4EI+2rsHnO4UZ4F/MnjvE04HBwwi5SRHvfQp7m/z+AUkZb0K7ItfEjZxHW+J8IR3qr0JLDvE9m5n
t1adLEtp2RHG73CkQ+bTNXF16chyjibfTDhc0XYuO6rKigznrw/p6Cukh1AHQRZKYLPaVzHS4CRb
AyLrWPJQCmxDjyOWgpyfd/paq6+76Hlu4LboHe3uc8Y1opYFjYFPrq8zfEtQhK9nuURbig6srHVi
zRJPkKs9nb1IOGo3x6J7aexMQIxI7a7k2DhAM/sfjXInhiPUvEZ/LTxXcmx55v9QKNx8RAzfH474
X95AI3xxupHHAcH2D0e4XGJxguNCGzGa8YKZHodBGa9JVtuUCQ80+o4WSwBxxfaZR/dwwvFxnmI2
Wvq2jzvHwZwxIrig8VPZZ9/nLtVtRmBh3rTXPwiEtWUmYLMHTeIKFmO4eDuzVrZZ/Lbz6u5wmrEY
iMYFSWv2q8LNaFJlqc8Nz68IHHGrirXA2bzr7RfwVoiby98bQUIpRh51DcKsU06RobL4fM93/jHM
ePpaS3q6zn54Lsmnpkg8siPzl7NOmpWlX45Zs0lWsbdxDKS1yBFZ9s/pMeI9sW24IAL4mYFt7xYK
NubU4ZXLO+1PK2PVgIv6iht/dSWWsuk+EL/gsxUIiUCJmUPoq9fkW+nfvUiYkcmNVYfT+bAZ9KnI
d9jsMXb7TGc9xxocpbWg5CEG4C5jV50caf6I697NKIoSdnwVBiXeCDDN+zVzvQcYLMmHU7NDd4SB
gHZsbCfmyAp2doLWsA3uyDkQHPVX+e78X9bKqq4WpNIMEoL6htVUv33giwfh+k68PfqI8cmef/7y
6GEdXWstJQFpIdPSM+f/dvtt6ZgyRVNJpM3X/KWoq0+wzRuWSydNeV9CQgQb8/dM8egNxcpH2mch
KGsP7i+wXpPoE2YYAzRf0H+KV1DdMBO5+Be6ASYFEMkuO+bqi4CYJ9KMJ4EDNjfjMbGLjM/dwrD6
OAQC9jWbwFtJJxVSjLlNhMalUjEnp8saMLvWdPq8yeCef0+Tcb2JqrFjX27SNX8B11hNJoN23UPb
xj3a64DCizB9J0TWDNju48b8rMadzvJfNXaDnrpxwPmA5eKJlg8KY7UB7V8go3D2j4wTjFrQfg0W
DJJTNucB307C+st4NWsJuQnfEkEQrQ+EUxWFFJgoN33cTv8kNpFjJDOIYIFgJMvUnU8FICHnMYvL
3KrbNQMySSN717goi4lPBkTAuRucxgZ4Rc4/lstAHCweJyKWeV/sp8Hpw2u7A+1F1irdsIH2gCtp
+hDiM1MYKyfbBKWi9Km5M1jzwOrEK8iOEKFQHgTHtCN/NedQR/WibyHLb6mZXWmZhA/a9ap52LO5
xiN6w7YMF1/n2zMLgztDjyZC9qS9bd6zWCcXttRsm8Eq5lHWeckx+S8nXmBexDLbNgLxpLpVbXRP
exkoEBk0xsaOrk3AXH13SAmn2GDNrpu0qXXXAjicmf7A5NwHSlYWC6W2WHfPWCcbJJ6HUpPvOWeW
PUQVFnzkwgX4drL8po/yVI8kP93E43frsDVo5ZjkWqHixRhfAofydyDuzgaoskp14Q/hUm1XVEDg
V6NgKGcyv1KAenfzTGb6Y1NEzYGiSc9gON06tvfwUppHmLkRtxjWuEyxrw/CPKJCfsY9aDbBamhd
XvKoGa5rRJoL+0tNz3JjngvV2ViK+KNj+b5nbyE8yylNRgRM3SJjW6PV9D5Jp9xzEpik+2wqBMMt
CQ+OxxilbC0D9nL6ahcRgCQIM7vBwKRpVRG+wjzuQaG/3fCV5/1gWafezjKgo2L7VV3lH7J6qPgB
pY5hvKWblJqgASkYZIWRQwHcqB3hLC4H/PkgvqnMlN1ZBW9nsjxa2srdgPpXHLRKHpfcKlJoN4fC
8ScXQ9dpGi7rAZw7bmzSQUHimTTQN0O3s1mtZqv3ZJnFmJGKFgAeiEoU+o4JwR5wxa5+naloHLsA
JvtBDjvwwFiqq+IUeKmCDqjhU1MVybbHX4z6u/xPZLwJgd0WF0FN+B5JmvH9L+JYaB/FJpExfMjb
rGjAgtdwkyae46h2dxyDTfUNtUwuD2tKVMJDC8+SyYdnoGdef5vnFsWLIuImdOfkS2QePyxbZ9Jh
1A9358OOlkLTz0o71qESNdadLBgz+1g5oC1jbYK1IPuQkRRCkBamqGLJXmSHMF+dhVdSHT7UE73c
T6SJtrXIOBB2zM//hwaTex4YbFGQL00rJ336BlKV273SzB3XyAiy1fDpMYzYKh0iBLCYNGH9bhv8
AWRgXMk9AuBuoCc/Aq5A3bvZ8QB4qNxJj83W4MfqcxnOvtvbxqY4a6zELkEla0hMCqWTgY5DkQpT
18+O5IsOm3LX2cPzegowj1SbfNwt6k0/yBSgynsZyMkFCR0aeFyaA15bNi7c+xm5K6KM0s+5iP+q
s9JWIvmHvnFRbs0/gN+wJiM9EIzOoxjPJNc8QQI9hYUcpRZrm0TZTy3DFmQZQ0Qpg9XgBUyr+bFL
ljGfnUM+aUF9XERU433zCbFTqVKzPQsWiBnXanbH3Ek4cW1DDjpEqGOPcnWrt5bKsMmkSgJKrpTj
0aOvO7RIaWstpfc2IlV7cfWOesX14j6vvhMS9OotXwb97GAtiBhs2BFbVeWEcbFvCueyAS6Xg14G
I1cCjQDpEeihFoB2PLGOBeNTtPRPl0O3ogH8ULKrJ6OES/bYD5YWtoixQ3GkIpn4/0FCB3Ko0Ady
bTAFlDZqj0OgbCaV6kmMewj57gYbCs5tW4obnNQW6/VgaNNelHlDumEtyaQNwZfaIKeaPY2bYsn5
2MDxruM3CTdBH7cCz5h6K0sz3JwklAZ7TFTATjg1fTlahVuXglT9MZcgbaEqXagnly+OE0UDPxQ3
yXP4QqSVI1amLvmgWNaDHqpskB8BnoEUwO2YfSuZrvyS8IVSbHNWK9qmnVxW2v+0gP9szxJ66zQB
QEYM88qq2FmbLi5wZHSe38G2MXaQmM0g7VX0PNaCd9zsKs0rTWs/j1qnskcBele1oS34hI4IVTog
LJs6CXcm7KvNTbDeHR0fO01jVZ5cRslrX/WHdVH2f44m38cMlMfz8FfvgfSkGWuFhA+okIEKuXrM
T65RPK9gQU3eID2rDfro2japlueEjOhEko5UxMuslZm5JhL68LH7QbFsiY+7heekGKqRL3iFN8MG
fBBPIIm+FFs1f7MS5zezetikO88MKVNWEpKC1Uiyq8IRwGV9OPaCIoTaRhMRBzAtQIMGVG0yF4KR
c8bfB+KF+9aeRVcihLCJt1Vu4++JpDtLtyRFTSjEd+5Nrjyg4PGpN+bAxzSttfX5jBhGLgJoKdhd
5M2yk0R2k46FSDHpPsaRMYZwj+QOyV4rpN2xM1ZR1wIjSJsARHbQuwgAIGyp7Yu3iJilNzat7rsl
mXFQgLvvKjRgWGkIaDGPRvRIrO3/BEbzjmTEJFnQ6F6bCk7gKFo9vmqJP8mrB2zJVJJyFymv+2K+
Lqf0CUXosiGjCubPNa+fufE5+do3z5yRqBXsogRSvGSaVtjXe39//p6mQp5TYhFMRKN0swX81Cer
cXRlPh317vnASHKHIkneC5TWDX3FtIV6t2idi2GNo87FoEQXXloyumtLC096wOY4NXGyq8SNN/S6
VD7C0qny226awT4RbdTQhOZSd86Xb5RDCY9G4kOE+KVLS4iKZhEHsUjJep/swKa0eNz0G8byfUks
7G81OlXZiNkrSivu0vZYiSaYag3TeAijZCM4jZmnpTnzYnDg/6A45jq8iM79cN7qsB3M0lqdv3AB
YPu1TnXtpjhobde/naeHSXpgEfA1LAuK7QBZCJ7mfw4H4SUKHzYkPxKZfw7bXpPCSl0cqef2KaxQ
PQY/MJBjOfHFCS2pgG8PlTkVOFgBwQpo9X6HMszGmcgRw6hVFYsZGxOm4lJc4Zh85+gKYNrbSACD
QPxZz7IeYfC6HpbGR7bB1AN+EC2E5YCLPyKLKb+LQ8UsWcRYrUmtNcFbbq3DAD/XjXVnEZJ+Dfnw
1W/JbZzSSTxNYShlPftPUkINeF/sw77Br4nDPBmn8RuVHO8AESOrT+p62zH/9+pYiEiOP68rtWxV
zDzqHGjG0aXHyk465CixEHwISynO5T+HYnu+tuU5GiusXRi0EN3EBjRmXJHQMfYphqfVh4UeI4Ws
ofVaryv0MuH+f8J7NSzQ4LpwLqmMDnNfvw1II/xmJh0gq+hp08PeD7T8jaAPTQmp6j35BswL7lhC
dQMAtlIBOy44MDokpR3ut5EDympMAGRF0dNKA5rFVB2SqYzfstsLc1JWdfBubX6XIWq2mKvRpH0v
XOjo/XwtvNZL9z2RA+LRK+K2l+zpXsHXapbRnmQL68vauJeaE7lsImEqqdMTduVNRAyxXj3bfnH5
wb3hGWUzqIqFS/urEBUph8VVna2OmMHSskHV2TliynisxlwhwpBj0VUcnjZ3RwEZL8s2+CYebk6j
UZlrPmKsvv7kZntMtXBlhS7T0b/BFdDXzYW6KyPeiZZEtGkR356iJMyHfltQiOnNBznqiDHuRx/s
4B6cY/4Rtboy1rIzOf+kDMkrGKNlxNQw76S481OmI5pI8Z6bLVcKm4+Tapy9eYYJwg1wgNJ4nNNT
0N5wG18yJUBDdHmvvm8+csfPAVZZPv76Ga/0ymKmfoQSvw2vZ10nhGU54FG9R1qsbXojasNDX87g
TitPG/p/Qmyeq5dX+2AXVYAfQxr9nZF7nDkW8UiR0acTBfLo//SuKUWsOU0p5ET739dJvMF+pmls
6G00EkRcDmYQAdbae4OmsqYJpb/HN8Um9v4ky1/K+YAGiLi+O/YZm80okiEsnwzbc1wcGHBYVsbT
zvKiAyMYfr25q/LCn3J/ifPqNfauyODWFhuEAjoqRPwMJToGAJ4E5wmDesGLzuKakOsUGN3RfJ1B
UzNUpUJhwNxF0msG4/jzeQBKTtFN1Y6zp41GyOseujNU2gNjIx2cWFRiL24qNphuUDny3zit7KwO
Jl4UY+d2OLcFi1ePdKbi4JPHyOOQf2QYqYnLq8fVOMgcwig3HQcGJmgTbI0hQsaUemZ4rynD77e4
aRFztdayvq+AnRLNTjqhp+OER2MJdDjH77Dh+Cj7yG2VHgbBy7jriy9/lsukTuNMC89QWhuQZSTh
ZpGBIP9cID1y/Vq6Q0n2mQSNQfnvL/tFOz3bA2Zw9EqGOR0CQPDwyXXX4gOnBOtdvlL/DZ9ORZH6
eUMx+I3j8+7hjjYwzKNwBppA62MhjVMFs8Jk6g8M9Qahw3aBaYCTn38HUk8v+yQ+XsepSLXlQMbH
9gfVntoeAS5m2m92K8eaUD04FcWW75s5aAGAUeZuM+AcLCtWLVQ0g1aERBJkF/ghGfKuJxRmAgjE
2UJ0TNRUp+HNxUR9TzaEvDxNL9QsojnWOpt3jJftEs3WyBph+n7sDgVoOzbAy1aLpiEQoaqoNXQO
b/sdD34GkURWp6yxaEy/B2RRK2QrK66FZAwLL1BgVx1kaGpMNFwxTnyc7qC6LnSGJSKZEqmdzEgU
0ag+V3adcHzJIe5snxcruV1SgOt6oxf2gwkg4RyWNIWQ3XbCA2CuEC73U/VnPk9NGocU/GkFss5w
N7qJsXh9sR7t1AKnfVYYM0owkGDX6Dj+yXbPa1m3eAg/ohuywqMOOE8ZkmSY7LmMLe9UIlKnsgwf
brmhjYUfOPql+FXWteF1zPi5lws7ujgM31jsaS3ObF/+mDjtmOHAe7KTE6ocJkhdOZZgp/edtHqg
2M0Eux1BGTQhPcuuXk9otiT8NL70qz5je6WYtqBGaqYCfjX9SzOLr0Pj7nWFnNgvZFNsdLYCqhjj
gyc7l+4laXqtpvBG86pkuBTEM/UO3OYx1xWmUnY4KsMDXxGr3SmzuYmCjcSbz/+OVJmoDUolM2Jh
WFMXTL1onPjqQcnZX4+YX0Lp8nfwY5K2gseLF1S7QdrHCAzu45UCHry/ChF3w8tSpeNFDZoorMUk
fvXGdq2AOWmGBl9sHtfu/4FsVaVh/huB00ZxLSJY+IcdUDlLoiGjWkqsmhaJLmHZ/0xQ+HEUJETL
xVpKmkkQchYN+UhMjDWsE3R6+YRB+XpOMwK3d+81AyHX/Rr6Q+ikzvym5S4BPxIKOwzce+tCAGJv
ylLSWRysuIbHX8jE4wUwokC3wtpzvpxlCEvRW4cnGRY4f9ZF381NMn8WTnpihAwQhyh8Wd4Hm4fa
RMFy7DUVxu1I/+bynLkQu4HnWD+4hwYMPSDk+c+gHsFa5TaRbEKVKOr1CHRlh+ydGZhELxtIIS9O
Ur5QlZGGBIzq1dpt6GnXN3z4D2Gz1mAREO1zPcIT7EFJnxVSUoLyrxhHivfM9hR6Pt9QOA+ZjqyL
/775jXwDlRF9Bb94gpVUtwa/YiPl38NaH8PI5JMnqkOhQEHq1Mrr9cFqxhzJeXCFHjQhkJHGUUv8
nUgGlWSiuP/kcZFZ4lxtwYEPn/WQIFgIX8kJ0XtSf8bloRkUjeo8VkWi59fOuvE8SS9M2BQmZ1wY
TQ5liXIfSIdsYYTIiJZY8CDeUFGQh6n+8zbwquoVKSl3A86SBg1AMp8BIZf5I3gOAI1J+BK55E9y
ilAM1kMbjsiktZwjbRMrhNpwCkjQpLqteGXaqqdCU2B5OxTFotVOiIE8zs6MnKVTL8x1vgwKOLlR
m+VhkV63cYXyw9CQEVWSQuJ+jjdX8p5DDn12I4Bap4RTujfZczv6FFFn+Q6DMqIbB20VFmtZvVFv
BlwDAncGZlBm6sPNJ70QPOAj+qyoGuxik2LzBKDE5sZwZ0gvYsdQNDfEGAApf2xZiG14+wWIsWKJ
SoNZtctDhyB78m3tyyVWaIekUBWbI6hwmlcB4Wg2ZHWh2y68i/jWJP5+YedUdEJnSn/gnmOgqV9E
vcRdw25xmm/Q8PoUb5eOjTZsPtsZqx1B17xNmgz/GEOdOv+1fD8eQiTUUoJi8z5+sQteFVhof1UZ
ohR+EwyV3TsAYf/T/oVEo5RZKTR6eyesyIyjEJryTx1aHIXpR3+KpfD10Ir7hjEYuFzNH3XUsuxn
z6iEwA58XMFg2kS4WnKaQXSymJbs++SR4UtJ+1UPBc6mKfNdgzSgVnTJdYdIeAHilMd/oj6mkcq8
hjsMUN1xNRBUN/S0FqKhSot/aI5D1mgT+9NLM/RN814lNmE20A6yYI/U3eThtSgwVAmwsfJzV5ll
NURnGTyycyfEhgps+dEX5Bm48XVwEsZjUMKwuGD8SWOStgYb2MK3Z97rNUT4X2rqVUkW9aKtycLC
PJDQm2ewfl/AJTxpgivOAuW4OxkBvJjuErcEzEmXYPpaP007CF8DTBpB2yDpcUZEuxtlaN9Yj5nx
3w7OC/HhTXpxzcNqNGRtQ4pSEyMcL/40uhr0rV6YR5PEH6EfVUebPb8eg51Qbj19KzutzyMnK6Vs
djyoUxsYUC5xXi+2amxTocXvdnb6xizS4zAIG1sI/IPRFL3RvhK8kKoijoOTm7X0jkCBrRcJAMiU
1sruJ9mgpyWQ3hVF7hKh7MpstnzvVLr0GROzmPVqbvP0SrKyn9Kn6Ru9/NgfwYJvFEYPYlJeOaDb
HYLDBaTKTsN5og9CPNuTJWvbXXMeXgLz48HC/99KBQQdsJkeAmwuedT/k3P+HZxdzKpWR4SCtzzA
mRGTybyaAsRbRygqZJIY9vQE2aAI0xlHE7ptosLljeIwul5YJq96MGi3+M5292rObsuI9P64ko/c
eCN8yjMpeDnCuvYq6MUQkDZB7YQGZR1aU07rgj0dxByHA7AQeXgJ5X7YNQUYSYb4veI+voYJIt8l
SVN8uC/6ryiK9BI6VrIbFNhMjT9T6yhevgBSCiSwOidXboqHSrMN0fN84U6GszWIuu4V1qFFZ++u
P0g87bxWTVSJpPnJDKwRcE2Dirgs3ysViYf/SKoginHTQCNr0lXk5whGMg987WwcpdrC5PUjCuPp
K80Jr/DEt62HjFZMADO+shul+9XrA8njKPVblJYqAEZ1GdZV6Re02kbcrXI+olghKyAh22qSFCL4
XvNQIEZyRrs4r7nvFw+aXAv9e4XCscYMEkwOh5w5bewr2Qns2hYYxMzpbnZTCTb43D4S//XIkqzw
PvYER3DTLFcOO5i6yjaRi7/xsuVbd+1KBlUug4a65k/ZToWrAtV4Hjz83jaikGkU/cWKIL3OwuZc
ePGhOsgwdj5D7B5E20Vaqhl4UixRkVb+3vzaiiSQ8j7jn9cuqBMYrUiBAx/sTaK3gO1PxThRnX9t
1VINGZJ04z0katgeN9RhssvnWXNOY+QG9CFSiIq7soN+CQr+5hQN8DmD3JSzanDAA1JAsIovsvQc
AyuPF1aBDlWuHEflRqBfB9NtiSUlvnVyWYU282WSTWnA9a5RjsrpK151ZNeh81Jrxuuhq20ZlifJ
uPcZ0xD794NLG++2GBR6912jcq5IMDYbCxzNdN3KXfG9H8JgaKCW7JKk84P6z6YZwgx9vhYckU4L
goxi4aHFrnG0TJi+F9oOu5SKcl3pcVWXk+ib6NDLpRNOTI3W7Iktkqslsxud3B8qReNBrgB4aaVF
BbmDTDwT2IicPnZxEysyydCNgBofEXdU0hEVtjkk4UiUKa4/8itVGAnwp6H8LxZJNtzvLNQstYmF
VCW6+NBSeAvFG6rrf+Wk01pGkvagQ0N95AwmU9naE7j4zbknLlnL3t8VpLJf8EzA+7i1Z2wcHELK
WxtNbfhqjIJCVhDm9d4k4DV9T66efmTvJMT3VkbryC00dbNv1ZakVXAQA7jGqI9qFG20UWqlIZov
V+DN7oDfqH4Gc20DnHwI05a27kQSX9aMaqNgu3/F9IZRRTA4wAZy5T2hEeFbanxZxel8HNhNVDLw
SFI1OE70E0pR2W7rfaReVGRfVeXrcWSccA9YvdMHymD6feChxgXYsr13bx68S7UBMkcmrGFm/sdv
WZUKL5i1subizJLSyOA+75hSS++uMqmCuCWGlg00Jg83kfp7UJyi6InkoNriCo69dMm5RXAyjcpW
BkVYFNt5C8AzvqOHddM/KEtTvTS7c91k7C9lhCvSVl5NMa8UMoB4YoiwNsZ4LIHQ4fdFRjUj92lD
6l4a1k1BKtBP51h9X3iYKZ9io6qvNBCqotLhkjpd/oGZoCwZ8ShuNYFiuscT1s6XAB6F8GOkTBdq
tuZ4N6CjrPlhWsm6/BKYPgRwVacYeVPtQlX7NMoroAMdgO1xD3No/2GiNZrJePiHUdm9r8gmgXBO
8nZgyyLqkg7OPrpUIAPbi72CQyzfPt25ROjo3030OjySjijXyK1dNarTfObK17fLDTmPhyybxvV4
MeQYKcMFSa55Pbvve1EkCMcK75tWelh+XL9fBBe8DHPOjKyJ1iKe5AU927ghnNDYfA+395vHaHbi
NomlHVgWg+5vcEFgMkJiqkEgPeSh+BgYLJxk8Swu5xSMrc8fUi8GfGsrTBLOYEW2JAWnyrrFwbae
xd8xAIjnNOQxeW8AZBO5m42gyRWz/z5vKRn8LTqsiUg9Uy46JP4gwS4ZdNh+nJm7o9s87Dpfuca6
yR86soHVPG5IdHXZonpCoc+B8ilkiirC7qxmt0XJeFyMvr2OVYBDo1erVlXf4261nHFOgSytt4+N
u50gm5qs7HjLc+fFgs91nOi3i3Fkb+sDFmqwGcGoaRX4bDQq+dBtCQr+gQ2r4XdfeNzo8Y5XR5uc
Iwqugxey8BTBU9KCvD49M9cT7RiTkf32uh0km1FoEQ8hjl0yOpMPQcQRZideXbX2QZzCRPCD7kt8
L2qopxo7zy2b2UUu9ACLw6o7sn+4GQ5k4VuzHK3EOIWjQBLW/LlSgiezdssHpM1yzpYc7VQBHSyp
hIatsMs1GEvuiVbZFjAdqAY/F9x9ep/oWcLxoKKHXdaSGm5rFygSfifVGKAecit57zyG+ma+2MMl
YTo6983iKWW0RFCdlTXsRONWCtxs3dMr/lFPwcy2vB5u7HP6g0q7ZpLooZ3hAvHzTomHb1r8ZK1v
PU6CL0YjKYYuxGQJ2gMvDw+HmrNmxkddNS3eQv7gin0k1E5m9CEMNmfl3me6+KeAzT23nGZxp4Bo
qt1HAQdNmMmVQe2o8npd25TuZRfFUb4NAwBHTp7MSgIH27Ey1KaF6QNOuWxAdqJf+s5CqTyHWWw6
UQqyX2w7rTIR0UjmWntpJLHujAhOKwVdQV0Ap4xRvzJuxVzfMKMJksbl4kRLicI86c4EsqryoBap
zidwQRhlTgIXmrD4DLya2pWv2B3i+dUJzo12wtByd5PYdaGeLdbfyHrHRMlZOIpD0H7vSe4QJu4M
HUb+yU0XTJ9XTfsQsM/TawLQ+pXfX7L7/F/1FmpoXMX1OXigFLRrzne7uZ1rKdac+89THc8j3Wgz
hQ6tkqFQIDauXlWLN2uMZiPsuPP+JHFu8rjvIYJu97oNALrSOOAy4pg4n/aLGpVSTmzJvpy+IiDy
10L66aRTU40gmaZMDkAizDXoh8Bqd9igmczKZ5sS8eXMZ1JWHM7YD2euQg/g5+4nULqdygLQoWBu
jVAenK1znTTNFDmFWZFiVn1VXgQWJgeKOaH6BsHSr1N39l1r61L9mw/onRjS20XhcFKZsHX8gCpb
ldxpFu/e4KngHhyoV1tMMB+xn2D+/FM8YguxKLgZnDAyO5N5cD+V20IXrFdYFGHJ3JR3jDVstPhI
CKIyEGsS2aoK/R46tRN+72Z8pMGIb2WW6QnLFgY5Y/jNQBvrwk+sKtlGfjkl0owgrmFbkgYnTZfo
B7uhmd+CIlL23ByOx5gICJOhm4kMknCc82g9SWizoJiLYUrydWOih/4e/IIozc/ilkkt9GXyaaun
yT0tdBjkYkHzYgmKLtvHchK+HGQ399iedStAmPFk1qoQG6+P4Rfw+nZ578aYjyilpZT7j7tyI4rm
g91sOqiWZcVKrfGASHv82BW8Og5kMNR+4yF9w4RjgFJ5t5lxKvwNIL+Z3osLTQrx+DCjUHO6zI7J
pZiMy+V+IfAwX/Ms6dWqLscdgWPZWTZLK73eiJIL20GKG65qp92XDamJlst8JF/9Oiwvg8ZZvKB0
4gv0uToJMNXTIo0yCOSvhM2vR3vBtCXWMimJ4kLHKG2bjSueOyWUi1MEqfmtYM1SNTUbcTMA0QAh
0fFCkEAMg2fE80SPgB+ZoFqxmy6ihSkuxemwUUoQc+LhVtQakU3eCb4T2l+hE8/Y0+JNg6S2QDK6
ICsyW+rPse2fC0mel/O+t3sHNR8QUYfoMc5diL8DR07s+bCuYVkTBnPxhvyBFTi6VYsT90bcTLSh
BEaCQDu+n8+7LHlixe5bPxlnAb0rw4p0N4m24ojX7Ze8GhSlgKDGO5c33zYAy4+nB3Hin/9Ms2Gx
gAiiD1twuz5gfEHgsrnq66ff5eqmSBHFcTrlFGWDRtifk7m0U5HUcQBp7eLGdNCiyZSkOdy5qMYj
n0D/UJK5+AhsM/e9MBS7QJZxFFSeoo3VXxwDudkujdVX8+WVc/9DMR4w3U6hXBLTuk/CN6k3RGJ4
6PIt+CtKLUbyfhoCXaFMyLizr53UOm4hxxshFSQ43qqoilzCH0rZL00qmYkmIwqcW7PSZcbIGs6o
nK+Wzw6X1kDo7usyjeSaCH6g6HkHKPdfty5BLX0aWlQqyjioqs9Lm/VS2SpaoNmEf44XmYjz5PAh
EuP/9dndX46CAHPjj6+U203ZJPRcFV7lqzeQt8ky2h3wi/dJo0hYCd1eREoZLc1pTPqqHhw4lYhU
e/W+biyQTnOGO8StF/iJGug6ZX5rdlzNOk7xtaPotYC++zNA52PhLTndA3vwTJUFG4RkJfFwB4Q7
RmpEueSsKJkoVaiJzteZUN8+bKMQXbei8XnoGrPP297aGHdGP3+BDbFjvKadp1RXBz0TwhU39FWq
xvwNg3uroX82lDmUywQnyxpJJGhB2Ps65kinqwULvsJtz5NnDZhzUhag24aEb6EGED7ULFo5rHfK
6RpiSvmOmehuZCxfcrVQG7P6RKwrMKdiAL2ZysmxHG8XlS94Jqkqw6iVCqdf2KrTGU2HSvGhWabf
MPtDXaV8EJyr95cOJ8lZmE7qopvLxfSu6IXF4nA7YhwVwxZ1ThqrxMzsJv9bxY+6j0k7Hx+bIAk2
LI11GCB2zwWTJlEGolitaI7aSDl5mxd28kEmtY91bgu3+JXFpULHTfwnLZdwayAq9MfbN6Xo58So
zogo6atFbTGiqh/PVU0xgAWAxab6y5J8/ZiJ+0yAzEBl8SCzdboLL78IFqKz5K/+ej20M8O1MaD3
TVhAxGQSdHTiHCQRfQVMgpJ/luY3bCXD2YpAvL0FEIqAuHJzvras+hk5VXiolfYPsrV/B36fJkOn
61ErSo+8kDipttQXW1pKsZYAMP9jL2B2JMeSIojoerMzpNuM59Ex9e43dr7WBqvC9Qil/sSo7jC6
4UWhaFY5y5qroIUKbwlb22LlkTAJUvXzXRRD9ddAI2Hm8PX+muYyeOD4ybQ+ZD8Zm3MAF9OAe+aN
03xlc+TnEXfsd5OfZlfq7HmyU+tgTKdDw4xR2pRGTNF7tKD/YQWM/agaxXl4f8xKkhCwzBQSxEm5
BDMsUPFFPURLK4r/QFaV+jf495q9rOJi5gr0C7b+QjtzcyV2QK4D6u6++C04LtkpjeuAU+OetQB8
svElOi311UUL1yI8k3/RN1IoiQ50gbSpyu0+8uxgzNnBIY5ndWec3bA3Bp37T7efOfE6za2GBTpt
fltIWtrbqGkvRbVlEyu6GqIjQSh+ht89Sbmz1E7ivUNdgV2m5H/J1CuuVCxP7wrc3H59VsmCtu4d
94ad1Y/33DQBQnvQk9sz5/kwLuwk2llR92KXb9fRvfpUwzEX7CDicIhmF8kgJ5QnXwKbSxXKcsDb
ev9aqchmN8LBMuc17nYGq+qqZ1Nq+V1CS/CK7OOkq4ivW6VLGeVS5yiamAdXiT5kiW1b3PIE3S0j
hrArTIviXIxxRNkGwrGsEjSVCs3vAnOgHRIJ86qtUotPoLJ7LGyzlWrv/6VIrkGsmVwNYGBXjt6P
TTTgUDCF39x5rjqMZn2DgAnyMvPJs7+PwamauFurotsgZizcAM2J4iCQ3rgt/2hi6L0+kkF5fb5j
zogXJuxXx1v75GjXFepwoGjH5yfIAioe7+hO8sbJEUVHs2s6VKNqzEygAfxSH8ucoyXI0hrVZ2Q7
xLEh6HMugcz+5zcHwkf6tS/uyKJTKY2FLm0jDr4Do+tHJQ8JcsVorZ6+SlBpXFPUunICkuJ84mnH
Tp7jWpA6GVQjg9oZCsVRAVwK+ansWDjvGWwUVlgMgxkBjjHJjf4k2BkwLjc7+qDIImQ0XR19VFEj
K46UFzhzE+58ECBkQbUYiFc+YIw7F3Q2XUrhgKKxAekWKlCaV595ot74ceccafGeMs0DdUYQJz0Q
iWhcQGTjUkXLA2MXbzJB41Qfhsk9935OmSHIEgQV8EBnbrXQMs0NC25PcwqX26cZtfH6CceHPwKy
N04cyFNIiYQlsdsZLqG981eVbr8UU6ol1mdmlDfsRfPxSqw0+EaPJRHktI7p8Vfy+/IEU0w6AVZh
QBsB4njuJZoQkfCEeDAvhTrRqEp86lzZvn9eT4LCKHpXVmk1ZKfR73qoUuW4wCe4I7HqAft0tq7e
s/HFqL+X8415so0hlPLLW5C8+QYF9qaTQJHeOAwMsomolJZNbij+lJ9jlWwLY+Fexkc57gIvUwfx
PAEFLyV9BSTWCtYk+TorQXJ/jnmicaxcBnZg7CFpOo06jcAgQBpyqevPUIjpl3XA35KW2LDKkUZG
S6kz2V6MtXwv0JS1rz8RuXIBQUs4a5ni0oib5qYLGjUuiZgraUrRN/4b5V0lBN0HwN1k6m716iu6
3qwhwIqh1Zp9QPa2qhZEK+50uEULSJVXesLO7I/aOjENGWmILYUMArwpzM+nwzzDIgE0ywkje62F
CHQXsj11kstUGbfWo+ClEKn6JMCJnc5MVHPLZ7/hQMiFT2bI0xrmXloE6iBiNAgUuuBFD6i0ik4E
R/pOv6+S7l/9A4UzXz5i8i2rAxvv0hI81ETaHAOIQBHxCSSKC7G5M4LTNcCkprsoCAY29353kzJ4
jenP8fYq4xiTFQwnAOu6MLMEr5+YQQ7ydIYdHwtebOaNes0g+g3dC1/V8vKehduT10+eKwVrXfBY
IQ5vxxmfIkrGsVxWHmXMf03NrVlUhTaTeHe4ggIsJbbcpIdVLJs0lafgZBJYIx3ImHN+tQJdA5uY
zVgI3UBm2t0DAQPkxqN5S6Q0Hvz7SERjTb4q6CLlD7cELqyFg0ndAEUtylgFEib4PQxOL82IKLxS
1ns/yPlblMrtx9n0X/YtNtastcNdQ5JK7HIKBcf/rHH9ZBMUCPh8t0pOEmbAjwSVSroyaW8nupR8
sY7wfCIJAP/wwA+OGzF8XVvWgEYMCMOh7K+PN/wwNQLQ2J5eDuEftbVcJA3GhX2i5Kusw6iiIOae
HLkWNEGboJZb+Ft/y5LTE/uV2o5rMgPBWLOcMKoMihSukis1V8uaHd5zZCNB2ju3Cq8lCtM/D+++
GCPaxziXsB4+k3IQ7H9ABJmqbB5U0XwqUg3Uhjw+EpzhNTSVQXiLsyHl1FG0IG9hp++of0z21wOT
Gu8nZCyfkkeDUVzbN06QbqVbRqCG4gboK7LID0LNQuKPr1I+zx7J/9pRfPlPxOpjclLy5PnEwxd7
TBxHvSP9ynDlpr7xbWxvRx0PpRuM6VVL5w85+ws4QGSa1zGbXbyz5MylHOiYZGozXdaF3saPlZP2
48UPPNmH5swEU+u/DW+cwk5HZfFq3RvYDvK6CttVGjC3eYEOZrrP9D9vHrmvP6nRxV+pzuYA4yRQ
8TAlRS3ky6jQKLpzf+Odbl3jGkp+1GIv00rAnuu1dUnHqn+PHQH3WUQ7KUNJkPGjCSAPbrd4oMi3
+Noz4CC39jIPwJeRupsO/m6A7lNDGP+4tDko46rzRQapzRdSMzTQsdkWTm9rS0+IlV489cPp6hgf
RpbIxxy9phJDMaPuD/A+os/KGaSkjz7F3Qp3C0KX3pyC9LRM1Msr0OSWq7hBHr0Q55BXBCKN5Uub
k2jbMKfGuOWJLYzsdawEM8ZBdAuP6i9X0bETecAGResIb9zMRI7e95ZSKjREin7aHe8AIebQ9hT2
mUbLipk2EXGmgbcin6GMY4sN3otVBbRdhlYwalIXNnztuST/Q63Kahp6sGIck9qD6Q1BdzmrySJp
SKisprVKM2m3Y8ZUDQlE6FDS8tE+8/vd02tHgZpc2bPi60FcWoo6glCms5ldtxoUpEpYl+DAE3ht
sCuFHAtBmxFyipCN15M0L7jIgkoFwLbZUWJxT/Y6GEUs97/IJ3RhkXCUDOrnefnRVpAFXUEk/8ZK
+UnscxS9FIk61RMjH91LBdmpPT9ORdszHhNUDqDH+cuXSBCl2Ihoa7vctYYscGEdH7ENO2QNxZEN
+v9Aoh4yhGUCcI0oQ65K8/v48b3pfyVVAaBF72WKceDIIYJ8z6+2RyvdL7AoWZBzC9C7ZuFwIq74
A3cc8mvoHxNwuapAACVTURHEmgHrhJHdYI2vBpcHjsUfEzu4tLEVlx01uWbUvJAOwGyHnuVypH85
dWT2mssqYM2NlCU5QRzmBo4x7Q/EH89cf4acCsjzuhMCPMSjVJYcxMdKoH5sx/iO7jX+MzNYt187
ujv0MLEhZupMdaa6SJaxnS0M2vJgtIANMa0HeVAZEHb1q0r1kjPN+yDTHLMxvvvDynE0G4hQ09tG
EE7rwnQN5h//smQbv+PWGdGtmg9yaG3lrnbuNmDcNxg/QFD9zzu6k0iOY6MJlREg6KsqQL8nlNKr
WDjVImW8TTXcjwmuBiwUZ7W/6/sQU+2oeZrD0vPak9UPN+jEHTAB76F8u28cyyMr1P3KBcsATEEW
OprirDa+179DfFOJe3I3ZIIeancp4kTEnd+dqg/6UKorkphu2lxvSlwVcSoBamXOCdEPS4SPF2gq
sYVbwraQcPV+0khcXyUqrocPgVrKnLByMQJLn1GzmgQXXo8tsjGAre8imfu0H7JF+mOs/9t5Qbqd
YYdasMjRgqpxZohLyl/ITkIVzSmBOzL4vUM8V3+vt/RXuGvS+BYzxsS0sGaxr+QKxpqUQDLvioTs
xY1ivMp8Vnw5yV7vwjYbLc3eaxoEeyV7VgZH6c9w2hoNXskQLupzS1F4OA2faVWpmdIE5BZ28egf
Pyc5aX+sT9sI6vrZExWHKjMQHTnC8iplwu03gY38Nkfb03hVbTBX9LhyEdum9LI/wC+ozcPWDARl
50g2n87GELJBE6Hb+k67l7HZOPIzJD3H88+QNizF3ymcye8hyzaItYA3rA40ANde63OlL9UETNUp
nNat2jI31wlQSPib20QFxXoo8c9yeGN47kJblXfssWqO1kE8M3dT3hewEfmOTIQuzgDAtC3Bmuf0
Sz4kNGycKeM3QMKaEc/9jSDpBm41+nFDfj/A/drHgg8tDy7ZyE5m+AjPkcShblQPWKLMlqqZ2WCR
o5N0J3jYMe1S91COYewCLEkdPb9JXdyqrOdTWJs91LeSV9LKxGIgCHKfusK/4sO/cxXS6yueXn9p
a5wi+iV3+1xRNNuRqkSvtdPuqm1HhKOk4EmChAhCRXpbS/XQzDgJtZl5bmv9CrQ+aM8s1MkG3Nsw
nPNMsQwCzYCJaUkk5ZkOObXZUHQiuCpES25qSiUmIQVKkngKG0+EHcJhaMCetGO5M50daAtDBQy1
YNjl8AiWjPt+Vjxc7zofU1KRzGqDnQopbLyST/VYPKte+tZdRlGZtUmFo51BPnOiDaLcgMC96s0+
VyV/UyvPzAXqkYtWdApS0Tkz/fxEuNTXHXyJ0RFwKrfgd7ojjGQ2BdlCKO6NiYyDpsBg0ouUWkAK
ampoB++D5n2ks9cT/zFJgFa0iBIf1cy+ug0LA6IOdMt3XEAF8ePenupDefPbnVknZFxadojEWKSK
ATOKE1W3Lv5G6gcVy8xEl0RExgV5pDjm+CdrebyCscv5md+05+qP7roXcK8CPzGDVAXFzoF6D90J
QP+EM/z/TS7GLaPU78OtQef+zWukFWzzBDD+URPD+iHk4C+9F8m3NISfop8djCcZ4h1fCXVUvMiV
dg8s7eqdfV4btraNNbVdGaovY6/A1rqRGCF3FiNa/sIu+8oohAjpcsF7HryXiVQZVXbb4aK5QXYl
riNOHlysc6sfyxpPB5YG0BUtIk/z6IFBZyAHUdOjTFyFjP+6wEdVD2mDKypGUgHfYf6p0BeNQIBS
ZDtCfW/HI1ZJatKJ6RleCRN4/qyDbNbP0wSJSwQheRB6YKBTZQT2wsLL+fWxUDx/ydii88nNpCb2
RvtxozCyfl7zqGePD2lgNVqqwrNGvRDrUkhPQQ4aGJGMJzN1tz0/99WL7BKA1j6Oc9wGB5n13rhy
yR+N8RkckcWX5KkorV/Y9lqT9FWLVfdt8VmhwxIX6eJ07ditN1MktPRZmqSevdkqgMma4ZRVigEd
a7tmrr2Wi7/BIzkw32/eUv9WRcZgheYnH2Z5Ni+D4d/+Gha6BA+LH6oYd9bXgfx7p8mfcE2K6NVH
g2g8kc7GFbuKmHHgwWIcMCJ9zJ/vj31VFzjPjk8qoFoe9V92D9h6ZJzdkC9pIEehRO+DmxOsPlsx
nSl5YMW+6D8/r0a3Fx36KcblSaMqG1bpLnfD2vqbij7nDoGbXuIPsspbP8/JSBSI1I5Uc0j5za/R
6xFIbfn15GRSBVJGhVsg2buqXBE2GbKvyaTFWMC2ygqoKCrQlFLtFm9jUAZnh+k6IWk30alxjpvx
/NHnff5Z6nfGycqAnRTeW2vTJqV5xDoVbTtd8iIdKAEkCu4YNgVYgqztIY/G773WmpqSH73WoEkM
2HkFJ+J1f4w8mOESyoENvOcsQ65WgvNhNJBsijHLJ7Dr27KFpVj67WbWzkzLLJqKmIsZpdn5vAGC
ZnfyxYzW3SSuw6V3+Qc/YoqywFF4OoY08ydwU97BDp+g76VLEYSF2ruvlgQTX11iwJFLXh/g+gjR
WHpG7VFmV26iiUxcGCSjPvck11suwSLxITO2hAkYySKoxZfV3CU9DAEG1lX1X4Ey/9qZSYTpZqnH
vQOPfjPS0QZMvEW3njZjEeJA5Ul3nFxMaJKjW1M7ec3gbQnSKvfmAloE1a1bmzaDDEEXksapbX+g
T9TPYc/EfpDffEKWpiV1NBj0bCwOam9QnUu3U+J0XcOiSzwH22ml7SOM2/sSstbYQmv0Sgn1k36X
SdqXcgvmBc3hcciXGrsJHacIVSWPZjdAqNyUU60PaNWf8loV49uiL293CLyy0nASJsu5Vx99CEMZ
MY/QNvsbfY1crJfjUtvefmV8Oa3L2YL3PsgV0gy/s5EAupdr9oXpzXOnr7EkKLT42QfcWNf9VdvJ
SoiczaHXzXCv2gFNTOOfZO8phNKPFguKL57ipo4HouDE1pSF1sW0f4PI8u9RF7G8epDNtf6VA9o3
tHs5JHrzpEE18jAumYKGR2YLKCO+yZ3bBdNIP5vY2V0aulsuGTzVD0MWX1cc7SLC1rf8b0iLT3ex
hGAsl9bSmJCs0SzgfBhnphg8jf6k1UTEpfeICaACgCZmQIqn3aSQkbyZKQ3FK9iVrhbgUr1NxHXK
q5XxzIf1gu1pOqBypGe8dfn+acuFAIJMgOqCWQWCYQ2T9bij/3jYTDpAEV0/5QM4rvKfk5V044C9
ub385/36lfqt2FNPU/id5FNYskkoKSzz2nIu8FSA/obSZYi3BWMEeYw/u2CzC2oUGBvyy+t4B22G
Pz8VtgT72sLuyVs1Z4pADNQgDfKCr+5NqZYeQEXeNhKJ9DCjFnXIrxe9C8n/t2xYdftpkd2kmyLw
BIxZ8w2IaghwAw8vUzUwekZs51o+L5WmcvORyvk9NTn8gTEci8YKrNmaqKY9lUoVQmiOTOytFMA6
IcKPrYpwr18eMQjaAAKHlzVDZjja2m3vDadVWfD+lH7XE9GPxOuoCkFO8nQS1JLFK3aJpLOTXhdh
DIyYk73ege0EZiig2cQ8gPivf68N5HukjjwphTZh7fJFvvan5VwgMp+56fKcbXXZ0wuTdItSQEnX
27cxE9VE4Ar4w/Dk1PxqEBiJTp8sxjzu4PG5uA+53kbHe8kiYZyEu5v5vVrvphZiZ+/bxogMXQom
Q87A68Ki4bF2MjCTb3TvDuT4AJ208vkFKhcGuHf9AbP5lMMKO5hHlTEF6a9XvfwJzuTX2gRlR51D
TVK/WF4Ap9EmlWiFmaiImb6DUYRSKJuQp3265WbJyyxsjdWI4Ap5L6+11ixVBJJocthAt6eV91+l
jfRFV+30Mm9KH6KJ18isJovxUYCOBXoMyKwh6rwueWZACx2pEz2tMKSzlxSo/TrMAi/TvBglpOve
2I1fONdmVz9Pl0LzuI54FHXvi8XMpGn+S2eSE/QV4Pp0f9nfuAesaxA0LxC2qOqq2stT7+eN0p71
YH18+owVVTMlb9KvOjhLidSaZflpIhJ/HM9I1XU8dg6y60TZR/N+uS1Zrt8XvLpEDfq7ohZ0AhL/
ok9jMwD4m61sea7qaIzSV+5SN2RQTH+aGoJEvjpOLR2nzDn/SukydRkpi/N3r499XbKXNgpS1Rwm
K5JAJNaMq7xdOek2MCUMJ6fUcb410F+n4Og6V8ve09ImxdvUqg1bAEtfTaZsHmp5WDcrPayTrlLQ
3UA3YsdkvCs8OHJr40s/RHB6QHR00WiCuamZ9OakJI77PzBTuEF58tcuSZ6lN5GtOhmHf73QKbYN
NciYYC+aGVbCJ+FXEZdrJyTbBaMIW3bZ4hKVxVRfVyfoHT4WsBOopjrPREhL5ZflgatLFmfMUiZu
21nKRdiNnZeSexhrfvddLd3cQHbxLb7RdorhphhCa1E5EVniSwAj2vKSYMzLalg3VLH/HnjlTRAp
V46FedqcDsNSqCaDD0obsslRORcKX12mRMFnFsiD27DhBvWa2b3RUj9CGfHwllefgQh4R0MRYQoN
VyHE7Y/pDMFvp7Pav7lQ5rpcsb/SH23itv2YxqVCyNCsZ+CetynO03CkP3OX+MokEbKyXl3twzIM
NXpgGIy2YhW0EafkAoIdklhEkzAZtuAGlDFV/DbDd0nBTeuvk+1fuHio5cHK8u09jbOrTJC1JKc5
lIvb6RPFb39TTh2q8RuuTkqLp50rTXlmxIvff88cdb0HSJRq1jaKtN91KBdSPEbrg0FP9TYLGXZB
sb7zNwqSVl/sm0uRTzav3tLbktT8b//VLMcugH8r6RZrNIDwKOXSG8JVabE4OJ5rXocPIm7zy3/o
YRHViRAbGC80dq3QYq2r3fmikSTYOTCZLlcaHUXQKBK7QU4IuXRJgpBzZ/qyTsRJPF9TcMRu4dWk
/h5JpbH65hTQaClhf4vluCyf13I4VITrLWJcyOGRSuigTUn5ejYygPCmfY9QLPqWuWhPyVYh/Dd5
S/bJrk8Q/VeTX2GfaYMkbfp3yX0SuP0GXMmzW8qPW1juctnMpU/5M/pHrdutLyKAOn67KvP8IcwK
X3xdx9c+ZN74uy/RqrMXSBE+gBfq4sU5/+xPFaRsXbteJmBP5mkK4AOER4zuzUzudMRxfZZMRym1
RAmA9jT5kT7D5tMscsHVQbAi+i8rJ6VSivpZ2OaTqN440YPz8cgvnJwgWnacHSEeRBDiRo0ZhRHj
Xr6E51i5Oxrc813jrLyZoSYqQfZLpEt5a9qJCmKl1J4isIa1qxW8WKJ3O2G0qF1rvQKiO+TJy4rB
wA/xQ6WD7xj/Q1I4DCoqYxwEb3UwMObdTTeM7sNHpesuqWHwTsYCco4P5fWXuBBRbjCeW2sFkNig
Ut/RSs/9fHqJVJ3L15cH5oUxEN9XKpGJBcyygSGkxQenYz6QJdYEKcsZIRORRNZR5GopAjWYQZna
HRyCnJ1nUIY8E9IcAfZ7YNgcZYZV1GaQfpqvvHmI6vEj2w/7ltZVSs/Jjke1rWPz0vLNJ65+m8GW
N9TZJ3SisGknUaykBsOXJJR2q40xzsy3H4MEuXfo++G7UCNYP35U6lXenGINI3kp7F3eY20l/0aE
Wha5aYHM1RCQk2wkSlArjKYZcV74qvdrkB4mKphrTcIqxP5oo+vmNgcv2lRJYBwEnJVmtmO5/RRf
YyQccdtRWYrspZX+LXOTwyv4Xr5WFO5i/o9sBUy2HJP4I0pJsEEkohPi1kMymDVznO/dtPNnJ4Si
bTYADR6FB8F5OAytOnIRY6DGfWqJ8/N1uTAlD07IwnbqqJiS8kqrXAYj/6B5N1Ol8gxVle/aQfXI
Tgn2CZrgr6JXCMdtjMzGsXUDuFLl8kyjiIanGFCymExsJLDz9s2rmxwmVj4kMrTJMPI4dug5bfJc
wAbye5X5DhrM/aVFBLXza0pOleL3OF2tIATHvk+uZSigiCERLmd+MlhZJ71/f705kyMF781i6627
JuRGypaKH/vhXt4A7QHfs/bTHa39ADAP0P3MhXaebbywxubxBcoRA0wraZIlckGfONsI+zKScwim
UsBHb9QKEqan2hHQDVTTl/atNotq6uU4B4hsPWkXw5o2DFkg2JrpurWk99NpgocV327bLmXM0Ory
vCMzmJ47P/2JTAY0pQF3LybVxljf5rRsLiqcOD9KedErzVGWBDdlImVmjOsSJKTg2y/WmtFadS73
KX0PrMwCWsOq29GSAHolBUrM8APr1/epiffETqot5Hp7yJxGOFglpcvsbUAP2/5AzbD+Qqjzkqf0
2pqW5ME9xKXhx+u0WW8kZAoddsOZYLqkMPFsOc2e5/LzD0mQumjm2sTCg5UgjxmlGy+cKzb8tzVw
1dwUdhZHeyUnBkY1xVtYVPDYVaLsWwNQrVAEkJyR2kqJ17CZqbu4jePnOoMfL8eShukRSzX8g4xk
ssnHPcCR1P68M0D9EMcq6IKadKlroIV9cLqFjISLQtEkXqrm5xTlKoZ+ptiooJtOxKOT/GWXmY3x
0k6c5UlIS3DJ6gb1brxHQc+CjkOIYOjtsG93tKOGyyFjS38QGyb6BpLWizDUY1t8w22/rE0nWg4C
gMxeU0wFHcglXVIP3kM+HEPedY1Tz7SYIuqVFY1gcXYs73dbWLFV7siMxdpnfwW3MGKrXga3EUhI
viQN/0TQNLgjQdbDWM0rKlvYUoGibLnxHFM0BOyr183tPeIGoonsSrj85HyasdIjwQbnYEKl0lkv
5F4UHHSPas6sPoRAINFZ90VQwoLpGfDtFw3vVC+RdHUqUqbOmVFtRYE8tMz8wYcO0/M3AnYmgRpi
O0+OEG2Fps726xdAdAGQGuAdjwiTdeCDTHk7+fGZnmlwL1bxPpDnKp1JnfOYm/HxOo4azixXx8a9
G/fyMJpW9PknSuhzKaeBErAuNET/FKs9pmugeGxHJx/dJAuYpj3p0UWmEmrthndkevBSQ+Rxt8TV
k/uc33gGy3blkT6yY38Njy7hJLRM4Wc+amVReyFQw6AYValcOR2kzzM9huK7bj2lzV+Pa+MUaFyd
UO3j0zv3KaqQHGAAxP9338WJl9aDHUYXwB8ixctaVXnt/kSycnNALpwrFVwxgp1+InSsoaix5j0C
d1Rj+jf9QJevuoPZCDPCrlTTrFA4ccNt7WaUThcd7e3uOhmlqB2SnxTw7VtjuL7KAwFQH7Ar63cv
miF40LcHX7IneeIh8JTEPgOlyqXRKaayHLJw0FsapsMUdU69A8alqg54rTaNXI/7/58zP/9WAVh5
mUafCIscBjoWFyPyVQmifVG5upkTCaWHAhT1Afb9eLFYfXgl9ER71cM5xN8ZT6yWTVGs8X8OXfcS
DC+Q6lFFAmuqR/Hd2uW0XWyBpyfu42yCu+i5oSyZ4i3mYr3mvOoI+79decfQ3QEStjSInfi6fPxT
qMl9n94I9JsshMkuEKAup/rbZ++OMfpqmUXEVDSxVzaKQB4GxuW5ukO050G91zfwz9xSdgiOviw6
p47fzexAqRjijlJQcfSgFmLE/C03xXXfjksr4aX34DHd95t8X4bYzHaVuHLmszZdZPAU8bkgg+v4
yuNGeX5tgwaGW3NDOu+3Tj+wDMwjZWB7VN0ScwJt47754y6o73npnoqmYpIw8dpFAQvRNRo4Aydp
4roZ8P8hkJluSuELRgRX/n8fHT7EIx7gdyukjKpTRVuDPfCHP9W6wz9Y1g8FzNX+d+pbFPV4RPls
M6FQOrLdSoa72ESW3+MR1zNljMKR7UtfDm876MWD5jUmxeSZHCt0XsPQX23jeFU5tCQec+NQ+1tS
TOjE9NpFor9cNBEtN3Df/hYtnxKurgc9VhnGtsVwFOO64OIdGM+ruXaqwEIFPitMbug5TArRAM7X
Ho+6dmVOk1+MBx3eO26lN9tcjw56bNxe3iKAXNEobuZEQxy40NLd7hbSoqgIaHtl0z/Pr4EH85oA
v5lZjYIM/xS0uoYIl03Qcjra7px5voiiaXZcv6NAisrv9t6vtBtNKLJOTyFSSt9zxHXNOmP09xtw
SNStz1CfU5+Bdhdi2YoNQjKGv+xfkPXm81wvH6n9HTxVTweopmo2GQ+wRapwDS+PCv6Yq7b99CgL
OV7Y1Dox3uU2UkIi1/O3O1mA60okBZC6HL8OOHPWlEVI6M7xDnPeMmkJQ3sL6NORSNP2RsICm1i9
qhODfYpBGVsbjVI1Rp2utnbylcKSwV5NwporD0hrcC8lZk54eiLTz+daBq5GOXNCaKb/AZaxDq2U
F5Lq3vpB2H3+4VX2J5+x1HzBppgu9WVJ35zcH+87IUSU0dg/kPFFYlySNd3l5Ng/XKwPVPGv/Pn4
srpIycRUzdn/9iFzU3lsuKRY1x3+86hMTmYaAG+vSLAgQShRPdnvqZQ9vxeW1pysmRm+urRjYez0
t26YU3N3pM2TF2pxXNsdzTHOcocNLLjQJCPmes0t7JDE5R/CINdeQgqI5W7w+Lwx0gbF91aH/9WF
Yagv48182X8+rDEir6wHsrqLPAkQbC1PiUCaVwv6oOXuXQ80n7bnj65AtMNAwV4W+sDAZjY1Dw3T
+OTX9zWmZ5VOqpWFLsQiDeVSn0Ut3gSxuBre4g8TR2x05zBzGlPwuUBqkHzxOsxiKxw3xQixOy9+
yMYfDTPWW6zliypfyKRq8u0bBwfoUujQDBX6c3tunv9OgKlPP2OX6qu6gd/7pmfmrW6THZXH1yXq
n2zZe3jup3lYaPkSlJHzmzIp2mJwKwN2Z8cSwpZ8YErMzyWXj+sFE0ixBQlf2oTUnR+F1bPWr3R7
iE6aDTYbXMX/pjm1QcNc3jBmfZ396HMOUeI6j4H0kHjzf6L4P4WShYPyOcEnDxjGp85wzkDhQnO7
8V3EKXsVWufHCSv5mzvUdXryseWxFrbbCiE+0fa5M78JIrulqfgYdIC5mk94dJ/Xvt05OAg516BT
62JuFDbcgo7mhBebeeP4hCmP1i8Cw5ZdUDO9SxkZGdymQZ11i3CxtWCBOZ7XRD5f68LAYZ+vFTjg
qfKovTsn/lX88BvyR6vxyIOLuyl0HFG7X1FAP8HbUy2aAhgtVNs//qTW5Mx45IgNlQPs/PT2m0kz
cx/B6yM0t8vHZxpYocJtM0fKbh5P56jMrCLJVvHDnm2d12rqFjn0yEjCCv0R3Hftty1rw40Ic89K
UufMl1C4YrthzahdxAEuJRYA/lVKdlTXS5jl5PStJAgI1r52i35KaPmSVOTHNYadr2gmWyT1vDq7
KjYyXz+8ushtkdQTsEP2nD37jLIAtn/5vgNvoEqq6G6mDdWL4AO3a4R37qyJ3loPqev1b7cyPaCz
mQjx89x0Onhr3hW6Z0PMVll3QKADwEW22ce4Y1i3XZGbC/Iz/slVg3bfKyoFZDPdMSfpi8yO3M5V
iuGy+rKlGrOTUg1IoHfSXNnO8JkvtlI4MDFvcSTrsooV/46SoXmxgJ7I6f159ZJz+1PpOsmK7G8R
3UOejD4mp3S95+3ameOjsAkuE34U2PoDK0V8WJNCB85msElkCRqsYUSzfVUKVPALfWK0SvBdoNqw
szJOB8yJgG9ZgNo5RYYoLr2wjKhRc6THMdDyDsjbICZQOvV6EauUcKlN61J6Cm9Ucit9JApFVmT9
9/KK5JD7TRbjDwWC6PnHt8L9dZkocJXPRWQIFK+Vd+qwdmRs4zK3ClQ2rKN5HQlIvJvLX1QcnIgS
jF4drX21JfqvDdNTcxDj3MUtZQg+Eh5w98mnNeRfF14savNPS/f3ubBYfdJA65Mcqo2w5itHppp7
7e1To06hXlICEFhztSSNirOMSqHMV47QV1/HqnNgUibjTNUywywd3fzgTMfpDhriYqjWKcpEESNg
rQ3o6BQQF2fLl6B941fTken0QXFgshcx+QdgT3F0lQHIAQjUkmb0B4rOelXh98bw9Qib/k77QOru
e4XtD+6FN8zUS8cAtjZV0z3h4ulg5evRTEoicM8Epj66kR5/AAADMlF/LLjARnKPKGIMlZffDqWj
F7cGfDiqJNFSDiTSDSTI0qSSIY/WpQym/3r227YxcW3kGmLkT57mAU7Yw/HgEG7gXjmD8S3f3SQN
5WCmpLzKUTZgQpzh8N2bGTnmvew1nUOceDGIpYQAg7tC5wUI0UxEAOETdSokZlq+IdMrzaXs19u1
1rX8g9dH6AHBgrdCBcZ+nWy/LLGou+tZsINe1QWkid5YDe4pltNs8d8gtj2asCkWpGk6Hq7/gHuk
NVh4j5ep6OkopKaNk/DyEzxE2SUqXTZn5ZJeXr/XGEYXH2+mbXLJr59XAQv5jJPiJnva4g/cFDgx
DkKgEeTTlPAn6XGO+xgnHnft0X/6RFlMckjm+4FJR8hBO87PFOP7gGCFbSOKqWqSUI6Bu2Z626C5
nJoDD1c6Arjeg4IlhsiAIvQ345pFmQ25k7sRjVb0ubHYmWCj2k/Rrn/3IOJ9R9sAKIX/UgiBOkpU
W8QMxrWurNjZBVlp/lkBCsgUZSlovGe4yg6wsQOmxVCzwzrW82s2+Avg2FHd21NCY7UxAZvtaULO
Nr3S5LhmamYkI28tALmRaZWnwyfTujc9wDwzGP54paqsWL7PFBdao0BtU8cAlObZYyj+Ytec7jXg
pPWgoPj4lujXsU9SnpYK2sOPChK96neqUksSM65Aj3JYygCvVnPnYZcMnNMBAhPnOCaPlM99lH8G
SxLjATU2sMKNX66XP5cVbU2Sf347K8VsBJZJ30n4e4YUoWQMVrsS5+CIr8OQuHLtKcoz49/hQokB
Vm7NLUjBhX5Q/gAKudiLkEmNJe1GeEjABA9oFO3nAD3B3XG8S4jadCrI49trr0WBrfGKbBoUc/iw
RLJqpJkoIc+1mD74t4r9xtd5yDai6QYeIG1eKKfx8qpPjwLwUjheD3I2wO8MoU0UabL5zACaTTsK
j6Hji5k3IqFA4INg2MhF7d2RAz2Ob4+i1merwAt188tJWxYDLfsbYoQSeOaXoSpHGNzWueVLj5d1
789mL6CQJ/Yv0JCno/KFM2AVsqRgatcpWtHjtd2YSxcSizQYc1Ky5ZBg3WTK11Qn1vyrKzlRsQNO
/yhzzoAiggWEQMWS2DsgOtYIhV8Zska1GMwgsfy137SZ7znni8cmlL1Av1RbBawrnenewhbU9A+S
ud0N2MFdWY1x59QdbnYl1HXcPN7cjnDTRXWee3WdOfR3wSTRItvG5Si9IRmr162f62C6A1kF3EWn
J6mbPeci+0IGqiqmSXRDCBB8SCSQ6Mh99DaNbTGNR61z1E17o7mJGIW7ajGLg0QuttyYsEpM5/i2
tm10AdoUNq8JJ2jdoCS4rPUU2GdQuakruRTaDSy134F1dZnRjemLv4VhxIfONatfRFXN1xiNmFqs
vCiGzfF+WA5Q0w0RyGhSNHXEfqTYox3zsyqiogrP5J4j9imbJlabQ5zqpQgUFAH6f+FTHmIIprtZ
7775jKk3Zx62d3mjtUocR+v20cPyNtqAvy8DJiZ0a7iXNmTfUUoD/W60iJYCeo0fmaLtv9tS5O/0
ff8MLLt2OQBwHRVyUzmWtMS/ViprZV4gwhYaRFg25zpSK8ISKW0sPmWuejCt9w/YTc16IsLKTUX9
lyRklqhjyl3HTOqJOEL0KQoDvrg+GSaLDeoevtuVe7dmgdrr1ZaWvMbaD4osshduUjN6wz33QMZe
RXdxzxowd3vtRsXjJY2L2Tq8jzHxRSYQ6VA6+8xK/CTa6Px/f5+P1y+pDo+EKXJrfPSy7JjUFJNf
WcipSFPWpt1R/KJVXVWWNj/oYS8fV2IN3GEDP7vAIQRTteVy17ON3CsIhloo74Yv4GAR/+GdAA0P
nnXvjQBqavtWEQAHN6l16tG6Tu2emWWoqNDGGjxEVANrInOKoznZ2r9nS0tZuqEKc6STwb6MNVxN
ipafJOC3tcSvphOvlS2ZmgwlCZOjPbZzlYkPMlGMxKGNwB5nFVDWptEOWrUoKe0h07EyS2SPoLuA
DEMVJlMZjL/NY6tfteiygtKISeCSqg84yiWXnlxf7odt5KcECAD9IvuM0XbV5lXfWQLnO4M4UAT4
Idxj/iaqELPzsAOwGIPMzBsjcfUxGmR4wWE5QmBIwsTx32bnQQs05m9gw1s2oAjdrwbZvGuc6Yi+
NlR/a/z+hCi4492mQ9VimM14v9Ozd3GaKOTAy+MLiJSbyOOnTZSD3SyO+7UftLn43IVBeDFdqmUU
BK5FExI3gTPv7NF1ewQo8Fdz/P4IRMuZLRjXDD0SoImN/A/tO/3FJ05RYAVwUWcVcL6giqCZKjR7
2keG6DuWe9KVYjADdoBcqs8ZvYse9S94BWcxYD/OGMtCnjk26VYSsQ1wkXNOZu6rSnWQQhxtWIzu
Az+4vD2D+gMtu6GI6HoRf0d+xYJsQc2GM4zEv+HkAecup9BGcAbbLQJEIV0K6B5UstaftbiGYIuS
AtbNa5k3D5YaFeRa2SGzTqTQgs0zV180hLFuYNndFV3ymsxY37nBqCDiH6cr4hyFW+uEjwNYFG4Y
UDoIgtTs2ri6a+Jd/IdaNgo9r+XV6xhHRa7Bj/HWOJG+7jEGTkTdP+Schh3bDLwODj5fLMj6hCQL
S3t/C9o4z4DHawPub5dazn2mRaVbasiq1zdZC36uanNPr9jq4TzJY2MMasjQYaip/8arGQJP6p5v
FO2xXM0FTogPGBNVRpweAbrjWQGJiO3jzRjoP+HyjLKB0r/FcwpBC6chprs3XlAsAX8jBvHMcl+I
6mWj/oJpexqbikFbmfMm+9X/MPW63cPUHB+8UFPf8zi10HCJbrCpn1RmxrxFXFCPorAmNCA3X97F
JHqY7WWy3tfblmB4xRPglMX15StNZHgp9bvNrH/d8PGPLhOxsxgGWHgh6ANOTcxZbQTEKg04FSfm
R9eL3M6HbPPkmWh5Mz8wTeXsgzf3jPmPqXrxUmCQl+PbJzoA2KcBJxXySjZSvTj4weW+0iV9ytaI
FbCYzTGKP3Pk5n3NcFuws+bfb9to4LE0R3iskFfSg7qsAbHZcSLNDlbqMVqcBQH8VLzoJRImJCKm
0+sdlHiaBJTQaGTC6rySJT10BpB63hwzli4TwT8FXPZVy6+RRSF5Xsw13ThdpKLiVf4Zt7daSALC
hpb11bUfx50rlvsp3y1VObQIphPAKdJpBvbOM2n5eunfcKV2C+BT7LQgvQ+/ZQkq2DkYB/9XavTk
uC0MQyLvL2NHRyinCH019FrFQRWntLG9qHLlyiMeH+mD3cUd3fj/mf5XF7dSB/m0L61QNrklpQ2O
ifm/nv6LHPer0MF9lKoS0OPsI/3J/oHk8rrNbBtuzzznzjYWoL4Z6XMZ64IGDc1D9fiyB8NlK4TS
a5VRjxuvUgDofP22WXnG+E/zUN9vsYTZIzeKI/Jqmf0BqfjOQDOu8SyT5irCAZLfoGLFV3xyjHOF
tm4aCKEuZEoxrWWEfph2jgJ7PoQqWlb53+8lclA+IYMYeKY84UsbeKrWsu0wj8Ylrz02UMwwJUqE
TgcVf0F/J03KCi4v6XckfH0GjNLAzLGjwc3Z1E2/WZu5D4zjlRmLGkbl8mLV1X3JFpdJo6iQGyjB
M1n7sKouJSRU0tcKY8EqxLzk+3282J78DritFUXqL/4aZLE7HXzppcpCGRF5x391GeOkr2ZSF2OT
Ci2XXZRb3C3UW/Z45Ykm9cPyVX/OrbV5GdKccPZmR0wWS/BavQGi9ciq74RZtwMjPB56JuvzaYw1
PBheYpmpHJXTasrVvEzp0/G/qpuQ5Cxtrd6kWv4Lec0MgzvH4Fjpufs/b9tCJsJ2KAGTIDhn8cga
qHRNxvtmk+daZlbKCfHl/WyzSNA3kk7edHqvby8I6bqyNWbGdwGm9+jpVsATSgTRbFZrOmcf8xJL
cemk6jVYMW3zYRt7N8BYscOtlBe1+yCLq18/7NszKgwq7vNcm0Tq6GhIrr1kKOQGpCYVVztNYjEv
0GAHsPzp36ZmnlmFUpPfU4nepmlIse3rPv2/WbpQMWxfRLpqcnPIpf1qHWdqgFkFixZC0ljT35Xj
h3cwvU+6MeIPQDkOkFZiNRlMhkCEXFvaw9X8Eo3Bdn06283kwfUpNiRMhiAdS2h0AalVSATNdESW
Ahv//bbGmhJuY/5N7trNzU5ufN/Y0o/R3OL18i5DlDekeiBKqxSYT572AocN820EvBSyEEHdEcV9
QVLeUmR6oGf+8A3jmdPa9U0mO4Sb085O0/U3sWNgzXl5mX1FfdQx8Zhe0XLQfj/riVAFtFmyxzep
uvhbnQ8LhgKek65vpBrRa7zK2alr9vIkY8UfHTrzH8Ojy7+UsP4SQxdidTsavNmMY8jN8wXNCsvx
YBnmM5EdY8C6Dmb5wDCds8Yq6yH5I0q19f+Id1gTvnrsMXd596BYovgszRmKaFlgXxOhduY6cu5v
NcnVcbBvmdG90hZY7J57yKKQ5gI0vPhfmtEIhK0F/8xtrxg6/jiZTgz/h0T4CrU3+kPTWlAcjvUZ
HmCtCpBPoetN+j1WAPD3HweCe4QDhNr7oTt3abJ9KYJ9HFSyIqDkTLoV2CivOaeU7hARbFxEWpox
NN/55GFibJ8L13o0sP03bbKE0InFwF7lEDLDiwadkufNmAIhMINhUKilVn8xsM3Ylzk4q6C4KtMI
KW5j1b3AL72s9s12Du1m85GHnpA6wzGd4rEcggD9pXTZdeswR/q7dp7RIkxjWnMQpEEtJjIqPA75
BsqqTgPAp1mWk+q8YYOPzuHGYC1KuO+c1cwrODJsfKJczyEFif+aDk3o5EWqrs2Si16whFTQSdQv
68p/nezYoYXapAKI2BwMUzE1TRfpVVl9N0cnSqxg0tXNVbkbxVPLybMaxnhRRf6bOGm3K6kRS8oQ
hctbizMyjKwPH+giHCz0OToZ1t9YymcbnWwYjYI2ASRhStFL/+85O3RfFV2rQ1Al9CV3nQznWtfy
HNbfzFsLRbv2WoWSdGn9eO/Y1g6Z5+niB9DQN7513sItWhq9pqwvcMDx+frtxBW41zX45MqBb3Ux
IhjZabhwqYhB7E/ylY6po930nG6QiMf9o5Lr8qnMb1wsAUhBxLDwcjgCpn2ElObypAsGnt9nGoSR
WGbIaXwReNrd/Y6fkP9S3nhFde8bOvRXRy/XXvZYjIEJDziWWfZM/EMgDe/E/IhD8T7B26fCcaBa
QQPXog4xG9FmF8WR4Kxia6H6BucQbY6gY5pVO1SlYt2OsjJR217qBq7lfXRn82uJKb5V/CzNyvPY
wxq9h0Dg9ivwirMaLtkHGRMO/a6uGv8cURTuEd6w7h87sUuFnfGwNJJl6EcAm+p1WRe9Mi9PI8A2
Ggw1L/740mMimaLsy5plCQ61lXH3U20bprKWhF0YdnuZg1IQhylTi3f/J+WQhesMuWYZXoOgNuJG
3TRxSx8y6TcDFIF2bONJ5klLyw3G0LK47opISfyvxt40w7KcKc6F0iN+mqipfBQF6nTkir3UbN1x
sGsj0jM0QC8Q/lNxGopaoG+hdhykJON6c7f0oXUHfzwkNpy/6Uns7qposZAyb5QFm09ZCJUp30+B
hrkQMXBA8RpVyDaaUfidKKw6ifYCC8Sjzx33mR7QEU/C2kbMYY7u3UdQHpZkxjZV2LQ9zzh0PJP2
paSjxXsFv2AHlmu5CoXXu2nM1HRTykYmIJT0EL6T+wACtE9EAGVYF4BNxDV1aykoOstF8JXhU/Oj
7dgNfg2KfafMNW+mENzNAwCFYb4zBeZCPPQD8ThFvtpAW/EYIfaih68LRdA+tsPXqgq0zUJXQIyU
KO+Z2JGzB5gCaNXKC0YIUsD3RA//KZt9ItfAokV+mZpP2pp6fEps/zgSs/I1EUflk8r4BxEM9gLe
WcsdQzCOaKwXCKp7zPuFOTow9wxTHOaD+pHxHsPU9NZUho0qS5/xG3zzDzlNb+6jeRdDSN6ti1Xh
FMpsxMILiC/3RPSctcW4AFs+IaJy0g/5pSR8UkotN4CvuJEO1GZHfTlisNSofiaIE6kKjsJCoyqr
mBE1obG/oue1XIu2aixjcKLCEitH+tF9SkdO9vDZ1irf50lTb+gKOI3WHV9nCOJOQMhP3O92GNoN
umhTBmWElEjj3ofDJJ+o7xbwh5KeH9sgZKaz4SE/zRQOBzPQ504v/dm0mBp6BxqNhLRxg4b1/qSY
E4GZ5FFoZJALL5HpiQtFX1MiJPeb00S7UQatvADZoTSyvKLnAeVuYAsMxGeQ2YCHdHU7WU9HM3oh
+BHD4PEUw/ZVQ/U9vuo73hCfhfiB7+uw9F+OD8AJcKs86HSynTSPwHxWQ1vppcYgmrJDDogFmsMQ
gWDig6xNC03kyxDQjJK1pQkJQ5wdr9I+ulbkSVgAu7w1RE7n4MOlZxKJK4sBN+0vVCOsFMy2GldY
XVuS8CREfjZh99nhfPEfKGa/CANu0kJRBDz/QkVjrI2KSVscFy342b/7NzwU9Pzr/OXOM0Bp4SLY
DoOjnRLf8Dg2nXkxvGTAG7VfNmGFZeG2K7y4YByiVu2uP4vqXaQ9DMhK0UY0Z14fzkkTdVyO2j6N
5aZ3Kk4ag0iaWqFut/lkX5PrB/nGMaCe3jwJAyKnDhtvPisDDzGSnRmPKZ8S9O2dBpJLoPqVNpKS
elPkyPi2boPUwtSNGSvTZ+O0lrvU90SAFFLLjpPzgTeMQSjuc8SToWRUCZaOGUvL6oWuG8ZbjIRQ
OZ0VLJv3YdkNS8JR1Y+edLHfn0SgY+rpeg00lzuu2OgabHi3yGPOjGPKLjQr/yjKwLCimy6ufkUo
JDQ/6RZdjp+sui82UMvPemdNYqvsrXPCjyu5C8yHygt7zWJ1g1LC+do8KYSp3CWD5wTgpc2i3PTz
Cy0K321oJVfR6KGVY+fdJrqj1TDcKyTrATV4tuM6EZyr4SST+lUuNB8TFiJLEPAyyclL6tSlq/mS
PdfttIZ0RJPbVD970i3QXlR1K3ndjFod20nY+5FWablU/kq/UpgkdptLDJKoPtdtWP6N1Ve1+wg+
55LFBzzNKbbW4W7W+5vtqb85qgnihf/3UF+eV2VsgN0bfIu/JsgW0k+w3uY4bPo4Um5KJJK34AJL
IgfzVPGz1KMmc7F8bcJDFgQZPdcOdOVhj64XaGKp/q2zHhlGAzp6WtOGOjnNr8pZp+0njxbbgw9t
td0dWEf3qXNrXBc2dKd6vtfwfuMVj1tAmlU5xmYxP5EbVflykdxwSoL5n1QscFNPt+V4NXTIRcjo
CqJQMoVFsicbfdH1MiRBdn38i3FzWM5NvLdpzBwwcFSf3AoH4Yp7fvnlI/RMM7zsJlGyfsITtCU9
sRU8EnAp6JkV+67K5B6tQjcpWe14X5x/0FzKk1tsOCRjlqM236Hx5q4oK6WUluYFiGUi6mXOja8R
qPY78kgjveO2wrs4iTcnmQQUXteNdRPha0gL070rRz6NGWpXAC9Ikql/B5mgZ6/pBo3i+/f9MgDQ
DZeVRmv40f0bmCVlaC6C5GYDeLHjuyG9it9Y7L79U2MQr6a9ZLTUbTS7TqX9BHP9e0EjlHgCigk1
8pPEewDLuqKQnQWFihKmBBfUE0wdPrXQ3AzCgn2PdyqF8oetBWHjG5YZAWPDNaEfwFhFAX4AhFjW
pW6XoRwCCeWIr6/CtAaG/IY1KPGS5osx+jtZ5yvecj9ssQBZiNetz4/n+smyCphCqcO8MeekDpaZ
eMi9Uas0TDDNO5SD208MLfw7uBUqKMlUpARJ/Y6lWAgtiBWuS/HhTOXkMcJ80cLxDFLz5ZubLUjh
4x8UVl8e1HYnP9sw3bNnhdiQ55uzMZ0tWqxnuAWJ994YBI2Y1+VUKPkWIgELoxW7Z5pXXMbGa9MC
zgemCtf9SShm+ZduoFvgY/JKoWuAfu/4KFb4g58W+nCy/vMAyoEkZHArmBYUfrDbH+ihUXTIB+xw
1oJd4yUnKO5QSIDRlPHfkJEv9E1pwygi2VQgUf0/etaZD1BgtQAC3paJ2iNB4P8fO6h34VHjYyUQ
rOv7PYFlQgb2O7IaI9oMzDaV9G7TItepzQ8vokKy8Lu/0w19sON47oGXtlBokaIaKxaSn3hzrj4D
xFDuq3b06JLGGX7Lhl22WXl6NdYiPSbXNyUV6Y2oypzPqcutHEtoFYSrD9sK8n3Z+3ETDFUuOEa2
u/1zLq2urxk2vkb86AM/U+slcz628IK+YAgImrBJN8wKYALSDl2soamKdJRmtcB/0yjuCGYCVqvm
KuIAhclI6ZJixb70yXcSud3pVHb/jBKFTWOXVY3AwpaHgaJQSKsZPSryklTdnv15l+0v9BiTk8dt
Kn2xB4l7d6Mn0QdBKIDugAkXPFgxeSpMOkJ8Ls0EUuwB2ECElMLx/5NVdoz157uNLmD7TrXionmB
RIdC9fzgHCsRCrYuyWrxMngDYKYWko/V8KtgdV7xz40AuGRKSNBJckHlcqgW/7Vr0JxFT2AODVm9
mvPoUzAKuiEUw8F3NWD7qCTUpFpxyB87IA2mMof4765Qc7GY74vrLdnp1GuP5SefYGIjisspx54j
cby1X9NQEhlkmc47XVsIND8r1HFqS6tjLTszKN06BKNW046ck+4bQrc6QxdoepC+922ec6cyoNRC
RaPQqE/aYb7jIyFOEeqd96e2Q8dCgM5rNsAscpvo6+EVj/1GETuyCBfhFHFyhDVn7lxdSBYoFMOu
0+VH6sQRUdox+T4NGr+6GeaU2ZFYxmL97qWDjXO2Md9tJ/fRWKOK288vAQP7JZ1qx2jFvElk2BLj
6m+78/FjM8vERZKKWq7Unq69bjM9e+THUpo3GwWPcliA/NyMnIqhmSuP5VYpHdOScsP6P+AGlz7d
/Uh1qHIVNC81GdCSvuVhejYUR8hK5I70y2qERLvXhxXoKNIkM8afRJNS7o3DpqvZiKDF2PXJRgGT
yCYk3vxTEimnwXYF9dmCofPbKlbl4YWNeAS1jyCkYp14tluf1p9rRa+e6P8OkuQ32qh1/bu+L+DJ
JkuLdQevup+mzje/pDdUmwGBIilCC4X1paUlypN/iwYJIWrUjh3B+RLBdXlkF1LwFs1bpMaS90Wk
OnWP11pk7BmpHlvstr+nOzt87AVOZgq8TBMP3wZPtUrY/bVk49KRYOa8CIFZyPqGxBYW9TpJQ1PK
gF+w8ItXclcLaobS8/ef9ZfeR2/zorvN+sfAqWSX4f2iKQOlxFq1Hfx3PqpDmv/OPJlMo6oAcB+N
lZtMHMLqWoNMwswdpVEWa/jWGIAQAUx2WFtN4BnOQLUZwZO7mb8+KpdSKZ7YBWHou4ycPdfk764U
tkY7qkSp3xfb6HZdccv0qAzIBrGsvSDexf0LPvo0YcrpObsEdY9w5j45QXxu2tEFvzc9ZP6SrfgH
p9krVU/Lj2OtQrnz/ieuh3kgss/bRss6MT1NeqoCjNvtVD7FPlD3nh6UJjGXRsaOXUpfmv19TdEs
peO8Q9nxHpNyBrd3qcNq02SD+dnHq9YeNTJ3B9CWw14i+zTmFzxZakYsQ74InMFA2PLx0pB8jgIj
tlHjlx/8kE7gMxvCZlfgdYrKYKYjYSIbRjsFZl0SOIIZyDji6jGWpnHRmASFUtQ0Xzi+hgGWo28f
iEDcgN/h7iQrZ5egGTe8rpOD51rO1+Pj3rOHXWt5V/v5Hfbvg7Gdu8dIfsogNvQLrql1NmMH/ziR
6R7Vqp3bEnM4N4GveiOhlp+nfzUHEZ2/iafMMoUoJklzjCnThmtJWLOr7N+eqFTAqoBV9xVS/SiX
gM6WpU2V5vbBqTXOYAzPqA9fLpYPwBoPJPOTj2o+8wAg5pIeFzOHbUw1Sne7Crad7BEbz9sBRFoP
tigkZXWjwwpdRNXAPkNLplOWRuOz0NpT0R72ZtmYQaeDyTrPZut3ZmqWeaMy0uQlYTvz1avTO8UY
j7sa+st8iNZilXQI+e1ZK2a1Uk7CiCHIcDljFyC8aqxtrkreMOlTOQvYPFkSMA7VZRevBGnoaveN
R2iZURNOuXSZ88mKsWOYv+SZBGMJGyW487AvaJFI/b3EX8pwNbzY+dDTvpiiPnYQIbSk7NlUH5Y0
tlj8oB0AgwQn4zi+Q8r6+JNO2sapbNz+AobH4CldxjSAGg2RWCXehEfsuxVYwu4foYo4PLGy4nEU
L0hObTi8JA1LlfXd/VYZWmjxBNPCGvvbezKN0StrSWpy97aPC6rsicd/n/JhGopgmHrka0R2YWWM
oWcKoEiA3JxWsbVDLxylbZJsemQQd+ah9sI03lH9R/dpsgVPHXQBH1mde92f3vCaHV4kc5NlA9PO
vlrI8bhdgXP46JC6AjstEmb9FvrblSXN879CwpHlVvjNhPhmhRnuitrWIpAeRta5qDIKxhcZxIu/
lP204eCKSjtaz/a8UO9qodO/oTvZhyC6cMu7xdfoHCcdSq0pF+XhyWTgQXB1yDLv/bR4DxxA8Hj6
2vImS9NSn9vfu/i1YmJLmSpYbE0fWBwoMDZ56RXkkN1Y9wBIDclcUyfuj4l8yB6z5v+FeZzpuhZT
rGwIycY7SN7iB6zNF+dpj3lx/kJvi2zu9UtQKZORWVjNkLt93+mLaBR8IDx2Bw8cKBi9Xq+C2WEy
9RvvSq9NcevXFozlceNyXCFketTfX3ijblfPG5Vqwq7pIiekz/4/85J4PR4CbOQlI3FdxTj1OMZP
9orjXs2NW7pID37iQVHaWKwJiXtomonhODuq1ik1cfMmlrTjoKtYnbPxBPGMud9S7pfuPzJcU0Np
S9mz7J01VgltHvDCEuKrLTZaFxO4ItLsJ3F6isZG6RxHCleBnRa0Miho2wKbK22+nyWfdl/UU3/H
TL/Wz0V0hTO8c9abfG5ggypvnJz6fKUDsrIEmiuY8dRFvka5pcui/X5GUOJgYssJHweFqk4vEnuP
Id/01iUBNryJv//IKWpu+rfPkSdsrGs/EwNu4JcLko4RB7izy9Gj7gd3nmb6XmzulIWUYRClmFu3
uAYv3la2plp1Zsv+DGllGU3h7+z2egxzF8oVYnbyPKZisImK5AoAZCvj+aQvcOp0q4/k+v5LKk4V
SXJIgMOD5y0Uw6hAnz9iDDkjaHI48a2tbK/PbIA9ro2GfGKqgPhFK7ETYjXI1jxuTQLzg9pT3PRW
tRp2yrRruqbeukdH4X46yrNPtb0Frk4LaLsZ8ZIG3H3L9gYv2rDQP7Sd8hEH2JXkwl9/bUbGKeAU
nTgUvnDElcj//ZNlpvVSiqVQcH6Lra/tkzP9jOSGDTbeyFcz1VypaeQt/iCzwHGtqv+LMcG/l13L
mb85z5Q2irOGk3z8OWeqUeQcpFnDe4R9kpbOPtSmlJy/MHzc1CSXO/tq0KbNGC4mc+DjHMtQFqJi
93OU5c0cGTOfSnl7HnXuP3j784QC8IiUQ1sXbJpHReXLiHWKNEU5LYCWTfo/nyE93FFOjdNU/OvH
jGJevZ1iWj6gn6CQsAvCxwT77M0CzOirepHWIg2nasp1eWOim+2PhGkJd8ykiWLQk/wEqoGreuw3
Um9dnIZO3aB6WrkcqsNAhLW2Qft6YDaOpQmSABuy2tWIVP7+BqkOfw/nbigJJydoELi3JJgDv3a4
XUZacvpDZPSvF9xnLaKbERUiO75TZp0f/RS2oyd2Ssc5k6pzU0wjfMHSPmzjcYLc4M1FnufZtYGa
IhHCU0xbH7fOhalI1my8Jwui8S6vTmmP6Y3j17zqAiOvdcv45yIdMMtOhUQJPEWOOmnrhn2Q6F8Z
Cq1WC14Bq+rrzF0dlxCRkURfFACWQAK/fKR+dTtO+wEhHgpJh3+8bA2w80C19fOxjVHGjXEfUgaV
u9XmJaYTr5VeMV+4dy/6h2/52RUVV4qm9lkyvtYaO3HM5Jzb8seVL+SvLI0C6m5b6r9ZNs020F50
aOn3yPwLjbdQRZM1HoZeCyWZWPjQvosOYsT2EJNL8E4AZl2n6saNFV1pNHS0I8utYnXgnXDVzdM2
o1e9I2BXVXwpBzwaLA6PluO74Mq//mxUgjexdkw0uLDEFBSRCio6dq3SJuPlaAESNq+D37wNOehI
45T9VNm4wsJrVMGqe1sSlHs2ez9RsEheWZaWuZ85eIvw6r0T6flrfYQ7OIJM558fd91dsxoIurQF
MrUuRlDvtEHgzJNFpYqiisHv1GXr5mip7oOR8kFv7Im9L4qxIha8nrnoMYG5kUZZHGzD5EylAyix
w50WU8+/SUkO2lQvtG1/QB3nQw2DR5ryP4xLOBtbBZdFF2DSYqJTebRJJXzt6VKpQ7bQRLARulWm
zud06Ja5oaa6HEAIxhTz7i3EjC9j1si4ob6S7zXcTwh0iH295GwEVmXAZkxDgfqgHrMaC1QiWWyN
vvzbyy+heH1YOE6mB7CT+UmKEkqrgdTkydexGW6Zuol2kbl1FaC5dfXp8tyA3XxqA+9z5zdeC4Yl
s1tpfk10tj0IBOYYUBnXIFkOvhEXnCyY7POLAX6KLXJGSJ2g1TS3uW90iYuBvdmcFoR8rTPz72zQ
834aalzDis0/bSFFdYFC1uNf+F5FWMfuWJ90d3B/RVcZ0+eRORkoHPizVyPf6VC0MEGXWcyt8Yht
dtIc8k42c2jVPtiRjUZ1bD1S7uENRBCEUlIQZYF5gJgqpfip6iV7mU6drx1wXhRab/ImmfeQ9C1u
i9/kxdPjfGM7wGv0q2qWOMVilEKWtjhFad1RCvHkLgplYAORgROuSSFkq0cgLlN6Ar93Awg5jVBe
SzcdxqNaH9o4/t5KHGiNXsB5fhQI4w6EFSgl6XF7YYdw4hh0hmD3qZX/Smp/0stDgYVq4WwiAkPe
ISNakksakOjmrAIDZpz53nYghPXS8lulJKqFWpKzUXOoRp2rfApTIly83pDl5qPeiacut62uiQwh
H4Pml9vFCYHNWd0BW7QykUmX/JAy3iRUsEj9D1/0CKGNPJjGIqkhULVuhozetgFrnWjt0aqb0uNl
pkEYq5maHQHZG7h9HrF3SDRD/oVVhN1uKE0Tefpr8mggCg/kV/KM4RXw4XDNcfUEo0DLBoJm06zT
idwSKwQa+QBsOp2QxmZ4bfYG+f93YF4EkRkitvKe3FPT5wObNaSSO9SK3ICom61VDaDHRlYN5zeH
XPDhizg4ot58xrnWGXNooAbYrCjB4R8t1wCpfs946j9kwWtk8bGChT8RlQ8tqTM8Wp6q7kzl6OfK
cKGBToEoZztTUfWuvujECDbsEB3+B5oAKuAxtvtfPpTPDu6p9RpvBky5ZVp2FVKLH2czzPSJkaJl
fNBi4FxOu9CVllgFMJPhoPNvCH6tBHP9fWq89ySTnnaCTzdSEOnpPZvb/vv7hNUq46doCXBS41tS
GHeyphw+moy9tfgj5zWI3AociMIjhMFFWYjt66x41cmSur8hxP+7ucsHhnsPCLBgKj/H6PYx9xQZ
22HuspearmVE6aTwS3JYiqtDPUqKLTRVdvLTDtH/DbDlIatc1Ruc/naw9cxLKiXtIJ7ktbZ5ag/x
CA5LPlEpogT3P0JXIXRqkkUcZx12Lj3G/Iw+bs+nwyZOmKtElDOoJF0h7xOb6G8qI/OsHwB2O4+o
NKueZm64FgDsN1HohYNtc0QYn+p9sT+abmJ3+dhrgZf4FPRpsZOvGu3n2qk5N12DJOw+2RFdZSlF
HCgXwysvUbRVygV0iVxZ/s0fRHwj4NwJ3L3Qi5ABGT98BALEWI4ARghUyiIZ+ea8oni5ZhUwUAYx
xAKL9jkqq2lBXcQNYIj6vThWrQVjd/SnJop3Jn1QNhNKNPfhKFGYc/azitPpE3SZ0Ha9GdOkmJyy
AdWxS6XFbbmnXKX+8IJX442dN2y8cOwNZHKlOG/MP1kH9kUbChgwLurv3ONHn33qSQYswnaRdpw6
SFcErhsG43oElt/MLiWFjtsmcwE3kL6x1ppfeMn11dIIh5CZxtwg0CRJ3h2dl+vSFEjtsen/oj3f
r6efXRFjUzJqGXW8tNWzbjAXMJsttUTrpdCuhRCvmuj2I+3tUYhETtLmMZcnM0nDV1doBKE4AAeu
X1gftlX7H7PcCyMTjnhqo++2p+RJkQlTiKPst5zKrmhJQLabh/yqlSr7fQ/cYOO+s2WFtgwuDUiH
nCXsiYlKyBF0Xw+BL6TYTQhUvRSbPoWqUXUAPhkAj84vDIQYvOhaMDVP2CY6NnR9ao+kVCgv3uNQ
WAwHfV+Q1Elz+kfGfa7GSeUbUdKFltufTOhA4gNwih5L/4XpYKObOM48242itFgrpMdl4SwgwnD9
qKCPbCfAe1H9TrfA5NUu6KnD773PNWJA9PY2kAGFN3mi2ZZ5/v/1WrEPnuDUCAk3AOkUiO8/IOmc
FFKw3BSvQOzniukwLudzzRZjCjZ95u/nN4OOVzklAC32QEhyJ6cWBJDM1o2+vlgtTCkQW09Wogep
grLDR5lmIumxZPknPrEo518CO2bDYKXAFbXfihtVTYtv0icJdJ6tdWm3WqCOCdWOLWWh3T7+t+HH
uYsB44wBw8mGUX6Yu3aPNhGX4ZRe+PIAKfGBkHzUD0c8iXNjzqyPUNoODlgNRxW30p/MkggxP9Mj
AdtesqDMwle2BXZkF/lORDbCK890vZ7Cmfae+O4Rms3IOt+a6KbJHdISK0pPzwRSCa1+3naeKDFK
O6QfQuAV3eFzsxJBKeKlVQIWaVsvsdec4P3wbLozg3AnG12+adGt9JXJJKl4t56OIw1mk2Q4bI9N
yqIQxOIXI+NHtbKoPSe1uvnNp2prdwixcORjLbGsS+2KNpRhGKsmzCZOVBytzaHHdtEzmZElBYXV
s0iOiwR60TgrZuvVA3Pbx6QIpvowjgILGUF0hr2d2jKAk6ovwP/+piP1aagHvcF90Sg5rJ4bUkmR
vybRl2l2RGI+cstFcsoO0wcVoqreLCeh7EiJUqF8x1FOFxW4FXM5v5Pg07UXkryiKP/Xw/JC5YUF
BwiFMO0RjMQW0gIEcE/EFJBw34LXH8mKe+DWywsQQDNLEQqpfcQIXWXfic9pWnLwxlkQocMZkuzp
FWR/vKXiWAfU7Dtr+VF7GN01r1AHp1cdZpf7uzlkxpnHd/Mq86gCo5/IEZUaJEva/Eay7QHmCkRo
5McPJyIFN0lo9jV9LtML2/S2qEjhT4vt9D8+yyOH5yIfrD0dK3cPoYo3EbVRhbNIqSHk7OCOei8L
vYSdjO8yOQSskKUuygMjLWxe0jNaYFwsAJ8gon+sAdRf0jR+Y7vxtE6CQzrEZjKUeUI/fYPgJDTa
v5Uqz2OAtw9lnIQUopg34AiEah9YjgW1WJde5Nu84OJ6Q2eIErzKRxZO8/QonXmnmu9wAySYkzKa
dRM7c1Zbux5nysc9l886OJLMMWOxFyd5xDoZZH6uxAphNdQCbBpVZ3MFc5dUpahuANF/6LUg//wY
XdKCyiz+f3E8PEB5iprIUqrqrtiOv3XZB87nb7rsD67x9D5RLTLaAkyWReV4xiy4l8kiZ9U4o03n
aOp0szCP9XOSfNdI5iB4YRwvczQe9Osu2+TlRszuOREHXIp1iWBGcGmdkKOl3wF5NmeiyYhIHPRC
KpLqLY3W4A+FsFWzZgZxRouM3K3cv+akjokXnvBOIng4xxDu/zNkvt2D/R6pviO02Av8UUwbTeNy
aKnM231gAAeSqD4nQ77fsHNDX83tEyUqp1DFga19NfFB/DJD3CWtVvTSkz2xwBsaW49bW0ssCYL3
kJAis0HE+msUBx4IyDqAFnEStHe+JKQ5fldSwy0XYP9rsUJnfI8BKKMXDipBtd/NNpMp8z3L8BTB
7ECLJDIk/AIeibMgKRCK8rGW2X5tnvmpmas95FI8dfs7+XNGb/KuIvsQUvThujItlZDbpDcO/4+S
WLF5c/PgpY3doq41UXjdjA+CiZHfg3vy5PG3LmjoFoJgCAAF+OhD2a0QtgdimltXMVZ2/ddaTw/w
N2owe97IjyhqGFj7MpFtsEiIVqrOBY4zc0sxjungYiy1MZOiYHEKSmwXN0eM3E10stCWl6VbSdsv
OGt9w6XAidoHmoO8hOHey89JoqqURvCrhczcrlegvTof2iaMzoT0WxrUWRU0fxJjN+xQAkVaI14s
+Cnw3nX1aUK5Sklvv9Worz/oW/u95/NCwD2DdImYYfCuJ84+fdN3hvf3+jLxlrCqiKTFbtL6qD94
gDTRB/D8jqkQFNqoL8o8DIuHVRFkLwyRiJ7yDiXGU49jfALfzYP8PH6f/s4FK/D7yZs/kkuIziUQ
yIZaX3FeLJE3JoCKSQGhQfqQSoaAIqnkFYOnT1T+BQWtRFXL8jGinPUdRZY+qeNJ13tqRf1GMMts
RKIpXcbswllOijXE0JIRvzg+Ofw0hRyuIu3VhSr9bdhPslQo2PgaNIJghDw4NSIZbb2LKYaALJNB
n3RpOqsPNVHEyFwIq2LaKyVuActKwWd4eUv2ZhdtMS7GMJ8M0qqRLcty5wUvNfWGtOIt3RBfl6tj
ih3c0PDlUqC8Ggt0hJCkVItSdQkt4toK3dHMsGamDm8v8S5K/0PCLjP0MbHBRu8DgP+TTP3zSQrO
Vj4pbPCw8Omjb3jx205aavzvtvl+8nUOU8cs8rFjMWNZHvmV9N3vTcDltJ1SUtZcSssiJfxcjknf
gIA/f0aVdlXhZT2lumx8TMPyxandF0b4nfbm6DNVZ+pIulktpFsQBOU7RtjORHGPyMK6mCWzU+if
4af0t9w5Pq28XdIUJr3Iplj1fD0aMUX8oGD+CQgqcxYz1dWflnIvJi4WJXsgG+QDPEs/9ZmFBX+4
MqAObzCxWkWwqlSXTOOQYTIyhcuPOjBmJRPYrguOCtzWV8IAmTY1t91JMVmScbJyF+JFHxH6pnYN
F1OUzGbaBMvWwUgWM+EI0hcHVVSYEW//j6S5B32a3eqLBSLNKvnHfJCB09KmQ/ulF5AQEZfEpdtZ
8QRKQvReay+K6A2PbVMvEUpnuyhHV038RYy4xyWkowPb0lxlbv7o2ishr0lxO04pPiupyTmeVfvS
KPxE7F6GmW0LE8zjOeT1HgWQ7XXDNFbFcldk1p3d5itXJ2V9fkgoWD1ArypN1Q3JV+5vqSC1Uknt
UNTuxBgjnq8wslKdB8dIWLiUxlPUHOduStExL0bHjLBWbbTzwfloS7kJRsHhbQj4VwixUBuIs3C1
8R9cYFNpssrudjqyTyYYqLBWVseGSJCu5EPd1XDwiWam9vBQb684Z17eaqT87ie1FIzjaGIjjiMp
l7pxt+ElndVcyMeG1F4t9hNnfqmSY68A/7jjW/DeFHk9EMewiu9IAjNEiUxHLdZ1K9V6t6Ybovmj
00HjlWp1vNbMzr7/h8F3QMXTThODnPUgLrSCGdlA8FJPw+Sc1YhXI3ULjL+fByPZerDQi7sytCca
Hp21rJd74t4EzrBpHEMjU+hW/dE1ZS8ZudF13zPF1OeQBxVuKG3ktpfwlLsRh8qIPPfU7pbcZ1dA
MXiJL3gv7MpBlVoM+fZ3GMhs3fwg71GpFkeKRn1tPNfugFEkBXn71WJcKVQ36BRByZ/s4FZ30BIY
bdiI3JxdtX28kbtLcuPvpZc8LdZUGknP6jk5k0xWQAsn3cdRjPNa6LRLq+iGOM0Y6SEnRyxcvfiC
JaIRpdqExGmWx8C5tppqWlbNg74xU8riCkq9ld9Om3C6ckCFd/4sFX7grGLcoRT9wwG2kNBAkc6n
9elX6HZcZ5gNuRuY4RYhf4CnrrOBiGywDi3o52a1fz1C/NZSlDMJ2aY2GTJF00Ni3X8AWhVV9Yhl
fYEImzOyLLca8sEQJvlTbL7PwwPH0yNuzTkCJ5+IeeJp2ElpyA+6mx6IFqCfhcwm87poKrDzLhkv
RBc3iOi5zwur6wGc6nkzdB4Ra3Lu6FC7F/c0t5x7VTVUvzcCw8jkEr2NZL1Wg7UBnBAcsPOPjFCI
u39sjgsYvyL3bx2eYDi//EVJeqVg/9zDEB6geeU/s4WVXlO49Iecem5q6/Nbc2a7IFcHL9C6OSdT
/dLZqu4GToemIoaAdTl5Y4Ucg/lQRXgeZyTvrfb9LkFI1NeF7h2r5YtEsNZfkOMaoZ7crKTQ62d3
Xf471ucV/gx0Jaa3ZdNqRcV4P9PWiAUX74tw8QH6NhxvzAr/Qx5AxOSiPZVqE2jkqc7iRnnycS2P
sBxsaaepTtbWy/1Bhvy3V/mQ7w/kkRiWjLv3fT75itglmsaSP9MZ26RL9QxOnwz2PfLpncCvdXiI
DfviZMKAH0paSgPvVhysN9XyC93zgTePRjpyGZ/H/nY5jcIiioN9U7a1crabxfi9QkxzYrSXW4Ua
qKrghj+4JGHrWixc3DmhKE9CNPNe4kYsur1SVqW6qQZthyILhcnSK34YzkX7o5Yd2NwS+s3EF9Lu
GWvgTsyrJ4UYRMQAscoN33jE1Go1FSiiLPZH3XIHIxX0YfJDg+WdfWLV27G3KJjEuR7Yg+gM2b4X
RpeMqngfblIH8fHDNpfxvfKSLChEd+6evVWRyLMHBDjL7lgK6uKRSGt1TnTsFJ/jkqfnuH9dsxQ6
VWxZiNFfaC7PCrrO8hvy/8Gh6yNu+iiChBVWYsXDAWtkljkRqhazNzuRBWdSjTklU5ifF0G/opDX
qJ+NweESNHIYN6+ykz36ssGaM96aGtAVfyVBNKbVGUFQ9un9R6qeEV5HkyVZq8hBXTqvnvFlnAMP
gq/W0XNjrVRKKij74RZfC23fjcTLIZpJyaCyJZZq/3Cx3lRb3SGmxHJbAVo556bDhdEG8YVyxzCs
E37THos3tGeJqsX4HJQP3qOU8JQPT1seKABc1a+KnGqi9IIkR0E7p+r2HhqIJ59byKDgPLdBlo8i
aRTqS0y+eIBlCQAUV0ko+4mBk0ZERJ66NiwN3AbYfAYDYRx+fWMCqzxcrBnHLYPd7LUQeoWUArF9
3X3JOxjC2Xfpg5BanpS8X3N1lIs2eUMhn9IUO7Qcg5f1zWSZrHLGsQhWnWXmUiaV+xGrtYiWd4uR
MPBgH0sR5JpOsllIqbGDy5NLM1lvisefbXIJFasy/HpYG4iTaR8Rq7dc509HAXvqRu4WvcO/61J/
xaRwfqk7xRtXefMM7SoIx7gMIgci6d1qga0pDZrUWakhHrGCJiQRu25KM+y+tHXRHnd6+6dMtp0Z
VkHt02x+M9MlIhf255vHkYPe2I+zSfbcaXdCw8xyZZfaEsk83/xqByfA3Us4WApzHXJNCsCGtevc
bfptahSRoIQVoq32QTXk9RDu5S6+N3JiVPxj3fLUn65uX1Un28tmrQqPRwzLDOANsls9GhM+JoXb
WsDwFO62GtHc5dBnwfq5gw3V8xWFssrunW7Kk/Kayz7GohPdPUKIh1ZWlpwKxgsZAk5CsPTCogAd
XEO6u6QXn7kZLmWaiLc9xsHXZPjnxiafJdmI7cXQpGbRK6PeMQ2gr0deoSgVnYnex6Eym4qK+YAV
J+h+zuErRsBv2M/fiv6Lumv1Q3AJ8wAjMJn5SfOwr96gVNY5RqFWrdur1WY6uyOgaLUt/hSTBujX
QvBdeDVpyi//tSakQ9T8FkeVGxdTnInU+iU9sY60KN+/0jDF+bSMGNCp3mbQW0tTPEpwiohlKcKN
p/5COLARU6N4GLqONi0yDpqvMgdWBFm+F1R/kl+PLEeLpTBEyeSOqGOBlVN8o3vWP/bbbAKLpbPe
Sxkl5w8PnTlix62M9APcO/y8P3huGsaomsQQZlV/mSqL7qzn5KPOFDagCzd7EoSyg14Jdd+TIcME
QZtisllAD6DrDJPm3o6DuPIy6sZtiECWR5e0jowj3qROQK5T9i2qdKs7gyL3KcKD+qzRVZsXsrZZ
vjZ6QfjV642SPd/7EspsP0QsiA0DvHfJjQsSCN9YZkVYCnPeJALOUdGRj1PwR68NvUkjAdViOn7a
0PGlyzFXq/9UaFN29poR6NAaGhxIeD+oCvPBw8qceQsmwzI0nSR6wtXhZSObPOk3ULSQ5q4S5Ikc
niDwMAse1kW9BUkPliY1f3K/O+DNNnLjBsNjDckEas8pUhE9287V+5aPOBkgBijils5SOxPn13Uh
KqzOMu5qy2vF38XhPbONPCZKNEnJcIQ+Ya65mDEhLyokBhRJsUs/8KVK3jcCwpn3rYdpJ178hq0I
5UKH1L2wCTd7SUyVuiH69HJyES55eLjhxp5Vd+uXfLAUt4xZYBKgd+zXyUH6csKrcRl5J3QmvlIQ
mtxiQxVhRxCD//h+8/0OLawbj1h3LSYu6NzqgmCYTEfM/RphGf7LjWv536HS02YCwCeawX3xaGgi
XlGlDG7BmPlLXTz1Csh4Ft4UCYldzDzsNs4fvSu8WL/o9nLYxZ0kZbcagDCw9kStvxsKeK0GKo2G
LZRLmi4CO8M137aQLphdarFpl6x9sZp9cNAoUSZ8xjMZ6Q5bLMYdIXywJavNxysrIpXRDyderoES
FTwe4CMQCVLDxgFjIpUQVdScN9efioe0/iJOZ3k2LXP1+RF7Gl4GSf35T0MHsI1o6kPoGEdGR6KQ
sRmMoSHnAUL0rtYYcya/k/wrz4w59q7GH8rf7uT66FyKYhF+2ZxLK5NSazatuuAAVCmVbHWgXbtc
4HHeIuiRaiRfaw7OhL5A7GksKsXKJfge6GzoPZoH5s4s8RqnzHFcadMp7KNvy2SeeFbP7PIX/Qmq
t8QLnss4fDmMatYi35pJn1xgiJVkmCZPIo6Kcc9cDzcx6TjOjcGVy+e1KwroGMFGhuzSIIHo/rWm
RE8XQr3dAj6AS2KeVKkRoBG4CBZM/Z5xxJ70fozyl8gdDaOChp10JMNYnaF61H/pS5aQ/dnbPduj
2LqKhxLuEKzklP0YdVKWpNsQ7G1RkTGOCdZKZ4BxgE7a7+aHj4i4Hy2ZzaFGod7iqOszm9mihd9i
NJlxG/HMno7I/aW9R6yL6YBA3RpDIyZ3Yf7oR1+iSFQ4n6UqLJTECquoEjPcE+MHR/jM5nDDkit7
Iyd3WaVLFteR6y6oBXmAVimj0QPg1DS9v48fYhu9VBj4DBk3ZkfMvrJBDVMEf/bvaXX9VLmdb3j6
JOUJclwJBp2liHvRdLdAoxtbEnzTgyUJf96cIvn7ChD4xl5U0ITfn3fQSI+WqqT+tjroZm4ZJgPy
JcETqBN2kXMb4TM4U1VzG+g1yUUNEzutFmaUChuLE/ZwHZ5CUOJMx2N7QJJzRYYsigRrZyWhObwY
1ZKKl1jOVT5r9INAYZES5daJvKS1zNL425KZlGLiZHzEttCqfUlqYsgU0Qy9RzgbCWG0qv/WtD5z
rD4maOfXpxMavaqfn8+mxwiNcsnvLzgv77sSzQ7ZdT/OUX7T8q5pC3rMYYQHIea+bE1YQ2WNaeQU
VYzGxjKHfEcpElOsecq06TwycWi/K5DFa29yX3fvCn6QYWRp6Ww4R+zU0SczpVnBQDEXovRaNAFI
CMw2OCWrNAWQ5vQ7cGSKCG6+TWs4fDNRK+zkvzGJS4LbhHFRXS8Q9p1Q+yR9kcpdZZ53WzZOq+pr
WB69yJFTJ3NXTWiFCP3F3k2KW5upFamwIGL8Xyj73z+TVrASm09yyUUXuKB9o70ghMcUzZZmOhp6
ROqc1kPD/WOvPUkxMdCKVjEUiZN1NrdFE1x+f9hsd2gpjAUU33Igfa2CPZOcwgfNkFn216BvNe8r
ZyDI/vYy5j103yUnUv0I3culrNJ/ekwvgUsJ4OOXOMw05bJ2rvnbv532tpeSMDPBM8A0ZV7pA1dw
AhuIdmu8qRzMUdjCTRRlYxNO9MU8LBID1UPmk0fx+VOdcQfUk6l7SOWfjL0uVQN1voLnylPS/DQh
ysc2MVX7yhfB0D3Vrs6JyqULw6ZyoH6C86P3OeHS7TVGfnGd65P/ufgv3jblOQfZovHYx5SvbJrD
WAngDb32g9ORUK8u1Mdoga6b3kZnInZDfaToKgLyN7mWn+1qO315xYysxvXhWbfi+/H1Sb5s3Bz2
bWvxhxymAGW97cZw5f+/h1b84NNaq3ir6O6+bXlzh/jVAH7/3yMICWeumh27jXncE0GwOYXNubEE
B4L6FKe/LF4A1Zw+Txspvd4l8qPYX8zekoXHsvPWR/BG2TIlSfrAk5wh/i7M59OP/DRXbA+ThWoq
7gFMOMu3Cd3+DVi+NG6t2vQQBXsjiPff7YIe7fCDQzzu6BlxBl1NS748E4KwRWUT3hgs2O+6tBXs
rvQ9JLWP9LNosJu/YdyZsQwsSYvOFSjxuLF8pwQt4587xK53aKw9yPAqIfVwEcASF0Ra3UN08Gx8
7RrNebZffrBquu/39uk1IAvZknOlca/q3VsEmPYwlHrjLYh1f2bk8atPMIZA5CVwOkEusMNp1SQq
+tgRBSBdmMyrcgcssjOxmBpzr+sURcYddumZsySe5M6jH0luBDwrV1/lG6DXCSKr19vxQotCZPk0
komb1U7uGWT8f8+4pi4xKVsvqiKt1PCNk5UQPELivEzU60ll426La708meQi0CzNrO4fngGahKfg
aGFSnj51dHRmJI03hNBLoIvMRSeiMeUqMI4R2h9A8RT8Csx8OBPcNXhvrDNVKxDhxhRLSV+2SKzs
RUJLZZD2peiB1p3vt+kXViojpHmgh9VadWjN19Nx9y6oSYq05emgLhLyKMhyCCHnHEGwK6Fa899S
F+IUhYucGRK+kE1deqc4mgXjWz8fXX44jE19HUEAPrYIckqbQJ1FHSnTbrer1oMbbrb27rRONLZS
sux6IQYKGznNgrRh8EKT8gSvDNsn5wcLhymtFgcyto94Gw0yNfxckzV6fJTqaeT1jtSa91PyuQjM
MahcBCnosDo+lqaEgXktP2bbsDExVhUimFt2QFb9OqdtHSbgs91a60wRrOH4/F3ArvErDVSfjA3k
TeYfeJu98wY90uh8kqdzJjrUt2A3+3YM7W0PS77b+4ljUrN11nJ66NDANoUW0Rns21+8Ue86A8c7
XZDhvGxuX4ZHcv+e4SW7MomgwSmofrSNZGle9q4f62W3IYSBdrY/h3xbAdaUyCHWLiE68mliUtdP
rYPQN1186OM9TsrGZmofentRcCSvlcpGMu5JeRdmmDxc+7xMQgyElKw19mgIeNywKQRFMXxcl0EN
wudtIqJ7hnQ9X4frYtUbOKhhFy51lDuO9S5yJ2Le3byMzwbBwi2NPZv9RJ3T558ctvehtosRLhBe
qs5sshsJMPR7n+5Kqr4ZD9qgIzSFC+cfTAQhif4xdTp87/1sqOVI5mhkO0xaPVGYRQQiIueNgWZf
PD9YHW+mk3/WDA9FOeTuYXInbciSCX/FtRxTOYHsXfIsV2OaeF5sWGCucYb/jsRDdiq+aPGvEn9t
7vTlgINO8YrSkHsSvOPVLFZOe1ixwWuU6KyLeSxqmK49Cttp/m814SaPmcYCHCxhtgOZhZHDfJQe
lo2V4G0cqktVyqlmhGLD+hNDWTOF6W5TX2zvtg4Y//AAqAKfAVaaymGQ7s7k29Xmb4+JZB07W5MP
5u7lKCyTV0aVS+I/I0nMaZ+gx4TmhigVvx6qhYpAiOz3y/MTvHHr4cPMyhGdjlE8pRW3RwFhMCWh
rrvNQ0B5rQpGYWKk5XPKTsqFPC6gVm5nkveLXC22FYmcw0kSHTJ+vvCyYjIqwX7A0gwHckPYq3Ff
L+Usw/wA3fyPOKVds+CNLg/rP2Y5tESiNrxHTQxZr14l50PF5qhG8R/jf8Jtm4ldpH5voqW7qJiz
RS6TqR1EL62ngTRS7QUVwSkurenCVJCIFoGBykRRBUP5CmrlKiECoZe+WvwjMtUXyryTVQ2WQ6/h
HcPc/972ddNCPVtev03lHTmDAUZDsBPnGNnn5v9WiQQBiI4hIY7Z4I0osBGwB2p22yEaYHFJ0Z5n
Qt+ndje0zi1U1b2Cxq2PZGITQEBQWidbCUjRbnNC42PKiR9INcbW/Sj/WUPR7lE7oRVLlWodv9sC
h/Cwcov3ijY3lCI+CwvSCatYUHkPy5MpTIU3Ghbz9EMDJPv3xVWp4It7qaewrVDoRGvpjMVO/IKa
9X10pNhRIFpXTY4AwG/ROcPqDj3RfXer+z+9UbmOYqJ/WFuXloPoWU3EnbXSdTWYKD+NI4A0Ksu/
4kuryRU+wClqNFJ48XW3I8y9RzWSTUODcO7ERp6BbpFru8sldFYyNG6KlSfnLr/HmhhMvrOoIvuO
jrpi3g/SSSLSmqeVUDN2JZP9DuTS50XoY+9yMojl7HivqORN2NCcLVfjC1EL9IU8ZA/DQLELsUH3
gajUqylJSYEvhmAYG9rNCSeE9uImUO31+Cr5qWjfnIePe3vFPWO11bkxMPgcodiKDkark8s3WQqD
19nZ5cFRXAj/nfklggFMtlyVdqZ7N3JQVwv/1/SVGRwRaJJorOo6bkGPjR5AzPz/ozBHmgzaOihR
w7KkFjvmjXezFqJKqOUGSvCuSfC4H4xWBE0bbngCCEfGWAsjrfEol7Jl/23yXeUwoKLCMM9tHVt3
RMGdfocHMmpNG4+q4b8u6JjJ2+U12+7RZnBTs8qm56rKur4Y8YCiShZOwm1RcDljgwoa3ihTtTMi
BFx0Q6ukx2zQd9z7kIcDFYpnXOrGIxza8h8zicp08tfm+yiubXhLIcelA3jLMoHUBBFOt4rOJgF3
K7Evm4/O+3SqpK5hGwDbQjLn0ZdEamq3QyJuuXfbVJrSLokE0TXGUjUPBGrSCDEleoMlzfHNnVhk
8hR4e9z/snkozYMZNWrnYk8JFrKS/up7arhrn0BDYvSmk0UXW6iJGpSim96XJeXxxGaMNVrFgKrX
FIQwZegiuGPiN7evPZmTiCUCGBI+4Wxf0u0huRAs1Mb/Brv40zJD3z7nVxp+DVfvpr3SaBU3KS1s
fYBXZCemJ1NsLs6b2LOJBUsqZ4altziuMUxq/pjY0L7sQsar0T2QhO1JKJQrJ9/dt96D7bRJlnXu
+a3a4cpnaklgneujK4rQwewh78QRgR1KT8vBhdzglsZiu0Vh9AjngxTUeDvCfCrJ+8fbI1/PpAdt
ao/IGEa5LoHbQnG6RQpfgUb+gf9yvO8kRSrl7EsWOVLzGcYVC8o3TdoIWKn9tpsrHgOOtw2URQMx
tOkattEaWV0x7sI2EEOq0IKrjw9Q76avUPPDrqJBaRsir+1RmKZD2D/glOnB5mre4LQb82UM8w6U
HKIMpFBJt3EujQGcDzlh0bitUEKsUj22evVJYED0A7/VZKVrC4SxVCzUV1W9DVzNP1LGpeKx8Zy3
/VVEtZUf1OUjecIhvzm++sI+e1q+RrwY+p29RqSZ99v25V22xFf7E6Ij9Eu320AEal0ftM7YGXPo
rZG4bEWf9RldIhjREp5+ABBsdSYhxD8Eo6+YAy5qFh0Rl6sOmxyElhTgPwE7pVh7tdbcNWMnOYuK
RA8OeTujrLDKi8VzRypSCsFRxQE5UKb7H33Cm5CrMBpnYaA5lMgsS5WYdzqAdYLX+sWnNI7KwTPD
G8fhyMU53YKE7QEN3ihtMMe4q+ivw4MGOiDCibobPgUiuSb7PPRlztM9V/CbRFtUUDMlV46T/6PX
PBkh+s4E6+WaZ8ebk0n4IIJCrb6NcJZ0HOaXRj4i7HOl/Rv+wzF3FswGS8e5qS0aVwhW9loV+FLl
vqVQPY4mKdvDIqPmQL2xKg9+KaNck+p3HDxGfx8UB3y02MGMjXC024eGYZOtwSAXIi4GVZJKIVNA
hd78EWm5jn63sQEA87a7K1XDSrpKDnXKWzkLcr6gvDKsuPLxVhN/P7EyAJE+3+SDt8x8Bv9YVKWo
/gj/wIMSjNIgfPcx7silrBzBxNJShGwg+LJfs4iqk2gs/IiSovEhqojiz25sMyayG9s3GLuAw6+D
ZAhz53OC/+A7trkKunGeHVs8KW8YT8/yJpO1yPcVf3abDGiqfNqI2G5mot/byQzLmz/Q1H+aD5F7
9vV3srRHyY+QChe7ayBNcIgdEazDlgp5WA+eohdLRqw+BB//BvoKzV0yjszcdcT4nFiSX4QiaZ9k
Yj/taVrnT6iN19psRusjW8OxcC/ZaUKs6EkySzFAOGzXR2eqtJIDsEOw7mz4/k7FezmXx0uVjuw+
8Upo3Yc2ZCOFOE2U/VvC2IWxBfozI8K9XrP334LnfAjhp0RshWIqXOn1YoeDB4BNk67tJ0jVg0dq
F60Cb7JFz69Z9MqTx6oQkpcjZLNbmEdgrmDgXOqLz13L+ey7/5yvYaBuNQhrpgOJ2e+UQXa3+zDn
JdiuLN4T8snbjJK71+l4aaMEgjEVD5uCSnVAJYmaxjfAU7Zm4xA21GVsBS89DAdO4NfWNlxhDTCk
7EuqacyO1OfrNgAApIMvCArvcT4UvgTesWOCpHODoOsi9My7vu04FUR38SRk84/IdLnZGadU5UzU
gbXAsx3HMGTT5oCtQfGOJyosBBq0BI5LA/LNiv6TyaYmNLdXaO8YzRfnJJWbrVwtB7jzRmYQpTeR
8rca5GyvtPQWxIcJYHW+ThGV1QmFDy2HOnyGsBR2C6iUJSDAlPc1LI9gvcpII0Joo4xwVGBYLM+W
CODeCycNobTfMt5f3ZlFqbedG7S+me0IiEXCzQc4ipC2r6oT9tqPpytvdDoOU3yJpYLYKahGZsCD
h9Er+n1s0wuDOeU8+AXkzROQVtViWPAxtc1fGRwY6IoTBAJNfUsFY/FtEAArSAfGcj8ERgIc055d
/+h5dWaC+5QX5uDwkF1nSGbGm9O72bX1IxIRbvkM86DVhQCxAm6Lu7cpFYO9tB7bR/E3oV2v43lc
/LGc6R26QcZxxi7e3HBpnjSWnzID9Hg5j3AbUDdJ1GIt3909+a5ycPek6ndlgwgKJ73VibzAPxDF
MnJaMRYcurOiW03pkVX8glsVyPomzQaFHSU/NTA0pZPiIWTAPD2HC/lm8o/09VchL0M7PNtlHWVa
rvhcKuu52acuN5rW1y6oaRszik+OiIX33fegT3MVGd0kKduoP7rB/KtXVB8eCYPpAtxK/5k/3HpA
x2bVo+4021iywN9+AVuRfNp8TRxqRETZI0QRs19CVsaIBd5F+SFmePpA3EwjlYcWMdfQ4tEvh04n
5q3/PwgE3kUfwqNDQR7iw1KW7JXHrV7BmB7j464x9fVZfbgv0DCCfMgHj6o0vno6nzo0dinRd53u
Po2K4vE7HzCvNz3LUGx+7GG9MPFPsKz+AgLMMvy+dFuNIwSbXWdoTKgfZzREgXJxPDxom+bMFWqP
3W6kpMihzesRcvoKu8tK2WobBbH5tM+sJqE70EYiA2Edzfx6uwGCV+q2znx0B7rWanYIn/kLIbXV
mY11XNNq7tvj0Vzkkvi25JDjH+RcPVCF3plTr/qQK2Fc8AcwvtEvPUNit6tnBMjzjnXqmiKAo4tr
FHL9RviQ5WCNrjlpiQ+Zyk2g/mYyWuPvmkjNTV7YA+3E1Z+1TBjmgT3dOk5nTxsmHRGNmZwhh+pg
cWepj3NTB1EM9E5hF3SqHbHzFKbTP55WyBB2tN4JNLo5TYYcyA31HcsLOVKn9SU7XiDc+lMyEZ8e
e+73hpxA3ni/Z191uH/incd5xWg3bOExtYPMkZRlji/3mbFIe0bqCvhh57zACy7au8PHBdx7qBGr
jZUcPv7xIYLMeBKTmtH5jy7kW2DwNgqBmP3Fu9AToeHZRv8C2daqT4YFIW0we0hr+8JROkb+rXMm
6ZyiKMYN4QLw0vQC54MRrkKgardmIjYbhqXTCJYx9pgMjkvkJNdDr+C8qwJPzQKFiG8Xaqpq/YX4
VcLIaqQ4tAIXrEXqlLNxuFRtJGYvULxl/4ky37WPLkxju2duYFBN7VYW63mMPulzXnP86Lf9T3NB
ISnokgLMTqircotRWgUY/2lfGXoFhL7xoG/eg2lMIb5J5s/ddIM8uJXMookFeCuOhuCG+unFlWTR
Ji1ifgJNCBJl1x1WDY4joo/S0GAMqzKJpziJkxc0NMNTfJlTzhDvctcVYozELGneo0gZ6o60Aapq
rKqWYdpWDhOdF+tSN3+7k9Z+ZJwke7XjxXKxepgQtxri3e4Hvq2Pc9pkbjxUvxabckmMqL93v3zE
ClxtDkG+1OFaZN72fUl+bk0LxY7twKZVxFfdHQ4IagSPp+1gs8y0Et/JrdA8oGONqDgThZz01SaG
h5ZvkADP0htEOi380SuMcrmuATITAhSRMfb+5SsIh2HrdBqCHxvuoBPzQCE6xbXtsE5zFMHJfOht
l4AUb9qXsfjBrl5zX42cVkPCL2sgYeqj9OY/AykDPDnA18cuvBkdDW/sW0ZIOlQFPHGNQAo24XRM
YwWHwYzPtxJLP0VZCP4+8yzmUg82rUitSwQWk/RjwSHhfpPrNtQYTtApUu6wk/D7ONtfPS7JjLCF
9QNECEuERHiAJdEod7QIoovR8+Q12sIQPhoNevrrIaaK4QLY2iR7Xzk7GWqcYTKvIeDWqoPN8tTY
rg3Zq668zWTtQiDQgjllf5XvpKpkFvr4RtRD6gP4pC4Xf3M/+pwbqSgH6knlzKXZH446+iS9+BlO
3RWwW+Rx3KKa9EctOK7KyPvFKUE0EmdChT7OSqutgsuC+QVuMTe1m7iOLYF1bWUIuywkj6E5rSTS
TambNiJn3rbvwjxpRZ4LuBXPI1cK/pv/2QJsJwDXhhlUbr/ycd8naCHFZg5kSoY2KgfvmKcYdy3G
fVyOZH2g5+Nu6Parqe1Of3af5Cu6v1oNY7wPTIbWWQWrF/b8lCp5rI5DQaDDbTPJqxPRASAlgEYB
U0qwIwAijq+5V9tVZiwJ4r9j6TBr/lOzK7TtJx3J7bB5U/gnxPoN1R0DwZ8reRzHW5Ktnr8absQm
vSbO8r/JcOUAwq0A72w5RasCX5sCUgfvll5sh7zr3v8fzs4AnKyP7cXMcp7knSGSZqqfIM/7B6ZB
7tkAGeuznb+KCHss+wJHXbxGage5NmpKEYQzBA7JNSLXf1cEyaX+xNO8CQcXBXQbHfQN66m9EK+a
OMDlhqiODeJWtJFjb3cSz9TIVakW/p6g4Bs8kAcNRLU9QXCZ40vC3rGkaSYwZsfA8S4f95mfC2Q+
VQrMyKJBxFONEY+Sw4uw7b2XwATaQNK8cHsFZuHgyDxd5A5rlVGQ5mCX0kSED5MVcpne9cOpcaC/
khSXzHW/2Nn/65U0/WVd6RyW2HcD3J8BLyin4tRyVER+KaKxJYEWql67Lo8fYKtoQQuucsvECLC+
Tur7a7KkG++CGYklx9LgzLja8E82R2ipZQ7yvMPKPlsEh08WRjMFy1qZ1SGgKR2r1aQVwHa1Y5ys
TnFx/v3uE+KMFKVJ+oD+9nTZw/jNwRw/9L9lrnKIxLyak7rEQ0PlJHeJar7/rT9TZ+S2TM8178px
ZNPgT5pyngIOk0x13aR2K/itrbq9Eq3ibqVRcAax90HYjvKcb+Po/NE6Ajq2sUYj4Ok1PcmDQERG
6fclCNFw+DrZlqpRnp/zBO45E0+dqto7LFnXeG9irr0uklr+8METbFVnftq4mKZdnLkT03GSzVE/
+iU5J76sfw1F0QzcCgAw8iDtukz38p89+rLgRXgEGD2nzAMHz3TruDIz94rGb72I7KWa9w95nLfk
/PjVwVf5f0wgaXke5K2L6qtrgtyUxmfGNQyTTol48fdDAUNFmcXvAWxPGXhC0Zm708D5x7bBGcip
j/gDgpl4bAKrI2JekxTGVhrRaJ3omqtUzPz1AoYvmBMHflR5ONVjMHt3bsaBt+DUE5JU08euYlvF
ovWPYxstW+AnMlFUgYOJIYllLToyUMzAP4LPJhN7q7OTj/W5FOg81bL0YEQz/b2BHNTyepENAwrU
RKJaoE3zi9flJ9kTVGC+hHOGqoGgMhpzIz12NVr7MESI3kZlHrSyWyNA8kF2U4d5kUcVYr+JkmjY
qahTgnZodWDrcDVcBSTgraInMCWea/YFx6v0FgvOtGRWat9KblJEKZbsP6NKAvhLnHnKFpYn8YN6
lU+UxTSBhsw9EHKbTvNQISRRqQ3w0oUymDi2WQh1LdFGzL4hiLaDP+caU1hyXnQQa4BYrgqDV797
P+xNteqk0N+x6+mYx9elbCFutfkGPkHcXeQqRrxkbSp8vcrRi/lhtUNXNgt9abfps4PsJmo85Ffe
sLRRUkrouiSd8i7WRtmYoIQ34f2z5MtKujUihVd8ogSlO4tSjazg2TOeLSV7K8WGL0uFLwXsyiBv
0nw/6hjx3KZo4j14cfYE4Be0Y7yhBm4xHaQzRLMcQT6JIPwQN/KoWfRCHTf+y4dJblOFHl5Qkch2
B7qQqMIzF027xcUTYwmfOqi3KlSWuMre4mZKzc2O7wLcSKR9ZNuj1mElA/89ecTp1gqbUerMK0I3
2tlQGoqbEnA3422muCz4Sbw/0B9uqXmsPKELs/AAHuQaNuvzb6BrDV2Vn/BQXioxqw4wGbkwS4nV
SR+CS9c2/VrWmPqKiWi6C6NrXIGMaojuRdUvE9k+wfnEdfYMor5rWpNyETaDGNEOLSHfwUgr5Z4B
YEjVwCTy6uXySfC5NyteTz56r9/DI9DPmtM2gHUdHkAzJQ4SmJwK3eTez58y5VLxue8lc0QBy3P9
LgZhCFnX17R+RpuWeDnHNnSD/Mix7P2D8CoFekt29jkEgW0m/FveXVaSphVgzz2O8ERYog9Mml2g
O7BFi7fr8m4ftlZJA3Il3QPOdX4ym/Z/nXlG9B5uimE/5V4gA5yTNj0ihKwRsjeSU5g9hXSBYBZ4
736nh4KoYIdhUhTYQVHYzLCMh1o54i9YU8GgrzA6yUyH2ySOtGXL8tBfuCZdFdgILqAbrXRx1G6P
IPej2Zaz8ny/wlX1ec022UW/fAraKk8EJs8qT5MO9/ELAag2FeYJ7LFOgez81NX+LKv79D29Jt1m
aD6ic2IOjb1zB4xoj1sOPGbNOZK4UGe8A/pjpoAy/kwR3jATD+z6zYe20RtQhW7oGkkcEh3BSC0i
KJYYUdOTXsW5FbnDD0VspyWbvQc41h9SzJ51VHvDzneWvZBqAMzVsGOsH8qVxabDvPoAzRtIdgqF
xDvUvtVVG1huB69g0bD0FoNKXC7EBLgBbvXmLPlvA1cf96txDwtTwqJK2CTLZhWV6lf/Zr0r3dvo
GGg/T5fVb6FymgnEJvIIH2B+fkcFatx3P1IdnmkjYzKcC4cp7c3Trg6YcCBAgBJd15aF9HSXDu6H
Gr09kc5XNMk6oBrdnpqoi24TErrvMWyaSxamBMuXlZwTNaTd7zaofgzFEwwRyCPt8cTwhaIIqfbN
9GruZSeGNPtnP/ir5P+6ANENqfAjTk+1QRPraiN6mBq5KRNj55JUMZgbay6vIJkoi/Cd/g11m5EC
b2UPz9mZyqYBDn1aTbYf/dKcKBrrc4EPPYbK7Z+NG+NmLi4EGkl8UBVgBP0fYyzKGaCp0fZ79/HG
6xZBmbHknRg3hjOJ1dpqFl9fA4iMZNlZm5Y0uG70fLGEtqe9XuITsooRjh432BgoMM3OhCG1t+Rs
WynLvZH2nrw7TbLd2l+YLjFdhuPdwj7SKz7dCMpeHxqvJvKZi2HX6M0wdvYjSDkxM1Rwltzjfpzi
v8unz7cX3x8RYb6vXFnV+Bw2xDOIJxLxs4Fa8MNaF024gKzaLfnS5Mnj+ygKmeQCs9LmX8I3yTOj
gK/C61DE+ik1aWDGgarTbYkvprxNPjF9NrCkU15kvj8dua1NwjhGNGNCMUD4YiHMq9CSsGALlbR/
W3dU2JGigERnvbSKJYjmX66qitn/7VlDhvDPBOEGE1bQKZPV4gjs+KCwVdYimYusyP0a99d1/fWM
v9llvpsVO1BXR03+PQI3kvbLdfhWJ/e2QQ2BxKvjOhT9oXhsSQ6TZcKj3Hs8s9YjE+q2K++9oooK
NhFflRlEj4foOskbBsEzhTGcSJidXorSQcN4mFCwBgPQ75/dXSJ37/gQbVIZ2xiAHzuFzws/rXT4
WqqJFX6V8KWB5JhkXQurnfgayQ5P6171ClTL6gXbomRzJprhHpufEyjbohB01EM/ZOYoIktfOTSi
zkP5BLF8Xdvd4plObr04RDmTfyjbX6j1r1/M+1In7Jz5ur26VxL77ZFK4KJ5r5i+HtfGqoW9BkK5
sBi8MNqcJx/XlKdqNDiVhRiIXvfyOoOgao0gLhb0wqoVqlTp5jC/S4Gg3RcpVDB/vBzT5WyE0kmZ
/aRV5xxI3QZmDuBN2YTmMYRFEgOE7mFvPoOAzpdDqI2kbhNPNQtUYrQGnjClDRftryH02+w1Xvsc
0jzAjuYEotOmE/9N5R1Ofo/iXztIqlMiiZAcFrqGH6+GIzT/rnjlLfIZY6RKKLf9PTdY2A2Fi3kT
dAk+GODxq1eorg7vhldb0nkBoodRmSk7MrvaNEKM+CIYvSsahsAVa/1AMC9ZSGTD5o7OOg+fz+K4
AhR1bEz0lDxRM5DMOIejLTcLZEiKAbXzVupRSl8I6IcD8T1eaB70yte0zZ48RvMu11M7/Ikuw3e6
mKLHhMNqNnJCGgRXIpNt1g1gYg0DCEaColsIoDPFyuVvmrMI+b/Gjq23Kgt7Vh+AAk1ooSfohv+b
Q1wh1E8ta/aPQht7V9nKaEDPWVCICuP5I37uhsGEYznD989nbOTAlC4ZYBnCzScUOG8LvG18aL2O
yNRMSIp18qxdNVO8GMmP5/m897XobAGyijF/i8bppxxXIZgqoItylerTYPOBpBp9bHrknP+RfaFK
1jeS+cdj4qrahV1Jv+/LXGIgqV/dR3fG71e4V506oMV0kdoRbGp57cjamnZ7ZMOQMH0lspDgnDzh
oR6ngsrEuRoPT9z038jtoGMWt6iUCovaUYZdPN7EIt7+4foAlj45PCY5AMDyei1okPyRJeMtTEGF
on7zT3pMzDmKmeml0mRPGKgeP5TEYRrYbbtAEV2UZmho2+swvm+93TkzO3d74mtUMHn9cAC6TF8E
iPi1Y2tpSgUBpctgmKucoYDEQAaDSz/otNpZx5z7EEraK6x+OmA1dW9J/xgQo2DK9AUAsXvgbAFt
6JGPwWUeQ8xU3BFD/50SaZJpKtSY4d48ltjuxqbnE+hAwXYW/z1E6mWzftl6z7KWACIP5+u3iG50
5IHVrWP2IXszAIHPy2d1fcsK3WIbqA0OeUfvZnUXT4VU6xqToSj6bLONcq8diMt4tTJK8hUkqmki
T/Dv3nUFEMHLt7HMGyI1haXIUGXJ1im7F5RCp6e27e/PJzWKOMXPsL0yRYEdrUNIfdThWBTBlFtD
LN59VxMpMY7d/QZ2rIzbhxhnjnHXL9DpkcGlN5tS6lejcg53OeYO5tslPFPdbVZ+AlMIPCLJP7c5
6dyyAff2xk8Rz4nYEifxD0vkFOgyaJcYbc10/nBtoZYo0SMPsH1AKkYe7LwJy1ytdP5atoSM7U5Q
wt58qHSED48XiG4NJfyJOLNTt+AXabctkfaWQdvpzaPvhAiJa9hy6HiRiRFTixHXhdSoiI132+5u
ASM1EEXHFhlAse2szIncV7sc/cYBiwQlnDreQ9eycI35/XLd28ig/LlRiuf7L/dnmflp+W6slrya
hYep6Fju9hmMH7glwYTb14r35xHYSr3vh0rCvXHfvY8UCaHCaa2xNRqQlozEuAOMA7sJoHjStMLk
XawT1Qn3zmCpJc1savW02eXf0ZpQX+GPX2BKEoygsYlLOvltimnjrcSleY4YgigdNwqLo0hFxn/8
W0OsfBaVzRuxFUljDs7vSdh1yh9krOGr8unzD0G0WKCMXULYy45x9nJ9oL23XHEtsFee6+wKOYwi
qSMBOf/bmoIIwnV+Op+usVW+e0f8aHy88QYfY98t1hNZC5ocOt4F6/D6HpKGCKNpoeq3SBvaAJCi
ZHSF+0TKon9/Q2csU5UDu0qSb1LdXwF1A+Vkl+kFZKJcfSm9uLjLXObA9Dd0w20bpDwQVQyJDxpC
hBuKhRIIkJHwB6ffY6uILKlNmSdIz+6fdM2oCFlqk8FDfEHUzPwAehU5XntoxJpAQjMenM733p47
nFgGzlysZmIonwQMnllM0OX/SMljjpSsfcdA0RO3Ph7QNHw2VKu3AdxFw2hau4VYt1HwE86nr4DX
M6WTlVpBl/c/0PzNoZ1EqGRB0Dx2K5Wb415pGe2wW6ErhiBaY02c9Wqj7s2V+PFttahF5kcL5/oE
nNi9OyCvOFZZ8zIqU1aezJk1TreN2n4ON0j6Qpovrq73Q2L+Jk2b+ZCjz8nHJkZPBWCeuvbIV5M5
JTE7BoQgLPvRwBxjOdRHbPIxnvqkkOyUufQHoqREDyLIHyeDLO/Oq1elW1bLRmX+V3XjOUeTI0AM
hoq6B2YkJCbsJYmiEMBp/idoHhnku+93bNE/g8dt3O9necdXTKgde7OtgTHv6y030tjzr2jbF/+S
m4fqwtLxkZ7ntKhucqJwcVsWscgQ1amVwYRH//BhENG82GEDqwuFxiT7ib6BTe66amBAGx6N/8qM
YaIDDt2HkiOj7VvOnhoM4M5WfaTvANSnWLoz+GYB9xX/ewXSfPDvjzsVyM2dLCnVELGEHbNI6R0s
wlSn9irwruzEgOv/mcUYkbXQ4RdrPucj4Yh86U0kJ4FeO+pf0XPl6IRPbLLg5AqoRXmbV1ScePHE
YL1vqLpPOCw7HV6E4giVB4YzZbh75sI1D5yZ5eI3UwBMz8bv0JaLyDCg3vsmVjF5J8m4dzjrRMtG
JdCcvEowNQjz+vpFMQvGg11NCQsPBmbEwdfvbbdBFOq3vLrQwKQMky+YY779IhiUoltbk04TWSA4
Im+K2Ys1oMp+TnwEd4kZ1MJg+V16lqd5hxhUyl/Vmu2Fq3v6nsFjKJz89kppg6kuh/YIMc5hecgU
IojugMjZy9oZxj/Sux+YpCpYw4m8/giWy9v16lMv5Zz7RkeUt1YrOWnmXdcuE6J0l3/REXaOSpDp
iPAuTJtStcUqKl11Z+uofdvA1rmqkb4V1f+1ttvLmIpDugOoUv6UCqN+mjrHxQ0KqhTtYVtNJE5A
shn1bVy+MgC5BHBCst4/w3tTWDFIjVGEvlCdxuqFY6pTxs4XkhgBOfv7aAEcq9EM4wbQm6/tAFui
gkQLYuon5W7ziNNTfrGjNzY7wA6bKgpcDANIxXE6vM3ObNkP4zURJmuzymVEp3IpB+IUith4Hco3
3vak2bUsNOH8nQ4b3xZ9pd4CuqUJJtU3jk+0yd2uGbXGENh799ah4IsORL0+3Hbob0tEKG6aPpcU
4Xxu92U+pr6iSivpa0PSEOyGRXiQes6xEExfktBlwkI6mv6o8rTe3o2t7R6Iu+Bi5bXR4hWufwmv
T+AjUVYhuF2l3gmJAyyhUOIMRtvUesRyybQ1ZBVLg4x3LQrVDrmO61pDlGRHXOld2Ly1z3HJgFh8
Bhyd4kiJPLwtFdLNB0IOSELB806El+Ei2plR8JMzZMMesfolLLM30Druvl3yEhumc9P9orHMoarD
wc3cbkJU2AYuh3uXxu3Rddm+0gQINv6u4WHiX0G0Iu7BiYIjTx+F7/SII6ZHXOaHu9C3XVmNcM68
z5vTTVhCz1ZyRsFNhNnN8vBE0x69E5Yd0PlCNb9O35tJF4bftoZDUdnr6iPgwDSGkb7MVYxHVVIH
rt+1blGjDCQKqRixuLd44e++Fn95fgW0LZtMyf8y5kmA0KxXH0jVRjktKELE+NMsgd6/LC1Cf3Bu
0Uujv5UkRu/hCKLTjMZpmsN1YojMZ7M3AhOr60mpt4DBRFO0vxCqI7vz8f+m0DeFW3j2R/ynJwbN
36V2WYvSjA6ktKnjxhv+erZ/bBS3cien+qgnOhYwCiHcz4ttMkP+bI2MLZA42hpq05pwW+5Vwi+t
BpKmwyObU7nw4Sz/qWap+0OyMyDaWq9AXKvN5LxfxESYzfYtrVwck7uURPcLESxmB2G1ZxVubXDD
TxNxfTBs98zXL2eeMfHcU6uYnHwhjbmYGO9dEEr5AqBrP7wAYrKEm0ucOE7nH+pNa1692Wk9Xgkb
Xogb72Z8MVQlzM2uqol8wb2dmssFUVVa8ZqYeUso4fSNO52NdnK3KEP8quSjlrogEJaNk9ZItk8o
Sy8AHjrIFMbkjVpLd1kXzLRjFKKomYenBOyIvFfaCPY1xuXOSjOnfsg0cDEgAEZB/MTyyawMvaAG
m/3NucMopZwM9OK6NTw+wxYj/fj0R1Tc/lbe34K+8Qmtlptm9D/IvMpnU1RHoWOS/1GKlii4vP9N
Thf7QfGTgjSskw9n4vUvenDnIzqUgcF3AYtxdmze689KXZyawe44j1D3HAqjaMpwoZRwiSKi9Xrt
M3Xz/eVYPWUHp+JbGQVIX5ftVmDu99tgUYPb6AwVfeK9dA2hy0g4en7BBcgCsSNGgLXYwaozQH2M
zg9wJqLTkkW/NMXR+xT34beKrpGXjdrp6fIQppAEdYNQh3aol6+K9sxLw+v4qhP4JNhn/awLnPfT
0dJ2raC/+cUy5t403RnxELHRSAGlChZBYR1IRMOuiyxG40i7QO8Z8OtnsnQ3zFtsayZ1Sc/QxBxd
O/31EgI5+TbbjTSVQ2357MSgS6iYXNE1Pq7JzIW+Qhj3IwgiOo7TbG90qY0EdObY/FzZNql+Z8Rx
WFpYGjOKWikRxA8i4wmggBhzzmbjn7y5ZGL+xxGb1Pgov9xI3K9rFb8klMSsN/KxCpvbPZcY9l1S
dPw1cYkzrcLYEbeXlf0R89xdNyR6QyOwMM+ITB6E8jcmHpJ/5tW+K66+PHWdrVUlPofYt1nSJDVf
ydZkWyfRrwuvhiWfUqnSvmhym/7GE4plmkYqI+L81D2/1T6VXhz05mXiIHsostRifikqb+JqAOq4
qzztKWpCnv06Y5Uveivv4Cgryg2SNnXrjfxzvUEFjtpvIKafI2fBSbf5vqvgu8tUOrIbBYUJHw3O
HPGETDxjsCXcxkYn0m0OMV0/tBanc8vMQnSPUP43Q4OG8eiLaFi2ddUbC29h7q+nC789jwGRlyr8
KH4YZUKU9LUCYYfoUeo4cWxeJ1OaNr6ff5JK1ms3UGIJTJAX2DCvZ+1IlP0oH00oJY54u+ZM5mso
0puk+IYnTTWMg5N7RRsNi8dEXydQo9OoUuVMAW3eXGkzoQVyhDaL4HHK8IpPC5F3HnIZicijGj8/
MrEGqHszZWtuzdwXE1JPzvtKzTJeUR31/HgpKYHS4dUPK5mdQTt6KqApEJqfMBuHiX6/1vh86sqj
CselKKi/ydNz6gHGSVtWmidvEev/53bQVjyoyId79c//P+tze75hS5r8gZL+KXGSOWTKG43gbEDK
uH4ody3VYqisugNMeYitSI77ZWI/DsJgy5cEfQAIZ2Qx0WSNdlrMcL8gKBntmWEjdI1TS74FeH1g
ltQNdBrJ5shz9g7TU+sMbHrbIhKR75LbpvmBcOPy+GXQQ939sZdpQqccyKrRLIg/nvbNVsj07oco
6V0BhXv2V5bTGVH+OW3SC0ecyXK0OvEA0TwscyMcZ2K1edyRqAihQc0wu4zDRfxh2VJao/4ycsVH
HnTgVfKVHhKgAmSZsJCtJLBQ4iAiL/Q4wuObMmvR/n7bO9772c1aLYjcbNA6HgyKKCtf3ZM36fFx
X4t6Qbs3c3JGd/7sekXoyDV4EVnsgD9paUgn7N0FcH7lImx0pU/s4Jxac+e4imXRA+PnC+Rafmvm
5sz9fsZJV/uQav9Ua99oeDFuCViDRP3KJg+YDi0Nuatq99FreDDeaUA9OG6DSF5r3XJNGOk89KXS
zSVgVRFJ4aDvm463SoYtsLXOPTQP6St6cCT7UdexdBXcSeGI9IO5OtQLZyxTPHcfdwvgYtrhSPao
l6r9JOu2bdqn+XwE7XTZPTB+I8Gvk0O3RmHxh7fjbpjmrUaA26E9W9IuOapdqYO/Zj9/NVMfROPV
w98vMRVJC7eu4re0G0nq4DzeMlQttU0xHbL3y4RzL1wuY/fEdg215NPK//Z2wHVh8itv3ZWtSiF2
9j2lteW6+D1G4cYhefToTAqzLtTBcYel8wj43WxQqkCmtG8fRZBH81Jeuwa0BMA1Lvi2G7IzRmYW
VkuQyX6noQMOHvye1KgPgGkjjnmYUToZIUBgOIuSWI6tItlpvWyMkiv6Igi+WCSy8svJfrbxe1Wd
IcQQnor1/5Xt8IKgIQBaQVU0SwPaPItcHFhjhBQ/DPAI+yRW5fAEq4PCKK4BCZxeur6r3gzVN5f0
8+ZAhYB/GxG2lwy4Q9sgKNNoesP+1H0AHrJmn0eDqFagmPkDmut+1d/HC0UQJbhohYL//P1LzKwa
eeJzNQy86H5wlVqyl63F8vr05niCB9N5R9hrSSQTcy+Tame9gSHVXsBJkzLFxbDrcWHIn1hrYddU
if7TOeobwFEjV1AyaQXxyhWUJZSfemQSc9cFc/G4bS8p4cdRK1YYMmHCjgkbpPj/5Z+FwItpbDQc
bwiNFIC49U+ZdCx+YNm9K/Bh7Sx0jBxkKd4ZtNcjnWruIc4IjsAk73iWaHyceQJifp2VNA/F5/mQ
rdoq0fC+rgUuHkV/V4GbO9Qjmrktovz4jXlNAphYqaf/Scb/KfmVTRPfr5bWPYxxCnDOlur6W+lu
Bh2i3R9tWTHQce3xFMLaKkliZSPSgo1AfH3gmSQDwB2F0rdsACATv7Wfcb7jPvdsA187JPn3L6Mu
gQXPxSMu+mwwYFyCH1SQ/FqFjxrBSZICdI7k8XKvbrFXXPdCm/8RNAWnICLSMcabsuhZ7C4TkAOB
y/z7ardGFdnpNBNKj/6wxbtUmqvQbmWrrMplzqG2o1jBZ4Nil5WuB+ZTetKv8ES06NrrbrbWOuXW
r4AxaEET2qbZT9kNAciF0hxxRvDR5WpEeHFK4qAq4IKibVR4e6QEl/7ymbnwxSbFTnTfPtHPhvjb
iDw1Gtb2U/EUHXPUOvBKyE+BH1yeJSNWzBSaunSM6Tw4PMG6J8rFMubS3OMAdNbs0UnvJ063uKs7
LUkGtsrd6z7GrB34dJfPGgloq5Envio6ezul6XNQVrPOs8WNtbdeYG/4tqACgmTCMeAxFljJJbwZ
wMQmrs9QCEfeEtXKztmjvcWFv3juyZPavwqHYZwpO2VdmTj0VEC0liq/0VozUWKZhhfkKesQBGOt
+qNMMXSgfGAeYuWudUP+DBgyUESxVuwkGqhMSTwUSxTCoPiZNRPjEzFM2m/qk3+bo1MUvyROxl41
W4GgEtIbPf0+iGyw6QbAlH99Kn7cpQ6GRjDG/2lqD2d94+BLrdDlOKwUSPU32WoOswMwhYAqXCrZ
7PBJF3c5TZM5pVFHifa4H2r32WEWlUA/XDUB+rvPPZzSxvdTvG+zXtXj4jByjxbWIQos4DIaM1f7
X/+a5Huwkdcol+RcBBpeN2FZfiRoS2+6UYSkfUIbjRXotTfH9mbCtY879oi7zPdcq1DEudJF0eXn
eRpwRRZip/PHLwhIume/0warwu3HfxyPBV9G/i19BihHHI9Or80SzyQLgBBJ9C8ZzCUGMIjzX/9T
PGrYUtaDCRhNRbiph2HXFFlMW8iOYOqSyYwpAufTHORVMcF1r8I1VDbsDru+KbpEqW5sVxSX5iv0
vnCXz7+EZ3JOt90k3z+waYxcHpoKcVYNw+bnZ4ukYI8yTivAo4ZtBWi0bCzNduSyy1qjDGuLLiWQ
oZqNdnIu2JAqHLur7VpMRzGRP6HzEWO7hnUZ7RjUyc3gzQR1vT/RFKWDCkJN3kAV+AdgO/HWxwwS
ty0mGVbRtW3gisEbMaaVErzT8J646lIx8KjY7yRzHFbX6L2+zyA/LZU3lnHFnnnomx3+OvgqQPPC
i5VBc402PILK7nwiJP8U1XaTDkbwnP+i+nSLs5KZvzsQlWPZQ/+ZBHZGsDeEBRxoTJx+uCr6USot
X/3qUAkbKOz6lLrIRsLNg5hN5KsLRxpSwDOXxlw49yEcKv4NCB618SQxWOX4hYl2N1I9SWry6E5O
ZE1FeU61qI4IVLixKWcS8i8UumNN+X8XP1rXgxZNepRFfpLxQA6x6sYftYcv88Faq1yuT0oljIvM
sfcdmsWzlUg8cb4ni5kVSQVflDh2a47zzbkT3mNXL9mhV8Cietjou+LkMolz8wJvh2oORKZ1DmwW
MU9N6MFBaCehc4jtKOh40RJggof3q8zw3Ny86g9kS6sLlD2yBhrVrjf/MGF6hd62t6E6nsZD/Pd0
Zhp9j0SIoTOJGl4ldshlyDxFMdieCaKbGXUGC7fUYu9j/p1MiVQ8DC0VIOBpANS87Lk1WjbWr/qV
fBFIcegyjFAeFCjXJwUw4GTXRIR13uh5EbBfMHfd0xEwoEbQe5QuxnWTuDOfZTJkEkRHDRPChDd1
x8xWFM3xgL/az0iFWumwmshzmXGFFR8xXgpF5LJKVrFuuGOeTdVkFjzhIu5clokXRpSPzn31wc/N
1IkFTrU4OL2s/1kTgb0L/TrTzkpnqpn8e24mKY53LrOWm+dqNd9Ai/cMHuYVCI8qp7OwJr+yLpgd
7Q/kk4/p6DZqkzyo/Q7bMOiYrSwwVL1QLgmYDeH2871yXmlmmiHsqSSdKp0BH/yccNCGlh5VgenX
96HvLqo/Iw43o17CZktFHv33CUKh1611BprBZpwgMe2eHocLWr8g6bSyh/FKVdVJPfOlCKYT6uwv
Zd0S+tg9h+B9BeGWOlg74fb1cq0TevrgfW8a+64FLUwYyZi8S7rDVF/Ku86ujLnGQfkgaUXl0m7R
4dbUVOPjRZDmZ6EDhJIBMHkcCDKzvfAE2Dll6MRW5r3vI7H+Esolt6Fri0HmEcMxZGejCbIIBNSH
qIfINh2IMd6V+ybG492N7SVOC4qp1DoEoXIf/mPoaMwV5g/0otbXwnC6yNaGFyF0em7wSZ0Hps32
6BHP6obl9jyz8Ttz0yf7aIaQOMCzGNY7d1RFmuPeoZ4/FeQWcBZgWRWA+FnD4WzDCFYUGLWfDx9m
i+H6QzK3aqIr/jtUIzYiSh1oPbQiAhc50ZUyaIcVv5syFKgF0RWe4lV6ws7lJUQ9fXNmrryw5wYn
s2H5dFQoATRw7gKHE6QmLh0V5tmZxiAnoNbMbgvWC9D2KgOKDQfXNxlIjDTRIm65Ecv8oTQr66PM
UgERDTgL85mf5U/d5LP2WFHLhtq8ZvbmAOSVcZhm3S820abS1+yIV2T2tysKLe1tm14oE1gDtTq7
nFrx7kqxD6xtqjF0Lq6zomq68hzZo+ox5Pm6b/F/72PhxPt6OiPV+NbshwOia49UtEooejibc1OD
oTk2ev8mvnVa1qIr8VIlrn5XSGu3fJ/Hl6QwZUaV+pfxeia7HcLirClC8FSGQU7kaStMH3BUj1si
0JlGIAJLXUdp+hOOQAeJjp0/rRXWR7iQNCFHsrOL5ANAGSHdWvjwT82nbIhAZcQi7go0vB3ivNBA
iWge7d1TvN26Zx4McFxdYJd38mBzYlfKr/JSnsbh0hHFQhy3F/LI09LaXcrTllqtZK5TeoR+YAIJ
qvFHLEPilxyYtwfiWye0vC7kgoWZRw5jGGYuGNDVkKUaVlRch1dVFPZkpR5NXM/dDASqDhDBOaIw
2aQIAITNF+X/gNFfNR4jQGjqBvAPeq8BBbNDr2gk3PP+xEF8GRdpYa7gesvoo2dePlhwkGspeGLe
YpGWdQJPSDukkLrd2WP5kM8+g9cVZTaDBAwJuevm+cOf8yU9w2k0z34woR3Ksny0CEeFOoxFJLXq
gWwHsDw+ITVIGp+yBk+baiicAeUSTMNql4ha9CrCD3er2eXKIhQRDzGapKRVkW8lmQwCAIgg/PSB
G0eTIAuowrDpttUXDpL1kPaxScfTRbENrhkiy2OY555liDHWWg+ye3v0JPX9GccgMdP06pNWPnFY
ueAY/o5d4suDFjVoN0n7CpQUoI21517hCiq0QkvnkNst9BnbJp1NSWC2McagKD1sQ/6y3YWFqLKh
xFn/yhHq8j/BDvVtp6ky7DMBs/XbfKyhGocSbniCZ7c7I1iCn7gfGLHQNiP3bm1UIXmupP2C3v28
u1Ayj95Yq6tgXhA4271CLge1AU/MwZSWjIstZcDNLvT/kDWrBvEQB6XgO09jIWWENZVS9hCGcbFi
NSNM7rBRQWELU2Ge/yN/iQhG5yiNMAegsLIgaTpU9OQWE7aC2TmWY312pJ+dlPmlDe6Mcbp+FFNN
ztQdihz9+aOEg/dG4J5K7MoHzZJyoivj3fZObHceN282TS7ZnW/F9NQg9zhHeePNEYXqLoIo60O2
Tj0+gL6bp2ZeWcNy1zinWi+nLXiyUjGAnkHl8YEE1+/LihlkK34KjU82VIzO+7sPDboj81J93D13
SvYcwW6v4fh9xUYvDwXHcRXya9AvVj5ZRqEm47LCkQ46wTxiDjGXH/O2u1cxlfIDoRtgdirZexRR
FLgLz5u6z7J5HhWggkY7GoRgw2PhE3t8p8RDwbwhR/UBs9t/OlcPy0jmJwY6Yl8QbcZCyA0nlu9w
yeQqNjylRt6rXDx0r8A50KUkFXrDnMAM4RwmP9+ZGX+uAGJiLpwB3OdSv8H+3hd/Rp5RUyWMW7yn
os/H84d3WMzdBLaP6P7xE7RKQvt+QpIzHD4E4+BVhOYkJZhtrwswyNRZqqGOWD0rGqloz743w5nU
2liwb7nSxwwRAuS0wcGDJ7svqBzfugL2GlAdm2a/RB+WGerdqXnMWPxoHwM7GjO+NaegT2nrGCO4
x3DRECDOUNKrcWRNl9eheitxdUV9Oz4G0R4YTTR4PDrlomDGZ0SPWSt/HV8a0xaBOEvxwUIOqj19
HeENO3H5z+tXDW2XeJC9yBbtyc7XuA4FooIqjG/kEbkhTPzBLeIvCKCweYWTuQNlY3hzbttiqOCe
Gqp6gkxRlFokeyQIHKqdYmRqfyI4aG2H/1hSayMlP9FVK+R6UVH6JXC33cmgvNHG24cKIqNsO9M5
s/nR1niQFRGf0pgO63b1IXO9dW4opsmVGYfsndI2hStJCiDSKrMF7OP22ZAEHg5cpEQsjebnv0ZR
4LVfIbKWO/t08xQmDkRWzOzUuWLqDbTgWUjiIEUY/E7SNwJN/558BsRa0txMn4kHM4P/oX2HpuvG
ZPeYVb3kGbTud9AnDi8+XnFvBu3zk9DgupbzvLmbM3UpXdAwAqcpaJ3Ohq54k884b6WTTIMCFiZs
rrAdksAskTofZCl3VLQQT/E/GeJMV6O324XwG/Vtw8tmUYvR0J+2cHvqNioHSVmlQ5zwo/lYpsJF
2TRQLE81YNmw8pDdobw/a6jnEsYGQsTodYyYekhrNLIm/9TSSmDFIAzRrz1O1L+ASnJTEL8OFmJn
NELNmNaKfiKDOeBpFZVQgZrAzoSZvlONv59mBp0YMUFG+wwubS6895Boae2NNXzxd3ROllkIZ2fh
EpTCRgKiCOUTa1xxDW+K48SS9uk0z5fd+ADDUwcvvPYyGdRoraLo9Ydzn/e7tr0HFjUj/f+SNhBi
ziXqb+M5gtnpDbwIs7YtnPLzk6P7+9XrHEc+fRMIyyWHRiM2+Rvjjvn5AlbiW1be5VYtw6EBV9n3
XNfXwn/7yGofvN+mNQd+i3qJx1VicGKszvg7slduCdv/x5MT3a3/cyN5tvVMX6zTvNXYPzjXUt5F
wEp7Hdni9yFJOLZq63XfTTqA4XKv1Nm9FgylzS+6JiX4OJ+pLGOv7ObNRGQlH959FYyEijsYGr0e
UNPJCTnUJid3h1aj4gDNZfVT66j9Mt+GA73aUKIiMYcvbfFmh52Hy0MP1bSbi/PXw56u4HAOzR7R
wP10rc8cEHtYnl6W2pVdjY4chPVoPfXu2MULtuxtgOAZ+67UB0P+JwzZHxLmdNA9uZ1xU547YOyL
vLON2YBWbSCrRR7/sHzsuuEgDwiBoGKPDHtvZ21yCe1pqZRC6KwRIMb4UyoccpKrsrCJkgYs9p4k
7YRz8YekPpNeMi/oqHuXLFf2zVz1MbD74GH3udXc9YSVWd/BWM3FRXm9bApdEx81tCep4wIvaJNP
lAXNmqv3r2y8iXjq2X+Qt17UR4o0cO9zfEB4bYBHSMKUpnEKrJdkFuXJQsdPvg6ylv7ahVbkIuZp
KJt/7Qppg+fVsJ+3PvgpQcCxqP4HXP7CRakTlPbEzMnK4DdJwB8Rkl61uCIAbnD8PEXjVu3eqq1o
/xxwy5rV6qqzZhJlylw2bPHb1270h+4oLtJeQfN+m4FNISPBv/QkXBADozFFKqH6ov2e+aAQX6gn
f1x903eZNXwl+gHNJDFv8TR3149OnaAhsE3rLXNBGQk8bjUCdwTlZatrZQXkIv8GM0T76Zoj6rsK
oDVtG1kzAW6qWFjo0HbGWGss4WCSLNZZm7vCgVj2EkFxkimiB6GnYqGVRwmbTYY2Sc+eymUhGqAx
7S/FOsjn/PiH2TG1HHksBC1Kc+UkFH3Q+nngcC0/s6oU/T94OWjhN+R4uDTh/IBwHI7hwu/VNP1w
ElhhLEA6fMpmvAjPyiV5eBmAwFD/jWQODep5ZBINn8BRmVafmOlwCSo1PnMsnfsMQIw86nSYOl3p
/Kj0xQikRyEvxJNM8sJ8ftrgmuBEdCiBTZ7B5gvhVPy3Rf9EtsUIiWNiSwsC7GNyZUhz/WGG59Qo
lf7EMEVOIfJxMiSrDMFACKCyoAa10VCrYCN6lxFOJ7AwSPFY7m9biIE2NolfHT+Qltudcv7B9gkk
FHpadIJLCtskLLL47OluMVCpHnBx9ly3rcWHl9mFsicM6p5Uu2auwUMf9bN6/+QyvqDTERXv1Arn
BDJJfV0rZg6Ip5COoYZNGTFxThYzHZI6rVCxBstR2fHnuLul6DlM8mu667SsUCNIGViFtF9N0b7F
D823zdOGuZ28EszLfjXlRYqfbZlc6Aakcv9dka3h0POvSoChl5oU1RQLo94li6sgyRMmMcDVgFWF
Ay4fHEz5iRX5zXBXxnsdiXOfY2N/b5PKx/LjAFHBUs8lfCA+XGdb7eytR7CTpYudPBsBZ19vkqd5
mBI7gJe6nRvwjdSpbgczTHJ4ldUwvvUHFLfVH4wUMXfbEZPXf5tBgUlmw7F3jkMzlGmsM63iirDe
IIDgQU752c0DHQPE5EsrQih44L1Cke5oOxQtLsoAweOS80Iay3RbYCbtnml9gq+J4y36vo3wENGp
VdC4+w1HuG1oj1WCoYbN51vnlJZ/AplH5Nnk0J5G1YRWwQ9gQwm+A7nzhN8e7zmpydpecwL7ZJkt
7/5t3L5Vis9z7NgC+zPo5WRJC9w8J8CIMeHUt1kUepyFoEeY4ougYEqjSrxm8MjUdjzrbOc4aLiM
f+of+L45WtBRaET4of8/hulMsELqtF3EqseSaVmondUh9wAiXdgX5+lbGFq63iRp9PUojfKUS9iP
8fDARx28xfB+NBZL+3lyjTuA37QCUzVLyZ6E6aJLENWFr0/LS8aKcyc58UPeDF699gfT5aXRVwHj
ebRxLaabtLSII49z7KqoSjS0g45sx4AurrXoiE0XY6PahIGZPVuupRF/fmk4cz7Ly4Tqm55vB+TG
o68SNT/LdZ7LU9UzN8ze6Y4FOMMmifBE+UryNPHzTtAnLhWHdWrIZVuhBJfn+F6vmRPze/iXsqeN
fVadMFo8Hi3uzg0qoVsjmXh5j2jre0Yh+oY8NWgvI0bO+oEiOz8KP4ArE0EMMB4p4/ZYk1miOlJH
pBII8gA3p/gMkDYgcMTu0fOsh33IrpvDnTpvLfv4rpIBLDgEn+s4kTCZo2gKiXTsqzX1WsC75upc
diItlzIhxGtojTVZNU+2klFLQrEKe5vOvMMZWyXAiE4hgCoBQ49bU34tqEdUF/cLTpBnpfK3Qh/W
agmdwClAAOktCXSIE+/Cg13wyxDY4l03QFdbLaD87fMmBNO2Ljb1AvNSLdT9WjhiQFpDhytPK7RS
eXwDD0O8ZCFnH+naZMqbvPen2+r/Y6iqlIN270iqrfJDGzsKG1oschWwhehJiwWbmDu209LVlH0U
jXYbd5QKDAtsZwHNx8gVDkmz3xRrYyDtNgLv2kF4BAEa2IOn7tpeNWB85QiU4PgI6lJicXQfW1CW
i5jq/Xp9aKzigUcKtm8+r+p1pxlNLfzHx4QDV3m03ACRiOIGMY+WVnhS8iQZBP5w9kjhCs1SHumq
YXj5V/NCNQMgRw/QDjo5KyatVcpddIdldT/0en+2soH4zA+byj3W4OrKQg2/l7UesUwk2aD/qwEk
njvVJ411HsSaGb0FbgiGQ4bLhno3kjlGgEAfOoGfwtn6c8+cL+v7xPj7HIJdR7M4M4xNPXhkD9gX
ncqNJNuMezESd3zzFhCup5EkUzjvgvPCKtzA7vTIPchkibS5G4nrlxu9/W68aLX4xy1t4eYMlZcL
OiWquiJDsBklJUv4CC+IwVV3tl+T2wZuPRM3EA3JtS9QRTusRZ5+3r/r9j3FXPOtDcv7SN+XKSra
QqFcYGAfmBc3u80jIccV9TB8wL/UFS7xag/VWwPpxwfbtwqntIq8aKns33WRqwfXYxrwwZ38DnNK
rbC50nWwh23OKKDl9lBojC19Hu51Gk3NbXjKWxMrlcSBSFUluiOrLoD7qqxh92NqpjH9MLDuprY7
kjMSNM/FBwoiadQ6jL7bSHD/sCKEJvDBeFoFWygkZHjdS0SOXpnkcr+gh1xz0J19EfgvBlUCo9ue
ukfqYXOTVLZrtygxPJBiF5LX9rF1BhWbfCfwnmySiAsWnkYP2YEHU1uEDcKrPcBGWKa28t1aIG41
BthhxacbwRbNHHBKhNdmFuzG147wiFpW/YwZRroE6BAUr1oblBx4TMCq6vypzQ/Qm0RLUU8s283v
mAA9CqR9ZP3itdDbUXVhJezbCQocG1iCsjYq0dpQrP5yge8webMvPG5MmM2JNB5U/mOBxJyoKvKn
aJ1VicQqb9d/LznkPTJMx/xUGbiJgarn1wpZPur/l6uqczaS67xDanMaBzgBLrVlDBhTzJPEbvd9
0O5NzdxzTF+lqgutrSK1zRvULC1mjqM8lD0XaMnoxuTLgbpACwgsIHE+XP81fg5TFNCy3ItGNOnz
Q4sRHNEb2eEaiK7FMTkAClnVMkw0jtkZAaA67e/hu/tN9zWL/kvszNZ/DZJBA6GsBIp0JasproAa
EWStFd5xYcpAjkD+AWGKLgmWJe44uOJOj1q6oTZ4qf8KY4iJ5sdyF/tS/5rEbZYAIT4G3ymcTU2L
fGqeVnyPWK8fD94Vyaapjhx2k++qiFUs2VPfXKFM9pXsJVf4O+/aLxnealeKCxVV785ksWTEj+A0
u4D19CAJMCX9grGz/WUJzHIq+LMTSqDxgsWHPRv+lA0RIJ+iSwd0Tlgwr9usJFLy+26xQo23IiIT
Iv6BRCCbvRH5eeDfrBKNESMCHdgZoVw8PSBjFhGG2tPa9NDIY0Z/8/oh3TEZtIQjrMFJaJxdhBNj
p+KAgTsa17GDvdFxghSp9prWK1dl7BF4gB7Ej2IWlfdyPqwGakNyJjVFdd9bl3thO6bjBSH2E2yz
ywwkaEhJjhAeYbVxvmhn03IIFGbxnlckH0bOfjYCfJLssTJ6p5rICrbg3FTUCovGXHg3wkx4UzLB
cx7atXxzsXS1zWPKSNpDT63WOSHOPdOFxZ7zluEroF2hTmvwlt5f6ySKuqQHH9Mcc8ZQ9PKcuUTz
C/JjuCE3O7hNIiONFU17mVO8dVZL8q4sCSHbYuHfAQliSI2Gfr8RcWMqJprHC0yC6yhfiZQ8FyMm
wdTa2UeXmxaMAtgJ5aWBloKJAc1Ep4f0lgdji5TsxclhhMVEgJpbIYGlygKyR+BfP08TxFHZbj9b
UMqxXRWxxhaiA4EGIXNNgakSUT1eDG9/b0bz0eZgrWv+t1wI+1OhpRggWHy33w1RTnxd+2+0C1PV
FM7PhVpsXRyxQt7t/Kh6437w3/xwvRbp88SkObe3+fSwD4I82NFvsNJ2yN1tgR+NOGLHG8ayDxsy
DK4Q5AOvGb1SoI9VDuRpizSXYQqmu53ZSLOkhO3kuR7wSxvFY5QF3zS2MSuRl6+D3s5k4BDucI6x
DCtAY3hq/NPSnPP7pyKJ6paWdw9rFZuzy6f15Cs9cxlAbhJYv1Xif5iOqKQA2xo5Q1uruqF74Vjp
xKke03Quoz6tx8Kk+yG7wpdtObUtsYeqvU4KTmL2KL0NOEg6F4UvLHkHEvfdAf+r3Wd+cMfAzpbK
VQA7p+aXKfOh9uG7/DV3e24Sx2KL7F+Ti/p0lgEeOwbGyxUGeho5WsPa/n12NhOAVZl7Tr3VYskb
3S7j/0okyoBVN90jwJc7CZ9pjZIKmFJxmyhOAcUMzXoxdiy0PS+ON9w8uX8bM5Rbmzi0VsJnQTDE
ZWaW63jWSXRZZSDjwTglOEP7+kFQKzIRTcw8yi+/1+huh5jS+ULFYLKPRss6ZaCJOS7B+xY72rDx
ra+RqWD2B5dCs61Yrwacm0beegQTBHL7VrvF3TzpT6yGfXZOQms35k32+H1mGJ2SYm8iMct+xHLd
nXn6EV7D4hthGSb5WtkU2KNSCBraqbhXfxQlv4UOSsc+klKITqjHFFRLCWYugSNxH6IKQKtSDoo2
N87hLQ7qTcYLv9cg0e6GUckvcdvc969tG5ztB2XsWutRZetqRQWcn3lN3Fral/qIvWSGmv1MK8dY
Q577GwWbspuSufgB1RvEYGvr8hSNHWXOo8QWQRf6tYHhZZlkluqjWNl677muUG90RzGIVKega9MB
CSL96Qiflrd/sG8R0YTjK9r6Kxo/0vKdU9P7uaKRKEb8TUt5Y6sjD2p+Q+EdQnBDqtQqyLzRAB1/
ONAGcxpazHtFFq7S10h4ZTRg6IOoG8v0f2/c3hOaMm+xt5qlfoXpzVpMHdtz2uhJdoQtOG6HX3yB
/Xs5oGnz2Nv/N/zQlYkViPCZix/3SxuJjEdbHFWsXesPMKOUN3hVng2h/OROiJb0jWdAu/QS8bMM
7czqKW3jOVaE9+ocnkgCqxyLllU2ALSkTMFQedwoVWkrV43XKPqbshrItCVFiaG73AMKxAeOPlAu
QZ8UXCQgb/USwkbv9apG6loh3LD2Bbq1ar4s9YM2Ib0fbsn572vDQ+/MQAu1HsWOB0tV782CjtgT
s7qMrWtUwjz0esCt/rTGJ+X7GaLPGYEAAGdGerIE+w4s13CfN15Fy7tNmaD9IF72UP4IRLRayeB4
rc9hoWebyJaW3MkYfGmhNjEColGoYf8OsT3mzWdTCZdLt9Evi8Pj83nCdIgNo1Gz2DhQM5/Eknwz
rvYzXkO4Dq82rdNs1+kwR44Rkx0cmh4zBar6/5/O0s1lSqFjpaVQry1XycrxCPQJa6wVb1bSrpNI
/E6cDIGCjfYO9S8+r7i5bMlZfmQI2k1QKdqni7FD7ubFim4V8blnRJEm9ygtjMQXdxUhNvBDcqNd
EZNE42u5ePQhShLXtLx/aAOD8wXwIo+edCtOsuRXZ+k/EBp5fxiRZ+13GljAE48u/BFkS2+B+fVG
oTzXUKhfRtwuErzG+cnu38/ETwKawkdAiZoxPlcFLDiqMcr8IJopmilxE9USZrSSg4DIu8vRzMHv
cuAZEnYdCKdkbw+sxDYjcN0k1jVModrGRa6GYEQqylHxNHy/bD2WSEoKc5h+6h/sgbPa/MhgQ4CM
HZjTGfwKMedTA7TWXL72WJ7FfnGIdH3GCSA2f79praSGYc8vG4lPD6CjB3EZJtEYXlFI0+SmD+pL
fjJK9ANkPD8GNQjgAATD0g1kEbaeXuH07+jfElo2TBf1pal8GCOzU+W1q3/Wn7YSyb8hXsBTWeQs
ZcE61wZHqiXKcnuS2uzuc1Eq9rzrhKo81hBHzVPSmtZ7ogI4N3eVEpCc/+hCsjNC2t8oal4446zq
Cvo5nhIB8Idna3+zU3UmNGM7w2Q8Dx8hms+a/z40BmZlm1rP1QTaUGbUHV8cxKzAxuYjgbQyjEvS
zUlqZeopftQvUGccKxfvjJkGEXHmvyXSHwFmVWo/0aDfiiYuUvRZqNgp+Rb3noWkpY7RAQDTUZYy
zzz6yfmd3/IJvrq41V15Q74rwR26Va5vxTJglAPeOw3hY3s7W4vV+I8YZdZpiPv/3ktwuYr6/OLj
h3G/ZemODz+BTe0ZxYbPzcuKJxoWSFpImJiK8ih8g/J0yylKICxcIiKbj9j7qHadVteZh/sd7ciZ
i3QWna3pal2LYOikRSiIghxFTibI2S4MBSqLf+d0bQfjDtDwT1V+U01tDkStB+oamBMsHCnyBRRn
P0FzqrS6DzeScr6PeliOy8B1yeS3Ddk1KHc1DYyZzPuPVJwAJ1GTRvhRh18NC0Pu3iihnW2SX/wC
lgchvfUnJ76hZbxOiH+DiW22Fgliup0hNxSVwFhlYj8gy1U8z8JBZkHOYXqksm/hlyXSqj/PODVO
BC0AZLp5T+HKRlT6S8VQ3J+E9f2Nc9gCjshmMpUyNb7Cik2RAme4WVLsKwy5+VPzD/IPdgMPbafR
pWi2AjFPRyWWsLxZPgRVYmhEUAY/HnJ9P+BsN//3SE5gQ6Laf312dX66zWrLlcp27ou8O3ZNafGy
38YoI2Nl1/xSWA31l15dxIkuBAoeZCayuWscCqC/P7+UzIclfxRE5Zj0a7zqXEhvxe1GTLBqtZtj
WIe7ydUKteewsnkRjWd/xNxfqPYGdUNOnHZcb1FO0Dj38rX9zwnb1g82oBE7KiMU9AQ0xveJvqXM
eH4AYgOXCSX60mHmwYUR+AvwCbIZeebRmulkknHTokN+4dUAK97i68etvnNDEC1Q7xQHR3mixi2X
tJOr0V7TUwd5FPZOi1YeQif7gIJ6GqSv2dkPixTH/A9qbcNG1srMWh6yHEqAAAMOS15ZcFvlJP95
/m6kLtqccnWHbOFwz8uhQ6fqO6/MiAxXxjg9HooFNEESxOkZQQhYOcnQULOL6+SvnHfiAqSMJ6g7
HzMlvqK81qlxWBBVB/N7UzIPK0lB5AE6Wc8pzMfI0fuLUOrAXPUwKqTNXolAwVBC3JUEOSHk0pBB
kURZAvbYup+1DbfIDGQXidRHEJ9DoKtAvi2DkzELT1qFVei+QzUNs9aBJdGPh3Cx2McghfHzKFMO
8WpjV16p121455jLaJOCi8QKzR/XM+JZwZLjnv2j8HlLTjsfrXcreHOl7oEtEBMQ6KsQqakEe+Qa
JO+8dSIbBIwtpvoDS9yBUW5S89P4aFJVe1oMcwp5BlO0W9+cqt84OGLrJFeI1dfYfgUhFtAEtlzv
okaZFrV8vz/iWX/YGcwhUBg28uxyyyMF3hmlf4tSusk84aatPI/rqjgyAgjl2gQRFs0Odel0jP/C
0AnKqAyGQoe84JrZmdyBo/PbW2KG81Rw4fhn/aDk5bfCE0Zb5XCjDlMJq7hjpS/EQYYgbqj3FB+E
GX2np46x3ELq3ApndnWk9jE3IYjZVoju8eX20EfDeixvd9UFHdH2mNuTVCEHHdht86SIm17dCzGb
hkRugQuh/JSYiKhgods1aLlU2kS6kruPUJAHGwmPLqi8hf+kZKEbJFW/002XQfz1L4LmL2gbpqdg
JOrOczA9CbhEf9C8EtpYcCUF1dOnYh1Ti+UMB0zXVO89BxKd7O3hcsF2HTxui5tIhqmTJU8NzoUQ
3ojM4Kk98y2YW9M9auuUkY9jF9Jy52G0488iR7Gzz5EPsiot40/iUnHVEgs60vxToG+w/SQKCc3t
nWu7+1EAej6p9WXFcqI72ayE2CFK+1JiVZA2HklJZN3q82JW31mUU2aTxi6dis07anMHZ93QaXK2
DRPrKfs48vYv72Aj1VESuM/KED9NtC6gFEG2WgQe59UkuSTPz4b0mOqb1Z3HtyYejEHffE1CMDsh
VRGxVlDAJrqWzkeLBFLUToF7i6/U3dnqlDZmAynhOHq40ge7VGmVG5eYugbkrrDHqHfKsF14qt7N
DBK0HHQ7Ah287V8dZvMHrH3Vgnbl3NiaxETFxnA7XxPClgGyeCKPeQV3WnN6NAWuN0o/+VXmdKoD
xrQUcKVjniMXSt3Rp9SkZXTMlUI/IuigBW708NXLDH4xuxu4ugIGVNE6TuHFv6TKi+YA3YfI/iiV
r8H6RJjPKurp18GMzva1R17bVqOEPWOyoqFo8SW9pRzifcDKHP0kX9g6AlLWjeeAj9sJBNE/N1Fh
WMZcCIGzJn1O6y/Kja0fXYrB15JGqnEf61eW4Sbkm/XcxG9485YeI7u1wM9NrQHSHFaDv+wKG16o
txaVMtSELrd61Dig/CuoliQISDhUg8b5Y39P/YbpbDgpmU8EN/y4RaC0+1WF01DgsjgtuQCLcnEC
nrynIqJ+o9FUMySafuo9fi/ofmqIkPGwFpnc6kZWwrhRAkkKwCnHn39kunnV1vT6bUHnvGqZ0ZiR
4izphPeGpJ/YynGcDypI25LnavSOTsHoOQS3tNgNBbru2xkXGxd2SAL9JeccpekOXehwVwbqXngw
oFWzNzQPYaVNKDQnE/74p3MiRSznLdbBmSTaDDSqUtHYpMS8RGJyMScptj6QBFc4YDS4QLdcbqut
pvEq2/kWrvx251dJzAKHgFZcZ4isIYQROC7fqW1ghrMrFvPT7StViXex/6m7bSDznMZPAhtDPjg2
VEn5DZDpcEu+7OMdONq+TMv+ZNhfssIPGcVhB3ooJMwMiDKeV7fl86gN1TUWVuHVMIPpQEelt7cF
31hlrxxB1jTE8d2/GDncHtjTElutgS10I02xwKECon+Cih7tGMEGfLauqzc/hkfUa2n68rDcbMtB
MLhv3U/JJ1FQCcDZt9BzS1kv1z+0g7cjKX83/rY8Y5vLgWfUPw7YdFCzfzOR9o66uZ/xyAeEHU6/
kCyb/Pff8dQZ1Xeg/PrKfztv0lRwD6blbd3qdQhmTS5ZCig4WBqM57p6LKQfyTsDkfz7y47aooA1
C2sWXlCpzTyKb5ytiOLUonDGVu19DYl5cBisdrJh38Jh8BL5wta/xbMVDgGxyfwDaAKzsiJNuenB
wCMXlW2Cs2AcBis3tTmMiPoX3gBX5E8RUkuYPiXDtte4Ra9ALT286f7ZOm/KQyKHjWA8UyI/WCSf
ye2cJG7iKcDWMrlRagRIqcu3JXCUmljomediE0y0s0qSxQ8y/oV95MgWHrpPPG3SunPeuoedAnSh
q6nNVm2TkijvNUkmExu4mhyJvJYjoKMFHKBS+rVqqWpwvKHEL4of9AXvoxInxW+UntTGaje8MmjO
sS8YE6k/c7RkbuxztydK5Abs/f2X/9rC5MJE2JgF/umHPucCVUF76vCSyv/ayYubOEx68AmCiro7
GLJ6GRQMRkNqMt7QiqM6DlIrfS4iORVbT8UzkMc8GUGqYL8VXrVu3wNbhIGQ5QF7DWgbkMpHgtA0
hSVryM3JLtPNJ977GL8K01ptMG9lMR0HkotvoiJcteSmD80sjV39VDU3iQfmAHjNCIC+p5flZlp4
X9P3v3Tk9Qv7zkrsgkixQMf/hscO1wP6pVSJGov/zyPpHpCiPIFANwiGSy8QhN7bkWTy40rPD3gm
Sq/YoxilawI2Pdx9MUNcbf/R0l9mKBD/lLUXnr1E3jEJNUlLsAKtDNCs0L9pFFI9LtkdzcH8aai+
lTF3rG/eS4cGytIXeOgS8kPPHXWIASWfi1kksR3Eid4gjs266uHXQA7NdOnm/eIU4TjF8n4j692R
qfn/hw+7UbRLwuxuj6v0vNhQtJR2CIFN21GaRctlOkjdE3FBHA5vPtbRLZWCeVSvWFlsCydWVnqq
R4E7H1jbJo4p9Td0loW8JN474ycbWjRFzmBmW7KDOnKOCByEJb5vGVmCFakB5sRhJARQ/KGwUF9f
H5dmbmjdtQ4c67JCbo8UOG6bqKMbOMpVHpg3d/Tx48w2VtfGeOQf1S8iqZrGr9rskeaPk4bCUVG4
61MSVKpN5KktVsANIMUmJMuPucit0Zz5/l3frQDRql6Be/YeCOV5P2N0bbzIRtNvqr7jUJ+6exuT
ASwXTg8HyK6TPyrPVXrYWaIww2iwt4HmORU8tigeZ5CsCvpkkldTQsT3iu3GwE+prpswKep3ou5Z
NgOr7mLrjqCVkIz9025UL2SqZNvVzK572/pXbWJvRxr6Y1Djlq+PDJ631Qv70xyNWt0Jj/lIw6j0
6IrGfzqPJvQ2s7gK/POJebkqwjHS6fjkvQkgZk5lrkGtoVIyV8dB7wmO3mMSsWGYVEiHWkgzI7Sf
030urKUfwz+0cH40IzhGp/5/Pc3eTCioRbKNfuqAunK5YOKMQZRLB1D6FfUl7oUbHm2dXzmk1ut6
2Bjk/cGsoc0kUr3h5f1IvenPd7RHM09Z9JYylNZn2kMGqdue7NmEw3gvuEOCYMaa85q3MiQhkKoC
vlPLMh+hlduWRjL8ohp9RPR20JATafyU34FV8T+IyulB9E5O+vr+cbKgrjV9cYbX1FEEeKQJR14K
ort7kGjFnb/uX4iU3DJAjE4L/9i3WWfU/MuGiijtbrVo+Nl3zI+0zVGBTsFRFYW4GOzIFxnmBvc5
8bXvqIMCB8Nq3Ei52GGx5NWhQe7E/i6Fo1fyVOi2cYsW0dEujJCPZpd5yUYAwmx/FgxYKWiaWkFS
dTv0RCNRPSVUerm4urnWaVJEBPTip8D7sRxLSYoA7d2m4gECsAREJVRex2xt8bL3lDtrt+o54jkw
1qS6kCComRB/pZtQHg1pDdH0sDeMdyzJ9E/UUvQceMhkRbssZDkMK+tEc8acKm4x6cxg5u2TfNH5
SCyf+QIh7CQ+pm8YzRWdS2T8iRPKCcI36RYYfZ86WTOjhcp8EdB99l1CdN9OtfwCV1gPEIusw7bK
niZF1J2LFmFKEY0mdkTUo4G61BNPIofO8nG/zs/nKbhqqrLXUi/WxL2o10ozxzk/bMrB8HYz67HY
swOMriKWNWm/M59NXbrljWvIJLqxOKhNzJ1RamjhPguN1oHtd5DSRdVejSldnxfR+wyGs3vqkEcm
Zr8Ar5kZKVwo+OShc7KFBSIWJqgOzJp5lbOIBxZ2OremY8Zz906PZa/CHB+uGAzBoXBGvFpBXdZC
INZjBadMrGoPMbDYce32GkQHsWbkuFRE2wmvKET6DFFVWyuEkjQG1nKe0+99ggm4eSemepoCyBHK
nrnX4PNR2bl6d4nZ3hdIsJWrqxQPgRLg7ks1WnduqrzvjX+GFruXSZ2agZKGO5+7fHXNoPSOCy9g
d/obTKq80xOTvB3XoUE26y7esx21FQw1EIgYRkXY1OrdnzHjBBoLd448ShcS9YJuMm2hJomKZ4PK
bky3iahuxbuTNvj9XU33j+jH+YiYFukmeAaPJqTnWcfcPPNbfJMohfEfGzmZVJXyVH+un0PNcDpB
aiSTDV0b+YUlalYOaqlvmdQIfMmATpQbFOfL6AXRV6E7gzG42u1tdC4H7Gij+MWnCH9brzIS3VkU
lQsjl2DDdT/X2oaPmY/8o45VhmAppxWGuUGiXlXccggEocuYxqyBs43BJESA01W3Wm1BC0PwS+N+
Cjn+i0bPyhE2JH04pupTkVuaW2Sy9JL68kXVEvar8i4nQHwUiqODNhcnJSVaQfgowWDYDJkmqVFA
up/AjW8+QKmZKqtzOHj4+TY6JEIVp2uHL6ZpcnHG+bISKmyRTNzZYzrGhenxGlhq94YqzQxxBKot
6p+NV4r63BlDJFAg9JciR/65rtf2wDlNoc8rKU18jDz+FIaJIAReM4iAHsKiB+hdRjqi26TxHbJg
F5ybQJKivNHiLkJULhYjvlNkNtCjPisaaAdQisxmeTsCFQ/yBFYTucM/UACSPgJj+qZuQpokcRYu
DCYiA+J6FkKtHH7DrZb15NZec1O1358t5UkOHwVB6Xb1JIfNEstXEXKgtrJXpoCU0mJWFLvK+FVi
4WbN5B4/korTpyWINBMTTDAiRa7DRc3u6A1SdeH3t412rwHO8R5TR7dzXFb4g3rAhOlIwLXJsYX3
0isesI9ZNC/MvA5EZ0gU+Nq5+ue3g1/d/9JGG1gQPMmtkGE62QbHC0FtEdlNH1+ULp2lQfqaozrp
ERRaYgd3kV6P3RvrhmvRkBKAVuEL10C9oF7whsnWu1s0c7Bvyx85XRmbQM0yQ9iJ6iKBDQzXznnt
ngKkdPZo3GDdy4iuXCBvCtCzMff7KOOdRkdc1EZ6Qvs9XjXxr1Ku/ugz/X5I3UEbrWdGuMVYlUhw
c3rUtYWXOlesRdAT4oVcYkb1fbvTQtevm/RqArbsSLiVrDsvhwHIHpqzXKE2H0+4W2LzMpiCXaFT
uw1Q/Isul+F6GTVi3MCvEtr+pKCa8pzaRaohBF8lVQTMbk4cOw1wUl/gFpVVFas4oofXMLHYqmrE
w4Rh4kjjYKqKxAmKyjgjLVxJ7UrfiekJ+0KImVaI/MjA62v8/LTMnpdMllerPmbx3q9EBzDZC9BG
5lal0mUMiFSqZ9xg285cOTsK9Ht5v8JxCaM78KpkCAlLP3VG89Rs6TMAUrgmYkvugwYkbBdzsFfQ
aFhFISIj0Lfa50gmpt+m7BmEBiNzVAC4CwExmowyyfh0xMttOW+9r+ejKJzLgic3GTxZ79vVMJDL
2fYoHFmet3OkHwTsv2l9Bu+obJKg040LhZ8kuOMdStmyI07yI4u9rsIBf3PgbkxNSREjOX8KW6aA
fXdEQkWBdF/3+h00NFOaMU7DGV4nqSjYkbFiDvSZSfWf6vPSjgTIAMya4oKb7Rqb7rCB6o1YzRrc
VidZT03Tj5wbZJKNIOyDOwhELfNIxgR8RYNY4kenu4I13ZsaRSDryXj08kuXz7CdBM/amldz2bc3
LqTotnsPG7lKLZmH5oZ2P7SVg4H8dC00o8go+JfWt3dGCaV00YwqjUGjBMFdnwLGYn9DG6+6CP5v
VENQNroQiyq7+qJpdxhs+M65hc8IRD/3I1zYt1nb9NnwzEj6S6DCWCy5Ymf+LHiEmmb+ajPN8OCx
q9+cVMg+rjI+iLf+YuqU8A7XIgrD7bw7yu28sJRnChFDkdjKQOlToycnS7HOZqEusVCOZ/F31Nd8
x1+ARfOF9pranJGkL4Oi9nFdCOyxD4KwxGXCaovssRGOqLEPZIBH/B9Pp/5jSijx5W1V+nQnISHv
FlVfxoHQATr8UIjUkimDZqPVGZxK+kv3K728KD75/GoQdYGyvS+4pF9A0SMdzgGMKVm0YKWX9jYF
m2W3RZYCjN9CY6h4SO284A0Qal43gZ713Baw6tSxA3Oy+TYMjGgoXO3SVxLV31wSDzoWePXfGZ6G
qH5QPoH1knCs+J9qORViaSCPTmvV54Wkv1mhS/CgeD3bALv19Kc/AAtX0u0JWY/nuOLh/8iMY6xo
GAwFEbK5cvYn9OXM2hdr1/pnG9teym6tMMk3aPY9ZSRjcoRmfk9wPvC1lmKqxrV2DMFd/fx8OeUm
ZN+9Kz6PBZmyWesH13HFgFFBEHfNlMbh1jEAk8zMw6hSRBA7iu327xMO+YkP3KRiZYXACnuxgaOU
AvwUMn5C7syyrrOIQRV1F081MgKDbY1o/xXMf5MySug/E41VhbTOO6FGCBk0j3XKZ7+oqWmqWlnv
sP2aR6sGDKDOLZ0Q5YMFlW7hkP64bAwNwWX9DrzyaHPnQyu8HD81WaTDiW92A6p1v1ooJrere1SA
P5pkjNUG40vkrLmdcDsy0nxJeNwuXwXWXAKGbK5CetHBHtqnq2dLuqQ4qEenLE1b/nxEV1pYLCu5
TvcCpsMk4QXLkDv9nxU2a7JlAGl5500FyjTBOjp3FYk//3Y99EbGkihcLBIaSFaj2nTRWvI/DUdM
eddS8kNZPOUYJFUfBp8aG/aFKCbmZEg4wtdDN+RM57RwVEWjmEC7GWdjBiSNUJLPSmK5RA6C39oe
i1loChm8fzVQfiizHzit0QUCWsl8/nxerB6OxGQkOhTNOEGuEkBZ5rMi14F1hnN0eHfX84RJFm7C
AHsTzuiliHtIUISX5ErCOQo2t2fxAQJ7+ZCeDlaL4mEESw7nlULDA1NvoEQtDE5CUarEKx5fqU9u
YRIdoxGlD/xHs/QnRZEWQiprMndxMnq3sxdI65c/HHaL6JMmuo9t2KiguPLGsAky3moKBMmy/857
X73zm1bQQBv7CzKYgDiO27jpUj6skU/flhFrluCZVjBSnmP2wLO+Fx6QTzR9S7dOOqTD+vOH/BlD
PDMqIkm5Gu1IAayclgqhI5mv2Je72WfVkU49IVSfkmiThtgqjRKpmCCtVs0w+oaRJKgt6+sAuspG
6/7rw0ADL0ctp/TGzmPuL2tzR2fb7UHTvcJP6G0hfL6cdKrzB3Y0Nbz8H5U29KMykztG6nnQKrAB
6NfkUohP82wIKgWw9yJBauATvTWwiRdKtRICa2PXTb+uAfjS1fBHkIsMhb395mROiBVA8TGzWqTh
fbnQNyOOofz0A7NvSIBvJzO9j4uq68QXC836VLHX9gLksny4UE7I/XCLJc5+pYAgwxSWwBI5csoZ
H5OnWY881UZEhoOezIhjYgOb2VnOi3LwQaCowywK67/sSrrZq/Ja6ziZMFPTO8GpXsWOVzQtQiUO
QayIiAdGAjpDsZ6lwgIc0vIx6tRksfjz3tu/A0sFk0+zaPq5fShq+yxb2DrGV1zSdu7LGALp0+1d
7f54/YSOnPxvg9GdiPNM0ddYPff+Uc7NCQIByn42OrLwv0W64QbPsGWZlQxncqO8tbs+QBtLhUnP
uBT+NQ6dugMxdF5QVrFXiDdRTsqz0tTwp8fP1HRAFbkkh3S1cp5DUlObHA2/8INee2nKnkUPhwXt
9DaSzpZu0VYcrCkIZRawmDcSBhTDO9UFdbuTEwnadFXBC+1OFKNIFbIQABY0TbCdFgZcT+r20dkw
c0iVuCkYcv9CS0nHFYzAKvYVeKC1xspuqqgkLB4Vlc8sLnd/R4I6bVBtduR3WNoHU9NDPgsVPI9e
h0lZYCnAtK0+BR/QhAsTQ4h5VaNmK1XFI45J0C461UCtK2h6GTyUzn7+pHnLJLYT/we7ciIDGnTz
6RK1dzt7RkYHNKdfyD3QB6bqL6aX4MGidGDfz4PH3yKEi/mslaQYqIvgmK8uwBIWLXkia3bQeBsL
wRZbCg20ZCe095luXGn2ba8hkIECUzlM4lvB+t9sCpErkmpS2Ju9F5Xvyv3ok+5AMDRBjORNA5Pz
DNabJM0T0y/RwNe74NMNc+2h+69xJ51iahyk/uwHhZFlnoj1VsDKo31yZ2uboHekktfuKx0uftUX
cpYRkHtC6Vq4ka2uSFqf20kEKUDzyHZaYnLqDOjdJTdn1ADVXxm71uPtHH70rJGCfVfhDliIz8du
ylnvTNqaYx/t88bqi7gSwbg38n18vPQaVcNEtTx0oCoua1pja+NNYj0oDnUFsx3ruYp6UORYEnUV
wOsM2lhwt/jJYaoC5gS7W6avfhqxLyDfIBvMPxGH/02Uf6xeoQ1ORw6JHm+LjpX/wgnMreW9Tv1o
c595+sC061RU2gbzIe1mmat2BohHWf2CNxtuWVQGax7gCfGRj7XnUxHu7vwr/ZW938Hz5Fgr2P7D
Xqy41/sm72xyHez2KACRE+GhSsOplK+rms82EMBOmTdVqxDkvH63O8NYy+2mUbpEXc1qW+YwqmwG
V37t8EWCQFicwjzLQDdqw/8aYrSmcz4mUt2yZTeLvTfctJtKN01zBa+BenMq286JANaYMcYMFLu+
hOYUngSk5MRMcGuEbg0d+AwCU7uo8gTZdt0yGt/ZfDaajCY955r/VWTe/JLip7hwfVlX2lSWQkt1
A4L4XkOeGpf/IA1PXDIj/MOkP2k1GEO1M601ifsBlxJ8U3GBiCT4ef2XbY2cWNNtE2wYt1fiJ1uQ
SGc546uVTTboJqguRT2yH/4vvJkgQOWtmI0gPq3eeWGurrVWtDv0PiJ1vqYmD5g9I3e9oA/8nQkS
3uDuwXiY02W7hGLZ/rpt5eTtXVxSWnR+BNw5thVRX99nQoR4KWkDfTmG9yopyhdrbOh7GQSYiJQK
u4P8bO5damIjCKiCUa4igeVoj+vICN8eK92qkJV+bwgghM1/CRGZ5XgKktnR7AkZUo30Zzc+iLJD
nYf1ki2Fe5XgVrKzLTXZ9oxlxpudw+SzhcGrTpV4KMkcK45GDlMn7L7DLOdB8xwpKMnABGktpEri
SFVgFUq0i5oVY35gIGCS0rKoR/NIJLid8pUEHzkrHeQ1A9finUZIt03YTikkLXaLv7ED5w+QJ+0l
mWxpSnFQgh/N/Zb0Izi5JHYW0bwWQOjO30huvdFMyPBkDpbknxhYiVZxyqrt+GR3sQP9KHkle6Uf
ScQqkZRg+pYNXATFP0LygeeCWI+SfcKlhz2FvUr+OVopSE7cSOAp7oqlwm7pwGu7baMO6VBhSq48
YIv2pJtkexDGUTHCHaUI2sk/d/pcKGDm6AEI+xxAyiyoMEn0aQ6iXv+j5ufkjT+7eZ++ulSj1nNs
EQLukCDRYniNalm37iOxJDG5DmLx3ph5A2oHS6vt80Uzo/HQAVkAzFoS9C4EHtH9VGFCloJdReTg
Nh4jGOkSs0cCJCROrBYAa6Z1KgH8paljhKlY/u/YTRdwaTHv2mcelX9Z9bwuklR82aTY40Q8WbdN
QlLTZa7dr7eVIOr2Q9c8ziJYgYKHeiUDmC6Q6VqX6cHItu8GjvWm7rw8dzFcDHthPpLvf4d9PN//
EVL18Pds/jBRWXPRycUmd8SRilzskTTjuJpl4FYRksQlrP6+95d+2+R3ItJ7uMzKqgFaoHdZ4c50
oOWsTBLyPCekd4pMaSbhorre8QwtFB1fo2K4S3GbbBg2I60pOi92bzxtH8YFtzO9Rl1ZToxpZek0
BvhrbRQIm64GGtOYnt1cSokOvj1JjYeF3lOzAGr3cTFcEMQkgtILpt86qNqaxdq1buORkt4Qjc7E
QWsQ5j/9A60l6Duj+LktMsNFFb930bxW1EqF5BIlcT6a2hn74sR08z7AwWnqg7rqmpZka2y+USIT
eb1TN/INFAmvKlh3KIc7179tNbHH+V7P9Ceb4+VEnV06+tzI49fKcUDrJAHVBnRWAtgtuRd/agI+
G0Zdfo/nTDZjm9kQBX7vE54RJqBvVdlwiZ6KBOUFv8kHmWrW9G+FOtR4XBCkWtwMBYoS2r94iS36
FvFzDKKexwp7Lz4TIGaJPVNqR9eKYmI1CtdF0JnoMKKsv04Yvp/hFzCLaXe1ff82WuoUxxBynZ/X
NqU51lmBibbN4ggwynz/m2nTfSMtre8/zltRF9GnJD0H8WNYApJzmUrtXfcVQyhI1PASHbxxv0zV
DXWIVxmmPFk610vyRvTkmgjE58cbIiuDzP3iLZ79C8ljQ+kiF6Bpul3vSDs1h+cfqF/NY5Y2v5Af
R5N39nqq14040mFyDgqlq5yQ/j8nwLKjvSeTKjmum7e5maYtbODZAVccvqZaUXxlA3NkJNLYWQDY
8J85uSyQuLbomrlNhJ2TeKMPHIf39UExYZUkueflkQTHIMTn22lNPzCAX6L3CeCx7I4/tQJl2nAu
UWFpyg7aLeSw6dk9qf0CeuAcNrYH1S2y95eBhUy/4KDdgXGI4TdfQAnDXV/G6sS5gYEaGXNAi5gI
kPfxuDoHortgg846Yu+Q68fQbVLVurvtDyHY1Qxyn+CIoR/FDypuiAoDc2tP87wYLUkXkaZ6UqUd
RpODQJb0IW7BR45pHTkLjYlgjTKJJqilXKhrmP6uHL1P5I48xPgtWoj1zcid9RpFNMgy6/7qxV8C
YxPKmVRtRPF+uLd19uWMrh8JbUC//3nItJ+uFQXpCDUeT3WbcKtCfJFIH5UlJ12QOzgPTBPDYEos
njQL6fuHED7koK4huKyciAzqViUnmhGBSv5XvvvYaV44iJ043HwzlZ2+oAyARBLRSSjtSHK0Ewdn
9LojcqOjpki4uu0nJsiLRLGRw6LSiMwE5VNx3YEK491YPqhqKrWW4BM94jIEMCCyQDckkiInDDV+
Dbiu59G412pLzOBUTijFscFsVafNEhgackXv8Lr90zrD0I2tE65ZHkeEGVZhHoyOisQRSFR0PQ3n
wSHw5yeuiFXJcjHgCh18DJMviNxd4vD/YT9/SHw3a30u8rLk1ClqWouvahbiDLp9gkR6L65wvpJg
lOFIfNl1Ua6eX1ZKpRNbqI1jbIP1WNJU4UqU7rs+dcSbtqTLstf4mlPQB/ufHaB1eRWpAxbHFn4M
2TZOQsE6fo8I/L9Buek8CmjFfnqQNiF2ZnMuRYe/tiMnjV6ap3/QH0JPXxPF+6ZoGqsHKXNGvxTU
lGYrstmEPPFPm34+Xz53osz97qvmkmTpJ66oKn1Qhzl07at2gRjQJ2bp/GxIDCUbEwL5+fM34eo0
h8riJSYAUNaadRuW9RhJPzmehiH/NES+FbkSzV8cCY8I11mSWLRVw2Wal4cURIaMWX3Scv5gutHS
CvOAr7dnQA5eYN2XzbzGtyFgT94vgdY707doDF4Y42m8Is7suLWVUsXw8+pYInx+V8SR6PQ3l7Le
pYVzu0N4ngdd3523EIw4odcRrwMIainBlnZnA/71xvKP0UVrymeTJxMQ7SjrvLf3hoFQZOfWiZHX
WRtbdfk5h+IiBOct7OYGMCv+ciQyKTT1RRIy7TXIevsXKTkMWjLEVc+GOl/XcNUor64X7hDiMjqT
1M6FUBbx6s4JXU3B75aIIVgRuyMMrfxU15erBKd72QO1JXLmPluMAJAkXPU95UBB/ciFuPGLhTl8
JXZ7WuqJYiocNvBEmzVIWcBI/kwgFTj+I2ACc42ocTapxH+FzDeM6OqORoxY6Ptqru6MlYl47S5l
MUTm+aT+IHZDsrsm16aFr4AveMbKPbnm8dVulHYbSxQUE0YbtQaSkpam0m+vbg+EzPfmglfraEIt
bXX08ziIQzQKpQIz58vx6fykMK0yr2AncgpTaXT5gHzPUbdAX2a7NYBq446o+5KZzyH+Be8o1NTs
RXVhTM2KhUhpaeU3rS7AQWailKmYRABU4dB0n4+AMYMj7Sye0B+kQjW5uPsSyjL3AA8Li3l/dr6v
Mxa4iA35jld4nVRrjt0tipi2G98VRDVUK8HrY1P5q/WHTrNcczkwHoDlC7cGMo0RyAqqwnUZDBmm
R3BYGl+7ltdDTylmf87LfDy4kwwQFZag6OrDQ1m2gE73bhaYKmwnxfU9eyJ1bo1bks9fuRi8twr8
hvFNEkHzY81c4VWiXecJN8jG6EN3a6ZPomh6pOZalpIhwf9h2tEqxm9hsNJ6krq0J4NkX/npwVky
XW6CMVncerFJpp5nlJyKMTBjrhH89xzMK1Vu/Rvjsxie6ObDBwrUoyr4hdafT5pVCxEbVnwZxXeK
N5wYxZP4gj52LUg7Cx5UJDdH45QeTZRGXFBw2fBHuoPyu1tiMS/KvlYHw94RfA+/ii98whY0hK7u
/8bpa/HfQ85sCN7InUTRI+QApmm7nq4eRL7fkjkzIuGUTDcwgTQslnbdwLyLHwUegXycDGwwo3M2
TjhMrGthO4+2henw2b1N4Gsg3xGR850ooQvwPV2cz5iFzVD8oTs+ESz2QG7tEeWp2P++R4FGEVIu
ozl6gnRGAwioctsKs7lNaeTdsfSgzjufa6/qE2zIRMNCPHnPo919z6d++Dw6Zjz8/nLLTBJxupw5
M9RL1+gdhvz4RaJeoXR40qceNcg3ZG2FZYhaZI4a/DT4/dzL+DnJzkTexcw+3rh8U8JPHHF9U84B
n1ddNXtlUsLI44v2Cq237lLR+EPUxgOWqPwpLH2ThBg7UJx7Q70WyOcqA6mV/R9er7F4PDSu4X05
do9bUGOY5AA65HlHmIBN0AEiFVyObcczSc7YCtXrsL1C+XzTNw88+a9LsVIoB41vjtI+wmLq5WHm
OtoPyDEj1hPpeAxSIbgtkPqng7EcpWbZWhdz14MBGKH92U1B6tNME/Ct1GXpfTfQZ7ig2TStPUx0
2bxoKJOrYuPo69WYi6GLjt6269Pq4J90yEgLGHcSnP8VlngWw52qpiFZICKg9WjBna0FXuQFyX5p
2JwfKo1YGzH1llXdeCyj33C/QP6SIleEzvcDZLjM2X9MK0bP1Gvq7KmV2CQgFcWkZBBVGQ4Y5s6M
Qcgzp5RNhIJaEWS7XH51u7sTOOx0xpNIhrn2wuvcuawbRmqXiBa611pj+B3oAQD6HV78LkIGnNMv
UsSQZnfqAtpYnjdcWoAXfWd45QS+Tj8+UG5wCQ0EvFsEqOkJ6KLvJqcxNDUVm9/8TqSRCqvyDMF5
tIqXChsDst3YdMx138Jr0uLeZlan2OLgrRP9puLRauTQiQRz68d+G01t+fIHgxoo/dms2wRPfmte
2EHNzrIRXvOjoZDNiA8lIunKcXn8D828Fkz3p0ekJn23pjp68JXn0ipFRJ87GUaraxbetGaXRv4K
2+Stw0irOMgYC+0kZUHIdgl2LFYCMBazyAOYYrPjTpjTidFlk/jDcCrQRjjn8VXKg+Mv9tzDfY/P
Zgq33wzcM2TVDLJQUApMAgyA17a+0PzSmQ7JkI3AUt8JtRxfzE1SFc2fQVUwesqOnUFoOPd0lSFi
aVzWGAhmIj2W1Vz4807KgEpE7GnOHTXW895gsUc19+g9wAJWJ9P/YG8nHweA5a5lzd+pQcFciDja
p9kQoe3SJVTx1Cw3to94v+DzimOxkG6tGsj1sepRmgACYxXVIOY1n0eRkzOcp9k5lVmJmrIBWIRx
hweTyF0KR/y9mkwJ5wuEtFiPH3oN7apP+GczxeghPAQRVjd9yB5F8XugRpp2bnohmOWWFe3zC4Ra
nxxqZ/rSvhhxcftwbRlx4ztrpk/DngPWd/13NxB5amMMmsUkUvZChBjTS93IGuaBiMfkXluIv4WN
o8O4mIvO9BbW0TVwDguiHZT55UATgcE3halxHAHfZmUL0KE7Lha1zyiIhUDpVMD9+UPL7XaykdUI
QRhyuMOYgFgOrlrFMrHwWdiBJF+7hGNq0A0fOo0Xlg4ylbntsCRs1j5Z23LZ1Hlqv1cu8C6ucTjq
Kh67gnwpP7vrIO6XtY7wWI82DMVG9QG0CGvvgQ7WyonWKdCtfgKZLIN5fItfTaxppPs0vx8wLI34
dUitDEoSvn/tWttqdYrfs3Vqpizk5hcGMBQgCbTMyZnhWUG3NSyfBrbZiB2cTl4BItPetmOmVnUl
v/6UqLbSsROBGGBE075KgxdrkKltblwdxoHxX6n03E6Re5PqUOfWbGQrfh91amSEdlsHy9ygKbEn
+WHZBHJLUJc+0ltwYuyhQuOHxphg9S+lNRPJ+LlkOIyWF8G2h+j49p1ZgWDvVEnvREp3/lGpJQja
M8DUSHJiB4mqUHX9GqUZPaclXqizllJYBla3Qe78euiu7WaQE9kt8rsOJJCFuSGT3LOKw5sEPreI
XYnN5QzT2zD8IStDrAs4YcFmVDKUgwWL2sc2erc8RgSS1bwzTwVetRGBJfVzsNpglQN4CGklGRPW
2DFvM34RmgacJxg5774p73iOjSn0K4JD01Ueqre5fnUd8UXBMy4HGOyvt8DVlmDTS1YTnT77BITH
jPXcwzxDhm8jdtMEJ/kwg4o2tZ2XQUeheOqTzPik1gN1lmqMhZgZWT+KJfjOUPWfooGCKHdIeyuT
UTSWgVrJNbn87dcbYNaYGrGb4tAg+xebenYJQgrQ2cmpsvQHIpz2j7x00cHhxg6X5UuKkjkeClR6
AMq7iZvIXr7H8KUxAaVJzLLF+BrglsFMkSGeQBKcHVtOA4wMfsOBfB2fe5a7PF47TQAurSiqBnOc
91xGH06+7gjn/AkYH3IE6+HPwtB9Dc4IpQmj1/hxaIIfjXh3ZGUsNnGrcfWe72w2sKpsVFhmJtYZ
NeSFdCQLwceaWt0WXws9hKfUs+cUaZv9VjKXnmJYta0WUGZpSIuNW3gOOeUHdcJx1HuWcyS7eX+c
jhPyt6WivFctigUicNTG/9PdR8xB60QriRctyroFr3fQIBBa5To5CtrSvI71q3UUbim0WPsCRCc+
zeVEh+NSYv06+Z2tjD3neANYNR01JXmHCI+vMNxWtcFEf+oaCokoeTeF/v5343xPlcuUxwBWnHIN
QO9V0+s9TcbBuJ1es1qMv1qzyTM/jXWgoSBUcobUUpicV7LMK30YaSKPKWjMsbC289Tw5OqUwvIn
yttYbhaWCguoSmAqYrMi9sw4v3QGWZgizV/uvK4Q21Kba6ruvzSJUR2QRZh3HGVdZa6ZBVA2ENhw
d/oxSt0yDb8jDFbScwrdrCgFbVuiSkdU/Ixsw8B8al3R8iiKYA4TRGx383rHxrRdONrxYImibvLF
MDQQKAFTqDMDOckaCIUUZ5/hPbzgIoe6IG/u/JASLR/yIEUranOAHptBztv0YILj2xDBfpxIyap7
uB0qnWbH8ns3tCfrTHUGI4Enb9tpUbNfXv7NIgsSazkWCEZAEDmP7G1Mh1YImulUGPGRfBBg8rYi
hoeZQIy/3v2luymKXb7+PqwoL6qg9+/v7jxTMsg+qgDVBIUiWYcafmyAmuQCbREdEkKunE3t7PY2
gRGWxJ748X9uJDgbwy38rhv1bMI8tEKeKlJD7SCBGfZskcaX+5QrQ6Ksc96ZFb6IeDitQ7b1v6SQ
d5QLAPcaq+EnpYXGUQ57TwanUlh2BipFixMZPiTohpSX2I7X57Gj92shICQKig1p1ni1FGmguDA6
1csLglKTCMyGHl5L3jOm8jIRcdBfnQfYKL3dRcEJo9YNHUMXuMF9t8nhkbvnGq2pBhmnF/aJzCjx
/YYQCgsxVJt4Dk23ZPjpnzx3hE/O6xtUxCZufu3vGf/N9/aRdsA0v47OQVNh2ATAYII+JSxMMunH
AktdH8NDZyGPgfxrV/lCvuVwCozzyoz0mWv9Me1pCVuFxrh2khJTOeQ5RqTW3kXiuObJi5wQqWeI
r8i9YWnef+wuldYgZcMAAD0ucK/KzkOrbexFS2ple2DA5O2L4HTAcxOEGfQK0jw/Bc7OwS2YXsF4
i1wZlR7xbpBRHzKTVtEINgbMJybttjSnrDG1cA2k3QnkOoK7ICLoy+vrEu1goeYULpEtmg2dnQOJ
7cX1+9ofWVVE7Eo/lelZdNQZyuUF+0JYFF8S7P3j86kkWZYsv0QIQkJ4V9Ps5NGJCm29f8TVc/dq
Lz/73Ryo3Tkvi2Cq3sXQ9ZdIY/sgv/c3OAGGd3fglwxSkMh5ic0+zaBdlOqwlbHRgRQRUm9ki1lu
9XbJoGYZvF/T16HLvO7/ZFj0Y//d9sMhFpLoOK4TPKX7XrBBjFJmtnjDcKcEC5eIIyd7gSsYycBs
r4yRSs1VaMpqsqEszesvEHhr9czTYwCk4yIzjDARaNxvtHsMuDLov498e4DV9/vYV9aAZqx0dQB6
QUAq4G2Gy/sO7B/aUbcFwRWzRElYY/O2dmnHH2sktemYN7Guj0RYOl+FpPF7xsX7BTgOt0/LorI5
asaO2fxNJdyD5lkiKf4h2nmV2pZHgZQHdvK18Mhf1rAJrrH3CXO4WIlz3osTsOqZ9VIPbrCWosuR
u9lRXkSiFgHc19R7DiDpXQMw2jORv3lAB17EWf/Ara/ebrGLzpnAuXL9MQ/VmZIbhuRJIskZmXl+
4dgLs4xGln54Cb6/qemPF/bDk1oHfTAO86neNmfynYgzIXIdWPlo7b3jScTvp2bJ5n3J22ONUSbR
0jjR2rNvQTSbMqDtTVPwpu389pOeKXwRj5Oluipqjco6FHuyOhFYVej7UJHjdr8rQQ10rlGPQbJy
QsjRRROTM12V45hceWcB8s25lNL94R3uGVFtLVV1j+xW5+WM/OMy1SvjiJ8HG8aFYS5aCeUAOtQF
twTx2UPekST5fYXZV/P8niDyUSfxLrcXcFjXVTs1rIb0OUrpGji5KsePVgdXE+qDCeQFYDZh5rXz
iHNj6RkebZo49AXPOfVE2HU4YBGtoQFBs4YTQV8hEbxb/Ejs6sLoLfeb+K0QVqykdKqNcuBctp+x
wJ/GIIXg/3jw3X2WXa3gdM/cQRcZsnPJzsDppLjmP9FdwIRqQHrLXY0HqoBCH7sgeHAZg305bd00
Hsjv848HOfTEtE9IaJL4jzeyM5KuiIvojZyknFgtIaeUk8OBG5qHMVyoF2MBNeg0JYoy4V/x3uOy
B3VJmvee5g93F7uivMGR1p+2IhkK09ZPh/oXp4dYL6ptHTpcL01QLUL1pBw0EgpFNkHQ8gtZyIm9
oj0A1vu6taG7XXTmk+gjKiF2Y2EZJmcwe4L+Bowe8lj6/21aIiqP5s6h+ytHputxbmFrPOqpmzgR
ZRBH5kGGbGtq1/iuApMUzIOY3/YSUFxGVpavH5H3UoDaxAM0cfO0WnocMUUzBuOlq/6/5TRFW8Uc
vnp24ILycCF89Ef6qhJI6EPfLOQKUBpca2BXSevSKGm6hWh9KFyNgu1YqeJ5B/z5FhBXjtSeMgtG
iA+hFY0bf7rrcHKAXcN56zzLfT+pOwiOIeRAqVGEG0bsZh8JcTyQPODaSFrnAe46ghKyLneYJvUg
B5wlgt8+yY3WlJweNz0mgNJQEE64BdbD/p5a8n/WZXgJ5h7ctcRvQqW1wMX6/ZniO1GACb/fAabS
nMT/PaBSOgQ5j0wM9wrXijYFzFMZzLTryAR9sJRaj3Wec9xNDQQz77mMEJsXNQ3QavETQZXlmL8C
sdVxr/3cUde2KF0EsQl6QnWkPhrgwXJLyRUCE6E/IrMMJTfV9D5DSgvMatLDHRqernJSM7Bsk7Th
MXeuDcz2DT03PcY+uPhdu3tIYuXYLgfrdVJgqvaWbwjJIPSKnFK/tXYSSUotGZGqKWufULq8ASWe
igdvaFb+dEehclWYJJMFXAD39vnUWRk0GmgeXrwJ/WpAsv8EP0/I0kNfPnG3YfA1KkEBJLUkYegL
GQgH2kR8hdLfn7Ntw0+i/JyyjH+2pLqLRHJMwdu+XQ/6ARxEnYGJ1bxfX1N3vVdaAsz1OQ+7L9Md
Ep4S69vI+KzOyNmjGW6zZUzJ/MXHgvFTaKOO/VJhtg5uIO906jzNTPGkShosRcEDas2dzCZUsi7q
dvEpd+tgGI0M57z7a3IB39qe4EOLJWzc3o5ANcBLfh5oZIC1SvBspKWCNxdeGAnaWGXX3XD5ViGV
6Z3mHKCoB+npl6bO2LWJ/jtGhr6Zv/66/0XtzWmwO5TsIp2ml5ro/tmMF5WkBIkhh9NI5YA9xGSq
h8UBsQaO8n5FMJ//yiINMjYRYOw2aHPZNYubtIBnfIyuzNTcx2CqnHIWrY6ymyhZ43q95HnEjyQn
0v7EyPeNqIo5QuGFIRzDA01Nl30rMViyAPvoZREYPr62b/aY3coFZpDnJxuj9LQMaa9NgY3uh5Lo
MHoQPF0cMXL/zvD99T3UXh83ddQx6+QrPXfc3/kTKzPsZJONJg49X+Pfk4vv6Tj8lPy4t42uPCCJ
989brwV28M+S/HDg9WAQy/V5a5d2W4d/NeP/hmtOvvK/7fesyYzpLrKVbmHIl1S0ZeM3M+5IFKqW
v5GzVLYWP9ULfd2lGhWHC2gmcaYyzWH3Ty3VbRjs0eO2gboqyctgB1zdI8O4yQwhTamZf5VmREuV
frtKqCQEV184WobJ6GbCJmMBPnvo5YXPTg8s/zagvQH7p4BS++oL2LoaXGSUlAcJEvCbRGwYmi60
pRmUrCVhr9L4wXvAN5MkMKjMSW9H5NmKAMIKWB7kZxIyE6C1KEp8oCxAeCumaeRCp7U70VJQrCrU
tQztzFElkP4YimcIWrfUPjzzWn4Qp84e9Zs6tPke6RIppJiA++dbaE2j3tFaLpIhv8+tTHYE8DyO
O/bSs11YFMrfJ2KvUszoWyZbpv+sixjlrI+pJMBqVCTgLULfY0g1drO+sU9Aq/Ffb2BTLV8SR6+X
EDBpisOaafcBK5OyD/Dq4D7z/qs2fLNWP92oK+3/WPh7u6im3cu9pC8i1J3GgRPKAfjCjDiJysRD
U9jj5KrFJC5LZz6BVGRQpcfS0n2cHxFubDH4fhI30F3nodEs391xl5WEEuPMgxcEajLawscfbwUU
Gv1fjEQ3PMzR4mP8aied/wGERqdh9jZYn4fJ/maHM0KECxV0kQtXXNnzMwBFe3M0r3cvLUilyGiz
6bqWDLb7VXujzsyx2ICMv2Jj4FmWuFG0ByvNnPEcsaToPDuHzMfK5BH+OXA7ITL9laKK0f3LWMVh
0WjLMv8Fvsh29OCXHxj3a/vJPiJKYu6e16TBByPFx4iYK+B1Hn64sX2Vk6QlMq9TpE4dI+xF/eg4
cS5UV4WK53ILYGaYjv5niKRai67cKZw18pc/1O5k+1jEnBrRlmO0X+0JS38gBfBiOOgiAj2xoSn4
8uSrVulf65woy5zUukgytI37phEhju5T/vhkePsqdRK5eMDXWD3cGcJVqBhpQbJzzY/03HllP7zc
Mfc2xOsWeGJMWBFAUO337qaMscdNhGwntV8kSbd0qNyGpey0HTIYAeP8vVai35tLeYr4uj+rlfNP
VHwporHxPlqaMvLbZh0VdlitW2HLbkRCkT2N+ag9R46RWGk5H4oRg7krGLLid3bUk2WwIjlVa+UT
UmZhot3R6Ji6aI3c9venYbKqSG8gpSifPgZZilFutnsT/VZ1PjCGiFZY/RAny/Xr3/s0AYWCpdv9
N4DOoq4gp1FOhNvIgFvShTFclM0P2tTLqmIplqZidIkquE4hgBmknSLvN7ohADxpND4cmxFnaU77
E6Hgo+THizvS55LwXDUPHD/uuwOvQdb3juVfHoYTVX0pFF9+6K9B85l52/gUFZuGI5pULlZfTBJ0
usDEnhxk0Y18RIpoLt5X3QL65w8kW5LIvtoMHkDwFinNhB8+2R/OYc7y9EkjmpCuUH5CHaaRCqhB
1yFnmBxZVZ3r9leWbKyuHfmi4qWifWo2vZn1a7lr88/HfMlWs7EE7COVF6BmYIs1IrVUEfMwkjD8
vOV3MYEZvNc+ev0cwooSFbJz7XforF6z77mbPBZz+qaM/oiOLGuZKnxKoBzzdT+Svf5rLnOw60eC
as1c/2hDqyh3OQpneQVRfiJxouHQcN75PxqC3mXisor1oEc8W1Yibz99SQNvr9SY2IcGPr85bn/w
HVscnNf1la72s/OiYYHLBwIT25S8+CcZGlkVUofG5MA3jXFBHhzvZofrxTzGZmeyEPqRqsK/WS4u
c5moBzJLSsn7ZSiz1wQVnNnfYNsK4ogUOKRFU1yeUA4+2R4Rio3SeoidVV/4Whfb9srdP1tcdvdL
3i9kZr6EfcpP6QSrKYERUpqg55lF/bN3FwHBeGRV830wuMxS1b3/ow9PT3R0EWj4DXSUUahLOABS
B3wW3HcJz9KGj+QOBlP0gnJYQMkSJNsK169LKnaDoHrfvT9yy22eMafRtGQrZ+Eg3gxMgDw94xSq
YHyEleW7P4UpCKBlDC62knmUaGTpAD4ntr9gNSQVZlYwPqXBM803JdmNNpeZgvmnITWLZvUGEQgq
oMEBY/4bC+pba4AJlw9G/5XiBUUDfQnSBLoo21uQsKQVCRdvOIz69yrkVXpOW4EI+fPFFNgG7eyE
P/7enqbWY9aQ5DyJD98LKa4e5haUlhYAV62EEx+Tfjzcop36L3ICQxTnRIPWnTpdLgo4FXd9DCvU
ZPDDG3gqD5vm/mfkWvaW3A82HW3hJKgsBjKaMPiX8EpMI/WkECjonPekcEQt0a6jY/Np2pYj4fRT
EbhVqk//GoarvQzcw9/IZRsdVfNP8J8Ars3OnUMRZiLd1dWXB8wjPqojC++g9jqPUl1QNf+n33ER
2rbsWrB2aQiAn9Vd0wsN9zVAc5mww/PKbSEHCPD19rdOlEVo8uEulEn+JXtNoKHEpnpPZL20+8t4
cKSeldCrgPIAeD9aX5+ZOdEhhX2y4/6uRpe7bCy05bt/yTdsUOrDRSkdQq1YTJoU/gF9yUXidS4y
VifkIaBN68UCTjScJzpJmkgCrcVoQSM52Yr+YJO8EscJq/s88Zr5KxuM2woNt+bB97+Wpc5MNT53
LUqmyFd9qJlkcslwDPvauYWCXPk280sbw0W7SNtw+mqDvyIMi22uO9cjb4r9CiArMoc7E1h9GA6x
5Sc1z6Xem7Bb28Cv/GTam8PYSF1MRITgcc+qEaRLk5PobQoWcNUlO92bz4TGhYskWyj81Vyn5NV1
bQFd31znNHHSgiNunG22CTPU4PGrHoS/bxZR6lThqldtlAEmWqqhsTtWNz/f4K7pnA6QMq+TQ2XK
ePtPgd+Bssjn3lD4zotuMRefGpR+yV3u9T7xJxD2QkUQrgNgz1CorF4NRLEN5bKGuK2a48rA1p3W
44qXTnznYQFAO2xyiJ52RAThBNq3Z5kQ458winhaSQeswYpjS+4pK0Hi4EPPHJCofJCvSvkUYuJ2
KA9pS1A/OmgKCxcN/HVeYAm2urRlAzvO5cJlaeJrZbmUzSZgBQh6yysgIZGVJRkXW2ld+B237glE
tByYJXFprbZa7VCGiBQsi5jue+S8P+EcEBe9+c4NQ1vpZnTayFvdEV1Aqco7N8S4TP5giO94FLj4
pEPS/Q7ghNDYzCIkbOjeAIA6zVshU1TddDN38nJRkyOxpayfM6f8yr6NOxnLQtuKYdWE/GYYPxwz
HHeLsHPigGX06zuJVEf+WxE2bDKYDg9X48Ep78So+M9AcQ7/mAGELthoLdwe7jwqSWPXtkYVIf72
ymnQoECszdifNkqh5+CG7ruKnXC0oJNUEwRQ0Nl8qrXyRHf2va4LxSi+6VvoXewS9gQ5UetVUljz
JXcgkGhACkUbmQpSNrPwT1aq5s2AmIwKTxzF6Ib2Ybj2W09qa/qGpqKJ8LzMGy4sZ8je9BrL4C5X
7wmoCEil2rhKgCtnG/kQxFjZqLe75whqTGziIF/8KxOfHDDq7sd4WHmsozKUGon8WM+96dyzRZAo
1vUDnTekoWAxq3keajqgXX5EQHqFnn3sykq8J5jxlqLxYRav0t3YFn9h1a8wXjwzT2apzINoAH1D
hdygdrtbH0CmJkZigcypg2uy+91Ey/p8CFzmS9OCWOFSG24zs2ZRixGd4xYJ+njRFpBB7Os/Ow/l
gvzWndFPs1oZr1V4Z2IUnFHa6uI45I8rgO61NH7LacA1NgoTq16PpDympewyrQty2LFvtAVBIuOP
FrsELJhTNvNX7B88WF+QTMII9rcWE8YOogbWsMKq0Do+96pqEMPbK6UHRK6omIqIRuuDQTaL+nat
tyckSZj59c1Oe1+NVWtEnoJTbRdmV1jewzOITTbL/NA4iKeLl6sTUDfbLmX0CJ+S9Lq2ou0TpYpK
Iu1/JhCekKCe6MfodvBCbxh1PtNnT+2a4Bt3WaIqa1QElq/FXet54Sy4iklq1sihYMQb9s4fPxza
iZMRJp3kUs0K9ch/yZ2LAuFeK1tPwD0ECAQClZw/vM7CbeslX651BXoYqDOIgRCJw4r/FWKQ//YD
DRfElaTc97R6ymnkEie+vJHLtk8l/YeR1S0quGZ77VXzIdlhx7qg2HlICMLDp9fG5CJy0NTqk+qG
NJ+nSUu/mG332P0DXs0s0lgzL8JGgr/GA/rK22wsAKs16kYFLq7enFKEIlLMrXHiP1vDKi4WbzvF
BjwNB6xiD9MxY6vxKqvhG2RkUnU+HjYq6FXQA0M1w1lVoqDt+vfsLJViKvpJ2X7+3p3o+8hHCBkl
6ndmvzrXLFSr/xRT9kldxdOdZYmuBSJi5ooEmecSg4TLUFsreK7fR9ekKUkZa6HKLUna5kDwrzCT
89zwQPAIG8oqH6owRT+mhHWjKFLiGZcsNjoL7Mk7KtcbLjGDH++gDao4XT5+3/Jl9gxU+2LXUSPr
Sttb+lSJADs9b1UD4v8hx7uS4LHXUPpQpiAc/G+XSerP3T8Sd8xY96JTqbdw4IETLP9J/kwTkp9n
XCtKbbzPb3LJ49zXn65LK/zpkACVT8ZSTIGn+oHOF7Vo3yj2uaYRxUtVY+Z/xAvFyyntSInfvYH0
oDSwd+5NIdwd8qr2cF7ygwFQ+nKERyS7wdLRfqzMElitdODHgkX0tokJTwu1zdBE2LTpeuoYJW69
Ws+H0DbehtdZikIiZJ60P9Kda+u05naBV99jtxJj6W71xGqG6E/8Kd2kQf4WQ1+DdE2dYf3JncGN
W3nVIoQjBSyMUp2u9ozfK+QDW0fB93OpqbnRN2mhnh4q9CkHTRvI8gdVweWLkzbHm9f+MEh1dLcM
H0NEffJS7Omkuibk+TrsnmKBzWbNlFEXRyTcqBy04v4+BC2beNSN/DeXy3alhjDxCBmoGyU1Apla
chAUeO/YbY2C9L+vKnKIpsJKrY0BdlhEoaHBk/+8bm5EA0LeWRXSgP476J5CDc18z06ohNLQ4e0q
GdOb5k4xk16vOEupKZIxHf+75ABtrACDUcP0DZtt/UGBwXaNitDuC1HOgCeXqiPS/3Zf96cq+/3Z
rM0APJ+zmr3al21+dQXs93Tme7ccG6p0jNGa4r3vk05d19V66wb3TFcuZ5jGrWBFbqScRvRqw3uc
WUZNDTbOHGzpIrLSL5bkiY60XMNj59ysJxlL/9SHKnO2leGz2rDniJJmRYjVn0/zWoDE+/ezZ9ir
VMWp+WLesy5WVoRX0PuC4Mvtc3fBKlLQ9KacXd0AkWnMRmnz9o2MET/+qY8/I4YHIFewfzNZR0SW
+xi4fsq+0DVOhuC8HEbeAiHXCSackM6kYmAueRCP1QPjCvZfTtUSaNyKVrRZ042Sl2HEBPfT9fY6
SSR46JQwQDFDRYlCMG8AxeL6mhqlHgQskgHQPXk6sztZxOnUIElJJYlVnYrmG7BHaGDU/dqEr/cS
M24Uv7DIrt9iOZXoZ2kCVwPUGuPIjFkGAFb8kmiFrgdrBv17lzTGlTjc3tnSn7Niuvn78FN9YJz4
91FaAP/l5nh07d0FiC7dp6rRI2jFSAVzpdnqJ5WO0TLUV2qYA28/6HzDf/e36hVDYPb1MJ8J6eOG
uzDpneHakoztgCnmFcAp66aLtgXC2p9j2TxB9XGX6LUPHoN7U7M6QxCvXVMzj6sxlvWxrJgUKDJS
3UewVGpkCNc/ooTubV6jc6QnMzPhXice9DFq2HrQbrQtxPv6K/HSwQlmt21Z0GRpTZfqxTnxLTQq
qzhSP2826kl6vidadD2N5lFzHdBKrcKi5WX3ljI6dM1YZCz8iU1fnv0LNo/s1HeX6UVH581MmX2h
tphvepI70Vn4xa31AGC/obArzp5HeEJr/yT21RjCwylwdDm70By1Dsv2feYLxpqx/YWJeVWTKcbz
8r6BrcBXJK05Co31NZfh0/Qmjv4uu472qusBuwQ4wqHwwD8WBYXLcaVXxQjEyPHBzupFsqx8++/0
3IjK8W6lqhemxrRt7z3cn3ZFWsyMrEW6bB6WfmQqdtFqhJIIkratbo+gJ6D9srJEVv6qL/AurDZq
qjNDa4PD13Q8xDRiEsYZ2ySq7oZBoranc1dYxHYuCRkhRd3RaHsd37pOjRy5nXI6fLX0xP8MGv0V
lylHmBby+5xi6muaVvlIiZppqwliVrC5hn2FnH4HJKg2GTsnRkOOHz/xJSMQqSDhw0j/OexN+Goy
StnBZyo5vH91pHxbrysMDXZaZ5Wo+qj+9lKj3IraopAem6Pj/zVlZPMsjiy2Wm9yHXEMs1tXHJuR
tFhzp73bbe9HDLFK5UGpJj0INgmBXLnTJBd1zSRBDkJpBpPAFJa/kbCK8OZcdAaTRxxekTYC21Oa
V82wHNpCFVQKV691VqnFyBoQDVYhV5ziGDpB7FbvX6YkBF9HbheXk2cdHXsxfL5QoIDZ+Yj6gQwF
ROjN63YP1m6PG4u5GZM1zLyaC5f8tyrvoWLcODPift9mVsDXr90TxhFMzaV2qsOMfMBFuFSAiQF+
j5cLog53NYiBh0+ulkyQCvw6c38m7HvkkX2ALF1UoO2199sh4izh0DAPxp3kLCvDVihsNwWYDID8
Om27u13N4NHAX4ldPoZf+FKQ1Sjl462lPDufLxlVYMVEDT2i8c2VP/dZYjGUNuVGeYKH8jXw82iC
dXtTKmt6+vpyaUnnNjXQj5o0eavdD3tBYPFaSsJqW+BamdTajSNcaxAAGoelVVeEhp8+PtwwUtQg
GXKAEnYTO2Tf7f2n6J1QssshvxSXZztbPN7J+QYu7mokhsjGlVq7tlGQDlN0XCva09Z48tdceiqc
5ju925WFbjcDoGjL0yGzgB+SyG/u8kP3i3NiloY3zHd3stbzwpijUkF9EZ/qTSEd9I010iVX9s1t
XeDJmPHtIIE+Am4aq3tzDJrnZP7O294OciJbCXNIG7fluyp2z2yUBRoneLjfIqwaBxD89utmlLtQ
NphYhfp7EQXw/B+NMsKTHDkCzoVtqVSgZP6a6ErMZ9IukomWed9JzL1mM+DHRAplt9XkUkISYi+A
IDsGBpgTwdDoynIwkVsh5QQpCLUH4NNdNiz/qx11Eym3ERR7zCA8KhtYTE4eAvIKh6KODFqR4Tok
ifX3lYEfvEkL0atqcbZmvZheJEDkQsNezJZYYwwsfFuHfGP1ySK75wdvPudyq67qzSusj5cFPwJg
BFJcX07UjxzLLNHkjj4foeyUBc8S1/N4GjrIg7zrYpZvCiqUkgMXbanPvmaB2eIHpZwxOTxathki
A9xK35MOh3HhgCRpwyyKD5+lc3JH+qAQfERsmu6EyevrxA25qp9IxvjICh2PRMxvzpsG/q6F7Npp
XdwWNDizoxyRwhRBwWuPx56f4fp0tZ7tMdV0q7yMN673xdlSx/hSNhUcx6iGQNqkOM8TWJmgdkZr
K2vi053mIZCCQpqoLb3e/40nqfvRZzwrwf9JnOzojF5SkBkPh1RI6SVnxv4FRzAIR6Rv2XTlh/Y1
Dh9emlXODD7wdPST3NppZacAvZA9c4N5Uz/808J1qxRXdV2bu8k3/JBSW9WA62hVeLxwR/sZesLn
Xs8McsPTZuHtXdw7mV9fPoVvDUY9Ox57GUbIy5WJ8azOFq2xb5cI6/C2ylTjwoBBC3m8fybOjAC4
zmejvd+dX58J6B3U00t7YI3y8ZVhYyAaDAgeZThsHVErwoAZxTKcB7ECu5mhDeL/bDWilFdczTHs
hlGxmaNiFlLEPuPcQg2wGxdBglx1zgu3nt0vJFeBH0IaVBdyDVHduf0xi3HOz5UpavCUGAWr+MfY
r7V8yvWy+Fj6ra7XhPO/+khJEAvLYovpezRbeZawb1REs5+DX/55NOJ8VsY0e4mtLBReG78hWqvS
YV2vdypFIA/0Ep3ODX0cr2OYANyO43idT8j6wQmYOMNmEWV/P7xH7Kynp/dNG5c8Wts1UOwsExYC
nsPWRGr9Kf4ciRQb+9VdIQTHE7LfShxoT80XVCnP5RGQWUZeQD/o3IKqbKEIQy4TMD5DdMp9yJn8
FsK8c96pety29rnfLrR9lTkCzgnFeuyAKaDhbGJIz/VyDHtiSncrbP/thkdvFM40jt2Hmhz7LmMI
DzKZxL1Rsp0qpsO+q2+19tIBIe4+bbeWcsI9ATLjqpU1o3mCb71xl4GrXGfhk9Ovc8XxYcuyto6G
6gCqIr/4WobqXo9sXtjB42J5rKmENve9a1ir2YgOPT6Lhc5AZLS0An0KBEmIor0X7ST1ScDoE4XX
wrxSRAxygtNMfNddT+HUfYQIC1mtH5Is1d19pAamHJjcIjJfAtZ15tySNvhKImy2GEHSqV5WOL8i
Kp4H3xz1z4u/LIpYEuHs40UaQZLdoYb3g/jORWyO5GIGAcVvFRCAszCRRfwk9z+WVfnbzHl3rlaY
eVJDDqQ6OxQmZwnEdyzVmwBe4duBtK0XkDev1RSD/mkWs1WcDApdA98uPaI+iNRHvo/3YR90Uius
Y0fTFQte2Dlk6Rd69KaN/JqwKV76oOSK7jU5wjG5le8xC8yxst/neO9yatHfu93Txf3V04Hk1Alg
FM9ARmSzZWCcfVFlr/56ywktFx8uiLiR1CuyRhwlirHAasBzJFzmX6x+Qacja1RENBtkEdb7bqth
q979IXZ+56LCt0MvnPtZgortp+0lOaVs8Tj1b9KmTm1zJxCXsp+JQG9upzQ13QSvRd4zfZRWp5WF
Z5g/0bpslZTgHFSm+QBwk//jKzz/yoKZjMWVNMDnBAifNI13rW1QimDX193XPhSm8K0ceIgnRlKi
xOTDBS/bkvQLCMf/jVVX3Nm2u/rV+n7xYtLaCWQAn/mTSQRMVtVnj6FiboErUUNd4VzPmdiOV0pc
WTeoYEVxKx3+g8lka/Iltmbf7ivPh++eWLc2RltNu/47IhLgr6N1iR2H3SEHnZ1FOOBqFI5+8vv9
ejsXh9Mts0xJoOKvivCAH+FN2/QXzfEWW5Gkzmp79s1l0L3mxp9PguNpFJEoV4cXAyj0ZwFUMADU
UY7rLLVF5TjnkUbZAT76omM1WAcEoMHGWROpwzKOGE6TjCgyya1TGNdowUZHE/veENst9zYTEJ0l
We8+5k8Nc6c66qPT2mAJ0afW7BsMI3a+GzFW+qbYp1mpgqmiHNorAIGI4jICQhp96ef9S8+UXZUm
smy/9XpiQB8VN5b+RLdcayZrlXqKKafoao1Nsevw9jWe/oq8k003/Q8F6x5EYqUtXcnl6sQ3kgCG
X0AVR0cudnyq8D+xE7ZT9nSIr5/mx7Xm+jTVc+1xFhyzdxbFGXK/KU54OPHq+LIq9/xm111BX6ji
VqSWcZlaNd27ZbjKnwV1J64Y4aTRQOkoRxjS09PBNKFe4ulSPZlvHN7+muhJjcNMXH25XiwPM4WA
RRO8AB79jTScsJcAyCVwh86n5nIhV/8vX9w+pz+w9NgPyOdJoFITZzmD8EoDwaq1s66TW+0TdOOs
BhJBXTLhbb5ptR+ccVcZVoGZBUrsnlFZpTOBNYZ5QU9g4exP9fFm/R8lUym2qEje/WLeIbDh2TMv
qSuknZSaTxyZx2C++TshQnDuS8MQBRfY74AnXp4ST3wR/hX+s3KqsBerYxpWZHYXqXE64LnYhfGM
xHPXUNgsGTvfxlVuCcLTUiKV2uxW05tdurhrRnXVSbZBJcG3r2RFKOOH6kiQo9kmpWlBgcnseWB5
RwvbgJpjEbz0zSO9yZvD2i88Q3TcTYnu3mHZlqoMdDzRyp/usGl6m1mzufscO+jU6tnndq0Xriy8
5MJDlnK5ZmRSnG/9LJEqiGjSn0407kr9WWHMuK6dnxy0Gd4T4yWS7JIZ8v9RcQAzkUtgWmzlZbp5
6eY707UGrpTYkC53mWUrLuVg4P2jKoj6WWaJX8RNybqhYcH2xDWzGD6gp6zBs2d3/Ns5Aqr2llkV
xQFgFD499ADMwWf1e/TFuGE4y/vcKVSYWF78rxBerO1tNMw2/gepsFpdv0WCNmMPgz7dOqjfLNya
VOLncqvml6Ff92hhFEBeN20rbedzPGce9yUH+S1Roztgu4DvHrLb8i8ru/pgmIQwrD8dx0HYL5sz
8WgSCerGkIQOyTJNupNDkh5AybtyAkTTyORNgCEIZN5Hp0grvCV1/2FoWvojJXWXev9dqkt2Jq5o
Hs0Vm/N0MrnBQM6yjBOmTtnAs3Bs8OZNMq7qhkD6nsRgxBxyYQ3qnCa+6lALAvVPlHDSPt0rbsf0
D+SOIqpCe0e8z6QoQFOH4eZQguzR5vF8M6NqvMTrxsVK3WUXUlf/OVhk2Zal1PUeMoyVoncS4Lu9
8m4N3BtTUFydJpmyNuzrMeqEbIlzDsRHysBexWfREdjfFmUdyYx8WyPjOXeOwaGQ/eJwduifJP4T
CIjGycuvOZxJ7bYyCF4FFvqCeEqzCIXRxB9aXMvqUOxYoF66ElvpNmJ11Ayc6AGFZbundvAa9gei
CSQlsrKJcyXQJfncsPHnyz6kmOxSzxFD64K3YFysXFIpTBqfmRR2S4xE4dUMrA+XppI/i8Kaj3FO
2NLwOrTsPLRV5arlc7YB5LShXABR9cEK0YVGZd/S49ccOENcd78qEjaiA8u2h0B2m4xZ6xHdkGRD
q7Hv9mCge3Z2fWTZOrAZyxcgdD6Fv1kDtqJziVi+kICdGxAJFK7N1QnYPwXt1j+PhrA6WmxxF+1n
bN/sjjsliKGTnl8Mre4e1HzXYpxLhj7r7GeQxyQIhkkx0HklIbuJACq14PEIvQZwlWxREBz7vxwU
ZId6lCYEzNzMr2XsNrPHUTq2oNSR9DxOcviTFBoJU3hJObBFCodY4vvOI633hN/JiDIGXI0yDXLz
G40iw1gYgs9cnjvSaJbi64oAsmuPHcevxatzckbgfMTyQ67GChEv+fmJHGJlSFaszWPskigItadK
PF0VEZ4OpGEnin4S8WdTVk2X8VzvAt+JGx3CsLKMALqecNuQ7imvqcmIW3qe/LzqvbZSnq9IuUw7
X+gg+RHGufdTabTa/TPr/RG2qf7FlCwrd/NsOiHqBm9/WmOerZ2dsvp2YJ2iqekNB6fksqvw4cbu
oMO/7fFnb4Dvh6YJqg6Pfg9SHV3tuwYpPwuO+Amcg2qw7012vmtAJzeqzMVENebZWRkNTS+sCgLc
uZ3VGYNqvwvktILr4SlE6WokSgcVnM+XZc4hQ9anR9d5AbV9ovqLVD29IQINmsUf4b/vSyPhdR3c
BTl16EY7wlgXWo1gTnrz2vlooOh/IoCo5EripSI2yPpBAG8hVhlWFbKgkGrYMCAlIdN4XTWVQX2z
G4GGOk4ZGzNXbqQav2v1fs3Fu/38F4TP0UTGWZBPCnqZUO0g6o65722ywfQH9jL7rTGoxyV3irNL
b3WPgj9/c0fh5ClgPTDcZ+NKp0SPmErvpiUxSkzwR1u7MbaGWqddPBE+pcXR23fIfCl/Cualr9WB
sCVKwBd/ncpT9F24ydgo0Oia7tCSdX683oadTEBjlYT02Lt7duP3+hZKSFqpMVqwZnXcAPnbJtrn
Dn1/IfBwooWZoSxq1GyScA6t03IjZrePwe2zrFn7XADzl3k90NNp4L67qQproGOmd8wt38PYAYAj
ygQECMpf04Ai69ImYNkEtmLoqUaqQX0sMANwxE0fCh0YY2Zan7URK3SI8m3ux5tDvkyYbukUEe62
iJe37cqSq5G1+i0j+Dz3tpgcxK+msrFIHrBrVykc61DDMseGdVT6kyqNux+OXW4EhBvDi7tMIIKg
JZGyirUqBIUj7ULpMMObnYkqPS8ddLodgTDQvoqkK539JsurqRsuaNoAv4M4ZO8S5zJaPTCjSCJt
qRn21/iOjkOahG7g+efLgqysFoCzpj8vpxvE9CzuV+sFUSa8Uvb6MHY+aalIY0yZdebP+lVca5Z7
aMggq0d/6z62AtjKzTs068KZMw0MdCV3cTDlp6E8sWRLt7t6XpcnZUP4r0SrtAN2q1BAaqxYpR6i
MP4brVGVcEQYj+y5Pdis93vqkU912FSk6aONrxu/6wAiuKqHWubzH3sr7VC+1kZT9zJTz0kXqosl
LkfWeXbVPzfYos0gMJ4ohrKYToc0cNsNpePb/BjvQBIAdHzvRNidUQoRmvzRWQwApilziEusVRrl
9a/sbLRiT3YrpcYeONMjcqCzbDdFsZvFsxvBrSG5oKrqWv1hiH5CSz2X7giJVYqQG/U9sw4+lL8U
LchQy5JXpKwWJqcw+kIxIxfRSUVDNUUpjVaboZ3v2RWaBp09a4k0HLluwdgA7E+JQNrZrxbgsETb
fLAAtg6ZZfAbcdTUZYLwLZJ6wWP2UjtyaM9+Qe9z4nuMpBKw5haIXYa+743vwHdaJgrcRwhbawUJ
ZJ5aNujbLOhpZscODy5j8sMlkgAkgRGzN9PE3CyuTGJRv8G69a6Y2H518+a+xuf28QPh3IqiB0zu
FFSM327JCzcXzuDu1ZrAayVxPEbSZtddlZ2tI0NB1o8ztPySj5O1V6hOIkZfAQPyX8GW1pCoadtT
PiXl/2YfuDTYSNJRdJGqCG8OLeGMkf2aHobSoU7g7NW6v6I+jKVeQMTMOQuscgG8CN9l2N+w95i6
0Mp9uiJT2IvJTekR37Sk8FLu06GFzkkgl3qTxnCzQIPneWtY8VSnw7Uez5MhZzuf+eqS1MJvZ0PN
ZCInKZLP1ugyEiyOQIo7l7eTQxQnwLZfX9iSdfS0PFYOdHe/mAJ0jELvw6ZapwZI7FML1SNRL0vk
NV8ro1IKMDORK6P2sMHNKb0g71sumt1Ve+8mV5kNncJq+YGyYJlz2rZLTZ8ddDW/Dp2EMmBC0H8z
dF2HZuF2j9DO+DAkWPXPGs7ecyQgYAEV2KKB4vZhFf4LUajS2ghgbGFlpfmLiBIzw2NtIcINWbjQ
pq3S2II9x1+qEHin9gFQUPtOfOfyxTaw9lE33z+oMZMIBP/uZyLAWmafiSIQngKVRzyk1fOrSHb/
j0URmVUlEvh+SzbY6orU91FUmFdmvkjfMLdLzTPP25EiPyrucBQ9qmTbqxfGzRIFf3Mpa0Qhuhn/
CgC4XS5cV8tRcvmzlULZngF5ngxiMp8M0YcA3/sNnbEPBJNsW6XllguIAhwqQY8A5Aph3ZKGTq5j
UcVx4t1f3olmxZfBQX2al4VOVUXncrT3YIacUnFmQpfLF99NckXVloWTVjhGHrv725mWU1byDsAH
Ke24s0D/ww2J77eVoGlQ+5MQsZqwT332GiQTgY1hMOULFNZTsG+HtAEXzk9ybNejBa+F5MC0oWXP
x1QKDxWwvEClj2UjyZRm4s3boQTBWtY8/eYuSqbB/sof6tc0f7yFpYgmhDzu2dNdMOMhrH8CkvIh
ipMFdbgzdlvDIjToc5Sih27qaoB5p+OPZDhfzcnbF5aNqLlkOqL6uy2GP6p8+dD//97ylOBmeqd8
ptcQWsVESJqVv2cSHivIoIRgOLuoPWe/0owqVBZoqWbTUArBXCnH1V+fm8UdllHVP8boly0YLU+T
wOQjOx8ydsEOADztnuiKEzVRmDVZQsukzzU/ItAia93WsUEDUomZ2pdlfCWkSnu21ym8vTpLfYFL
1Z3mI1RbGVpemufsGO/dbf/g06rgLBfGO9azHZtAHHj6niLrU8xwompUwmounpBj4zyQXbW4tHuQ
f4GhJAyZoqB59U4Snxrgbv9BY16MhawEP8xK2Ei7jpakckC5NVVJAahpv2zjGwN1DcBksTOidcao
OJDgX0ykbx6mNdQw0kPgcWgJRy6h1M1ba2lK/GP+6BZHGN/Hfg2w933NIDXBuF2qKqxC3CaV64X2
LvlisqcsHGgfakDxhs/YskrQguY9nQdsvcEVYfYuDulAdXkgxFCMFBwE2p5nCthAvylfmpF6EIab
LE51d6WhgylzxGXyTSoMNcg4oDw/xhuyxiEcM8j9bz0qY39EIBqu6hV6+olgzClUsuyF+dBVpI5Z
6/4muVJwaY9Hnc5AsTRqK1tascafn4wm5obR0tLIBUtzKjztfTO8tuW9MQWbBPbThsLwKabo4wtJ
gWDLOx3v3hC0K96RfF2OjgC35HzV2zSqdSaQgX8Pyt+M8uBnqFv6zJ/aPwBj1iMlSkz+9ZOpOcxf
NXTgqnC53bxKnsb8RYo6XahbjzB8s/KRpKmVacoDtBuEf/KmmFg7CT1VbDPssTCK4CrYT489f1Cf
8mg6xgs/auaEo5FxqpZl5vOJT9vhKIyAZzRJPLV2qLYAC0+J5zzdfZhcw3FAyNnBJRrl0tgeDgLh
odi5c7cnkcFwRyGIwl7DUBCGJXzWyNUg/2iRAos6WjQncciJuVtt7UiMpzDDnPSl5z/QeK2pN7mP
l5ooMHpeaf/RdUnd7QuCEj9VZr5l9XSytPRyjfpetfV+nRyxX9MoYiBZ+fGNPTUsZ7lUVK1j4CjE
fyYACQozJag+BGkWUQ89SI9FmoAbIBb+lq3MFxHU741xsrIz5MXYZ4j7hF8bX0KKr8azX3R5bG7X
L17TAkWfgxvdE4y3RrMRdw270dI3lNti8FeWSeCVk8LVnTK37uTMe9LTAl8+UMFYRtr8uPGmURA+
i+aKl6Ccajy1GhluUjURBIWQvEy+UJupsryv4uQGRWZ1Kl9J/F1cx1kMFZbbfD92Qmj8VFJHbNi2
v/7y9wcg1PIRWUX16eT6cZ9+JWxnHFbXSwSfdPyM3YnRdQDlVe0S8UQ5nHkxMZMCZI0otgIhYVja
gRN86Tvn7EGsZ63cKAM+xYsPrVDxHY31oAx4fadeBtzLe30iykGNwruTE4wfY8IiQsoFtAFaKWGS
KP3/ypCbz5V6wWDqwIUfe9Y4B9Oe9jnH7hTiYpyx6L+lZnDDwnGS51oLnPJFrsYakudojtWnb9wP
r62cpb6N6uqJHz+VGxdEjqMoYaB8ftixI5GfeULzUXyTEly7FpT9DbrI64EIcF5ts6ALVK6mIYpp
2FDwp4KbULQgTrZIk/2AljmKDJ3/1JuBKAQzQrStoU0WAE6KlzcgBOVV5y3IjSciSo5WdwDpKMlw
4mQAHciNFEFpfYZ6Z5SMYxQ3UTlG/VFq3MEyBolMJi1L1IIExY6qwEVqkMxoVKGSR0JIm1oVQ5JQ
cqwjuS4U4xf4h0T419zQyppiz3szT2If0s+plXtGiN1lLdtqCFIBEi2IPlMHpZZxPaRiRQsRf8L9
sdBYSWhDCQRyqXTgxjJ4+pXYnwSxYaCzdoC0PpgP+T+im/b/Gnz+TTUPOMUDzZGpq4WRxZrMaoz/
GEUrV/9eYtNEH5ikWTYBVBK+7i71uiBMxiJBGMWRZqtLu30lluM+fiodGv4kpD+qOcR7ja3eNs4G
y+bZVFaNY46oSsyBr4GIJLGPvKb6FrT6ilSD4Sopygmv0UFZRAqoJwBNFSv9FG6pLdhU+HU3LPif
5iXvKZBIpXe7I0F/x8Uomaaby/rDNPP4/D5WG+mP8qH2dLmGQHvxayYioOveK0oHSJNrhufM+hOo
Kns4/i+hOzYAYSeYJ5ZDoImABHSqBFwAVx/i1g8i245pXucNZZL8jB3VMDSZWA2Ef8P3+uKzoVRO
x7TZ36uwlrl/8P4gWG0syUoDmQAhgGxPlYRcBQVu/dxDtT06jnNcVH1h8z98t4Me3lJuI88XLi6c
SughnYmZyDQz+kpJ2CuUWtnncfMkeDW0ihEr3PSVtXNvTZhuGuwqY8QLGz8i/4lYzdEfSYcA9pun
oYwIr1NanSMWaMKMg/DtEbXH9QtaV6DWWXmGnRQ2zug2zQsvyWghnd35fCvTnE5PMr1W+HPsfxlt
yMZQqXP/GYL/UMbW04XMWb4SA51OSmSjXme/bUCu8kK6AcCgnrgR7croVnNoEwqF01qeslWZA1pt
/JKsM9a9fvMHlkg3ADsuis4mSCfFU2RD1pKvIZFl42vOZtZN0K4I8KVfJLvXdEyw9AP4iSiGPy0g
cGbhFigM/LPPLrD1URGoKiiNfRmdpZ9A/7ANL4sqlprNQl6aC6hd/chT1REorx4q+UmaGChwe21B
txp4159khCHMGwBaQhcuEnzb2sMEU3ApUvI4d/MsXPuLeyrsID2CcRMi55NC1nGwqIuWMfueqOCJ
OBwdiFfemsmjnOOkzgvcDeXGkvYysuGEHSw0IolR+qL7IiMy2daaSdvYyxAX5gR1xHY/MD1nhyNL
BWcn2bAaegoCsSxU2Y2UToXRSjLLByjUcmD/lt7nuny/bZSOHPXlADlPF0W304LERzGQVJ8GOXuN
ppKR2V+xoNQblTzdCYN6cKRFHwjRAocxzsPJhjm3Kz9O0duILlbsW5U3y7uAcprs80MAVV9K9G3Y
JKtCCKYXc5mt5brTt0FfOdDOGcFMEJVvuol0ZriykbhFDz+xj3B3t+coVC7Q/iCrk7dhjzs7RlyT
D8pSfLtDcWxHTDxB0M0E1eyqUWSCn/I+AESqCUdCYa0sObtQOlk2NdWjK59NtQcdyBHXM+CVQO29
epkDD/hZUI6xnDFA8S/ZKp4R60bHGp0Uvwul+HG4y/ytuBts59GtWbRXG/gZLx+iU6pXuG61FD50
qHnVfM5CGIYhdu4HhxM916aT0zcqw6R2J86JjFjzoEBk7g3jHJ20e/SlpQiXBR2LAgyxA9L/zLF1
xTzFC5At1HyllKuv1hi0+hZ9n3Mrurs/wiX2uRW3xvWvhTj2AOrX49pDK5tcuxUqZ0ZjNfGs0sQ3
4TbwJeV+Ve1wk9J3Njega0FDka0+EOJyCSDa5NKLje55Hpxf0SLqBHLfrRVb9no2v/TUvdSZvB7t
Wg0MziM02Oyokc4PCpPgWK8IocUBKY7Gact6N1tnko6NGfQtNYMf1a9fO2fywJQs45/HIU/YtLhd
81mtE6d4s9nc5eOQVlvn0jX9hW/ddTLcgRQ3GNYvu5ig2eMRf57YFtSfK2S1sB0+0CeqZ1l5AhXV
FV2Sptvnsesq6fpm89wehpK+0azbAsbIgzux1XCgxhrubn2PycpuVKb+EhTj/6ArfkjweBZCE9Ht
ZOLxvQHTfQayJG9Zmom+B4S1w2b3yfLxQZV9QFw/oEd19HAlQF6V5sWR4Sm6RByBwj1nOnq1n53L
3UYBQaZDf0aPS9bJS0A6WP29qeAQyYjoQUmiFb69NvgMFD1ClkmvabEjQ8N6YY8S5hznyKl98tuH
6OMMYIT9w5A6KLBzVIPRyntdFrpvR066hmZLwglXqE5lRsRWBrrynMtgWIL4fWonPydLGS5R5gBB
+huw9P+2BUMjq4nwfPgfeToL+aECxAC+NFGnXS3W2nZ+RMdE5t4Qi8TGpAG2f7xwbaELbbbSn9wa
m41S3B8c/xG8xFwYQ/CcwffnM80phW+jAO5Ak48bDdlUjJV6YpQ29x3nsXPa2Xo9l0P165rWGz5x
qyUoM8WzNlf40VEUCHLOfRCIgCHC/s1w3vrdlG+ncjySh9jFW30CHkRyR6NlK/oyak0yL/e3oPn9
hJlaEqBT0UM585+e3yhIBdSLFjB6QvssGQhlKxkjLuf6ggKfXu5lmLFuhPNnHBNeSTsJnk/4Ht8S
hwRDV2WlWdGtP27SMXXOatt6PUwxiBpO4ISX8/EZJOZ2NH8SGi+4nTUvYH5G6CJPRzGYcnixpnCy
9AUtJFmHhkBR2D6rKiVJI0pYBioV7gWhIVSoLsaPd4uf6AefKQeo06fuYxkQo5TVL5WGuFpNi8R/
fSULFBAMA/DrPmSaJjuTrbm3ByEO7yl4FZOC2u8bNOe/jPJkwuJwUr7aQAT3xtE9noYe4/nKBCp2
oOj36oaxaKtJ/5hEr3F6zfOVHjLKOEIyUc4EsuLtAji/kXPIdiwbEztzg48YcoNgDKleiy1A6qPn
MSpEiVDQ4GfChIupIf5cQO92jaeunmt+gW75apm6+m2F9Wk+ONg1l982CX/NxpWX5l48mY49BSes
QLdtIRrB8/pNSu+C4Y/c6USJLNpvx2xPS0fGJBP39+RO4chlj2XMNU6yCcIimadFzNCKTfCCAwEm
5L3ITpgCiQOTqnxO1yXDeO6lDk1Hs1ZAMncNnah6plpK2QG3GZ7DMTYAVioZO0KovN//yWjvVl/k
zCLAduxdQKGaYrMS2VHW58TiDx0xMjYUFO4/VYSKQV41+REEBh+a2YcJAIYwaNCLm7I9qW6ryACD
9MLFNL4dz5fpojhvP0pEmYV/hLcxXMfU/VwZ8y7PpD9B3JeztKcAsjPy2iIZocKNtGduanhviVGj
dTBzgT71I66PCp6daVOL6TcGbxiDJ1dFeeUz3MeQuCUIs9z59h+DegaDceUqYYB9ptTzk/m639qR
BthCeqT9PamfAmyIrDLJSHu82RvIku6suAOG5j2ZNRfUY/iwPaDPutBvYu0y2ELb650DroJcxSv1
zWHnFoL5HSOybXOOWY0HsrBJVhzpecAZ94NwFTRIxPogrZ/kGYZrFNIDNrmc39YwA0XjJSV+GcUh
cwbvsKPvtYRZox3fLOdDpkOQfPrJz2azRDFZRdcunz0ZYgP7s4tCkW/tWa1w7/niG3q4xk5R5tuZ
Pc0ouOZeQ+0mD0v8VEHm5TFyLJwdEdNERfMb3AFBhqQSPLZsAXt0RbW1WwBTvkgMcxds8rNmoO93
slCZmdqYqPvtJWUnJpQA31pFZEy2pgNhry6EfBe/455h7PFAx1EkjocKQXeuh1U5V2NpR2n+gMbe
RIEhraItTVEdmLeDLOwhFwCaK6iv88qIu2zbofo3RRqkdegwGZDZZYrq4STKeMbIVsRgiVUo8Nq9
crjQrY8fNG4F17nGN3+97rO6Fc+JNVGjJrZhTus4uCc8uMUCsN3FTG4GafkbSzD+oVT2FETrlkuT
Owiz0joZ1spyskBhLg+kzg5Sr21LdM1VSSRvKR9xzjr7MvZIl3TMb5ci28GiqQKcEBBKK8z9Xyri
qm62N5G2xeTQFjp86vuJMptpI85mTTVhDgjk36WBoOAN5z/G/ToMLr8eouo3o9bZmhDHz45GJ5Er
KT7iRHARG7zNnCySd5gnFD/OG3F8cLXPdphD1iLNCLj0wYmksZKvPWJAqPGGNk44pO9pY/6MAhbg
F7FhQgPJ2JSfTHVjlrMPSyjt9n1p4wpOS1fW112f7KUwOXu6s6W7coTWfwmREiaaz3DxnH0UwuL9
H6Hvmv706VZp3hSCjqowNEE18Q805CPDOC/7uHvqNa3Y50DIu/k3up8/O1md0zDZTENy9CnKnm7l
gB7DwcCf2RRI2WB6VYLdGfjeZuUagwCMXW8Wgqqv359soOFvP3nzH21G7DHuw+SfCtfpqLdGoQMM
kp/TPrSoTgKZiErRF48DCyGkPKZkw1J4KAk/ekV4RJI/9EPgpVlSv/Z9a3tQOToWxdD1JdiWlqr+
GbFJ+PRxP6xSbwk4BwIXYUYqb6cnc2FIZlCXMjHF/ED/aS6mqJoYCIpc0/Fw4M+72mNGQdXy1X9w
Q89EZYP+EBoe8a8189MYeUThE3H8cy8v5WzKiuO+RgRSo3r1aBqmAKbBdGkyBPUaywYU3n/86D4+
KQduupCkupIz49jBthDEyfs5L1ryXIda/UIsTjxrUpMvPLquJ6OIUHeotlttQSQ+ThjR3yHppw88
825GRi9oQLhl+14LYMiGVZdWRr/ZA8UYWxFWWCmLOJya8phISvZoWFxTjPekxO6UyWO/70x/odCu
SkiHbG5wlSLt69a7za7ZckT6ywO2EPgvZY0zbP4KDOFnWpRdm20stwsgsXRbcuOXvQSNzmXPTBTX
2vr4qS+7oiHmsACzc7FV6EhyntbUmVQRvbk71fux/0hpS4Iu6s4jANtcpuTSQm+XnPVjjDgU1Xb1
UIwhNoVUfHRof0FHEdB6rOizW6EyvggYura9/OuWq5WTkkXlifgP+i2F3Y9T1kU1FUTjY9jMY8BI
KLz8iTuUVk3uLfZTrCLYlmNXqT3wQN8l5aOe+UhmPkLKnSLWDuXJCmhNg0VAJrNLmeZ1i62Ap+us
GgUf3rnlkC8PB1R3jiB/4lLEGQQN7aQjEx83Ywq6E3dCNvNRniyiM6ItO3ezajClFxlnF8rc0g8e
QItPnF3VXSwjxbuT0YUIzDEQnzRCSUkOcM1RCf4UHoxo/RHMa4P0wU3G24iUsunQrIq+/OpIbub/
YYfaAirST5d1XVO4OjeJwLLOkq3YvTCy35BBZ1TPJe6VB2jPItsMSmVS76fRKeSBJaV0iJSYtiBb
YNhg9cWh6YqA6v3PQaznm6082m3ZqZzF+gTkIAgmzMcNwCWERX2jKkeOXFa0lGOc59MbBJHzQCb6
R7EnvmUIk79JOmA39ybfPSpgZw0wZNQEXMplU9WrKX4aBUD/XkyO5dKcNEbvY7zGsLnMgX3P5BPj
HlGCBySHTuwhpAQTb7oKKFG4TqzM6+HgBwW2mRpZ/QoeZpi/ABoX5+7wYcuzSk9UydlsdmslUCTl
oLkBowJz6cCUZEaGuehbsaSmBfxweyqESYjq8m+BejcXRqQoXN7zaDBtCs6bNMNxqJsFsN5RzD7n
RpQHsz0x9pdP5q8nWJmwORFTiN9qxePeqQeqzoCtHmFOF75uOBeZhmoL1vJGEh+1nL7rtRk/i4N8
OSS8zttAE46tEKcU1Xhtw6Srva044IoGAW8Zl6drZwY9iWd+QCsnXpu6S42mFSeaLDeHFjlESCkN
3wH9t/qM/jLbuWF30b815PjvVxoEy6XI1IKoDn5jmSRNjpHfhpo4GtJnEZlnYzPHgzWpXOSq9vDT
GtISFgHhQjaMj6QPuzx3qxRAIpxPv8aIlkZZ7tda71UEzp+WFW+0GCsg+pk8VQB6ZcPLHYM8ytCt
9MuWE8x0SSKLQfs5Rzl0/+Qt51nCXK6ar2EHfqqwjl4hmHR6W68QiQp1uU86pZRcROsT46boe39L
6PcJ70LcQILZpu6UQzJCvli2wg4WrvrXFQ4pk5V4rvq8zqOdWr2wPaAUgxGf0khhw0ohcjNbQJtM
zj8IJjLW1erF2im9GZEtYkChA6YfmraAH+wf7Uoc9NMNYO7yHPY6QG8dX/u8mUza7HdfHtL7gqwH
jP9RqQWtRzxNbVVtDUql1weCX32oKvpPH0Hl4NpvNik/NPafP1IuivUfcaYvkQzsvN6DsJXz/iNs
hA9kfmkcOCE2im+w2xnn//mRczT/Y5Vm+0+5f0dDuBdB1jtBKxdZxZ3QZVnqqwNClNA+k0yqLTVm
IZQv4U1Xc6lu4zmecxSmNYyBKJxqaM9nFdPmpWkAoTtBKcXB2PxYmpRjI94lxO5kiDfnNJZUGnfi
Vh81KZ668rNWp5cU3kxmYf4eGnBGLdpkrKhbnmh9TYs9GLajS8nJlgfNZdpS4PFM4u7s/abmowdI
ZNxxlZ1DAGh5eZk76m9Xh4CxzOeCYiYcrYPy//3uznAiZULediXRmdMb0RxPvY+xmu4fOcRzm4MY
YcxdxmkVT1BLKHQdCHuwWcLYnJnMAjwoD7qqiMPPYd31TGvZ9CupOsSPgoc9RLTZGB+fzRiYo9Kk
ZB02qxnes8e+q0YIp8+boq+kB1H2Rna+phqx/fk99MsqFQwdX+5IamYnz4R1c3QhrXWkvEduUxK+
ZJhQaZhUo1FlVSvefCPBqHoL+1MoO+dRaW/S+ghoFIvXtSO5IgEvQmbX2R6zwVD2XBmueRSRNQNw
v9dxD2jc0lxpGkD3jMS1PUI86n10DqdSQywB3utbqDI2AgydHYfl/PFbSAl/QEGlyxG3vFLQr203
opwlQ0k7Cf4c9ssoHyME1AI9USF943WDH1P6Rq9bJ1rbt7CfGQOfgpPb3XL7gZNRcjBUZDlVt6iU
dl297MCFLcGTUNBQuAJeEu0fRwe6U1hEk3rbvz7T/IiPXOYTCUfmoZyHG1kJ4j7lRYfYxboSxn80
NvhqcbCzsKTOQUQNipFsUv3RGCIqBbldP3HOmQHVYSwgBzn6o8IIdpr//Cl4J/QlLEvWh0zymIsQ
Rtc2qQcp9/4A8ZSWtli+VlDvTf6mBjjMHuDOwKaf2yg6g7qqY7qm8iwGLNe4LtbqT5v19as11Gqv
EMNI0FdNYQ7WLT1Iqd8ztF1K8je6a2IXFfSUDolMKZQTSXe9TFLY+eARoHAKRHCLwBJBKq3HX0ej
WvNQJMlPbAivPQ2qlND2oxh3Xp71kf/OxW9Rrvnc2bW1ESMFD0Abk+RUp9/HmD4i1ZvchP/Cpx/F
X1H4EKaaDx9lHCURJqkTFXCjr4e21KK04YySTKPMXptribktnvWWfPsw/cH8EpYZ0v3OdCUMQkdq
wu75yfr8CndILs3DpVcApr/QTcD9GdZ/DWj/TZ8wRWo6NpQKEYkEJTJoROpoLiw2/n1lLArrhlgH
FctgjLOTxtO3MVSgCdC9gRn+NRaubyaQPz6GM/aYChRIaoCa9mvE2uNdPO0q/Gtl4rKOaJv/XUXK
o7nFa7U7cJmkfZyvdtol4LDI3uhspumfghUYhgFDuZoC0+wnEOTB3WvLUN7YVeeDYhKYbtbv5Kv6
Tpox2YC9FSmeYKDHx+zDBx8Y47VfFO+CwOCXvKhth5ickeWOnYyDhlVy2Vxt12MP0sqjA9c3AeBg
A2lXnL8oNF1gjwiCuWoH4wP13i0atfMucdVegZ2FdwgR2J0lY5wI/wwBt99Isfsop7nNWTaCXsPC
pd7Gc1DlneIrftEO4ADFCX2s7kIYgB6Xofb+bIqX4vJXXJLMg22HH7noR2QpvJgL7Cjz2GKuzW4C
FNkzCD+f4L/y+vTx31Twan4zz06x7NxLxgabazblvlonqkDP89aFfkNRBzhvqBA8JIxRMXz84D7M
a56wEsZRhEdJqWob5t6kvOTE900CSkMLnTiiQpuv6JgevuzomxdFjdb2svtO/Lm7V+p/IpKfeFwx
PR0lB8uyy6unUBOiIJQQzI8ba6RYlWfQU2CaGIfvbeWqGQv5Voi1lo+5sXtYAOfQhYrS6BG0IRzB
Ix/iC90WBq6wtnzyGRZcjt8EUOdwu5uzBPH48L+3Lc7++vGBToKOKZt74Q5a8YpG6jLPSTqeG9jF
ZxzybnKdlIEObUuucYnvLG0Bsk2c1cFAMPpoZDdKIelH8NVFWVIFDJ2jnVVOtqZvehV3KC3MNZ9Q
GsPtwVvLV0rQhamgW/u+3pemvEJbFSPGlMJENhcHyelk/4cCocsOwSDS2OeU8b6Vmzpavn/RhY5s
aCZe1GZE3LmLGfqXTQyiHNy3XSb+ScYu8ege516kaKLfDF9NMbjtW2S5ehje94+SidZqzQkRmaUY
w7j2MeuwmNmDZEiG50yFUbCB+a90TAKdGI7t1JUyprDeePlmlJksklLcuYq2O1EpVsMRN0xhhHgP
BlYqFL0ofEsMXVGEjtobw8UUSHPTAcMtmjv3Po6JryZly1bg88xz00+w8B5CQaUtkZoJeuXlOt4V
eRUnJrni7b+/osu2BBzl+2PRJjT+g2AxjK1BGjbEKC2ikl26HnB9fJ71UxV16vRUPt+RUPYza2Rz
/jSXhkW5CQR9pGDk5KQL4Ye1xAiBA1lNGR1/Bcqf+eDFuhqNVMvkCN/kNdDYuIbJviIuqAt01MEy
VZBs0OXMs+lL90tzAcEuBlCfIguqnsFnu9rlsZwlOeUVpS2NEw2AV2NGTSfK26FLs4XJlTSztZkk
fC5hF8/T+TyWgT/IlVVuUZuulGMxwrBvaQrtYwv1DWkPUJNR2OE1R46sR6LwwnJtkzBk6y+1esaA
GnIJ7wy5sgoNIWkKxob0QG6x0U1hSj7/S+2XfY48wlIk1b/jYoh0hW6v7suyMIQCKYWR/ScbO6tf
xJlXorzSDMPuiME4F/cBUJZh7FsDCnYQ/yTtmd5boY8dhmGP2wjDFOHRw4x7NkZF/5D3GnnaIsoa
ZWBHsK8qhJu5VLGv3ugCeKHNIAyrlEr4uJad6LFYTL4ZfR6NEV05ay7mlq3xAC6BuvErxmOf2Bg0
5KTeQi4x1r1+M4e2zNE4lQerBoGaVOn/64/NNi3Vjjrc1kCSehD4mo3vsGBAz1ABGPlEiQAydcUW
+IpaLd0fMaH1JF1cOZQMNUgx4cA7AkdW6vELsu+RsCAl2Et270QMx/rV33kMW3ztx/I6AbW88EqW
w8jl1pN755g1ZJAmHC48BIKRURV1SlwmsK5fxnwMmF3OSbmGLKQ0zx6P6RyUeuuYVpG0iMH3Jah7
qErmRp5S1y4XQ2MeqIaiW1jzP52J9gAnAd6PgOwBal1BrbW4dBb/mkyffO4dcm3p7xDe2NPzscUh
31sqDo7r5zc12eZrsZ4jhPvu0R7/yZohhD5Z3KrXqgoYbNGn2eCUGQdGg8Ys9LEORupoH4M76lvl
xRFs7WHFCBjlS1MYZ5BDOgMCEC87pakcYgGcAHh2gD2KuVRzDkyPsh50HcIOq/qoS4x0RnE1C4/P
T3M9glAW6baUE2w34h0J+eSmnTp6gp19LzATR7wC3zzzB9kAerVC79nWJBG41pLoQDd7oyrdHb6I
Cb2icfAd+cW/8+kqTaPWE9VVAusyJI87z4WgYSk4XTPz+qGO5TfGEdz1cu3yO3Ogvt2yLUp7ONmT
sus+sgLbVI4Df8W5nJYo9AI6s4xq8LQSLwiDBeD95SV6s+ZRY06mgFziyh3qtoDuBW9GOEODUCYZ
i+7KMPJoOI8P6m8u/cjAn6ERie6c+V31ha220E7GNW97wScvoPeWLFq9CY/UTTQw2dBh2XTwlajX
N7u4i34gF+sPMJTOcC8y83c903N+xuZQPcPSA/pZb2YTeP/8gX0eak/DkOd6i9f5Sun/J60B9fj8
las2sAXRlr8BoycqzyId3Evyg3Yy+ijQxyQviREuJgs7mU6Cs2NbDGHVwbGN6uBkHzPPTATS7wQN
qPwA97H83yaDE7NhF9gZBFWdBWCqNbpGd1slIWGBTuWELPmqFYV/9Ru4oyO5FqBM2cCxSwm8Kb5F
7hGYw2cav06N/Hn4Umq14NQmIFn64GR5d/HRGC8pbW1OU+wFt33qMxJfiGZG1cstOkcF3by8QZ8K
vzTvvYt5w98IwQt3Syeh0Z4eQXkjzQvgzhul38k6CgSEW2GJcCwPPgCJrLBQckKqoIdis8Aest0H
5WtBFDz27teF9zEsiDBMgON6yeoP0yqSDyz3nzmT/N6u+DxGaWlVUjBTcCqfA8Fwv3Fkw+/uwfIt
tf7JWSERTHBT3plE0VPFANn3Irvl/fEj0iwu2L+37D3JBppdJXsvk+CeMVNQgPI8Dfk5NzbgpogY
/1yYwx7VO37EJh9qg7CSDCBREkUejnjcF0pIEFfjtRZfKeGdUh0RPRIySbpVk9pKtCFiuUlqUNRc
6xvUiyVgskTRq7ZibJ8RxIZ8OsUAmaYmOeupxEX39i2g48TjoLuhxNEjI3bnZBdUodjioscSRO9I
/9hyw2nR/vB6PHPiiItyiOyk9eoBmwk5ZG/Gg6Ley+iFueQz6KoNf7lC2GNxllUKQv1WziiQJEGY
8SmbZisgV4hbtuH3nfNHZghvWuBvtrjPzyi/bZPAnz2jMNtL66mpRAuR2mARchWkSF4/Ghfrs+fU
rOhGS3na0EbX/ZkfNqrGKJGfZTACag5nLflM3NUdqxgZxcxk6aU6Wyxf2jegeDOXet+Gl8XCEpBX
4po+ccS3JV0pgzvdCxaxzV1e9ZIwEvk5n0blxpTOlXmjWiJ/yZne9oyRH2qkRPAL9XzkjIEhK22j
8puXGWbt4RcYA7n0ikSkz/K4f1+z0qBrymZco/xq5JQrRVdvyAFo+JywpVSCdriSchtfkFoPgXRt
mdhq1MFNQYq4QkIO1TprlWV2CZdJVBtTex37rJrJ53mJ2MMaXx0MZVuJeeG4+GFZGXcZW+jbKIoz
NrSgfWOBCIpsfhGdNBwmfY91gZ8rjTuMtOPRrqsMDGHmAjZbwUu0jM/G4BScGHjDrd0MJZJbNxWo
r0jYHKvklJrhy7V+EShRGe2HMYnt16JTqhqmlgjTreYlwSWxxJsg165MiCP/3GtCcDjZCkdheBwu
7q5sJDTNVxZtQ8XohLTiLSbjVHKbyLubXFNuSLydECIOHPC6S4KiWQwqcRQfKiLtGF0DZxswTLWf
qPR5vfxIB0y0WgGHh99T8KCNGMqafq5qRw1cuMF+8ytfBbyxvtYMWPw6OvUj2aDICyps7s3+Em3q
TXZOaJibyZHDCz8yqgfps9q9Mwjs7NX6cLAGNsft8N/hj5sgK/BsNrtrSxHEswwSxS6/b/WOG+Ki
xMaavLiY3hZzIJnkRKx/8rhjfVHm7SlodBx7GGHq1XBCmOgl05y7eaGg1B10FE7dZXHYlHtPXaBc
R9rs6fImboW9IK5xn2r3JMw1mxsampD5BbTT8iwyzDJBbV8Vpyo7EB8NyvQJ+dp8Hpi7GqGWHRqM
Sv+CFtAot4pFl9dd48K7wnPFsOpgYTNeo5gHLQM7ukI0IKQIFxTbgHCW3RsjoXYRJxHrbxqlewi6
2bOm40RbHr26GV/ySjMP2X8QTokeAXzl3yyVeEO7xVZcOMuFoCXCdKep+Xb8kpCP6YSek5TD3yO2
0QdIR1qQglQaoqiPLtXUIRE1kje+D2uQTxQKs9w56cKFWmGnq4c5m0/872/8EZu2ElS/7c9v945O
ZWaxk5eaAHLGEqcjJAFbeaLZXzaVtos1En+PrZfieYRpm3PkdJedm02BN9tOQqTerUKvaJovZJMG
HRn54uNoZg57iv+rVbMoo4W2vydAjkjhFRg2ffri/tvkvo3cxmC6XcRQv6EGr8DPjhMLq9hg/G+l
ZnzqSMhOQPpSoLmr+JUqenLVtZWwFRyf5m7/aotD6jMOTZW7WCjONKfxZX4XZkLycVcTdycbOP+j
R9QAhjnZv+BI5K7fNWKlX44oz62QLD7kid4Nzt4KRlcn8BOo+cgswxmZQnrRqYjvoo4b7sTrO2BD
0skifxjcef72iDjZdlTKbMf+I3V1OrOb90XXIRJRsha8hAJvPH52ElV6f/u6xY119HAiUbk7LSm+
C/t589X67wx5D7nrAkvrpUcm5+8zZi/YrFgKMpbcW9/O7rd5GyKpU2pIYZftZBryQNjAzOSEHcpn
0+94W2wXa+L15ZSqsK/S6X4/KtXOhJJ6U9gLsAZE5DfgGALjjxZXcbiOXt1HWwrkJM+Ck6WmAMtW
9yn/S0CJbcnnvkCh6D9I/4vvdP+yh8d1eb9kd3A5vKRWFufnEoOfPZDhI3AVMp4oCna+BNJ6KmJT
uQBKB9fC1xvwJRpfYK/8Wz3gZ8AtrQrfm+5owdJwpq1LM3tmJZfhFFlEv3fvEL6YC2kbWk65CmJH
DXqDQxZOLRTWs8P9/lioLUvI/lCFyLQhWfKmgZ8SOjGsvSfwPVkgjOlSnsKOAqHqoAZN/s5HrqwG
CVTmriouuXJeKM09SFFIqpa0gfasOfSd3UIUFTjResls/hGYm+EN0xuZZ0wKCJHyjjd1fBs/Xq3F
2Mrhm7EglHDcnCwSYxjZydiQruO5uYqt7r3XB33KzEDe0np35yx2rEHN+5j7HfuuuiKrL31opOBB
afPh1E9iSzuSPdI0x0mRsdI/F2xbF127gyFcEuVo6VUW3TAQrzlUjqjfWysylEaV1GELgGsJS+hV
51x7/6FmRUXmn2O+wTgzK4bRHaPJ4QT1xifpa2Yv2gLbL96Ngrqxhpi28xXUnSmTpAY5Atl3tJLS
DU8LiG3IytJ2cIS/pAQYfpRaiXlTIYV17djn6whyPUTabpV8WlNzzVnRbD5iud4bMmKfkaBqViIX
s1xU0TTGOLE+JYMw+UmEXpW/rqGHAQapY9EWNUkQsjxD6iyzKT88K9jAJfVwL9CSI9U7xlgo0DDA
pxLYPvxx7laiNRMmj/nswIf0T30ha+7tBNC+US+yV2xt/neRV50H4i7xRC5XDkEj0vRjSqDXBxsW
ASbbEJGucw/veL1jkZhmtTpVQPw5hjPwFclPYiltAW7hO6LftS7Evz+MEIdAjrVGV1ECZeUzUr8c
9tdCmCPdmuyTGGwRLav7bb6XlVdQV0HeVw7CyGb6aDzv0JUWw3we7hVCVRyOGrTD8LPA8iVn5n+j
xhvHMocJ4T2NPTusbFFf+qlq2/ee4spK+vOw9QrHDidLiP3TqNEk5K1SrSQD9jvnkvemz5Ja1U4a
QQkEpq0VO+KbpshrnfYs1zQiGg5BhLsMz7wMGlivlIcnWGzwmBOZHwDaYOXiypU2h+vdp4yPwiXj
zGb+2gL/tl02aHDRkFPE1p1T/M2n6sGLbekzyMOZKFFrWX/B4meBAuqewMTWCqEKvFVMjC6fAAir
rlNUcBliRkkTry7WwvadslYIyKjHtXy7IkRa35WwlXwLvhA+vNq5Zs+LitBCtY6ZxGSfMJv8bU88
8pq/S8N2IdLEuhJINXkz+vxAouugaDTjTUDNjZXgb4XIiaroBsOei7Bn8ZHN+CWg9uaYZ0BqEn4K
hsEi5JFciTR66FGHqJcJYbo3wZxm5VvsLvhZv2shyguosRtwZa4c5TtNupQzX7iB2WkDdLY4oJGV
9koBg8yh6VpocAMqPmfIqLYAVHRwcrBmmAVijCtfHowRlnogrY6CTxfbdkffHBqdlTLJ5f9+2OKz
G7GenfxA39hCrY0y61Xt/7P/rVkdHbETS7uDDF+JVVwcdaFkIlpQehl1iUhADA8bEctqmoH+eJ2u
26SgslUbCdN6z8pLVkR2SjeGNl9HwFeGKM109IV0P45tZ9Kn3O4zYULN1ew7V2YW8CXKhkpsMoPR
VXbj8TGJ7mZRWBD6493M52ZwAyYLyCKZvQGtYVy3eTDzDrZHYP30nd8oHaEBFMSnODH8VHdqeilJ
DFknUs7aXLvUKUrS+Tv/UkofgsUa50KrAYHh1Nz+Ja8lM3NBhJzB/kLfO4Z5tUKXPZvogqckRoZt
xhJu049arXxnsdZqWBV16hazFehD+ek91Pvvwqj5LEXnMUdcbuM6Ga3S0LV+PhGub2R63Vxpc+lR
lKtrzjeR6/1t3xjBVatomCwBz5yX0Y221ldIwo2a+0UZCgmcacrXvm6fh0ix3f2sq8dM3TqoRRaK
jqFDzJN/5ONQenpP+KwQc6cy3epSRR6blsiY8pLqqCEXCwnOh9QGGTlbLXUvPnF+E+xzku2DdvXj
BaOFj7SXxaDN/QhFl6cGWozlUN/1YHfyUJEz2tgJlEBCwhXL4SBVmlJpU0yGoJHPQNm0XsWfzdYX
E/dfTomrpPoPbSNIAjeZrqHFG+qhEKbZ8nvQL7V7Lk4nCnN/YHwMAZVObsI31ZdYLp8+JqGteAmN
RFL8SSADaw4Dve7yhjImhx/QLGrfOZ9pa0lXgQn2t/raL0Vd//vsKJJfX9ATsTIuUBfoBctnx8Ak
dQGaGeq865iHuytkL/a63DWFtcDYXyPUyGMIldTdnIrrVwbiW+V8fTHLWHI9F3TaqOtV09q6DFiG
fVSkbNRnt0fWV5HOyqQhk0DdVkNOyszLO73fHgUjjvDD6ylLJ7raX53ceByCwlxrXjlZu2qG5FSo
Y9dQhr9m2+JZVykNGU08H1xb+hB3WNsQRFozEA0eKGywlYOBRINtJQli0a2uOI8XKlrBTom2aiaA
+r2hRCUyGjGK8CP/z7ImpGipm51NM3f1BSD2Ge7AXQx9wijV4kz+RlUC+kmibuC15Kf58DS+U48x
XAaKGju9GKB56e3AO1So/0oR8JjtwjT27VEC6Al+WVZ+Oo6BI+zy8wmWkLNPch9xK/2HBySXenAU
ARz536sUnlsp4LfpN8ZqVdnOE9KqqUIyZbVqDn/xILsisI3Ncx0VpCSzs2ElKW5H90OW0dpM0bjb
oJS3dvcGNnMw1kv+4lj6Ruq0rGDhYJ2QJVxbGsjguj1shK3/jYaBsCYkdBBIJharv9vSINXNNnLa
15jAndy/+pt3gZiwLzeKKaC0N9NMh055ZKc02JjxksZ61Khr0UEOEn+GFMvxiUbmBogZP5MKCOK2
26euGnb4pzEr0TE1WrHoS4VW00qgIfDejpjlvY1g0frw7WeqV9pdZbxGdwLcaxyE+AFuXRqNhjEo
cQIwbp3iOK43niTffcBjzLvDXY8jkduutKeWbN154P5XcJIgdZpNG8snoyDmCqS8Ljku34CFzxm/
qtAD3rr+LrYLUpRaQpAcRpaTX7IAJaRL4qNqKb3Ag5vFeHoBYnLVyW9CeQTsTBRUv2yAb6Dzg0TS
LS6QP459v1tSefaiWPUP36TAyDtWcv8YG1zslWBQCzNr3seT9WAPhMa1Y9XWUa8NiaxzVsMlfbeO
U8n1ua25a0tiV9WeWbM7K1Pwowg6RJfRRaHhPEBuUQNe0CnIeAmk2l+Xf75rHS5VLGtioE2CT7fq
vp1Xd4uBNZ57DD8ZpTD//xOQ6TU5rCuqsJippza+oDqqfShme6YmHde2bHvYR7g50bBt3kNKeIqc
FnL4jwfsx0z8Cs/V1zmk3+3lS9t3o2j826MKFkyW/1iJgBaF2xDdzSEyuQkPlKWuPNAHCImzq/Oa
AfK2OBvbJc+L/OYf5TY3al/emzWiL63lv8qWh9L526iYEuTSnu4bw5etZOPe+9ihxr4z4OW9icrW
+CFd8TuQbopD7in5X7ixmePU3qFUr73CKA2991go5KkSWifjPhtr0ESijPDCOaAZo122gGTF/jI+
a0l/g1fiktZrYgNCAE+u8oMrKHxh9SsQWqxg1lBvER6jxJmWl49AT9g1brK5J5tecEkqRw9kaXh7
9dtfBTQJLDI+p5UPJaigMYYxLjahZTo2wrlCMnwh91AE31hppzLNbVwgWicCMzPix7UKTL/Q3Zxe
3/AVdBG662V2ZLmCXBZi8kNMKaWKaFgeApEaMoEL/NXhIT6SNOlSOI80BhpcLIdHoBIPR0zt6VQO
Ic2GircAxS+PvT3bsjMi9qYPPhK90ENjMeEfP2oc7jFDfDBcV5KdgXpQnIMcWQDdsNSBqiMBleV0
6Zi5pJX4AxYEAobS35x98Zh4u/EnENlCzWI2xNCAuVBdneRW32794bkKGYTt9GM22EO2x98R1D66
ApgyYgi1dPdKjMgYmZi5aqQzw0jgiCtw56Vmt4NBAd6Cz2q84RdwFh7yrd7l4ZIgO1Nh6TbApF16
AgDxwFoa4zDx/eMN6JI7g50PG2qmZsFuSg5uO/axYqxCkktHBQtkPSdhm6hT7c0qFlCRhqDOQ+f3
2wIkHDp+/nDU+mHY3g122w7+TDXAAbqiGMAUHlXFEqjR7sFsJL8Ac5mX4wI2S73O7VMVc8ayt0qu
fPt/Z43KcrjEfsQY1CgDEGEoF2vOWEEEhCwbghjYrmPJF5Mqhj4JPGjsBqaPyPXufnMIfzruTX2B
8iQI9GeWfKf+u/geUxAuKxdekOK6CvCoZ4o959DucO3MgHmE1uQIG0mDDrWimG3bYyk+SOs2VTIa
XExMbXhxY9E/k3C5dqnpXFeCwihOjjTCCbExkX9+Ds3Cha5Y4Jx8JAkuqINiVuIc9FDWZt74XICZ
FCaGbmnCOizUtY+Bv7c9SluO6//tsceMuT3CPlwX4cUXSeXE5OQsfvSGBzWCMmv7Hljj9spfsTIs
ahzSn7ON7yNVYXSDFZA+ZyhCeup8BSkQc1/PcTTGI7VCiTJ9h/IoDMDlk60MsLWmI5AKKEd5/SmN
jEZ4jYNOOsoWHR5vEvAK1M3KRUYIqI7OVvejuuaREr+xR6TnIZz42fe/S+9rRGTdxrqm2n5d2BBv
U1mc+6ACLLlU0OV+HmWSmrTgRrJ4S/lbJsgmw0/W8aotjOD1Fr6FEvjxnktKTDy9QXhzxcxA/bD7
CGygmp2YWa0h36ou08IFi7gpoCLzBKDrOKwL1MHG18DkOXbvqr+4d5WDd3I2vO9nUQzXgdX6wDFe
8cYKoStL6pvDgSMKWgE7V7a5P9PrFVfygBl5FMP9Jnfk4ox6hpID1Be4FnYjmRu3Bt84L+0C1x+R
M6ygLW3fvt+shmB4VNWx2w3Mrr7LsfbcTXgM7tL3Jfg5i5EwPkXhIA+lN1NoSf1W3vmC+v+Q4AwE
YcreJhQuanmm8Cb7Fhr+XkhVvmewjGuUHxA6UGdZyQeUkAq2IKw+qCcTw2hzAzgw/KIJ97p/8/+L
RS1uCDEDKZrlUXDbmcMqky12WD5wwsZWzZi/BbGBj62w6GWPb8X0xSE32ciYt8V1gEJogmJ4+LWw
YXLzEE90isGN9aQuN9WszHMVQ/HXCX8kRQJHqrQ4g/XuQWTR2KBPes16aJUj/JEKYAO4g8oAs7Z4
2wm89bBznTDIVbBWkw8WivnDj0nIVUTWKTkA4l7g3Nr2kGN4W9JFnPKLRkGwLh2XyB1cYQ7cRerV
LVfgRAldR6NT1WpYg/NYyKkFQng26pSbzGZqzR/627B4EK/tJZW/UhmICvjcPCCIyTGJN+GWYy4h
vnNZBRU6BTAjNEBkN4c9L95CwwWc48BsxpCqeaoFw0RHkZAUbGf81DpV2wO1hFdp2HkEx6Z1j3Pt
xZA5nbvE/IcFzoH/vsHOd3YK4R2iFSjiTLROIIBq2VyIwdocAGTW+Jj5j8eH0Q/hGzaQ8l+BtEHQ
/t0bERdppceG7S+K2BGe34M9hGJts2a+fhR7WFCOeQUVqhsRzmBbP6bOv2xRCncmn5bR1LhwCBZh
4Wjd11csop/r51lQv/nbwnc4KLIZ7S9HmsLGJ1PeC0eZriKkRRHgqK0ycnCgdbqgKQ82Su6BTd/B
12IwvnC6FcyW4/W5N3cqOXGqnU4WgWfPGLMjePek/GnY0Qy9IGDKtmwMqqmnLvutCWKZvso824p0
FCfl5TKQcazeYspEm9s5wVQNo1ipq3SKNHSWQ4e3X97kVoa83HbqA4mS18/SsbtMJPHEwyHgyzC0
k+4PgwAA02ZwWUnF//1BKBoK6DS55zPXsYs8hLQEXBN6Ajimz9tkJTOob4KU+Nxx98wpTwHr5OMM
iUKcpFVShYMUMmW+KqjRQZ3Uz5hzeFziILMe046ANAhU1wP8fnXmqeY9C3Uobipmt+q01NeXnVP0
vxsOxT4G5rKjeSdq2VUaYHFpz1Bj0ddhXBSMn/Uwc3kzWFVpVd2C4mKCR1pR//dAX1on6pxtENAV
Rxo9g0/cCIf3+UpkxZOnXopUHGlIbSF6HcCDilnpk6rIZDZXimkta9j0js/rVRYHwExga3rP0eYF
BNdMbSAThuroMd7DnQBXrEKsMNU09Yp+1hyxASo4Nk/mFzBQg1p1Q7l4a0dtZ16e9GUa4ehGc04T
v+IsqSrNk53pOgwkr6uZtALQNAcH0R2rloYVniwQ1yWAabYW7A7U0jaGgYrBMFFIT5ceHtMRzTuI
pDFKiE7fC0Iv5bVFzJY4Oaadvrlq1AecdwHYYpxWgVP52WO11An0mU2CUSCRo8vZiYguVQLaTi0L
PzAmtwnd9uoang39DOlV1d7cBJXmO0HtVIzhvR1Fopz+C1aOwNrDpIvRbfQvKpq9aVuouL2awKJK
KsdljCkZUA3xC7CHf51z+NBJUrM58L9wfBPDhRvrZrQBr4titUKU8WOz4kES1wR++6cKVCCRLJ0g
L+OJ808alRXRTmPx+K62ALyVEmMzxeJSY65u/osxBz+byHfN7FJFK1qa/dQFMn3R1U5DLJgILYWN
gf7VzEGwR8TL6N6mOxmlFKnopAggLJqRkb7J8kSaoKTtCzg8W8L0pdn1rKrlQR7bGiYPp6AdpXDg
rBBGZsAvWdlocvgDtBqvSRfrkcN/1DQl7O0E4XbQLaPS1iwsCRmPK6DqAuSI0kSO98QtpUD/NYTr
uiER7vWvxCEHvaHqmzh4t8IV5utc3gND97vIVsHwcDR5jCptXPmteDF/f8ulcwNjPJfgQc5S0GX/
WIUFYlsoafJzHe4JZYyQ4292s8ks2iTrEr0b7S5yQaHM7d9Sjyq4SoIUSiqSqgSQoypoOBdHZcIg
JHMp9PFj2h4BBZ5SnlA93E1NCRZJ5bRiw2dYNiJwzOdiOAlxx6eKBPpC7OuURycO+mplnECGmJ1s
VpkqedUkqXsm/8xGoUv8tOqbPWOKp62Riwi6tN4QDMwT8ecgz4KrQnIDkM1ghVFprz6xLsHLWtJb
1Spp31lnbEILx7qf4sju4Y9XL70c3oc8gAPrJohRnwu6CkepFpKGuZxMYMAJKVCFWPFUFbDWD9Rk
y/sk58I7jIqdLsjqHvylOjIthMMDUwihG2McmP3oFMozwbzGawo61KqB3z5lFKnVNJDs/RYMnT2x
PCPqYnhJ1Gy1H4DUZjl62Obn9RS9cgx8xo+plpGsmgRKeHCQZTKSM954gQLKVXKEAvlPZ9OQDSDB
nNQCqP2wYKYCkeOOAP7aqrCgm1LZtobNSBTO+MzIPgVZFOi+3q04IEXNRbUtvRzhPMYT1zo9PbAF
h59CjR0HBrUg45cY29ulyNWPBmQhOpT6z9udYOKq1Q+PIUQI6sgAd5NcQHEsj/YfA6IkDXBBpbvI
woXi4P07IotBDU3Cf8dpXrYBYsGJGDgnM741yARZAbc9h05YDVjWQ+8lLRdnOgatzif8pwkK4NeI
yH1VXu/8p2/A4oy1pghr/RF/363UZWOH9/pOxiDascBVi2OO/rlc5WvURBWYqX3iGgdrg5CLgqQ2
TJZ6bioDqdS08B/gCzx09WmvIYmlUJYLm1awcsD8foXbJmB9aXISjqDwrHc+vu87kYvj9Rwch5J1
F41m0xmbOrby5G9xtJfoKeNmwJ3b8htQoqvrEpMGj+ySnMsdTEcNlLSfYqnve6E3cQasZ92NBxoN
m0z+08FwTQa79S49czIdv83zdBUAS3U3yj9Z4WJ94/NLsvBDTBKQasb4RUrzkpm8WL2/Wiqjyp6C
HwAK01qOHyS9MpdRVwg3VsizA2+DEr8u3UbeK0EMyDKZuqH/uGKmZXAi57k1c5Owrf+0HM3TBUcM
kwnfPy7gF9Q+7jks3MrH4Lf7ERkQvCYKs0pvUh2bGva54Xg5kFWwvBUy9csWCTPSFtQbSqLMwjX+
vh+kz/byUX+pVNOrKWLt/5ycM07t59btsAhe8ZaCQvNwtB54diiWzLI41CFPHeiP8f3rRBcasBSb
AC30ijbGk6qvs5rLigaezneXZNW9cMXH+AMAMrMA2FH4IvN9MmRgb4qD4C5MGPXpLv33GT1M6MwO
fwhkEuf6gpKnfA5WFZzIFow3TTAVcszuZeCJPxEb7HRHYExNxVSah7UGuZ56vHh60cWG2iWNGio4
3ho27froOf1302bedaH49zTV2j3un50KeMKpZHDcRjIj8Z405oM2RdoBkDon4caqqcuAluDEwpwz
NaEbDfvrOTjc0diZJmGU7F/j2gSyi4sgN7NutC/EGEQ/2Nf4tWAx+7sxFWg0C6q3RUnKyskp+zFd
dkXI3IWfJJ/c+9mHDxj4vFrAJFEY8wFtUfhnxWGqJFNTCD/hLoWBpfKJAaiaNx6nHJJnIFvsT5Kc
jzgD37rGHCVWEW8OsFZ8DN781lT5NWW5q6mZFQ5QpRT2yU7D13cUrYaWCDIlk7j82S95nWTcNale
CgdFHuH6IBw4FBd2SU54W3BTXRHg3DxxoXXb2Vu415QIoawQgpFNFUcSSsyLB9jHm7DqutUND/5L
pQKRPMofjyubVZImKBj+FqMOnyp+Uyaz+engaHFmB/JP9n5/vHz4maLNkEgFkM7w85AOdMnC7vB2
BCY1c/jC99ctdR3McvNUdlVP34lgZUOM9yvoO8k2/P3OIZ33QtvgBKAjJxTiOvTca8qXAVcDnEfi
IOTrb1qIYZLZDNQ5e66k/MW74I/wzlkNfxi8Yz25p5UiXVzKqYdJg+x1Q0RX+zdPnNsdALv+NT9K
vd0ws9cWePJaykayzrsWyfk/H/YTZJjg16Eil1dBahZ+RNYqi9gT3+HabIL+yMAF+Ed7LCmuTY1T
5cgbasrm81TkwDBCP0QJrCeTApa9azUZxf5oNSHpYqlfgHRxxai2frJdYwYc3ti/QLOGZsqzD9qC
Tm3enVHRFIpm3jmKxnc7/KQ2Pcai/T5FANE8a8HDOeIbK7UA6kYLlgJIqeCYz+tUniX1FSwJZUYj
3AJ1N1phKMdqFTcDfwJ10LCPp+l8+1vrplUOJJrj+PiMCoK+aop/fLqung6pTxJKm/zQ2e4wvtJU
Bw3wKxMWizlf2mmzs8sW7c6FQbAuGGE3PZ/vuf/VB7Ix0PXVAXqdVqAlLS0wbl0yLVt50nAsIQgY
FflAnzsthQaZZrCqugpKYjNxRlqr1BRjUygqaYgsli2zwH8l5NpNVAcdfJVBrgmTwLfxsduOASog
CFyJVKSnpBmcshijFXOrN+1Kzosz7GnJTigaMX7OqS2o4xMpvN7BsKk2K4FrA0piyhzerXNOz2d3
E7v8YhJivozrhoV7/vTRM/05CBocPM55kCNY211yQSD7LtOqnRfngdBkOBZOQWnkd+X11o4Zg8i9
/TzF7PxkPSqC96iUxBzQIJOMtkoEpolcfyhPwqL0saAtn+oZxAWeHp6opNHO1XcQ8RMngYth/SBz
aCeBnxetJMLC1IXTku/Nq0e+se96WJWaNhFPVa1JtLWCHoCoxS6e4PAkuEzt1d3Gt6XddkwK/KCP
NLBbt7GNUAqCeaSWyjYtFaDxV1+XlkljxHZsytmcrwqM9Y4OQIpGeEpWu7uPn14h9RZwRD48c4Pp
3rzKDo2Y+teFn+LoSJBZh3hPNag2AJ0OYpuYW64Sr4ZaF9riMQbYlPsPpZJEzXbSS5qkDeJanh7F
D2ptpUPn8wPzFTvTr4z5KdToIhFmsLoseTGtOeVD7AFiVMem6b2DUzZ4WS+5nThxIjDIJschK9YZ
2hdaLcdZoO0c05G8CfDgLfo4CTPbe0IWnsHARUnIJg45sroM8Wl2PCwKv/+XmSELoiiBKemLzp1H
5ovS733W4ejB34qhOp5Dg475kf6kZuSrsJ+im2UyAym5n5bclDeIgk3f3pxK+LA3qX4LeszCe1Ek
zHnGXabJS+Z4CPCzF84GsPaYtIXF6nqdmVqrhPTVD1Nas1VQ+TUQDGbOorx4y0SL8iXt5lnpVyg1
3Iek0bBNi+1EPMUmjRUt33nDRzIxCP9AI7owP65DDE90pHdIJ6MyN3s0WeHPTuAaXbfVcbjoA74x
ACeunsjwYF4O9vkwmdcCqFfOnGeOOXgoizbY2UDhUzCv4envT+7tjXQQATj+FKcEROSvPdwiZtfm
QlJOIIEV+QHuYVX32cPEul2D4UlcxGDpj+mFiwMuQLTtmXiWxXhJkSr088ete/428nH/s5e8gHr3
/hFb6Do9PCA2dvtstz+VAreouirRi+kx1i2n8FyN7DzYCxsmLmddnaLMCRwwR4kuTnBsiCwPNlN/
NVaeU98vB8HDfFGCvB0f8UEanKiXIr+8W/psngIqyO5ReLzU4CUAZiC8+h7zsPXDlbxd/lTd0CpX
XVEgtCkXE7MWnrCJEBE/WnvwzpemADqauycIQHsgA/pMFiyE0naVwWEcqskFt3HKlEglK/v550M5
JQF4zkK90vJoLtKj6wz8lNZxlwJIscWrrcCv6hmfgXeM54/I8ll7AZtbWWXoyw4tv8UTSrtOJv4k
U32aH7rXT/yz9jrY88ExHNGbLgfeyix3pZuC05DLw7ZDvOZxU685Jx1GlA+yiA6FIVk3d6RFfYxk
fN4wQeS0pKlNc+IRvt6qjKGQqmnRYp2JHVc6imSOwo52AOLZeJaWB0zYZZFEeDKTbJsCyaSjDtuM
mnsM/XEkiZysoUCJzagN1Xoac7G81Ew+R7HFQ3OIrevAQ2L0py+dwyLxTOHU9BPPd0trSxVretE3
VoFnxJp5ACs5jf+d2dNaCZJmMb394AHNI699DmDapFTMOtBL5xxPeTorprR6jr9qUAXEiBxkKTiN
hvIEjjUGkRjCTioV1MRHqjSBkplymT/32syBlRi4lkrc+xxYH0AyOv6Sqpr3sUXrC0jYlzKQweNr
TkRYoA1cUFqQfWTqMB3lYlcjMhTxRIDRKbuxtAzVuqcmSYCJs2hY+GHJojaEa/938PbPw8vetJtX
T1/uu/YvQV1ZIx6BCwhg1XddlazTEjQ+ZINrYkl/0mjXOOdyOfdEyp57qEmP0hnZed0dvQ6Db65o
CYB0sUxlMqg9qhQ6X/4eTFKVdmqkz5WveZeHwoS6ircv/HIOMmf4MWMYfT3r/4cqqd7WwydcNOwM
GvvCJTARZnlooqVSVwt5hg1X+MkxS3TuCNRRJiDx6Yyn2+HYuWv3qZw/+AZiZYaGFMltg2hhJAjS
ZSIxOTHEr2G3ETQCBV1d6eoK/DsAyWXRT3gVMqKctEX6jgSd2fPLODK5/vka2B3Vn3Mix+mwUQgx
0rWLrUV+A2HuK6JufrOfJxxU5sFvpOyNq0hFRxVTzn4V+YkStODuZYTG+lR+ygyyj6butGW290hM
ojVUSKzeDVH3mY7Ojccr+zcDkOdxW9KjT1XRCwDkoFRKemyZSmSQ0SWCH6krF4lrz7m/GJuiQtur
gihDflhKctlQxa/0r4gEahcGvspolJvzrCo61VhrxdhrAleLf1Kdq/AjpIGsEPHCntJLs6aTX5Ys
LE1T67E4rpecaRK18fGgV84V+K5pip9QdUGB82nek+ZLA9f5g1ropqnoAE2gEWa8stDGD36ZPT30
BxeeheCo+ORDso3LeRzeC9WWcYwKer1Tg3Sxe6gwkvFyMtG2l5nePf0Z5bJoBDAybLUgz8WTipGw
kcUWKqZVerFSrsGLvkP7zgYZ7sSoS7uX510vDJMl1jgWcx18H8zPvjVSQPRhqhy0QDr7LzfvCXWx
VrI5xPoaM2ZNqnZ8Bwsu6j3dHivkEFjsFp8burqAn1yMRmGruy72XwexCFu3UMlRrh1A3MVZrPJq
aJhYgrVx3pZSCHoHfQ7tVWxg+gKJ8zU0NLzM4zi6GzUgvOoIJv4ClLZMnH2qxhr9VRIpuzeYtH/A
PP+GZYFXs4FVXN+RUyQqTmCh36fIf+fFmkKDt/2xCP24nlbm4aCjMOr2wAdk2mm6An0OUDhZijK+
a8MxEBncuCmXaAIoXEgVoJ/NTIoyS6/XhGM9Ul1fqV7LR7ER+z82rk33htBALhpQJ2fhtGP4fFx8
vYrM96sr51g3Dl0p/neAQb0ZE0bYOFuSlqiWO3hW+Zu9/R6hcevXQtywkcOTtmHcD4AI8sSiPEMb
k1QQHV+FzeP7NJa2czkoPhF0gnFXve5KBW+mmp0SAC3Z8pJ4IPIX6p3wg/d0vbHY49j2rvTUCOPR
tucSofXOWRbdot7BQwJLbvJm81RKMfZkh8H6bmkQbsQzmObikzId5+Tm4aAwrEtU4nMtHyDy8gfl
Je1pJnwFijXOwhiPuLNDQgstruVw/X0tdN1+HPqJ/Y6b2M62zQB5+tbVgIGOs8maIWo3rdmykTOd
qa1dUcTNcjUNo/ulR/6eDeTgH7c7DTNnKbsd9Jt1gA82n7H1Wg5xl4I7Yf2VC2Zh0W7r64VWFsEc
0pa+xdvJEWxEkyQAUKMreVEs8tceAqquDeVHVgbG40KQUz0doM7uaC3NE5q/W2MKG6472qialjsL
tW3N4qoLyteIuJ5VmArF64PEj9k04EYLaXhCZ5RaYf+TmBkf+m/OYL8EnkMB9swG0Os0rqnEa0rK
I9u6Qev+BKBArer20c1BF26vYwUy1YiEfo1ne/iBFbVhfx/AG/QzF7mZYjLjwwOoEU4m62EW5BGO
wP37CN1f5BMG3+QbEKGSjr8Vis6Ms/mOztff/uM77yQmNkBMoLcTv4LrejpvJkjbg1IDUCtcol+g
7FkEJf4lgPOZ5Er5o96SYpqMHe4ucXxGiyn6GDWzLI9WvgAK3H5XJDQS32zk5+l3AVd+W8+bVWeO
l0BUG6mO1HQCNQeN2QVpastxluXnNSI4ISP4LeGYWRLPCMVLxsharxxnX/7ODFgRN8f0JAo5Mi8L
hTOnNkdtRU2AAXHPzj6JY/GLpByIUU++sLKrl5TqN/G1iter70w6sCuqPdGGWqlgVdU5yVfK5g5s
VNFlVWizmPOqC2XtsoKH+5pUJmnN9iUb3uSKWUlYsNoElqYlpzvHMlxeMjTOemnj/QApIIMLHugw
yKyU+W2unEB3GvjD12ztn3roJfIon5fEkGoELLr4l3gxq+kNQnN8lgcHdFgMoiMHjrFeKxn5srVu
mv4zfj/26xQxpbUjG/ZsKSmArnHucybSeyklZAgdBq6HQqGl2e7eDdVmJzbWObs9ha7prsDEYkqC
g8iAYIBhdPJ4T1o4ABmDQdP1Z15oPzzKPiUvw4rLI6DezN7Yi+ro+jB//4T3w4rGHX22vfI6aDCW
WtEJBbnkUuu2QJG/3TMFU1hL8NNGyq0tt/CgWeV4Qzl1Vv6yhdgkLo+by1Hk5HqbClAOfZ1gs8qV
oZt/giobSb3MVMM5YJ3fdZhfvylZJSSvSpkmblWj8b9Z1HzmWoTvKWojpFuoQKvHgYrk238ztlCf
KTx86+Qp5a7DIwt3gguSgeEV+sMPdFYoBfjs316+w5gXGL+bKHxAmzU5AXn6xB2UaRW8ChwUN6V6
0TyPy97f4LZESk/k2PgjkThoIMOZZbc3wVH7Bvv6aiqkESOhN8SnDlEUYdor27MVd536T3ZRFHlZ
BWTwZRTUM9VonZNpgJY4h2a4qagynLXXtRooQzXSr+P+3X3H0sIOlLR7gV8WUUsqAtd8vf090dX1
X0w3BOam2NNHtji3JFWTRc5Lh6NwsoFJqzu1WOQKWfPn9wdZk6SLI8qgkBGRRDevwsC9KsD/ZpS7
F7P1zjgOWgCxvcnRORMHHJDa7VAKv9bl5zXdJcjR1+sIFbNDikFdMWOFwgKiucPXtwmCPCY8UgUF
mX60WTO4Tv4tiZ6FLaN3WfZU2mopkzuAAl5IUsIVCDBk8JN2+YuPJT9A4ntpIFre/Vh2U7SvnRKt
OB4cBjjCxUc0i1GAlYfxxjBcBfK/Hlw++mHjBBryJ+ChfdvSft8VOM+xUmn+IZ3LzocFiRUeKIff
y4aZBlfNZTcod6nRbK5+bkjS1x3w3ekw7elnh6D39Gc4abU5gGa5KNBd4SsOUO4zDR2rg5xstCvH
5FJDpzAJRUeJOTlqc1EAA3FTmCJDIaBEAEdzIQmhGjDfLBkTy5qzv8BA/HwbLPqvIJUw5nSSQMgv
eEsT0fnETajbgHM+C8hzoFFOOxlAEhm1vEKNQcGptl2XCxn0dX8m4Co91+vNvA8RNibqzcg9SEBm
/7AeZeYrceNpVB8QzlpB5EqS8+hPBKA8BG2T8+9anI6aC1cb2BEsth0bE6/npuDVVlldt8qDa5iJ
PKiao4lbdzmkYKhn4R+3rGa+SDYRCXD5y/eeimMovG7GJhRlhL5MiXwx/wi3+oIrRkleXFDCY4wA
TbZwhk6EGAyf23Gnng6ADrSCJWubn2x/f7C0vuRCyO/nFAI5a9a41E+N+bVep1b9buhFhIW8wehp
ofQRaYlRvLV/Da3/RIJfbb7kovk1IrGGiIvzQjnElXNorxShq5aIfRbPiAAO62DDdTNldJdkRevq
agje1ZVnpG/EiyzjV7L+u2SGI27HHJ6GQJ3sx9CLgeuahXU7fajj6vAdmcymPW8CDtdMfkORaUm/
CllZ+e1SKk6fgM7OfQABQt9G0w5/D+Sw1PGz24mO5rvixMHGEs0NDJoR7hC+8tar5Dg/FkL5Nv/x
H6cN4pFRuQ/kDjCn8cQbPEvghz0wIcUNV7JPJuN+p1bijhSpv/GJiSdjghIdCV9Rw7+TgjdURCej
xniCfzMcr/nEzu5dztQpL+em3vId0rb1ahBOzpKKKXP6qqHnFtZQIl/Ohei8tiX8nV558XF6nqvs
cRmwSv3ZRjqqZIuswtDkGHgNgYbe/M626blbaTXXzomcKLn04WeFLAH191d9aL06O5tg1pED4X9o
P2tMJ/b056xAh4Fp+agaETDAR+J+70wjZGRyTVpxGfj6H0O2gUmYavZUMe3QZ/FJMKgBcUPWM13R
8E/Y5METqBRmTgGnBiM91ks93cfpQI/hx7vGpy/huLoVOd8dxX9jwdSLXZUZCxWtofsthSbKoLro
abzM+L2AOTBwSfUuWRorRp8mQKmvXx4fnbe+Sc77lZ4sWm7DTeHXVa9o3f2QwkxJ/lvoly4vKcKF
HPft+LrytehQtHoXLkb+cU00wnD+LZx9lj9FymkXBGI81c11ZJfrkeR2NLOK+4sd6IGcmnNB45Tl
M+phguVgDA03687oZSdBabaPREZWRMfVCT3rFq7uK1V2KNPV/Smk/S6i2BRZnoSebyOTfOxK6R3F
VQwqCR6q+3KDnzX9kJ2d7ptsw4iVYPERS1zXz1+/xnbHUFM5qx0KUSv25XSvqpmLe1AY49IsKX4r
02lzGocM3uHC+Wvqt4k0AOSA256m/+iTQuPY/GYSIiQ8thd4RtufVxkxBaVZTZSxxcIAn1T9P0Bx
ICKmmkIUIXJtPudExgLHAv0zhIjzgnu3/oqBfO/kqOa7ExOd3tl61g6+2uyQSTDVrIHv9ni7iH1l
Zefnk+BjKPpIFS2OLRw8VDI+VGRbA83VKJWRe7rEc+n3LN7ItWUvH8Ott9EgBmwkuFy/n6/gzji5
rho7m1rth6DrF1mgzIh/pitJMFdZI67WJ8zgXJY58w20Q4KjMG5/q7kN5MWmhY7uJ3QXi1svlXNM
/48JA4GoIdXDSpFP37XeLCx5zZb+lJb2tFg+3KaKGydJ0bc9iOl4owaKg3eQ69QnlFWOBHtL3tjz
mhLxh4lu72T4mVrDpzsoQ/uSjgcueZ0P3n1ZiGtd7PrkjgJdGqfcQwYKJvA9WK7DpCQtZbc9/M0H
MbVLGKvdAI+MchwZLFDANBf76nBoSG4AqQTiMRY+3mFb5v7RpiDdQL4pbL85AiHGvXL2TtBaqnoG
G8e1/TXI8wMC5gJNz6Cop5U2rnaYlulqkyiEdz0mtRundjtZZ0ajwPdzB4RGqi4QjNt5y7QjOOfu
ybq9RVE+nNXjdGBd50jWYAvQnK19beYBpfwhfnji0esXL2oGIVoRrK5w51cjZ3Os8twfNiXzSUAE
shfSxLQklIFctY3BLg6qCt4GwWw8bdzldsYRVub5t3oeOul6PqOhqhw7QisiY7zPcD2Xhn2CyDhZ
FL0pelcmB30PCj9pwb/mIaj3gA5YDOEwT8oCtqB7J4sL9Y77sUWaiEd/jd/9d7mQ0ZTsHrRiX2jh
ax7udFrQTxzlGgCmggiExUqrKR8mqFeLzwfZXtVCDCmmLOyO/iOn/mMvIGR2AkNldzIrOU07AYsO
sy57r0y0B8ZsVw7fvSqGjouWxechTcKcOJrTo5fIBsvEGv4P/nfeIr3bcCHr7DuUKJ5svKnNaNfH
sR/oykNxFOl+0y61n97eyI+URdYLHaOr7UC38JwCCuI4oFEDY2C2FDmdTaCz5vEgKA62rvGTW05t
QznDAJFK5vz2ScDkFwP/pSwnE6e62a3mwDDuL+N5XdH+xwQ2pbzPWGN5X+K/2bPnDh7E4zC5O9Mk
3JiJyj/gUw3AfEyqystwtGZksxEKcp+Qhk+oQzRLGpEtkBMyB9E89v+fp1xbbPPJBvt2QbLwyQhP
RZmWifZlytoWnyf2DZMvqwed9pggVTyBV+QfxquGEraN88zFwGWwqXYbNMTfE1aqp//kMKx38DZI
svwNAFdEh2MT0MLD4/JhNy5UeeD93QZ3NVHc9rGzzjNVLjVoNkuXGYWZfbO10xwSwx+UGSWQ0E5c
Sx+nDMfB2tolaq0S7q2MZCxj11+nLUMQM1SVGprFZK9jjpgF7OhvWDLbDnRJ80Se/8yAh9fVe3CO
aJheGEvR+eVkdTcd09tY9nkvGxdd5lHXKhuZVyYwtnfRTWihP7ndTuTlFaytnc4ai9F9f5MAmrd6
dhAmyZERQNvPnXnPGYsa1sMdDHDmClD1vAF1I0wd1y7l1FEAkOqxoa4RnHAMp4bG53kNnxNlLxXq
2JYU27zLpENlPmZD+I40wK2Drffad91BiGzyCsAeBHYNpHjGFWVBFHND4cDLXCRZ7OyrcKLyJpvA
oOxK14mh9ITTMpUieOZpKBTnObL8Y6/WacWveMybZY2JzIaOJN0isBLfUhZuEp6quZWyr2mioKYp
ibTE2SB6JMNkHZSloiPzZM/9/lu43EynkRqFflHQ6iC0BE6VTtBktQP5A5+/pE4LTt9OxVIah0W6
zmbg9Uwh2BracZivSR6hLesCvSqGLKb+R2g3w83MoPi6285CCcRjoM7MU12/gC1tiKKquGjlaF7l
lvjqXzRgTSoIHxVJE5coAEwoaYaNDJ2Gd68ob0pwZ0PP3j0LFroyVBVBv8n4rJHQmMqxdvdfshO+
0Nj7ExPzy1st4XjtjOicibHAY0ks/vuylgwSaqfcIOKB1FSRGdibKP0xiLJoc7BBl1uGXyIrOwJg
SPgbhhGzQ9/vHFZyFFgum8N2eVYKth1WD60CSveyLiTTQyw+Amz04qs4W/2GKL/qadu87M0fAPRN
Nfl5sVRDMyar4KXqZz3eHQ3m3kFcFB9KilijnnI2ZvD6xH+SfGndcES8dhV+iDhg1nn+6ySCKG/q
tahRkr+msOTMXSrZBMHPGNH8eC8M23rOUVAr+nr8bNCxHQbJINGminFKs4NnyhQTUqXBWHelwhlP
ZRWRBtuPjZKvz8W7cNV376jlCkgObDH75Nx00RD0GY4JOtceQsi4kumeq9RWpwt820HdPMottXh7
IlNyzWMR5gkaKUIJJa+WQNlWc7TrIDK9uAdFoFr4VOG1h53EKyOBIyXP3Y8jl2SlkbVAS8csBHp5
T8yGY6wYtfDZpic5XjyvqW9j0Z1KobC8CZTzOnVXMEaLOqCOyvE5ctY58JFqizgMHBERXD9tpL2Y
UHBeB76y0SYgo5zLJ8CyjXLUN5u6iMvO7sQjrFPbX6FRLGRuC97782wsI/8Zrjvsdi/QhxvgiHR6
Hs6MCj5wOsZ4vl+4CRKYp+ZMYX9sEs2qc33CxnqPb/WWTO4aGfNhB6hwyEOex5GiewXgGexg3uq2
RHUuzzoTvXUv62RG2N4OMJsosxyvxSKfULyhtoUCF1kLyUmh7+0AUfqkjWyFUDwhGryrpoIG5qtH
+/e0IqZDDfhooXg5yLdiVpWnFC7N/6Azf2nslBSwdbI3vx3MdBnzgUYaDvyRZ6kpJPENpsJdkGk9
Ubl7Is/i0WG0NxOaGYulhW9zq1Mis7RaGMzEId98nUtSMoNSl0f+Y4a2BGJHo4DmUbeR9ZwP0oRY
Ejqtr7+cH099DXQIjb26ZnmhgN6w+L7MF9ENZFZp8Me//wAvWkiCpffLO8lXKFkFZIxarE1vI0+R
XEnF46z6bHQmlYNNaDVA5tU/PDvOoEGlJEePIHLDRxoonXWmFHHCytagZMb+Odp5W5JfB8Xp4hd4
ZCcsbuG8NO1845wpjvJ5fN4BzwMUeQSKbXfVmGocmoaRsHP5n3H7t7ygOcqJYP1WtujQhkyu+gag
xzGzUc9VETQr5wp+ilYfVBFuWzN71ZWYZRjNMx5f/+adsvbzzZHdLghWbXA1pdpJA7T6bxwZVox7
HgUHpjAFMZMHRj5oTkMjFRURPJ/+Sv2+e/QqL88+4YcZa3pBdG/C/+SxnMI8mjlDZQyOSErAHDsv
nL/hwIp99MqkAObm/YGS9mOw7gmx/8RFpzsnrHVpMU5o2ljap3mNP6QU2vwnsJnMgIBD2/r5Ia74
MJMu8g6f2zmyFSfBrl8DQ+w80k581LISfJcn0TVbrJCDmTiXPShSNg3wZ8OQyYszzugWih2Ys20q
fxeoEUjs/WFA+hA0L2aFA5odkFs7Z2b7I4vdxDujGGJGOrsic0BGBSagvHD0YNepTdXHrjRaTOe/
XNZArAWaanFeL3A0vzVMHMaQQIELdj2ahfAEzHfdIOMHT1Md2KHTKIWUULSAbz7Vq7Xg63AkuAKW
U6awp2kGL/MPx6+wdfg3T4Iwcrv0yhuQpLGOHhZX7M5bBbPdDoYo749VqADVPcKrHKahOd4WIYzg
27yc0THoOvP371erxQhlD8Ucb9sc4X7BaQCSgH512MWziLNjaxaSRCmCPiTw7mn11j2EKwOC7L6T
ZwF1Xo4LgQ/M9i0VletFBuFDHupU9NOL8AOXCRFxEHEB4ZZ9PAP0rARqgk06109Nq/7cjChVmDay
S+QgglHvmrcGfRBvvMQbA1vpMVCqf6xUL8vbK2Vdd5FZa3U7xTpVcSKn1CtXRo1+9baZNMvS6nj7
z3JtT0KESDHIwvfewyuQ9oHWBNEo4+m4E5ZyQByvwPQXuk9xYCJcwnbWz0xOsmY4lIG7Ic3xFPaD
HcrePEbGCiUZ1pHxfTwtVfqOPMoSBD5zVQa55I1GXZcV13AqudikpOj6zMj9JLcfGl0+MOovg68u
GZ+2nSbMQI0ev4rwuMYEAIgTPMi1A74tMM7ISAKJPqAIgX7txZNgec/erF95ByIFnrV/SnDWUJut
bzcRwUFVjzUbwwHGTwZwl+3fgOrOhlcEGuIERp8YOd6vLJIJfO8xHpEu34e12GlJEZMnOde6+Jpb
/yKhfyDrFVV18IggD7ZzhkVFGXijJM1RVTMX9Xmmj5kIzePxWSAfhYG+VeqG/NDPTz/qrymfIUCR
INI7W5oYUuKm1dd2y7el7lBAbil6HsmI7A2nj8DmACAeQxRPFDHdcq6Dwz0i/AKyzJeFor0jhSmj
mTrkmwojarHmkGaatocwo8R3fzxElD8upDOcAqPwTujxrwCJ1E3RuiDmgw/Z2j/HWcbDNBUPiEP7
k6ZXeClfa1qIn1o7bVy6fYmmZzmJsiJntAXX/2vWJqBPvSufksqljMpAhHgyPpbeiFQJTl9U4CIi
BmwTskLca335995L7UMlul6PYJWpWwuq1N5H1UkCIQj9OpD8qAJAX7Ufkd8thUL29Bo/AiR1qwsg
6hAuDq7H+K2UPlnkIAnfy1mLMOpDya/0gbAUubWsL/kmoC7t+9Dl4DPVu1ZoaMZO0oTfTJ0KikLa
8GSUjIrxa0y8rdJWiyRreGENJ9XImyHcX+2GC40+csZsTHNeWj8cFDPBWL7wlwXd0p421aD3aPh3
V1hC3uwXAYjeTUbrqFSK28Vk+pTqwQjVH6kiJc/2w/fcLd6LHCKmBthlCskYxDX8zUW02NZ29m00
fIi7FlnzFpSkHi9Oqu3yBjyhTfL/JtQDbJcsrKlQx7T6EI+hSNQX3gWFVH3Zt8tLqpQA43p4KTVj
1+W0g61f42nHS3urR1fZw9XZ+I+BzK9anDJmHO6z22eGePDkT+fKlLGde2q1wqGKRmAFOokC/O+f
IdAlSDJf+ag+hJLSv7hPv9c8qIfuPOS501hTPhKWL7uDou/WnLfiycj6i8+RRzVIWLyXqbm2Di9u
sOZOtzouEcUzpCTiQCseEG3NAPoXnw74gVoqL/oPS6s36AH81D+aZ0MjpgzX1P/ck/kydteJ3QVM
UPNqFuFcg8jOTbmI1rAtt0QC6Ixw86saq0PFTbOVfV2wkztTSwqz7vqfJmcyrPuNqVW90RaHZVLG
4K4Ei8TgjODag+SG9e7Un0CaO64We0endxbs5efAKa8LM0gdEcNAVix0DcUR0lmnxMaYqoDTVX5k
BGKpg2zYzaMFK0W4M311RoELj0ATCg+qi7T5NUudIEMoOiCqEyTgbF3P8ifSu+uRt7oATNIT5aZ1
ufJnso3yZEjhTdOYbjvPP4DvaakVR5oqj7LqGanRxWhX/oFZlh2eHlbCeMV2nskv+qoV8B+wqCdx
+CL4CpMuu3ieOyFhf54SwaqzZ2iQ0I8hRjX3foDMw4kQij4vNTok4g5Akn2r7dcooKP4xlGAlk6y
Jp7tPQ/Aml+RPBiTHQ+XnsooA/avaaAdyHbadv/zzrlAVzPKdpkBAm4egYP0Q50rjK2v218hDdMf
Q1aLADKYtLU82jxonOv7lGpbYsCA3HpOJ529hcWZH7Q7IC8OH8wdmXweNF2ldMcTB4tY5ZhV7MF3
5Ms0VDDF7RKzxgS/faqHKQcVySs29waCv2S62txbKcuOZkOjQJM/aCc0LxKrNsVm3iL+XDqYP1mt
fP05eGMppUVUwMGwQNCsU8SwcuTMylATCTopFJejSGb3le1usNVRDEAUeAnfizEJwa0s+u4z59AI
MnCJpWiPMLIFphLXhQlr6CH5y53r1Mk2nSXD1GkefVAZfQs3TyzUY7+G3ILFgBD2m4KCVRvmSwcE
s0DuYpGW7Uci/QwCbs1jRxjd/E9Lo5ErS0pK/8AXjMehSMugQHW35cC9NwRqJjZBwPWnWrR0bJ4e
1DJF2s6kN6YC6DZ524qsdBzr75DK2/+n3b5rb3eU72VjOUxnDw68qm8ioo+y+OJc22LhPOLwzCCS
/Uhyod8Xy7vYIPsUZQ4YDmR7TUlqNq8QG36PxpoA7cNxDbCkY+vZZ/ffovRNE5g1o2Pz1NFbDZqQ
m/jR8RNkxkkKqaYSQ2pvG2WS77IVZrlEGkpuYFYrbRah7tvjdhrERHFrFgFYKQG2yquGbi/A8DSD
Cc/1H36xSA7Tbw4IC7zpqKSPBaK+6HEJ9AaurgyxiBiRDT3jjvrZhNereNpbVFIPZtDtAxkmDgqJ
csufeZRfakNLlla85GFlpZNXZ9bAzP5espSQd0+O2MRzeKuIEfLj8aOtG1a2WySJZGCq7MruclML
iksB3k3G4ZyTF5xeWrtpyKV0X+qcimwX/MLXpkWO/fX2VNafHVyV/af4hn2huTcqMTnqAAzcmckR
kG2BI8/jO9jNxmRayAZnz0N2/D1EVErcSuVeRDXTL4FWLMaVsCr4APiwZuADhnGYxYePHZvMmUo5
+dv9lTLmZyZdHcTiHtfMeOzsGxkWRch0Cf2xpGgwf1PvrpwnQtas6xQWHypvzSVP8BgYkidBQDUx
3f+BYOGY4EKX3Ml91UZyHrcnH1pG8uE7kG5TnMV057juVLCjFHyQ4cYYKXlrGP1OoUtkD/bdTcMY
F2NNdeHYQgf3BNCAx1k4RtnXdoaMcGIb6iVPpjtLT2XJDApCD5RZqxPdFck/5I6ern34uqAaZkWM
oi0MIVg2f+6UBYvOf5gLWm3Tfxm7ioFzfqJXVuZGCovXjHodGM+VeNxhoMQN2ud0Opjou+yfFpk8
5j5IuN5gS037/4FHsyh9B7GIi5CfJs7odzhI0P3S93aMHyGQ2IenpPh2lcOEZJSgYCG8auelMu4/
c/DU4KWWPUiA4yUoZh6J0qRaEm76SSS/WKxzOzdH1xGEpyKwi+uR/6z5sG1eR1G87287xLn3NaLj
RXpKQEDz43lGHk01XEsQdXGGI4Bv0qi+dsdx8/2DlCM8h94O9Fa/p0VN86r1kRdSR/yP3vGCX8pI
JqixbOTEgUzgDPvwnN/uYpCY2MEWZbSUZTmbL3U0eYdxkRRZweFJQPkRpKGlPKqnFcciyeAfjgBN
uk0Y+r+5Imp2Dc26zwUtg2/jDObpkQSUXE7XLNR2bnsihqOE/z22I76JZqh64+ltUOWWE9MZtK4R
bAkPbsFuuNsSJ5oLUXUS0mlNSATI9euSHSNUtUbejQMRWsa5t0Whou3w52yz9FM/IIwo1GgajKeR
c3d3/iJTFsLRE4q7z2FeUTNwpdEb3P7qvcTk6G6P8cvjV/WPT+YYpWz1ziq5oQl75k6fA0uzFX82
S7MTh5RpPIzx/l1osIQu56Hj5hTZ8jvVAqD90gJOFyiizE4IVN3Ww6MkpyHmwlkjVAHP97cPZ8Ml
SW9LJEwLF3sCj/RIR8VsaYdDJLzkgGXyUpI+dkaG0PDvyyrxoVpp9c9WrSDszcCxpCRBo7/X8CIS
Rcm9nH5b8c5Xvd5M4r/is8sdNPA1Yg3hpAKt2iW9YfXdKtyAWlIViqp+ixcBdwqez04XrgA0JiaS
AfR3Erp3VbvlyA7NRtwgiBuFZb35Y2NuAldm+ARRHq/0k5ebitkufvbudqxFeOkM6P7ldzKCJU5E
p7w4Q8zhyJ2pL2GigiUvQ5ojWr6RgqWqphah3HgaRxnsE7oJ2GPJWEXm5N7sB98vWAavcBDQNpiV
NKtPa662D3g0qJd6W/BzO6P+p8TNNp48BQG4CcLkEqQYFc2ENZnsMdBucRiRuBWgtMBIUGdyNZ9+
gqO+6RZuEfTFQB9skZvpMsf06xF/S4XprupuQTHmU2Yg+Kxm9NV3/TEQSH1kx/Yfd0v7Gj7ecDkL
vOVvPmh/4H6YrFOftGQKimB21hdPSQvjBjXKIvqTwMNyfbs3Z3mpbmqvBT6vfFo1rGiCk+21YsTq
JmRP4er/HwIMB1rZOLMuXttl5fbgjcpccInXxVwBkYIPwc9PBJWl3gxVXhKiVCKlfeSckuODSlSl
8ZkO46IW7K1Kq7RuoiijHlBkr4pQc6U0qc4pOMsE6Hzk9Y5Cy/UaqQlu2O5ywCxEJrdnD7WU4lVS
W/rafUg0lJhBwCsCbDbI8nuhP7Ax9GVAh9vjtMaHpcaASxSZ3VcM+FNlye/XbfNIZib2P/Bz6E0N
b4J+vUl9z5Ei1pyxgOb6OLalF4deY+hPD+W81iwA3injDFsJvZHcZRuoapyAhH0T63JR/FyYHtVL
gdC6yHJxGEE4BBHNYCb+KaeutSWpbCGfp2M3cj5P0zXXpnS8ZxsZq3NPL4Qf4h4qWv9Bh1ncvZcu
JOcH86K0jbO2jRGlLqyHT+wKtEYtHVMxrPieHyno4oWpGYp4Ab8zj4DMsxWQCqRbvF7do/FCcGuA
0UGYRrhYUmIC8YjyriZWuVi4kJvo1PYmLefs8M4u9r8V4Kr9ZljcwTIYjHw47HxBFDmHF443/r2K
Z3DYo8BxAmQHP7mi+7XOLq56Db6+brtHKYFyEsNk9V6hre+S9fYcE8R6cPQDy1cjJ/avb41Fq848
4KS5VIVbqSrKMfHvM8mQ0I64TpGPm2NYz4H1ZFmiO3tO2kqy2zd951u5yA5VTRXzW+xtu+pPB2Bm
fsWBWzE1Tc+m42Qe8K61SyFtAQHY+8cd2kv3n9n9rvNnEfGrloEYE5L4Ez4c/25iarvNkZRUT3AB
ugHD3315c2QBBlGI+3wL6tER6lpllTukXd54TnD6J3bSuAi3mdqlbqA7UvYtJUK1UG7QzAsM6bpd
WYmxvNT6D5LIjlyeK4VO7aY7h1IiGZtFABDf39ZNL2lzZtkWlV67n5qkBjAdVB3FH7D0nADXOZEc
UTKUiPh658aNzaZ+BNtkRRc1c09S5o6ZctSbyEoSa6vd0rHerx3dgbdQNaFRDjRxH1BezLRMY3au
EHlBRl/SuMjTal00Sk6CZ1lHqwztUjlfjzjLbOHG4NFDDKwj8a4BIph5KprO68IQ2MC/Tpspi95p
7HaXeiDMpWIPMCqABW9cRej/XRUUUUyAqW5qjtMqjcF1B7fc3L1YoVoaFODKbQDrT3KSkll82nOZ
39nz6lTOcGGt0OLdDg6qyMtpbMUGluIT7swcjqA54YkgaTOklciDwkLqkt8I6/Mtgvri54CfVdNB
yja8Dcay7DPA1lhKN8ZHHql0U1U+2hxheHageYtLehJD1JwkqwlLrD0X059NvJYby6zuKXgkeE/S
T9XwsC3oMYP861YkH2shDAm3/Yb6tKu7WR0nN7oV80qlyrEjMn2jr/1Z9LjszIDslA8ZxBJTxUql
GDNv2RJ3XaW7SBE/obEWfMyRTbHhFPv9MXaB/SCH26pgqfkhmRuZ4yEEJE9jIumar446TGoFKeLA
ux8Hn7HmLCxpPA0EcyIp7/ckWTBGSOdUE3Csu7M5n3Nje0+xJgGNIGM0e+K3OGupIhvuWyZbG+Mi
vQaUduhhM36PqQ2u3ij4Rc3H48H1u3fJAXZbxBsqCbYwXbSPBFdbbS18754/CKX2vD6hFmFXSqRv
pfhgZ6u/7H8NkfjZOEXIi++yRmEB5f+NUCdbHsEr871kasmcbKZtF11WQe5nJ+Gw6MTXE9TPS9M+
xdOhbQUfqts/HaS++EIlXP3Fgsmyrwu3ncfq7LeCAsm8kVeHviUZ1uufpVGu1LMh1IA3sTIp2sR6
ou9lDrSipPl/YVsWPGVUMN4Sumza1zP9QVVLlY5Gj0JjSohaa9ICqaw4NCFNGcX4Q2f5H1StnTy+
guWJw7qLbiBtn7xCQScrb8/dMQHAfNyqJ2yqTbgcUcQJngEWKNZ9oOFuqmaJ3rK5HJXO/qerJUqU
OSni86cxtIryQFAx2DkV8N22QLTwezvIk+RI6Vm19H0jXHjbyA3cTp5OUNW8ZfZYSGef9+DYIDz3
9BUpAJ0Zw3XoLLQgYuBjZkbRZKzO3XSnTBi6DhmJFUgzeg+eW4mGCGPqpmfDUZnk53T326SijQSm
GGCPzK5fdn7AhRu37t7lTcYR7ezMfXj7qswG5dIGf2/jFOlBT3bNPmCgYn1wsU/PdKYWQbjh1/4Y
xR4l8zvKwiNPrQUcrLeg/EE4gZbyug7msTJW1zdwcGTjKG08gvfK5RFDrbv6aWi3iSd1NhtNQ4Sq
a7J3XRYYGQeK0AwzqdokmIFqFQ2+OWz0ToMj0gAMhoD5pm+46gUbc/fnEWD3SlOhFpiftZzOq11+
uy7rdu2MSL02JBT3r4AeK8cRxrEjx9gNmVIlpnvjPAhbZzdJV1fxSidxVstAaM/UH8DsWRXhjD5k
iBYlyLRQDKzLzZk9wG5eQ5ZwPOMjJOPhkuIKn5bZc4mwnFPGdJ9iFQ3k/mL2cFOoqDxBTk7l44/6
X4QWbrl3jZuHi9urxLiOP5Sr2ocnYGklCLLwljJ4/uymAbRoI+1kkWWfwU+ZY83QBCzHJunl4SHS
zaUvi0cLM11HvUd1/D1xk0bhDCvAgTkWiKZ1YC++csm/9eC3Du/fm8svoII94neRe0/tkILPbVqO
0r5ee04K3LdtmVv78FDB52iFlzCUOtq5U/3gVgP7KFOEsbyd5XtbjVkCgmbUayxqZz485VEiz6Fd
hysiQT64k8LWPfyGPhiTIZxuYWqy93mPykMeuMxDejMOBCYsJbHsbNEZ1j5tOUhMprrN70FdFso7
TYLH8YKzAPJnaMJ5fg4/4zrg5FTyint7JF0lO+euJqjd63Ihrq5B3NEDBharmvG+fsFaq8dw+Nih
GM5svr8qV3AZvRtsqORafBybaiT1vG6RgVMdZBMyyxAz0cZ2QZjxVrr26YTx7bp03UB3RuBsbQNd
ME/FySRgdlatXzj33ia5JUhAWYvogbRktnzzhGmxjp9MCpkJHjUE7wFtEucTyKM8S36pPqFVAcrr
c/fylCR1fWDOkni/6Ca4ziEqvd3kWHIbuF8SqzanxAM7j9t7cE9UkSZqPm+TtTx6dzh6EQNjZvOQ
4Ow+fvN6/f32W47/wSe3+sL+GNfUJvZDuL/KlyIEeDMCMZMxe4ehNoQt1D0caq59GrvgrNVp/Z6A
ToIfVtfeNXzbsyp9JeBcc/MIj+9IYcQR8BGCLYujbuO+qP0nThhYh5VnLrC7VVeq2rddVMK4WVug
aLvrKdMYK0xtGUJa0Qzv6+4aL0momCs4HSji2V2DMIRIihdHzvVcbCBJN/S+NkKmB2rCCjjBXlnS
oxAARiESJ7hhGJOSdtPvqa3VqCC0NUu+JzU/Io1Ig8b3hRkyHwGkoDdVzuW0wKuEYkKliIYGE97a
wqLi1UWETXsr95gXEu3Bha/DWMkIJLD0N/N54pMo/bKzfBw/ooyzvC1Stf86o33cnMcXMjdHjkEU
bocEX3SmW9XUsF2sy0NhCVu7/+HEC7a7055vwe8QU5EvDFI/+gV9WXvPlpYVIOLBL9Sia6aH0HMq
3ySXCxlwBjXwgBId7+N201uvYrurpxGUyEWBZZjjunEPwriTLqSJ7fRWh2eOa81DYszRqpKY9WhV
CcBgNHXED16eX4gGdMelLTzzKGIU0dU428vdGRFWnJ1HZjb4FQikkXnNoiwAGg4C+RIWGJkKlUIb
Rfj/aW1aoGfkQHT+RSf4bo9BmLngNsjHycG4z6ElykYZl7yza195xEvO8BqjOcZX7q1x/r/t9TOo
L9mkD3t3W1dYDvwCm2iZqkaeh8NLOE8NlRo0x8gDqdRUO2BYhHlZD1WuhKu38MruxGdudC2i81Xq
TLeC1PoBrxPwxjy1KOrpmeboEaALlviiCIyNIzC1Fo15r8XPlMnEVRQS4nzvnUB/yxxmWtfDcNTU
dotVKRjhdkgQVVrtAp5z+fx1hkMs8QnX0yhSs5rP9MgDgP0BpkGL3GjW9HkObU1GzuMzaHGS/xv2
6Th23GR5bUYvLJbQh7EKLMIGGf6H+vgkZdNHE9ThISvM385hr3ulN9NTyJeKSwbbe9E2J8X/pJm+
qlx70IjJK9mgsSpaKGjnJefPDrOs5jFOwjwGgKIOUxZ5OCQzNrT+iPZBFeDEZ5vVKRJvgiFnnieg
O19LTRoR38x64j6VqnAAHPv2xdG7ySuNOQok+MB64GB5At1Wj/RqrQ4lLMjEoAdusQquNht6XG0x
y/63JlXd/Oi15tJoSw2bU3Ml1i6NltvdBDJ81J+mON1opWeDjGrQQdZWbDAGyJvCL4YvY2D2s1wj
KWZaB6gSCqLEBUcbQPBgRudZ68imJURLCQbRlNOkSlPOHhKkUOyXIdGxmGvP0eS9YVKp5FXw+XtN
NSg1i/Ps021TBdzD1f0cavW2ViXA837hoMs8dGk/TpNZP1Kblrb4vkSHdfVJ9XiaJepEfdhjzyY8
/jytKYHCjAbjhKJ6tcqqZ/mLiYsNoChXWhYSHeAM6dNdgj84qF/ZdJGw8ED7mpYD3o0879OH84B8
0X8N9XTT+rzOeS+S/0yd29qhfRSu6L4+qoRJPzvQqCJ0Ha8SMK46czjASM04NsC32YrH6PCdh+Rc
CKGwHXq/xUm564scmJ5z4AK+OZg9glMVufzjSxY74x4plTvIyn5Xe8XwKQEakk6/8mf4B0ssE8sa
+/8zBtQtx4dnc3EQKhXHA69ULdxINNGqYOTABSdpD/y8o25L5Sr4TkDwc0sxvwk40YzS1Y2jeDWY
HSAUUu7G/arSY/3whI4QMq25yN73d2KTNZkHW8tVFftyIxL/xpxgSmIDXJs/rOXVNDdy1oIFVzqj
wI+/rBM+4hAwXO1NjSgMQbwhvAfIqAKLY+h+WfNAGK6kTmJxy/3VF5euCQKDGSHkcA3iYSeI8jix
/8k2OVMHyONIWF4aVklm0mKraWARNZ/8kbIgmHHX+lFEVdYXrVQPXQv4IDVGhAkAoEGAp6dGs2Y/
0dUoMr1EtWa1zjadCfYCFDykoP6fDsd+i+Xwmtx5M9pxPk9osz/xB5QxsnTNWxFVsFnIxFAdhbkM
YEHOXIv6WUk/IVMcfXl3Xk3duoS4rOgG3yIKosVUKTtA3s7BCz4Dapy5qhdgIAutKp96Hq8XHurY
7ha+ozR0Ve7CPoh5Vzmi+/9fkD8kK6IbkaG8vnoXp5LzPueCP/0RtcSxzsSNrPGbP8lYNLyOEY+u
j7KNd0VjE5SYGvdtQ6T0d9cuvTKz29x1DHl993+1LXzV+RZdDy8VaibmyuM6WhF2qLQay+Da9riZ
UvmIvAY6nh3d20iTTPKtG3F+CbMicqSmg4gaYrmA42SVlSWCeTOU3gEPVDBJyRq0Hb+6WkAvyyVK
yjMT4TgT44a72paJh0TBPVUNzhe1LI0mkPYmuT+iPcWa/Mh3AQxJT+lPgFGVrU/drvLeWVdiCfby
g66YU9fH4s133o9d33TpOzS8jOTml5H7FQOyg9YsCtZ+VswnCGj89wdUhB0wuaAWS/Qy3QtXkfz1
AntzKFlyopvS0qYv12wTyqiVqZP16DpQZCSYcGmnuMo9Gwcj2IKO0wgwGoD/fFiec+XdFg5z8swU
jUb3CqhmxXzJTMwHtMMnCMHVJ47W5+Er1HF1FkS+AW3pS13xdTuOPCdINMWq5pUjK3uAYX1dBigl
uItwx0xkV+t7dPBYqZzel4asezho2ew1HVK+VPEtbeUu+/3HLuC0Ji4F8bYqNGREX0Ou8FBjQyO8
qsOo7TuXhaaY1+cvY23jiNFfVIMbkG8VQ6dmUg5F0O24h+4h4P1UMdOzm8IgPBYiVr1QqNyOdT1d
yXC7L0UWa6+n8MVKnZK4xJ+UIx0appGoQXiINYmBbG4jlv7n1xIZbyFLRachNQs+ZtfEADsa6TKM
ofduoJSEraiCIiy8RjoHxarfR7ERR/LbgHWpbR9wAX1cEXZA9le4QqDA5ksgsTA9vmYGYn/f+vXQ
32LYneATJEhCa1ltNW37bqBPPey+qik/dOBoE2zIiy0FvFq+2gDZ+yjGKkZRQz6ucKsdTt7uVMgz
i88X8JfIq2kpl5bkEEIK9fUnUnNiFipvy6/8lYbIgk5mDLogUA5X1om0uAODZtNYk+1EdiAuMvk1
tgUwEF+n0Dqpy6WiwyU7cE5HbT/cU0CAmQ1AWL00UUfAlvngkZTRLUpFtwg+te5Gqyg5VD3L8JhA
rjqALV4ajzQPDaLU5t800bDT04bzzI0X42t3nKa/GYGsOKnrdcCnG51I/WQvxK7q1mge5/RBsOH5
oM55mLthsby63jOYEUFM6Q1u1gxUXKd4bw059IPEy/Ad6zJgEg/vXA7BZQ9zU+xjQVc7aVVsmKux
xHTNgh54FDB9WvS40z0RQFxrV5CIZd8ZyzVC9kZ2W34PcQwyC+WczhgE4rPD5Xow+dPZiCUL2I9W
f02j7GoFfJl3Vr9ROzkedLQZTxbpQ6roJZ3I1uhz2AX0pHmc/woGvdZBKl0AlHVZ6XgTtOr928io
LstxuR6BPIBK4IpEC8aJlLTTtu/OHbLz14VBq6PsDxo9MUiXJkYLqBOYIJUaDk1LyyOSVvh6tonq
S4gUbnvaCjpozq04LYmODaRawldOufJrt8sAnnj2424p2S5PbHa8q6qo42HSMmEejHAYyPYYoo0J
6KZoPc9e4cLGizd+hnwsZxMwbDt3iwt/T7+WY3PUsnv3RbzdrAIATu1rArOJwk5s2/tEMgdb4tvh
05UwlaOIRSvmWALxerSD5SWDSurfU8mNnbXT+lpUeotxA0Ol6Pv5zfzvwjRpxcSsheoddTPC9T8i
7aDBrfbw0sQhdnVynBCmZpuh7BahtGf4P+fkTgW6jlA5uShyC9jbwaNHZ5UCrdnxwC78S0RPp7Sm
jBUDQWvFZ9y0GGpT7BJplm3s3nVNtbz9gRcCXx4a7RV51ZyIpQRBhSX7O62zl8M9luwJW06sIXVm
vDLz1xt95yENL6oukL6tTyfZQc5IrGPfdkn2k27Jjoi5VW0c8PafWyllPvp48ABBfQjBSsD6v3sz
TzE/4AQNiqSQKbvPLKOajdPHWpBtZStr0yOppOtPvGhyNPy6qxiVnHqaTwu/fK481IynRGLX8kUA
77LXrBQhf1NJAgAG6YlWXAioi/fhjQ5l6XofYw2J2NzASEse0vYG9wc8imtMQ5cjdAzVbmTM0JMF
Rkf1Wdg+ofSt/7y7EeXZMt6As3u/yTQD1kSVWkWvearOpzN1sXfUyLfdgwpxYPewBjjspnId0+EN
f3qjrV6RaQW/cJSV95LyUMYBCGXNR8Lu10g8NUcXBh9zoIXnBL7vTtSw+mKba83+6psHlcyyv/g3
apTW1lW3jy2EZg/WoyqBSBxZj033atu9h9gew5HOIwlpqCDlm22zTRS7flhiO8If13DUeffxAZMH
uUCx2GfWIfX+oBNgEwO5BolHAVOxFE4l8pvge720WTCYBbwN3zTwI4Rr3EOOFqH+DXTk3ha2b3BM
HRBKk4AuOFHhYl2f0dyokWVMHqlCnuUWu/dutcl669tDWPmufX53b9XFRbAm7OgG+EX9xTCibun5
pfO+TBGQqlp2lLIhYGHs/DoOvMJF9fime59S96Kdz7mz0eysqwSEktDJpPqBITwn7xQ14uCcWb5l
nj4ADwiQm5qORk10SKBClpPg2uRF85AH4YA03rmpGKl6HkWNixNQnSuM2slEuabhkapq11uSaHqT
8Nc8ebJEV/7fB9W0tucplKAhGmSrLVRbfPBlGY3nRFL7nsIQG2nVBecLPCQIe7J+P4sOTVZ+5Pbl
K3Bgg0JSCL+rt40YVQkuF8kADZ7xCIJUu9T1tEdWNmuG58GxFcGSzZi1w1tcxSJ/lhVIIyF/dOOD
O9fhkKyG5CVnwsmnq3C6jgPf48cqaystMf7iQ0bMfsZjM/7egfrgPfaKzalMdcRbzvDcSYbjdH7U
wWyv7TlU6YEloUD4I3cqDSqXIx2tGo1FSHT2MwLKqbWozeUN3PBrfGDsa5+10z29gamm5GSlIoYn
HP6NnnpNXsdv7LhCIRu0D8kfbOyA9TKscVUoSDP/J6Glk2nmtlc4xTr8FaRuVWPc2VGAIZ0yp3ky
4xGoNPwz+JMqkzMvSNvWuFREgQ+v073wGgs1nD6kNy9SWVHiej6MvlhrGBjlDqGjc2PzEdOuspvf
C24DvlIz3eRNRbabV5VySQJtA9m0XWvuS6k8SRF6fzjGYwgawA++x1D+7biSLvdDW3CUAl/bSe5f
OY72mKb8rY5lQ4GzSjgksQHENY/0cRjki00Ot6UY8aazD93NSGB+hB9Es4Hu+ueM6VhCkG93K5sb
46L3A95sUQELzpC/VOqVzM+PerLYUfZFZZv4BjHf2zfjXQSpIFqSb7149MDLcA2m13Q6sFGLq0XM
eO3uzwsVZtJYdFkUvMyb6lDXDQpWxO2JQNVIze9bmDHgY7L0TwC6iqB1ekcRzYlmsjy7OsMw21Qr
oQlpS7dj9WmAFCt5/If8F2DxLiP4f6lkAUVrFEPq8uXrNG4ytZMWtDGmjeycLqWtPV3QzyUz2SPX
0T1gSine7ay+zScMeZqWbfPYVqLizE4K6Nx76DDqUt3RaeMM2cxL7okVV4CeAaCrVij1sWv7b4KK
6BmK5ejNuT/giFTLstW7y5UhIp+i9dFy9hQn1K+jIMvUwPJ74KtRqFuuTqj/BTZ1c0ZEHcT+DFDU
X7yH1M2qkhCHFxv0OraaPtbAsVzV7+Z8LmUazehaA5G+dMs2VIhxwxtqsguzmhlo1Nu2kLK1WvVr
DM49BCVceQCQxb3dBB6/RLiTuU8IMCcsWX4k018CU7djt9iWnr1jhT0YMLfiPTJb0x42KvdBGV7/
KyMvg6xAHthzCBPNGDLcJp4oOfSGL5EY6u+JuuV7OFuipupQCzAsrDkrapLcjwNqWz9yhRJV296t
vNOdAdZjapTYNiUuzerQN7Htk+2j8Gh6zP4bL/z9v7EoZfL9kNbHgAiQbHDT7VD2WoFNqMkmeRPh
5vZpaRC3M89Re060m8T1Z0RnuT4tFDwplARoN1o3MLmhvMG/WuJNf/88y0p9IWocbjmlRmItBbaV
caH/gJPvtsKOlBnSvsucbFhVpTsuAZxpahPWnkG28bcW35eWb5Q81Wp1zeB8De/pu5fSG8FaNtll
052s5K0TLFlP9QHJ0Psa3Q/gZoRjv57ckosZSDx/834CihollSEwZkiyb4HzKAc5hCNaHqhY+l9Q
Aedy9t579RNouqm3WZ2YKIQgYiQyLDBE4HXBQFRa4g/AaHqI95O2sF9Im0biO3t8LK2RwXKVPJMr
l52iotnz2ebLXB0+YpvVnhSMrF99eJNxaOTm4Ls9P8J7qK6Jilav8yAZ4sb62xpLIP+KLJHuNvCX
t09w/nkqO/Ph1vJDzrkS1wcaekYea8KFDEqChvMC6pAR8pkqTwWel4ISqhDFFUdo7X/zU//eezgL
Ves4VR+SzsKn8Xhop5yFn+ztwzQ9Vd79HyTCxMw2XBbWfVuV9sLyEt9dKTuGfmue580xAgWMU+rG
HndhV4ZUu6M/v1aguRolyRsisQ4kuDBAoZi72lUwgvFIbRI6qn6ePE8gEaFkKw9qqz1DBiQkSN2G
fymAb021ObdwjF5eln9bx77HU9uXMcn/xXp/2J7r6FiPHFA5e9e3rvrNYoD30izkOD7ddHnnFu7T
MsLHgJ0lQY+5yXt8cKFtdjkVl4dC616In2TbyIQXjBFXrbpMWVQsI/jqrnaKMc4JbX0Q2cC+XhHH
mA2+Q5ijZ4K2qWVLQ9vq7JgHRGrEmhYGpay0UHi1xQJB9CpvFGIcv3liABtiF1x0PjxA0cQpJkKA
J3PlJb9G+d2tdE/s41/sB5hr0wgZVr7aBEp2b6En2DeWyyvxeBuQ3pY9yZDMaOE8Q8S5lKei7IPs
B1nnM1Giy226522F4nWXds3MW4KHOpBI+L2FrZ8NYUlUBcVlQK46n0UJaFMdGw12oGdKPcPjnUXp
6GJ5iiW3aSRo6AqkbcD6BmoEIT+uDuR+YAwtGbn+UPDA2+6y9LANI8yfgNCqfCQc0VcSMAFg9Gqs
vmPiQH9PG88TUiMiqDFJCT3avmN5GQm4s7wdA/wOwjMA928Y9PM3hWjCIXuvj/CLf5tYM+BhhpA3
l1jSLLa2xN3RLhlZZGHCd4oUhh1U2O6R2XQ0+/hgCO/ZOBLy3ghPiY8qdrlyTXKHkNn1nSx5AZy3
QAkd/HZ2BfOKYDD5nVFB8MT9+ueZw9+hagNH9kqmyNmLW6zig8vqdz/NXURpgU4OgR/+QcFpqPxW
EUWbdROv+QTy7fJOZibuMNiPhX2KsLgJ2BC9GJIW83uFXPUm3/hS2Z44bBq52p5S6U18MVFqjpv3
xy45UZtx/xSoowTjTFkqh/sQ5HYFJmnwNjzgNQdOVVqlV4ViaJE7RojcIbl4ni//PbfFTMbeFwEm
N4DCYj8i2vBIxoZ7+ONTYNSauCxViVt/LD6aoQbcU3TRiKnNAFDHtpYjEfHtgv56VwYxUjE7yMjE
k+r4FUBL1Li+LoIJ1cOxg+8MtDQA4KqWKIHSUH7JUo5HxnHRpSPfOSQoFZXK46Ukgw9Gv/ZXXIzg
dqzGmaA8HyHwy5TClLSWUVyyuKL2X+HVpkWawZHMS5J0tDsLCGmZfrFjSxYuaQosMl9NYq8yhq6y
5C5uVj85h7mCwv5IUCqXGkQnK0cQ6pqxdJlIEbX+M6tk/EYYJ0BA9+xNup2sJP69oe4yZwL8QZZg
Zw1jYnb74nPEnQH1JuNWJKbE8Qj/jCdFcDXyXK1+YXStL/Ldh7zZGlQf6aJm1omAcva6hdTjlyQZ
220gccJwi0QvlJHT6jLfPIho26aIDFCZSB+TN4gDNimk+3iQ6MOpUVmjnr+gYEiAPIGt8GdhwY1q
rn9CLJmw/NkBB52EHT5y0qsXL02xA5rFjoz2+I45wdmiAD04DgK67Hm6ePnyWRvDWkQ97GtraXNc
xXWN+nULHR7sMjVlMwFibOKtZTz5xW+iBgmP0OFZh7r8PIuih10rXS+BKqMZ35Po3rwdLESOM/yu
yKFSml5B7zi9diAUXhbB0dpz4dsN1aniS5QgFae92dqdteFZxhB/eHiafAgYWEekYe1e06jfygC0
iOFK4U+VW0JdNCPBgA8+BrJp/GZcTnR0wlfuscV7xEw2HJI7uuOMaVS3aTjlnkine6FIrHvj919c
aEdIJaK8LKr1Q2RoVyddu8kLqq2dkxB8HpSCsVjTvbP13tkIMRIOh2wNdVEPTh8hWSvGExvNJadg
q9TqhR8+9NSPQoBeX8YyoIko5kAnBTSD7YkparMN1SuNNaKIc1o68T4Jj5jkG2ZLQD7r3c5t3zlu
5RJUqDKOvob3gXGWTFZPJ8szlPumy1ItmQ4XHgo7zDHzSL8teAYpmDpy4ABvPfgxd4Cf7V8zUBjD
j0IBLBRc47iyApsh72z2/a8eYIVvX5UgTapfoitoGFkmdRruvIXSFq+uru8crKM76qllN9K+f25b
nYrLVaUSTV4aO/sdozqBX02um2FlQseev6fKqwwPlarm70RJ1QYz6Ka69eqqeCzieuvZdH1wlWKm
KFFf2IMT4ojxoxIUq7cZn/nSAGuocbRw3/7fzuu29kenuOOLQ0JEOlGNVxAndRw7Ue74VJdMXpt1
A2uoIv0Pij44GN6LfgndJMof3IEd+m+fIJaO/lgwL44LWpBXm/5tblDe4L350RPwjJcnz6OgXzPc
AebKb73yYR6qYP0ZYYjLDBrtTT81roATrbfMl1UvNl1EDvrJH0WiOpbKAZt/v6Y/4eh3t9piHvs6
ySNjlLvIC42Ibpzm39J0S/R5TRbZNy2UovAHz+Qv5dfh5VW5b+yS+5YGmCrRPwvyAAYyMVvM9dDl
1w9zg9Snj1CD7oUdvsinStLZffBqm/mnLvw48U0ANSMOwAgwcBLLBjiJoX9GLGNLHp6p78Ml7HNL
XMNxwNBsvIsqr5FXK9AB5Upls1SeoaHsW2dVqqUWYXKMG7mQB7RMS4E5dQRXi61nsfXQglJbDKkz
0HlscoFVZ6/K5FBqYIxnOHwaJZfY6idyC2/8S920g/nuyPcNM40l8P6Hml4UVmyDB6tdvvvsh6JV
Z6c6Et8YbNe4NjekyKYOiwV1RyDVvW/eJUlfI9p9ytU482xIcMP/wrKCDp7oUdU9Shk9+wxuV/AY
k+hXrvnyqOocec83RC+ej6rNXah8tQ/QiFXThqi9VqzQB1dJ975KCNvtBnd03cJXveMjrpIzWdFw
GxwEQW9fuHeYySzOai5srFyQP+IbRJnzGyLzsTciiJ0sCWKz+oIMnF7lxPN5FR97uHsqhqXf9RFn
Uxxxawe5Lt/OL9U3QSAiamZw59QpkRoXJKyMiqPSzBR2BayvtXK41OpIxSQmTklP04DCWaJBfHjK
i7uPD0alHxlbXJhfXbqojTRWBfs6GVPDJRcv6BFTZJmXK4FWkBTw6WP5hhP52EFnx3SI5JxY37y3
rndP6hYbOSWHzUUHPQ/8lGG26WT8WjVhrGetuzHickgPxqIyAaF0+GQFL/7Po3pYGzgtZPHoPjEc
D6b1oxlvSj32nD4tkoSKApXJc7Psk3C56wvX79tZzK6srX6SdOrMglGTbRJ1ZOiDot36G3HP0bIS
tCISxby6xMwxMvKNZqoEBCxaRwbDyZixAoceUdJdArnativXYc39DfVpuLS5DPmMuQUQAB0qtq7V
F8JjoSRBN7VmSQehu5khagK0zIUenuCQ+WK4AHYiU8ClxxGIFqumtcWAhuu8YigEAUWutz0adtl7
hAs52YztOc4DF5vEx+Ut3JRBMv24pR7orvhdYlRnMd8muM4r/Rzum1vCOolvEuPjO4wHrLrscpCU
0zxNlOYFWVst58Mh2IZh+gOB/utpPzyjPon9w5gTK2YIaFpREFZzNTNLJUFD8V9dUDFhPo86vDXZ
C4E21I+h3hbDVtjH0CIR2OK2qkFb4yhXCcn6qQseJVI75tbbBn54QmrWRHWLfuy2dlGqU6Hwwfup
raFFWKIpYrm2kkCYds0Iv0ctB6MU13u5HQiAlzXIvQVKN5D1q17eEhNicrMxPrYND9F42z9H7m73
+cwDZcLYtxszNd46JRfcmq/gG3+cpxwPZufDEZGEqeHzFV+/mXDt8lGttK7xg3yW43mE27TmcSTQ
qBHPbPlhfk9oQT2Og5N71uTATDH+0ocqXznQSoAw6A4iJN348Cai/mBNfReydp127JJjd1kk8acE
Ng0vrE27B5FQGo3wOVYRhhzCyhfe4vuDB0x9AirZJR77iJW+cXRFN8HCOgzRjUrWODHCopzhr7b0
tcegytSecNG3rcah9oZXp0KVrn1R/s4Dx5oIOORfLWD80qCj03XUcI2WwtKxtcoFc/x7vvGmrLrI
uPHq1Pm8o8Giy94/zB3lwG3PQxpby4T0PEk5zWKZbe2uYLtLeQ1coD858BYW8//cLyV8lETscmLO
PezYni08GXbcFVFJP95Ihbvt7uIeXznkwgFy0NJYQKlE9aq+8e8Gz98Z04oMESZUsEouIt5Ghu7r
tkDtuy3PqGE+N0glvREGqFE1so3ZUh2a4wHTA8WzGe9RBCrnnPM1fiDbp6c0XwZyGlAw4lQTAybq
1HqCK4Fx+Tk0rnRO77WOdeOXiLP6gNJMw89dHwVrAWhzGz4wBTJPt/rO7NLOCxi1f9C4l2C3vHon
Z/8e4s+BUeEoUuKvypoJha6OtdbAeiUNi0yEJUX9T+UqBBwFPgR+SInJ3A/nB3J/N/g9niDpi9V6
kjSUiMjXnP6FUJVLi0jU0pFlZGCq4PqhlHMDCM8hh6KLYUreFbm7vx5nG75cPFfQBLSztHE1B47m
x3+ttPnT4zFzYTIhlfPBY1TWwGTjDLGRGxIf6CaQW2U+FfTOEY+t/wUx7c/8vjeEc2qCXQ6wL7hU
osQp3DQBSEWmbIAXUu2BZMHz2sN+WjHy7AlNXXELdEJr0M5Hpq61Vbh97gg1UCTKYCvkck+jvKVH
Ow38eRBmxFbxWHPFZNbtA7J0FBA55o8Vb4ISm9meoiJc0fGo0VUDcck2hDpqGswZ8TIqWT0tMcM0
Ew1Pk3950GuqMQmCXua3G461JEaYEB48wYvUiIpOoDke2A949EjfP8KUso+yhs0l5ipKxquNZbuw
AhHCWyeeC6/rqw79RJq/8SAY3DGUeDpmAtTZY6T2RJayfDXNOJFcYFG633QkV8/EPUpQpgWUnV7e
4n20xJ7Otoi1nN8wCgnHx1WEeEmwZQIOqOo9U96qJqfWYhT5H8Dem/3qYtxCmYLqx19QCm1kDCSg
WvnwSpef2U9+Y2KT4qNfgr4KFCcurGtttVgvnQBVK9550UDDdQPxOwEA6vUQLbuSoElw0yTMlrU4
Ocb0XHbfh/+UQ556QZQKM5FQhxkrE1sM5SMSbeByMfEACzNPhpj6p+b68WJhYI2ei1ZghsqKZtKu
yiiFKCSxQjVLa3xG13cV8q5s1pJ4aEgjykmEXSGpNz72HJVl9Z6/4sjNncWuX1RlzkNZznVMbDvg
hDBd07UKqfflq8BazbNhdL1+bPJ6BtKvpOVw7eENKv68blbOAtck7ILHom28pLJU95LxqtQiRdEN
nDvau8MTmyRHHW8kvU1m4IZz0qRF7R1i0d+yTDRAv2Xeu2byC+ZMWq707kVcbest+Vdth9yV8ive
ZXqiwlie0TF+JClK7e7tBa1kgOA/cKQ5OrYGkK8TOXJaHCanQpXoxvKVCptRcmm5eA3nStzPAcpZ
Jnhi69DRdEPD7Zg2iZhYiXXcbte7YKBkTx8fU+SCZ+4Ddd4D3GRoxEKQoYDWI1+esUnA0n44Wu5i
9d7XypXuaKQkodgfw9iXFV97F8wvbLd9fWNO9IuvpDMbi2iQYySyZoP1OZkUrSVb6KbVlTW6POqE
IKZ2YxQdwgHwYnfKxEzD4s/YhlWOP6GYpsdaTOmE6NIhjWcgaSdtEfmgfPKPDzWSn65RtXugmAsb
M1ORW3zQRCeFb51Sf7nV5sHaJSWKWuHsmamdJAkNy6y/NA39AxjNpPiA8qdY87rp0jsLLVCeCsmb
O2QMpPKc2IE5dY9oNGf4Q1fxnjYosWMvAYTV6L8UqCAjxHTKzyG4fZNC/kScL96QzrrPyzoA7hNm
EWpdQRQG9BTxeeH3U7Od6Usg23iPPE96PSQT4yLc92xsY6zowPLmHW8YCaAR1S7bWQF/b+9oMzer
9g57cusXu6CwCQPct3bejlko1VmVbNUoHZlC/iLwcEwVXmCutrsS4Hmp2lxmaBHRqI0riMVIWUAZ
ZgCbDG/K+PScsS3Hu+MgzSpY/BFl2fkt799fZnMKx6zleHcgASIgXTmjZAvN0kq+oAqNr8ac8old
mQissDt9dYhApbAd2jkIgZqJk8j+G2mZdHwq1zLiReQzLefSpmmTO6o6WXtyyA2dUw5Jtj5LXlhR
NqlHTv5H43E25qf/bD3QD5Ks74HGiKobyBay+180NU8DXVZ9WTIE3+ICBm/bN1poqiNJkf2/RhFI
vzYCUyv7ckXK2Du2+QUZPlJHt/WypHT1kSeD9+CbTR+pOao/tGSIdfmNZaKscLUtesD1IHDybY61
4ONSrnO8aAa0njmnKsgJcPg+w48sOrrBKm1fpRI9hvl+hcFW4p/yu0Ohyuk5gzPnNWxQ79qAtJAK
KWMNcAEHK05rMiudsQ9s/2pS7ceyvg/8ZXc8kgfFfL8bRj0MBYBPV/g4EiZfuj6XTDXhtePOPfvO
3EPzoo4InkXjEr69HiSaCbElVFUoRodkpD3YaokzOMOT8PmzJ9HljrIJUhNaAiJfre7g7xRltu5z
NFw85XvDeLo8cZNr65Bt6Anxrv+O+ZxJ9xN3pZmyo6Ea8nEo5c3sgv+pEWof92MYMjCns4T4eMlC
QJFUmtjH0J+R+m8nrA+81XayxKKT3dgkY56U+v805znB/mBqZ4ugGI++rl7jQaUA8llQy/LlLPyl
gmfnOgZJK4AumqGn0rrQFlpg7XCeX8HadeZWaWAl1UCjfjsI47XXlSMrDfWDNAVxdWr1zDsU0tjS
xxFCogLefJy8+KBzzgrzXfDwaipMXpMFZjRvtPduh8Pu48NliVdXdWwjKzD0APzIVtocEnmiCIB4
FX1K7TJGWn/uEEGx69hhX71kySD40Cmmxsnlvc0YA8k5M9cQWRdmFo3FpU7+p4gER92ctMqxD/7X
NmTmX15DH+VPO/Y2T3lOoY4NHfLl4daXw+RAz8oEZUr0n4XsQC9MytNlVqhpmqrV4Ybdgic1O1Qs
/yT2kWAZWn2S+iJ8nIKA4w8iom0ZgsucOgARYmdj1zJTkM6UO6b4RXOVufwuhmCJEUSXqukXe81a
xdA4p0nL6PtpA3V5yuGSeevsGn1412WGHGF7S1eLk0uB9kCPJXEzfoOKvULzVGBIfhjlG4/hctIE
YrKFcVraK9EmDdQRJr+Y5FmzV9zltUhQ1LfGIvap2lImYpp4z8lZRGq0Hgm5j3YhTGTU46fwHq7w
ECWr3XhFJBAXAF5ZQDT0OgR+BpOKymJYB5bE9ZeJkhrqpLmNcAXbHwnOjYm1F5xI6C5vSdB5VLAn
uKp0paojxdzpl2bzR3pvG+nXPTl15gqbfK/NMrZQrIa+Kfsuamp0NJif157lmVo0QS2/hPSSac1/
ZDnzCom9zwXlm2H72AH5aK2B7I8hFu7z4A2WFJYkjFqnJEIs4U0lnhsRJ371smspZI7dzn6lKpvm
pP99bgWiu+nIIkZLPf8IbI42U8JaOQluJMYUMXnF37HiEFAyGekAyuj0vbs+7PUE7OQWSy+vsmW0
GQ0VbxC3idjXL67QZy1bt/4vQfAEG1/W5Trjdd1yv3iT46EVS/GQh41b3JD3+AKTMtxaXxXHRsmz
XQ0gp0ifTqWLvgc0kKpXKl4zl2uDDgKLcjroPYcbvDxNqcFCP2EL/luJKdKwytKRKEwLe6HwuJ8O
MlEbLjKJysHw8URb1AD+QH54UC0rvGCycI+M1f0HPNoZvPUHq48xiIEf+LQq3sOfesFItPaaQ1Ug
+2FqmDl3RF6LPnukWkphRJ+UeyPub4aW4rTWfU82pKF/4wCe9vuwatZoKOIMQC7IR8VQIIZeuKJV
6yF9wGYVyaIlkuZ7k+03vRJ2xYHVKaAg8R68XAZIW7X2CrziVVO7x58TWv1IJvI692quJ99F+pNW
3afCp1ZR6cHxLHtKKj6aZpUfw0zecZG7VuBjqEWnZcngPZd/40PB0OK9FvIRjtgqodgggRwvQOnS
/6BcNixkemdGrBrHTvOELdpA8hd0SX3tM35bR4wbKk13X2tPP2bN6RGbu63OQzYgteElM9FaVNrh
fZXPLMeNnKGbmdC5VurVmL+lkEA1nwC6G14Ypmm3uUEGkHqPR5ymbWFRTnSeLWMh7e4IPRNdM7i/
y2OwJCfG6rgJPB7MTM0yz6MJWydB7B72NZHy6+E9M93q82Ey7oEecYsP59MZm09Zvj6bIzbTsLyA
NI+/WQmkib6nGEraeI0rnP/RnwTBfDtzJrhM5mhvz+DgECa0uUuyOgamHZJ/BBQUOC0XdawC5zNu
atZbn0DEsPVtZLNXNr2aPLfN0I54Y3p76G7vzmU2LqXxx8PloorgFD9g+w3khkj+YuHtrlQsvyLk
AlEAKVrcVcB8iceW8nnufO+zTOvIoX1+oQQrdpkHr7G6mDWiCOGteO/Lzo54xS7bf4+JqrAlity4
ASPO+nTdCQCEg1r1rsFRxftEtXEq8lTG6j6HAlV967fuwsUDki3aDqg/e+C+MHMxXM5V3BdtuEVl
0o3lxD+hcW6TiPhjzl2L/JSMmUDCVKcf8a8/wOynz70GYOX95Tu5o+Ax/J97ziYCCJJUgRwyl50Y
HZi24qqJGp1GoXt1mEL0rl8hxJ7gy857QRgkHl1dDXj0czwSbV4u4usfgDIOUAkH7dwVThwxH8kN
lcjSM+sryMX97l8XrcRohNrwu/XF6mZap36ysWQenJfw6eW8Oc+vPGN8++Zg3uIf/RSLjtVG+2WT
6o8tM+HX3sM0CKAgxYcOTy5r1FaICiXWxTVK3/78+6WN2LJnA6HUTcwuB0Cetvhi47RzbOGXfGQa
aM7SUFbxwtobKZD0TaN0QWEPJIrGJ2onu4wXHIfV0CDlCDrw73BqEDWe479XQaRL8KQwAvnxRviw
tYICO5O3hk+vMo3Nk5ndFSHC0C40LeW7R6/J0b6/t0zP0sNPwRSxXhCLI8UQQ8szgXLeLY4A70rr
d78gq/Bej9dwFlVt55K1rXHb7cc4sP7X7RIgzy8WaddC8f1E5EMvz4vZHX0pbL29mkGsVw9J2dFm
39HwrUpTS618thx0rsdUfn9UgLeh5wfNypsZGcnDVaJb8DH050KCtiiKccuNUly6OihlKa/a/BlA
TCtCuH89B7/wcH0J8NqSX11M6MvGlB8kCo5Y9xickPRnzADZ+jx57jQisIk6yA1DWDNWHaB55tG/
245HWTJ7vJqgn2JiR9HBeuwpIPxyEsbscfaXp228EA2IUT9jQofJ5cH2/5x1C8ys4QfX2Xl52zhQ
UVoUFp/ABQ8KoxGfM153hv49s6zAwy0QHqBhl4VfeZ0VYEDG1U/n3qo7ysMbnss0vv8KGUXS6nLh
oAJIzM+mXLeaapZnUTr7X1yI5QCIZrg466Vh1UAeU+zdswSKc9Ln9XS+jzkppGh74kvs+x0KgJ6b
drkFasWLp7QWdzJUweCbUdxsRjn641xgfVm8x7cWO1Zob5pUBMa6cw6JZdWEcqppMKeIY3en55H8
tX+lfFeA87cJ6uh65Y6kxiB1ZA8rwZUtze370dtEHm+Qu1hf269hGzW+ah8fUmjlI7+EekXYsFRA
s0+CM4hQA2KbQ5TehgAQcw2l2IOPJOsaVLOhL3hi/xcof73XNKSjSa4pebAohvMk6WLfctJmoqWR
tySZWaovlGgE1zm/EfLFMe8QaYNPEZNAF4LO6J6a7GZQzhbxbvnSAOG69gsHqcHcCpIeKQYjxjjH
HH/RAg0Z963htnGV97BTKRkKjqO24V0bXQzq4sbwRNib+O6dkpskDyYTYJkyv6LXDQ0B6LCaZDW4
T+yaJd0GRNpCuBG+ff2zJu+ksjc813+TXG7Qx8c2LLvNZr39M0aXXJrnHdgfUaKFZx6Wrtr2C8HQ
Z+gJt0SqZANjVusnf5PDS3IuHEde9mW9pldcuglKuAHn6O9IFeFx3+gOSJhtRCkkzIfIazD4kX5W
K8dyCvLaEyxl4EHBKai0pFCs+0Pu1dY2+ywPuAjgDf0n+HgPJm8kPsd/ChPqKBTQjTcHcgeY4OM5
cfLbp57kuijua/9bELbaiwdguLC4XE1/Zl3fEIz7M7Xsxzw70qGm5/ylL/TgDkydGX0QyUsVnmyh
tESuoCJ75nNmhOlH5eN3I61v/BOYMMtrTH9pkeR7zElZLgGANdzZXZYc4swpG1fS2TPEI7pGXm3m
5RHltK+HA5kaCygu289FGltaLgP5HiwU6vISuTzffsyffmfuBCyc2OhvEpC9R/nREiiKIDRICqiu
ct2HHPL91XkJJQALxQOkjAhyfETNHm3ue5Rr1vkK8U81PU042qQx8ZT2lVLf0B4G2wPs6v6F1XcZ
sMKXlsXsV2OLys0NSgOgwwRVkZMPf1efkv8/hLZIF/geSjhTCwm+e5mHP+b6hHSVSxeAIku6notS
Su0eSEkZPgC9m0I8k36TMOGQFGjl0gqyg0XEn9WXPGbOrYD4E7FkCFWtzn6uSpJyZhlGCfZX2/Yg
N0CB3YTiYrv8BwvefaPm5SRGi6f8fEMHz997uX4jkChCC7ndltha/zWktG+G0y8K58MfH1mZTflA
iHiS0/oFZhVL6xlSDmO0gi5QfM+Ebob6gdfc5sjIw0Bj8z3PsVxZzZ8m25mSPuX75SF5BGhcUrye
39RuJ763i9xCtTWPibChN5R/FAUw4neS/JwSZNht7T6DF2Ldyd42J1J1fRJGzWeehyUY83xo/lYv
XbzAk9DzIl22QjW+YnsN4I3OYz2rYwGDoY39FnLoAwce+eEkOeX6H/9GacAVgbO5L0WmcpJHIw1v
DL/y3AbeXiy5XfBxOxKW3FUvu4PM1Q9jfQibMPTZ7/yOHwEOC1bXQOQgCs+xyvmR7b/U1we2CCEY
iHdo3HY0Cvh1p4gOkfVQzCrZF/kkHVlj9VZntW5SiGYwx8NT9pGzdmgtOTPUiOMNQ9tpiNP9IZsH
PPUrXuXpFK/YUZAKUbmTqexL58G7IGCjtDeKpNJoAGaECsQK3EQJip2/Z6m1O8XA0dh7RMA/pJvn
2xaiyFz2Y8xSi+Qw9b+7hP0yiU2vo8JyCSkjtoJXtlI/pCgPCf5y/YtzHS9mu/sX3U6T4bVtmjQq
n/YKIZuXb2Pc9SmoQRrYDwrjsXRxc7g+qZWE4TEwgjzOSzmKNbHggpaqQz1m5elviyzk5kLQ5eon
lMg+onzHyJAy4piDRVa+cKwDP4Fk+F9s4EZrfZEEilEL36FFy1bmROgiC5UemstvM8tjIIjSE8SW
lBvppGtIlbJ70ubB7zwiXHMy4u5tk844CDHqea5iLgMkoQGn/c/IFs6+M0nN9QAhS5id6RiwiEiG
UmkazLGpaICrEplqkBoRI09LOU9RPl7FEGNiWttm7voKuu49N/pQ6ukjnC0/gln1MeNeinliNkk9
/N7Am1MtncCysFzQ4C6FA1OLuyDw6hecWvnaQzv4rw4z7a7DZTdniElTFnENZ39dluO9tqvlimNP
kWg3x3Rqc5csaMoS6/JQpFxRNGTRRkSuWJJ3IQ5TUvfkWq2izqD0kUxn7sgUtr2CrZRgTFT265gM
eX5hWaCl0ZD600yfgJeDPZUkT4Swb8TdH8ihuMijm80neUUPLA0+Zr0qV+tjfb7syon4qc9tlwKw
yz/wUy5rWLSLWUZ0BGGvGRgpRO+aSV55CzoxZ/+Ny3IkvTZD4ZUTaYxOaAc5D9OkVmlEs0N3MPTB
id0q9PMmxaQ6+3ZqGOpcL91NhsdwI3fv7uHWwJwsU1IK5EPRW9XbO86V0ilmUCZbK11md+4wdeZA
rtM43vzq2dxtei0tQ8ir7iOOTe4uppCrRl69VlZPz+4n1tXl5tipDHC+iGeLzhnRgbjXdDSr8n70
B34ZAw5OYLLONJgrvoxQGHWDPIKwtbcXB/gct1J8NYFAo+5vRJuChvqPtw7/5dKCDi8a5vEMU8jv
tDHo5sn+3p9WpYI6AkCQpCGk0H2zBn6MbvP5Gffi8YjgxMQD2+nIrlDRnb94vFxNTF4bAj5wIo8z
BWNiMPS8C2UUqkTgHdztKsWN6Vx/FyVZAvSeGGk7oZoNuSPaVoWaVrdxR3JfyepCklk3IfP2Sfsd
a4VcYveJcq3RtNVP3Yh1r0YFaEzkv/RMV5Y1rzlOV4Cl8QNmmH22AFHq2HJ13yfPkI3dk8HkhM/N
1qAyViAReIE9z93VBm/6KfJCCcc3J4/x1SgrgLqU1Mkar3ZT5AC66/RDniZ0/q5dS4wId13THEvj
Buf4kdGFS950BAhPgFK7sA0t7OtBLOD26t/13mNRHXOO5xunh8+EmwNUaMl82zte5ero4WJymQQg
NDPZK62BDw8ZcR+bDDn7aXkwBhOedcTxTqDSmZkvAUpXMytip+GVXqJFJEwhR0KFGyGD3CYqc1pc
Oc0n9BlfqytdaLwqmZmPxij9fLd7ovNv18r+wXQ5IdELC8IpQifesC3AEKrXf7QRvz6KpP52hV9W
JCTU7WKWrEaITLGT0sthjzxnA04QlzOjpNku9xQ/zifATzGXOtggBhp2sY+NMm5UecJ5mwS8dZJV
qjPzZRwUfm0fSLdA+o6va+AQiwTI0CrK4uFgtk7mMlnwcDI8emcsAVUED1w7vLkZxUWuBiYTT/33
sa/x9eD0Wj4s+uAy+H+KkjFq9V4QpY2CK/6s+n6J1z/2e3FpEWuT5lwXx6ef4zOJpx79BIZ2ofP7
6CPhck7e9VT0fj3cL9ySuo8hykYAA+jEQYzWVPDKia8OhQvMywoY3Qsuo6uhvDNDwBXJoeoSlOGb
1en+0wTURIDrxNwt2xs3t88nohAb+M1nRucBRVlhG3V8jDGFsMEZGNRuSmkA/xSddvWzs36yekVa
e2rPhn1aNqSut2rruFn3TYMcSuXs+jQdCPSvVYJ7uwa6/hJXDbX+96r+8REY73tzngaR4477h6jM
6BkPCG0qI2P1I3gGCPMMYuMoTLnIexNadXvOWyNhyfDqspaQxRspdZH7hrYxsJICriTlBUwBpQ6n
ayhXezBFh1QKqW5OOh50swmZbbDCD0PpcwtVONjUmbDaQ+pkyMFq9ubOe5+Nom5ZigRCdud0Xl/Q
qFo29ycx6lCai5bQMmo/kxnOkZ79NwAiG7/Zn1QXJvrIomeENitllEPG+mvYNvf2Xv1GBAWziI8Z
UjzcL/56csz5q1Lf7gI8kCVCqsYEZB0MJ1gFjuxSLV/J/7EmjrTsPvymDW4mhZAdHFvSVlK1QMKW
cn5C3dxGyVzqMsAa/JvhlbyWzHhJROLe9xNgZrlUOK1h1KIks+joiOw0NY8O0IIfTMovy1o0dHe+
RLx3cIijcUAsXSZHJUPDIBnKYje4tFkGFGNJvNup2Rr3CK8VvJBGONYR9aqhCMKYAAdRf36fWapb
8Pa1HrD0wr6zYA0vMMTdtcBXcpfqRJ3beQgt+AD1R605SvVfppY5rrSq2zvMfPu+aM+OH03g/UuG
Lc/ceqbgvz1beKCx5aNfTykVMu8irFXjqdri1yBQOKRcDCJBVmCZYUAXQG7nM1jB9V2kLPV3NMCB
SI+Y0mCdcfSt9E/IPF+uKPIIGtNxyyoRfQS3m6wX6+gKvG4vm0bqHRIobj+O2RkTgzpyeEAil59Y
bYVQQVdTByNNUwwLNDz/tgqCQ4+I8KKYBgun/1UF/vc8rIKLdBUb4VDrLx7NdFfqpHPSQDWITziw
psEG57BBK6QbnQEgPNarpMwOlDHHzb5gH3lgpmL7RR0SI7g7eb18cd+MX3b0PUs439IBfplUQLJ5
eKKUk/WOAOBAvqfBLPx3PnfDav5IKsPseNRlaipV8WQltfNEt+IWUsBaLM18JdkHlq4YGUuedPpC
b5ChuiDRyFMZNRQ8vgUMflHuvNN1FHgOGsUYx7zV4vjq5vp3nfHzHKj9yuU4RRNA74nzunp2STUl
nSqIuTHcLo7fl5w4Y3a99IL5zpFlJotXwnxNvI/WgA/mKCNaypgW4owtp+ChDrAtaK4eZwrkvhgN
9RjxI3owIWAuNZX+C6aK/ejSPfTCciYK2Goo/W2dOQkh/03BJW+JhEO7DluuKCDSXVjeLpBlHE/R
4uTFbo1lWkHG2FXoEheP+SBfqxDCEtb/CdA21viXPs3ckzu5zSN9p0l8GzIiZz2edXhfeBtYcAbt
bBaJokZLTXhTxUK779+JmGJItwyoHBaM58DvMoEWKpmorge9TRSCLnW/a+hdCWXY1bDBQxv/XEPU
2hQ6ahepQiwR6l5y7l+hyxvS8IxAuDpR6sDO2tFBxBBp5DSSxNrzDEzK90fwME8X+XIbnD2Asb+y
AX3XSXUsccOy0L/tOCitrQk+Qs0WJdygbj0APmfj0y5HyF8ZGFNiaN9289Uo1vNGBUg8oy4rh8gg
HaGFSqiW8KgARsvfeDs2rqlAbao5ULqbtWFDMtgdLYVat+P6i6yTH3cQI3IN6jI9d94IraPEZnTj
gFYe26zswmQkAAY68wsDqLOqVIe8Jf2vmfhhfnhepdt7tyAz9FyJLRWpDxYnjjskZqd2vMXdMtMN
RYpqviW12K8bGvFKe4xoSOxpR6sIGtQh+i5eWsyXu8nVAuYlwwE5oqBYFm0/03quAskA/H2+TIRb
33AEKYFrjojbI34gpI24yi1HzBw2qhQPGOG104lcuDtzkWDnaIBZ1bL7M5j1qBf8dZdWvfBO6iTA
RJ9EZDxwEX5u4BMJ54LK0kQu67z6fWNwIYILBOWbMyQx5IYVEP7RZcg3RUDbTC+2j3H5S4MXaDGd
rphRCG76xj0G+sjVpSBf4XwhPgEGcSnZqOwlLHGxs/54L9WW9DiqNawwgAgbHJx+5AUHNPZLn4im
r0llsKQXx43xAPJTrMejh8JBAF2dQUGu7NJXWoxc+e56X/h/Ckf/GdIe6UViK7ClNvLg5PQf+Rje
3ptpIHiHATouKgGkRv/oSpr6CRFthPcHyNm+nb9b4bHR6rqfl297hfGqKJh49t1V8cO0VsNqZaK/
WvuyHVyyPRg3gfOWsX3++76OxuvoeBrWQxyfIg5qxmkCrHMHxraWrYh/zlwFtk0KPgr3n7iYgZcS
V9O2BvkcDIm5ZvTFST8nNcF+N20Jg75KO3+QtQ9uXdBqsHl8CYp2jyaL6kaXWBe5VNYAmdfq8XtN
jmZkh0y01Z/Ra+mM3DESYGUO6AtGM9geZi0xhBiKJzKxQCFpHQpGBOdyEs8xmrI/zkppyvS8tIgu
gcQQQN7Sjw3fvDkQrNK3TcjdXKIDlp5VqG776jfCQ+Ccp159fFb9g6JZQtusiIi7JzfvB6Cwz0j8
p8mPh7Y6c8PIXPqhnxtoBwLCyCxArbh7fdVTN85wT9UzNnZXR7pgN153TXbguKRd6pqZ3YRWns0N
BBYMJ8TME4qF4U4F9KcDCRo2eY+Yqa9WqR1dEiEwOdI+Uf55oQSgZcCB1sAzzL5Gwai3eEsBzbvy
4RZCC9Dv+0sw2I4RksCiPKJ1+Lb2XfvcsXLk2eJnjpVawdF6uo8PXz3VuCmDF1/EWsdgK8CbA1bG
d8TmDEpHQwoIwxSs/ToSf41quKf16FDX/8MvtmSx7S669CJI3lnxT1+9jYb9jg3BzpBwFQqSDjxQ
Rc+x0P8YZ9FBU9zoP2Ug8upXCoxRXDVlYRIzulD8/ifaPtGZwTMHcJfBblq7srXxaONMhe428i0K
6JPsNh93iSMe3tAkuDUJgfGefnS/qXL8e7cnC1nVcLboOd0/OivvycrrzT54dqWUmYoKFCKPbN8a
3DprDFCjbqzbrt2RxrXesDvoAlpLbw20/R1ulvycFQrYqEXZuasywSqCeJZegWP8rmT60Mivjh3K
VnGt3onjYJoezTCqRuFiDCHYxpRQ1WHrL+yqywkP4EdsZ8B/VxorbXMClrTLPOPDpF2KbCFZY3Yg
naVj8VVXEdtivf+UgGoP3Xx28BvrjdwajnikJaqCtXZA7H7gTrDzykYId+zrUi3/XIBEpZRBFAjM
Q+K+AeHXe8141eu6z620ZBwyJZElXWpJHr1KT9xQf7dPMP4dZo5nauhHKugNb5IeMXwu5h/JntyP
Udsx6/eCBINJiuyAF5GBqo8bRPmhui8HJe6xKgdGHHT15aKHHsEwGYYLEXnoryIcZ3dRHnaAIYd2
d86eNiV54AMMnTIzDB2mXTU6M23a4Z0ekqILFfHkkXozISj9w2s5afcYvbJdr3lqshRwncIdarSH
nRf2Hr5bazGrtc+w3dH9Gkc19VUMftEYzPskpDASjQJN/OSt/XDA7GSWXbejT2gs/+rr7GcRXWSx
5jdYmgpOYGxjEZCfV/ry58FiZHa/Z8RpakhHg6xkp8eWuvO99ElvzSTGqb12xG+4T4CUH10IORD9
0TF/Q2l0K8q0EiPkzPKGv5L23ciTRgkPcnvyjgo/qd6hnSnM4Cg+mz1NAkKGd44ipNsZ+IbFOCRQ
YA/zn518uSO+28V+Ld6/dSWiiJAoSgCVOW5OTmBiX8Nk4JIMxefSPIL0vRNTN2z21+ENW2SqDC5e
32ZrkDojdUa6w4D+VpxeV/06H+hHYWDKI0o6AfLbOkxfFXTcce7iw6Vx4ql0tWu5Y/PjDKX4x6fZ
sNgE3aOl/uN6jZ0v4gYVUxMhjpPFG2C8v5JqgSmIG2QuE4gMtFOkXzF04jpUAouwUPY2+KkB5gPd
oVc6MyCiPtAWB5vU8EKcAHLy7U36Afvb6/arer7Nc8b9zaeYyA4S/IJ4dlD2yL/hETnKuJE2FUw0
EeNFYN6fpBEqe3HRcGcDeAgk2k7PNeOuuHXCJQXFuvqN1c3d/OT962dxtLKQ5+7HGNrfRU08dUU8
I0v1SbHpBg+Qk8Tr4ahuO42cxFtkyepswIV3HsllczXHMnC7gvhTeKnYjsM8R+Pv2vDtlTIvTGCI
C6/8j8Ju9yFpmQeE+L2h/XJWSZnrup5xrtbpBGUfOcu03g02tdb5CO/XmrYc/b56TdvUqLbwfJ78
OOnGYeMOG80VOZ2RTR/T+jXOrlkhDtQXoyeJNG7y7iD3ew1HDLuef6iESKWctPAeURPRRIm4SnWy
Wt8FjWvGVKFu9r5aRpRjLig5G6q/7MGoJEgM96dsrjxCeOg3mtrfvNYvYZNq3uLdcrzhSxMC3xEN
tqXqGuYVPCvs6hjQHqiYiM6Vs3aRegnKid9RtsTtGCjVDa9Wxl5GZq5ybn8EFIvOnc8nJTc/l26+
w1MUDmXN8GILt6NoxKPCbePyTD9Kx4sGYjECLrBiGH1xTJhEz1X+MirYLA4mLjdBfs+wuqhdPhop
PVB0p7kcZkxHeMK2rmBi0m5IwiSw//0GN5sPVUw1+NWsylFjB8vhhjLH+gcjgpNTlZqOzFnmEUtM
eqg5TBoxY3gmoLHIC5gyCvIOZy0TRIy8/If65cdaV36tUAzq9hXz0tU9ExlYy2ewmlDS7M2tt/SS
AWZzFLETu33nTW8RJTfg7cbxV1VytzdwiTKw7iKmSDXAi35lv3QRfycFCOk94m7nNIAmvnJ4xeGW
/W0lny4anBRy3vkD1g+3RmP6xvKCi8oYRVALKr4xsNsP85BQ3GlwFJtYWGRVzJNnqchOkK6v9c0v
gcfNNjbPgn7jXbwSVaEYKOb8pWoeIMOytXo9MFNJ8IDt/Isq8Gal0/Fr4Vj3ScGiu5hzw/4LK486
pYUyKBDulZ5X6ijkk3JTfIiIzszoK+foiTZL71IdyhCvJOdaTYWJAWvGUC9UCS1KJKFYFSqHtLmg
LUvlIuT3nZ5sBoVJIbn+MS8HOwSFIXT+feY+JNFS9vJe9HcE/Lgl4QySHe3IEYxbpAMRbSUqeyL8
om7WjeOK8iXNKO90gdtJ30mzP4DHz7itL7KZJnOHqzcHS5CnRyQHw5wd7VxnVmX/z4Tp8MpLmjAC
tuEM8e1bsKutkk0tryBxHKgmYKnDNe9AQqq1or5w8KgreY+DuxPVkRweMbp4k4oXKrwqDXpGScgC
AZmcuvPAOp1vPmAwuxbc2anXDQJ8mZdfQWG5i9cH3iVLknnozIyERzxWTu/kMI1Rm1ITd+Uq4Gt/
fGJTiBFshjb+4JC/lRcxQvLdjTQd0zQllBx+YlB8vu/l8ZL3+FgJjYqXAxBIQwIbtaPB/wgN0hDv
6lJT4h9Il9SejhFcOCGPOSEAGMwXd2H9CkiDTl0oGkG6BUNi2Y9JGqCcM/YI2Yn8ya0R/di+2PYo
GRMc40blEgHYTnewKopzZXdHa2HzOjZsaXkuWcw/c/bbHYJTe2zaVg5YazB2QpK3RQYKsta5sz7C
msxbcTiSP/VLkRvCUsrr3YKhoESFaNMk6QXN7PXRwquq2ugatHKsC0djSyWgfNBhO5XXp0F95Eks
JZOhiftAdj1/BK4M+LyYpftaOI/Tp79Fv1U6ZzlWyoJJVD+1i0ZlAQgN3uXJa5KzTZrNDNnTCfG3
LYRgMtdcuPIjaRlKsDMtkxagjO2rVY62g9zxjqHRyXtngmQGUW/1F9vtZxbqVLNCZ+eI5l6tqFJP
D/ASqSHqQo9Cl+5XZBDlQZhx23KBXld3FqrjK4RMrRts87a1i80V3Kr14HzLjxFZhISL5U8IlDmp
0aaj3heMHDB70NSnxMVbQ71U1ydAUCut/FC/VtBbJGJewFfIRifCkU/VuyFtRSC4UaJTz0RwjMNL
ErZsairqyANTheMfsDQEO/73ddFp7TyVKl6hzAhFhPWUgF4ns/03SIYJlLprgcPBffu9Q7p14Rfm
uIC58qMFWSQ7q+ipyWpmMxnfh7ctoaRCSWocVP716Itzuqq3z10NMAaGlHGEnMi4nGe/nFlR7WAp
15tu4TloDYR9gzgaY8NpY7HwREbV4/R0sD1cwnOWr+kQW/aXwsMJ7cpKiGUDNUa+o833ITn8uik6
rscgbEBJVrxUjmTrvsnFto05SL3NGoShqmq4QeFRDUbfiF4jONcPnr5FVBfJa4GUZsd1p0d+mueC
uykY4Zjvz/otf/VSY3N/joX53lWPgiHsXxtElYiNHXCdcoGP6joQtseRMr6Il1JlomApA1u8j/sv
98BEygH15/bhmzhtKBlTb42TK90ISCd7mRgeEUrZHp/fq9E77dA+ssHijrk9IfYRhwmVhacCYySh
e6v2bYI4juiEySlyv24XrBV2jpAh7PJfSTm452jyGChQ/XXmtn1S9KCmMuVyYIY2EAdv8p74rMpz
+yKgki+BW92weYfJM6kGlYuyyo9N8VxuMh9ezN8Oe1lBrR0i5NmVL4kXDIURcy7smzzUP0BFNkT1
D2c/lN4vB2z0/i1uP1zfikQD9xV3/VPOp/M4oyHLu+iEAfTh/i/3bPkD597GtevkI+FXa3xoV0bi
Z6eMPbBSpfbu+89jbmHBHK8cCztQD2Zrzk07K6UtF7mg/JPMXV+U192lydY3TKCDUbtnJlWa7S/9
ZTFwCmqh0lKHlHz1j85RQxh6WjHSmNRMldHNFqrGcXmuoaZcBf8DeWVjt+6eC34C1Q9oPuk49Ab+
1lyd1Yr1Z+v4JIorb456zBMvCDd7X5k+H4+KIwxRpw6XW1XbSc2JfL1Y5Iz69ZaV1AmVOjtJyu3V
CxoUF1b8n6oyq/4G/675sDUlvqUb+zk+y3n8v3T+tVBLr36RVgVYkFhvsDYKhr00X6d0uCAVU56o
+F7EGTQwB7bTJDxjjh/CacYZM+mN+zxPjNfg/3fJqBcsLG2+Or1m7nKWzi8F0YFC9fKwx/zBHm+E
Xk8iZyK+2QHJox3yZzZOHesErh2n+vbVgUJkxFNyJ5LIrt/nhXM1BCfcc4/LvDC/MCVn1IDZDOC4
gC8RBq5wBEsjsfxChOatRjRasCVjyfYuIi0BzjU0vKEcJ/H3fXpLxO8Zw/2pXBTcihmnuN2RHtcF
jlLYPrA0lno3BVcB2TYRx+bhTeU+YNBA1pzYprSVAclY8BTCz51DK7UzDMF0RrCv+SBRuOWWjHCg
jdiTbgMBg5TsS6A1jujkz6h71U/4Y79+5vQH1RdVXm5wEGgyssxPfLKHmai5cggJerBDuDYEpAVB
YDnTYL5UsYW2W9JbBVNVGxJ21s/5vfNx+n1htz4SMuRez917w+bfyk+S6NDuc+juV3LSQXK8xRMK
/phkcnZ/X4KGzGZ/6m9Tn1drQQKWld9qQ/m91xEXjZoIBVZlST7cVa7W1MH1w3N6VjQv6nfafByI
oxD2OFyK75xfpYsH2K9EnC7h73NTfT9vHrj+obawCzL4pTrEZmiGDQhhx3RWcWKAS6OLc6SiTcZX
EVZigiaRL6ldmdvXdkIsnT0OzQUx7M1+5HBP4Vm5GVdX9WD9Xpe7vhPnnoK+wHsXWYUOyRswT6AT
rNZs2WbSpntwDIuNi4XxE4voGVwA6CM3h4YOb0X2ergM6jbWDq9W5xvyiW17TsP3V9FEwQNsiRAU
jMKT3N71kRlc9Af7Ib0ERryI7GKBV+6eSQ9OWfGRXlW5sugKobn4Pk+JOtqNqhnc8j86HL2DDY0o
4e42EIqt15ejqKjp2uEz9sgNTYYeD4ni/9nJFxrzQOAA6wLmrONHEIfb/iRWB6eaJGmiDB0L6FZA
QIIWJgrEL5hEm7BsBKhQH/jRgZbyrUpTql40mK7bdbP+KSks0HjrEkHCbWaJu/Tc4DgJFmjRJuzY
8AI6w5rOCE5klmyKlRH+WufvEykTehuRgLi3eHmbR+tsxvWzikp2D546T/YfXnG1cB3iGV6lZB+/
gHhTIQI/EMHf0BLq9VsLy4lEeuzk9i4VROelrSzb86Ac4XYyvKHaJ8iYuWtWKBzzQednwZ5/71OH
bSAZ8cdgNRMzkOlvWtdwZdm/wUoIvHqH+WzRUXkz/CGw7a8dzaOGzD1Qjro3RKRcz1bfWRCMoTAh
Y/7ARmis72WTITSaj3k32Xu4jXop51Ziu7yNnw4yLbkL9nmMY33vKD9mOcv4PHblcq37JTgkuPGn
4HyyNpxORULTOTkHCjqcfDAd2/lPZfSdTX2kpDs3Cxlxkz2X6gEF6ZNRAp4gWFICF1f54DGBR/Ae
BVsQ35NprU0itIrYdLGF5ek7j83/1qUh/fLi1s0f92UFfv/l2J8FpVNuXUIKwJWuvkSgukQP6/x/
vP5oLqkvq9HN41KrKtv7kwyDfw69wNtN2HxC37ujpyIfBUX2+7Qy7WBGX2Npee/Ttl6xc7ymQ0mU
5GN6YQI4O524VXp3TYdZ8ecYufE7uk/rndHwknvUwlrCAK2bZ9XRt1W5YT4ZJvwb19TjlepdNRTe
xkAVo08ND5Fu4vSTHlylU9p8V/1YRz8kJSrt0wEbc/bfIY1xgjI8lh3vKfTCw8QfImh4tZQD4aKH
GTSTRKwpH7MAplwhed0FthgEwNtlV0Y+GtvDs4PpBUWMBoUX7Uwp244zRlYbJnXcP/ZR1BXGShxR
zseZz8goRl79eEiFOEL1PaE+AXV9HDPEYdPG9SEP4v+XjjCx43w5aQPvj8R95O2XavufvLZ5tVME
Pn9iFC3/WrTv0Cu9UnrlgxnOYh70dIyNfPGiXMwbO4i+sBYK+/3I9O1gwG4l66zXiATUTVDatVsC
FzSNq97hhgDaY+tvfZs8/YZlfQbGVRukL/l9vPOePCOWfmByR9g7wb6awkmYMp8je6f2EmeuHnPS
lEoauphO+zuTkm/hkfSYvIgRN9ir7hMetfzcny6RgM7BLMFg/eCjqkIyZKX4ZRMiOVP8WWj2o7e7
RtLA1d94bwnOzwhDQgdH0tRo8BJdb7bgXFT4mWrEr8yWInNLgFQX8xkOgWBNEbh1j53TXU4bw3xT
iQRjeW88R6pOZrJZMB1n1+O4shmdhUD0WgfYn5o3jV8IvmumH376wD10L/BsVhuvHWHhw9C728Th
T5HT+2/cnHA7gK0v7iCggkgXv5+zkpJT5dKthnAL3jMWBCspwAthOw8o6AwVo5+WUKef/gbqnDx0
pON9I/ZHUWl1zUBkGxVnjsZPkQmwXDM5q7RFxvY8LnsscPYqG7ANLjngV+EW7WbCHOgGLnA0Udyc
QKffgm0/EdjlXHSLIIpXWxzCiouWgN76yetj3uIcnT1NMPlhGcIFRydZNNZsTnB7+aRuxLECdO9n
/ozTmQRd2MVUrmuIB0GfPLPcv5f07PAx3CiZvkX1BT5LWXKdevFjxDxfDGeLNmqldqYojTd13tfN
AomhEpqIcw/0YngQPlGaY/QMVLrikckVIfkGyOFHUhNZ3KuqBY/KYKzG5sawKUcxBlxWcBKxi+su
uTEzms8ZzKnGc3oWb0bwrgXhFgQ/MRYEs1KnPq7pB3We6eM1+2JRg2ZP+4UGp9BIE7R9wvwyRJEI
sefOL/RKkWSfcV6c1r5H3+f+vQJJhbbuWp8IGsRjdO6h923FxC3mmWINOwIjJJZvBDLGAP/m0Nyg
sSoTSJUmca6MO3Wm0ObBzm1uaSf91RtN6dW5s8xXvzvrPca9waCpVE//uf53GAaL4243RR0GpO+s
Sj/DxCkqOVTENlVxqD+3AgeG4UoPUrFPGHCdwSvlQZRCbMmIjA3nQpgRcyClxSh8NEF5bszKB+Hl
qsVrQeUuBZ3E48uSydQptkjzvCnLBuN4sss6DrsHZ14EkGbpObLu5mFGqqNwl4J5fJcipQzv683y
boLbh3nEevIps1eXCAu6fT2gbR3ZHuFT7yhupEGwsXcuxrqyzWU3S6ABTeBAp08Gb7HPDeRHVIhr
24Um5dfCcv3go1rzGHpv/hTP43hlGstTMyLRYHBE78lP5MPOHJ6bVT3uTgOznPTLg8ALSYbuSsF2
gA2b8Vxo7LtouZUCLOb9Z0Eo1Bi/yRuH4D41wIoxnkZNLs8kqbpDkBcwdDYPq8CGnuk2LExtQsdL
jBMv4Hjl6ILTZan0maNjJZRg0FYcWVfimiprZ8qKGSPLILi65c+Dc37BoVZQOZKuRr5iHmD4in/F
IYJGXPqN5QtrA56jQ5vTj0qeG38YYdUfl4veZ6zziyw3oXcPDZF15ydciHoJbftAav6PMCCAc6Fp
pe2faPfBQaZ7+dOAoLBqXnRBcH8XxxBddrJTqWH7vwqyi7GSBB+gQW6aAXVDEpZy6lE8/wi1hd/H
435L4fuMpCu33Aaamn4g9bP9wcy9PrwRXqlcmSbjnVP4tylYIdkkikBZcaIK/7s1ctXsQhQoNLlh
BhJCubvswTfGivFVs62zBB8fErMfENAztHps3+mRC7NW9MIZjtplh0UkHkquKbkq9dLm9JQhTMH+
gTt9akpBBFLfm3qnObxmGx52S8eRFbPk1/1gLJqQceryAAdmUaUcat6D21xOny+AjRNCtacYDMc0
rMYVusqd2s6nuMtgy6033iHdU0aINaqNabgL7BJGrRN/RobYo3E9DBeBJ+cpADcavQ18fE8w3MFY
9904gRki1Zh/F63BATWqwXEiKrzp6Jdl+NhBa4emoOMe4X/RglAHer33z/r4umOXeBgbvrqURZ1Q
xgU+0AjxhmYXjppiNAELC3m7tnYCE96WTc+VRdbX3WldtyQTSA5VtQed0e1fb39eAzOwL94jf/o/
fkWFlYQ6heyNgLlioV9tJ1GvCbcwyFKiNIYNqoAdE84WruhKj8dbix40OzC8JLTChlaKF3X3XfHx
8lR+OlT8/NQWxCjhAOujuZrvRPhBfkW8iB+VkPwHFwGVMi2sYi1DaeSeBomodBZp+U1hzTKTroLG
k5HrdD311XyaA4tZyxwpVhEAWWyOEzNUEw9w9hr9HW7eG8BWtwb6pyKx95wdxhwlcEswdwiB9uUV
I/xMW9eLOsY7/x+PUPV0LAIHeboZr1pfUEw6/RHEBETm5HiwccnclJCNLKwyb2P0p5YKcACwQ1m+
4qxXHxFxcaNIY0QBlOkNU3qJfzw9HTM4EoxK244Q13iulNE64G2j8OV3oPJ6Mdc0jtazl5TeYC63
MJF3dYWOEowp/vzuZIIRj3iw/p1UM9c/Oh4c9kTeb/wir/l6EKcDwnDtqKLG0BRGJl1ZE3dUIOIp
0pDLjTOGEYVRZGcYxLcrhDWXcDSzy+B6KYn/u9VU8SP1sdDihSXDm+Ht+HsMViAMmBnDnMjyv67Y
4Ak6guIbyoymcxEIskEZsUJPwhnMcHZQfyNghDwJUyp7rGY79p6twzV/ZU75/0iAnXkTItLcAvrq
CMlyRii1t8uBt+rRZyKv1JiglIQ/piJS5r4Mbw1gdz3JqTjl1XwenT03fcBn5bXcZZwWThOHgmKY
w6vY1SYEJJ4yOTTm9tp5LtkIKdnMFuSBUms5UxGt8mRqP+xn7dJ2fT9skNTZBwd+1p9r8I9iV2Yr
mI68y2bgFL1QgfufNgQ21jYsvQFZjiXYXUErS1SlPJcRccW7rPSHessOHly4F3k45m4rbdW6dIrP
Cz1t872Ndv9dvY1rzXyExhfYySweZ64pBnspOD5x7kuNfBn910TzHdUAGhitW6ZCcAzbhQ5cS+1P
QIS3Eq6XL2q0xn2+2lR7R0apH4mg/fnTSdqp05BMDC8HXMxlmYW6/QEqeSGlaKfdlT69HA9RTsl6
yEppLfZx+68g6NNf2wlvFBuHYXdSCWZZkUO6f1cUlAe30dHGZvhObu0KL7a9+y29NkGKuV2M+RbD
40sxVcTd/XBGNLeYOehQEjDXENyeB2vTHLhmIccz7/7kGWK6ciyK1dACrVLNswpJYhHqj5plo70p
1fZqxxxq/tqZJCv8t2RyCYNkGsVExwM21bVUnf5NHCqHiXGtIgC3AVC2Tmwq34dsWUwjmnJP8nKb
P+HzsIHadFiZV+p39PSBiWP3mvLisEBbKF11Kd7wR+kf1SW+RtPK41BtCVC61qcXzSEPlqKZqCEH
gyypkxiZoC/Aq4GJbHe6Itza+CB0OaFE02U4Vs4cIs3Y6pLkATspKBZEPrHqZGMqbRaZmvWcU52e
I6UqgcOtdgDA1j8F8guAjmy8XWVuZIcrYhDwypsgQiRyiWix1xB+WC/AnJ4luxpKLq1n1KEylMLW
FE137R5CtJ0U/xn6UWBG/gjDmFAsmfLOpz/t8gaSlNNYWq3PS41StJe6iXIKnaWOFFiPWWf4OBnK
pMLMXqI4S+KyT3xm6cLa0dSVumCwYBF3GcB/E5xJrVrSM/Z5y1kQ08SaA/088FSzNvCfG1LINVqP
+AEcZDGZTvOFlXvmeF9V2nKpoKDi+jfuM3MhMlZDmg/5KERsXpBrxru6i0zLrwxTRQzFVhMLxcVz
y1pnKt/5ViMYnreG06V/v92qN0vDQi4KIoeVH1xXZ+nQjYRYM772FfIDWsIaVH1tJtY1vcym1s7g
rJP0/vE19UVsj+V72ZnZRI5Iwtl8JSWHY2DfEgx1Fr5mbTf5eZuXXZXKIo8rssWzihLEdrMeTpge
7kvEDncuNOuqth5yY0GSahKwl8vEyqHsCSNFO4p40Ufz+Jd+5fk0zT3I3CNs47m7L9NbLnvKoyQO
OxvUT4OmABY49u28PkIxp+3rufYhGwVZofsoTVxNeLbDFlm+GdudxoLP6QqRSjceworaFv0jvczM
zIhxn7uasDaACx1Ti2zGw4YXYXeG/QfHAItrquues5jBnNBVsVNH5Da3GAabnoGrNOiyNRGtlzrF
GJLMVTHg8z14SU9AQ8hR3CU/WXxXYh7TG0+HS+/HtxQ5m4JwKXiumDLuTytnqJoNLHnR4MSRkZto
JnqIKYjnB9tUKaMEnbvEXgUIc+t3VheERXZ/DJdq3LVH5d/KQnWnOOExH246eNO5UFNg5tapK2Jf
AeKLtJPBdtCCTa0LoNA+hWtX69IAwNfOfB7Dsy/Kwf3TAZ9UM4HG7akzXs66T55WZrYvlSGdETxG
UUep975l5wM2NKt0riN+tWHIrxC24FipOjnDe3vX8htvz7N0JjcSgfqQifgALDIGRVxjr2vcqPqY
gh1izoasWaDnaIWeaHdBgBBkdA+F7hx9kZjFxDDFSsJ4n33O7XquII4vdopGisRSTJIxJ3FlLIWE
pCgI592/wAqXI+UPZPFbSk/hMI800TWQAfr0XYJV0cU55Ln6x98DEA6aWFvHE6082f9JEwj135RU
NoHxv0bDFHS/yQLwbNFt97a7896NUEg40vqwUkvsHYC7bW6EVy77W3GZt0FKCovJiJhMTQFK8iYx
c2mj+a5WWnMK8853WoCHiuDydQmdpZK4us8WZnNdNJ/eu6V4Aa+K56v8OD+YoSF9NgIvzkd8xMSf
0QGAoMs56hAyIa/NLujgdIUSjt/oX5So5PCVyXRj7FJEyOy5ARrMY3VfhE7Jul0H3Zzc51XJDZKp
Dg0Oz83p8OGKDGr+DhqPQgRbhcvv8v2UR5wdp2AJMKeTKyzm1HaRj124qKpI+VrgM0NchIWbrX96
UAkbBYjXPS6/4/ZqExdKML5sAGiUHFVb/gqqQF9ghG2yA/mH9otWTU4OD3QFRGA4ezdzHjgjYRgW
MEeL0qC0yvXy1sFQ4a3UzH/1C+agb3/Y4fbGC666F2oltTIA1WpDrv1gfCaU6gbsz3miJdtjYgQN
hAyQshRHUKYXTqrTwDK5oKXIDAY/+iGJXjGd5RGLBkkPDa/P7kKC8RuxFl67qAdWuK+OIMPkmcs9
ytPuhWs3x3mdnw3C6Wny143cqAza1Q8IlLAvIpXeyaYSSNAegqNz+OUjMphNR19R3hPC5KMbXqzB
QgK4mHlKVpk4Ey27qK6EdTcwgb+41ayfIFyYAgWPQeXQsZvPIonvu1mdRyxMeyn97UVUDfmniW7k
HH7Kt9Ypj+mZ8BfpN4svZ5bEy4MlWUlhk+9jr614v2FimvGGKPLZ06dy1dzdHDsObfO/DJ1z/K5u
71+bGmlAA9ikPBC0CskobyP8Bo3x9Tze0amrUmA4Snd7U9q7pjOPnmxjIY5/Fo1ulBwW6RkubHn3
wyZOnjbmKisgeaTTHL8oc9eD7MmilOoczK40cnQm9EuYvRjX+d5N29e9l6qt4fJ7CT35voYCboXD
X7JpW/HELu3O1pF7mUshVylnFjOkN5NhqgX/9RVAq6TzCxt+2PfPltNz6OdC5VngDU43FNV58F1d
p2GFbmoEicUAvGXiR3rgRkpaHMKAlZUNakDDw9YG09VcvwnfnNfX5Btl6DRVAFmW4vwa/kFSccHT
GuBbJI6IqJ9wQ6wIN16vrRFklX6RJ+HC8f8lsDWZOLMqZSgsL4LSLsjj9MFaynuxzXu7KP7r84s+
2VI7gADlS5CaCSvU1AnEWFqRmHO6gDXcORIxL4SDpZ6b771xUGHYfCnoeJZ20XaSXdOtFgETbAR9
e0GkFORLU/nwvq5Kv6P2pSZLLyn0lW9GcQyKXLh5e5d8ENOAcAUiAOM6LfeK/p0VFxgeAAuSvUUG
xdKRleAbJanvnHAGr+wC7TwodvSIj7pxezb0xp8qTnI6p7An7edGo+2+n5rKCm+u16CZ5jlSzXH9
wnOzDpELKyT7dJcydWC+JgyMvLwMrCKp4KBqZi4P2Yz/Xf+rO0woUQZSrmO6aMQZCiLqoGz9fqd2
8kZVj117B20X6RSEPv7u86CytW45DXDNmDlMNYMzxeFDmFaqs/qZ+G+QDLaY/bLsQbrEqmC5/0wy
hirEKm1xR/rmY2Dqyoh5qBKn3mHTRLAsSxrFViIASXQR1WVB/DdzO/MszUeZfaC8iLS9CZmCZOWY
8uVBurBpkxRAsciixLIHsgRvKUpwroNPSUgLL9ITGAX3TKZbQhA7EbBs3xWwI/Z7AGQb2G+dt0Jf
PSMZLT64brZTizfgJLpvDmn7RyPPRPEpXY41LW1T83GFDjeb2iExetqIbKyJDM/ljHozMCPwvdD+
1Hgo0bkvEBjpd/H4M68JXZFLZXmgh74g2p/51BTjiTKfSAzh9e7B2bdkkoUWEjRWPXxQ7D++++C4
h5oF3sASIKkcCa+LinWbu70UB9Jgv2cecgzkxLXpIlaQNsmsXbsMwGmihgdHvCTejr2oDj33Z+Se
t+fV6VfDASXklpDZDIw6uhOQ0n9l6gyPqu1Bx4LFGOkorPooAsRNdLvMspklWGoawanXHX2P4+im
8A8gXY/sllKYp/bxttSdBWu+SKkomJQeoTEk14k2u/x9WqxN0AQvAWem4c1JOa2oWtn+9LAPxoPA
53S+MMiDvjM7sKw2LU+tdZncqjIqZ+dT6Fz/AgaVG2kmiOITL8GWcDwump5TPWeY40jslcv/PqbR
JuD6BjKiEn7LYwDgxWffkKwMPHdNNhOfr9m4n+fZbttnmf0WqVfuu4dCAkJ/sot4Hd4OUGzTo9MQ
n/4GJRkZtjcC2A2P2s+tidqsZFS0qsn6XUegQygQX1U9jPnb0tLiYndsYbnDPwlo4MuOM5fmXn4k
M65vFS2kxcY3q13vtRQO+ctz7uPo8wNgZ6YnjvqNPbL/Hp0qbogAYVnTTwxNNwxvAQ5qolG4cTbY
fL1RiCnKiMXr6B/I3B5sOzx+xALPwbvRUXpU0Y/zq98dRtu9PkJRNEuLzThnpYKs4mPWBNVOLaZr
yFaH+0+ldUHHSbpkQs6m51MUUS4kfJ5qlzIpiUQOzKggjNSQWWX2RFmArO4lrZkqzc+yC7RXui+s
UDgbniyy1vJlyLtyFzlH/01PqDVjc/dTvx0uVXbsBsxSxIrjUR+KG8fzAvsx9VJoJvAZk6DcJ9f8
wyhDJwWteAFrY5tSOsMSSj5u9Bqdyp75VR8K0lE2UF+HPt7kNDp0FhSmF6hA1gMtEgd4excZymOV
SXsYgdEOWm2jCLpqC2cZtLGoX1DjNnMRyoZQHBS31ppJmTpAqb7XkTTpV65MAhKdrxPKJwtZWuAM
l67fe0wMgT5UXj4MTEHzlwBk3b4ZMLqgnUIeacOKtkB81DFKqD9XS8+10eaSzMnVsWVu+RF3Fpe0
do71vxKNh6Hf6lZWJ4txMj56nNj0O4KrhzOVEfpTK9kJHO4RxojJXZSriZqL0t8AVlTeIgW8iYHZ
xRQTOoTUFT/SpPs0hvX6b1kqudKieqWpEMP70+MuOB4t1xIxjkES9vKRmHYEYLpPNUNI/Z3LZ8nY
1eIPCyjvBDwYEEmsyY+ffP/icnIziL0BkGUAMPQjiPrjCBfypfWapC/PAlpVLRTXC/QHk0L4/rh6
7QDNY81M/H3bzPkHpFcwFtLRf2gn4ffvysbhKAzjtUwwLQ3IPLNipFupG/MJ/vJmO3KgPCMWw5yn
pn9K6sAdm4hO3Aj6vRNvEAHLmaSN24I5S5c/4aT/gqCt4kxIK4XSh+w6np5ueC9LTMN28Ux2qVTV
vIdZ7m4K2BSYQ18zTAo2Ej+Q110PJVtdFuUoSOJDm1DjaLD7AHIphlVb+FdZeuO8+4MOAz+FIyS5
Y1Dlb3h9Ni6yLwNmctHYv0le9zopDR1xkgMzAR5GHAQxtRWBQwto7JCLG8UiwozTtI5LgD+bHPlq
oynOrtnmj1KAp+gJEx4gR2X+K9dTSKypO6baadhb7ih3FYVbcNl65BV0VNc50xexTmKNK0bYrfuc
WtGyG//cnybF8zYevJcp7qNwBu6mfCu0on7kXzrJmqbSW6KA68ErcBktlFDET9N4+uGfhBiGz6/I
NA23UPglNaP2ANPUVbD4wV6G0ez/NHAU/5LGCAYKe41yu3LgQZMTJiD81K7950Mc0AOhjuIKvC1K
uDLibLYH5FTYPkZIgOvxXzcLzdC5aeo9VQWxdk7xiw2ZZNujTdziiHrN6DCkOasZv+IjldbzbQlK
MrsOCYaYLB50os1FA7LXBn5ePd1rpke/WVQKjqXYb6hDiM95OX3G4UAZnSZfRVJmCC4JCSdFX/oE
B+iavI605c8pxO8dBxjk4NgBrw8hHjFWiIOAnWbc7woAV8xKD+keFCAh48RNljdZca1LigSS9CW2
gqXfJsHVCLlLJnM30RX6cdoFASxavNoHMxulfHIlDBHvpTxyd7IgJAc6B3XCaA+DVxzH4HMB9A3M
pg+Rw5tNRMn40l0bB8V5xsFaCGv38U2KK3RTPjGFNq82H/qWNnNNOTm5eSHs9iSctrlmrKuHZ0PA
Q+3Y3yahIiHQ6zQ9PFta7MJGgZiSJCv+gxJ+lgGADimC6agayVXal5xI/7iwxtI4ChsVeUmrpPH3
LNS0tqQwO0v+n4si+q5v/Rq5DkSn4LB9SU69cf2QQUq51FJTjghbZohGF+Ld62pUYfn4Mg3fcLXB
PioNpjcfodhr0eWaR2A83URUr62v/kwDenOYnrCPswVgUWgL17AzKy6JpqSncrls/iO9AZ/3ivxJ
9EZRDzSWibdp0sxvPPb6vbJOR1wcdf3p442SKZOd+F62h4sb/khy85Wk4jlDUaUnfblKUSIBjmfM
ELl32DBixY0ysQRc5bULvLlMuV2xZlvw2YL5lDjKk7VTvneRRix1SHrzh/KbBfVblb3TibrHtUYe
ZoiwvkTLNKwujUN3WTCL8btpm7gWScb29ydkXM2MOljJyOCTk7LqFaJVuCAOnB1LHXtb5FYciP30
i5Y4mChc03HBxscwnn2nqokyxw+hnyYnRNA/H2vwy7JLwLFB1x4JYF/lbL6g9WYOdv+zQG9VU2jx
AxefK4qS1udoWRVKfj1+e/odpstRqYy9LU7AjdonUYgHKUQGtAcAp6MsMrp13yzpBid9neXZFCF2
jxrNI5wX+OjS9iOjHNbQlLUbRfVDEaEy9FV/Eurne5UvmSLW/Djqo+VMhjlWR9FuUD5isjHSBx31
afHxmiF5yXLjc6Ajbe1vcnLts2kG4Wf6fnG2tWUkS6OOohfP1BsISZx43i2tgI+BTsC7nlM9l5ya
CvbDGLqWpANlVLWOaW5ShlURI019MCwSGBV4PVtmwXhrRtVjcYdw1mWGAMtGoJQlrbyGxAnkVWqm
ZkOfUli+hHNcFtdIbpZjRMS2Na2QbC7b4P7jz2eKAPd/c8ZxuycWU3jN7BeIIfvy+IBLaB7K9Mhs
Pkoq4rfKDJzo/jmCpmSD6cpGfysdP8zC6PUVwngePVooJQ7o8dKVzUV3T1nj8u/Mrc4jKhK2hAQX
wCoSerNTjg42EO0B9Z3YU10txlHBSDaL6L5/5nQnqJSVJj48ZacZ22FJ8z4sx0o3Djrcb8e3+m25
HMeu1YOK26iQdwCVN19LgaCuoKuvyW9zGJoAspaRx7Kv4BoGIA9Xl1b6wJvtVdPCmzTLZHe7+987
8ABLbe4UPKTT6giD5NQjV4gErkQ3zNCBzF31R6VmYGj/Os1cQOlOQ+9Q71UYUuyo7GTSCCxUPvsa
uukblrR5RvY0/7q37rNUfzBr487myLKH0f6DR/M51eOcuQNZ/CYGds+4aP+yexi2Qm16bJaTOaTi
T9yIkFnkxNHo60MsssuOWSQtMb1TkBA8qZRyN3WhwWADTio0KA0HPVAxy2+2+pkdCGVp9ujfpFEJ
D0PweuKceDzeC7h1o8uyYnPIttvMLyelMppl+5lzzaHCPgrZSKtfzRq+LC9zOIb1QmxLpm2lQA+/
1lvRaJo48ZVgeh/0Pb0H/PzNwtr/yduzgH6V2b0IWoE6DMg7zIvzoq+dqVuTxHz6oR9EeaC6SvTN
kkNI6fq9POUIgfFXtipOkYia7wDeApO+Ioe9p9Hu6H24zaiiNDnZuFzmjoN/4ZVS9N+Dh9CO4juu
IJ7l9xat4z7gSt8kJoRWQfTwsDpUcNi5S8P0mtykUYdFf6obFKEAc2vu00oksf4bYRAux91G5qrp
ATrVZSS1QIVgPykg2upZTaenDcxOEVy9Ui8nNx4ZM2cstNjNf/pMdEJbDS7ku2f4r3VSrrrq60J9
0/b6SU+cpsjBMjwIGvIYuPfufVE/4iThOpz5hYHGe98fnI+lSDE1FCE0YN9aAKBJx+MVOKIEzTp8
3S+vjFZZ2Ok3svN7H5chmv0jEvTiD3DaFDn2E0IUagEZdwNjHku3a0hOPM/fQ6O/+eNG1ZEVx3J4
56Xfdpy0DAGlxQSqHv/WYshamedsmwWPQqAmKb3107U+work+F9y0DSt7mN41d9TWw4NoSB+/wlj
h2XQlfPCS87+CtUx6i18s3F3Oxjab4dV8jpQThpZ9d45lfomS99oVu4ks37SdErHaZ2MX+90crki
NzvWCW4NndOlSqhCBzbjCgw/AhRFt1pUhQy0slTfQoCt0hlKtrEWnZXCdIChpOhNga5wf0z/G6Tp
n07Tc5jAPen+mFRzHiGbQ0MNoWNZ6Yb6jAc0APcKyOmCIxbo8eNmXxMBSHKm1P+Mtbx7EumhUglD
kZhKGSOWS9i76h3+++T0Vj3qoafUY+SMk7AaicvmjpISs3a8vyPulhRlro/EJ62Eh8LroEFd7/s9
fKQPvKxGh1yGa0Af5JXZM1CMZoJbTgvCSJKMc2EBDn7q37zh6J0w0LPKbcbxa1RfVrRaVovfzUF+
8sJ0I+TUCxNErh1FjuT1F+pfdjypvVBGPCfGa4oN+wvCKEZcKSjb70tJ45HsgAWz9qqi8lOkpRrX
ONWD8auW12OR6/AUZI2fZpwojpgt5KsLdklCVxYmUfO7Bbg0A9UniekV65zadTrbBfyIUIfyuPgW
ojexECogkvpVsYTFveUbEroP1rrsIRyFIWdqKoAqbJd4aFD7U0GCKih4dSijhHVRywq7aIlKak6a
XQk07yFn+DLeXNK/rNAvC73ooyx8IRONDUF7/dF6+FSzrU8sZU8XsGY9xx8wkzb2MKevTfQJSbQu
ue4kQ/WfcvQyDaUTVL+82dq72SPyOtrP5/eV65N/dBcQ8dEx9Tv1nOS7udEslLRh3Em4ajVqTssk
OhlVNVb2fJeNmwbNohqqToIhAK4nMSJEqmVALa1djSw+e9/ZwX4VwR4mPc2cZJ8IutKMEzdveplE
+JAnrVSkRCP2NZalYXEaOa3OCOiFnrqoiL6Vh0M1YkGl6miXOy/xpgFGSyW28a7/JM0DoOVs51ZW
68545weYhlybzeKqPSMvdEXRkJi4oO8y3hcnGF2OReJK96vnvlAyXzCgyFfHwaHOrqr8Ltk6qz7Q
VtgwoZKAuECrYFSuHaWagN+hggIlLPre3Z/kt6ymfueKGBCtE9yH8iDZ5ykP4iz9ZVT916utzg30
7I1QN6IiwPUOWFtXeVVonBXtmeiqeJyCs5oAxSlX7dLiYPQ2qU1jVO3jDxrhmPBN5zIbcMfS9QfJ
EhTVIBrvbvEc8JVAGcvkgC9NIaIAknBde7xH2OxN5XfOEJkWkTkB4dvlBKFHzxtA6H4j2AIZULOG
cTzvBPd2dqH7X6iDJTfSg0+dY58xDKa4XbKoWnqTD7m/OtEeOl3X7e4CuY4dL2l4VfXdZdPFZIU6
PdJf/FO1pZlSUM9WXPOomn5HhsCgiMbSoloZ0ZOwhWU1te8RFIH5958cNQjQuN3lq6Zi1yz78fJl
cpvzYP1p8Rp6JQ527XsgfeRKcWEmmwP4Y/fi/87RH31x68MzKB7O9ve/Jxyoh9rsPUtva6jo2OH/
oYeQtqbOfXaPWNnHd0A7AR5rqvQ6Craqu90aTQVUktSpZJLjbXSxjoKVQVpPxKyVAPwL1nr3pqz2
uH920uF7OrpAyHVXpHu6VgpWCspf7ye6CUi4XnhxvxdQytihMSajY6XsvJGSkWqjcEYSLskrQvp2
FhXVOho3bLJeODzNDIbcRIjNYCr0tUkjFCDu87aw53OCKi0OVWmkI6zRTSTjKYEFtRftmd8qpLmd
R7+jX89KHgIuAlgmmCrKt3DkIj53DmfImMvRCyd7dWvSEA3XYidDx9MFGwnt4xYa/ky3nuPotbuV
ySI5rWVAvOcfobaIMWmz3lQig7yQlLbuB5VFvJk+9PwXUs9WdML/awj8WPX2epKuz34cre7o6p1T
QxSTLtkhyzZujK+HxYArLDnxjfbPKRnHSE7HgDxvXxKBPHYk/MEMpV+vP+8AS9irZ67M64aDDXGg
0RJkirE6SVFyinAsYTIKbxoshiLSllrDpUqhgEmQJ9OnR7hJh0cy1Ho3gLaWnfMecVuOycFnPiuV
V5K9ci0km44XZiOihgWNrSQiBPeOV7IRmsDERpriXLld1QUs6TYl5fDPaJ0TRboJoNA8mu99wdbW
MXwmYgFHZs03Vu7d+jf5t3iMowsWv4gQzZ70rpKWrLLpnyCK0f/QrPsJjK0sg5hEVjnUpSq5ljec
15KFgoSNlj6VqDvaIYmUn5aeoT/taQq/OgeqPbYuuemLMnA+xDMYNTz76zoXvRe5ushke/wz83rz
jjBLZCyn3+qXKizYiIvlmpqTT8aLKdix+I7s1yaJKCx1OjaHEwwzuelAD5Ddb5ip3zxbcOswLNUp
CfOaZmjDFQA1UEwlEThPbyLL+au1XBy2WgfUr7GCTIzzx8sSTP3VVbAzPdiIfKhCIK63G8j1i8T6
1CVEtc85pxm325daM6R2vfqSrOS0AAuNP6ye2JFB8BNTTZjJrltiRONEG1/Kc8HpP948QJ5bQYJQ
KWQa0tF263mnyLd6/ltT0EOFkHbQQMW6SB2r3WasxXVU8mnSfR4SnVqyOuQ/X0Lq7jNl/TYLN+10
8J8VQxtidByRVaVG+HA90T6hdVw2ZtLWaf7zCEA03K10fzo2We9G6b4Q3RQxox4GcDNdfUYuzJjS
TEmQmkFbDZ/54uv1N268979e7ieatS5F/A9BR+amcsC6nZziBe5Sxg6GndnXMS+WAnlqVxJlO2fN
9d7mVCW6CNTZoTs2soBbsr7YdC69MtxapotBZo5XVPM/fVSzNkx95zdXW52K/elq4HUKxv8FhvdG
tdwmAgEC8NPWGDVT7+OwR3Y+IPN7+/hzDf1V8WO6U4Njkp/BdQFTI71b3Ftb8jkUwixOhqsOKVGL
VddGkrGx3MFVxZ37/3aY5u+hnaiA0oSC9pQ2N/i0Cx8S59in82coDCz8uAYERtmqysnSVUIkTeYJ
uX7f4oqweael3SMGNWDj4ajR/1zG4N3Qu128JFHC4Y11d6xHEL8qj22dc0WROraV7bKmVptwqnuL
kLqo5IeeuvUfs9PITyRbBsd+X2sCMbOTA5ZYU2Lk41CLItzQc5+brhcdozo4VJ1k2nue50GRw1Ve
JsVXdJbSZyvA+th6Mrw6qFS8jT/HF1f4xV3L93aBgFIj/0j1L2x2qsuR+TRcRgNjzqdxtsy9oen0
yxA6ibmzPiC/irbrNyrHnWH3EuAQriX5/YAOp5p4cLbn8jPlnVWkEDeYvX1VsoKcT34s11i84pmK
2Qh4lpGhQPBn1sDr+eG6IdEPH5pmidWYtYp2e1+6P+MdmdXInsAmrhakcgE8iQelUos84DJdsB1H
DZwWWNPbDveXnaIsinjYC3xLq0PJLe2h+XRxueJ/xdzPJNm0FQsXt6sYaCjrIpr1qqbje6Oop+LF
uoe81uq7SmM9aTwmUgi8dFBFFDbENRWGbAnYIWPRZBhdPEy5e3Alb/LGxLXu98X2tpmuSdp4iAq4
u13RLdNfpmAyb6rdzTtVMexyTNCpPphfjeYSpr10mx7i/H4KITXPJjoXItFvjRgcjyX9QjdStoQN
UTlh0g7n8ooiegzZIsB6BaVtO9ORbZPlx4trCEpmxwFGaZ5uiicayXbGjCMpseN1EWT0QqBj34ZW
ubmAc43NRyRREJY6Tgv/GJnYLeBtAxUI+smaIWIx+YjQq/Vt7Zd9nNooQyqeHeACnPKJxK/uB6k/
SL/7b1YXcdrQyIwWrZmNyzeYdhL4EKFh7fXEH8vG1UqYXhZPgjZ7hjpwPjLUM76Or0UMGJmLEC0V
1O3yP/cIYqOumaL8jzzbfsVMqBCdbRnbJ+u+34EkKnOW3shzx9PT7uDY/SFdv2mCriO6h0Hs8kU/
AjQ4ZJSRKw/U7ntMpDI14Q+92PfvJJpTa74XnjZcKTqwqJRWwipPOV9IYAQS9ThuBTQYfLmZHDKO
op+5DYLIo2xWA1BFJi1Ofql/2/i3BTmrg8Gcs26NW4S2hhzs9e2kCWTn7ZxEQagwI34peAvQG6Y5
sGmbubKAlldc8Zm3Z3k45gh/zVmCFvwvIxNJ3hLE2R4lB9kAVcJJ04yC23/bCnazpJr3XzeLAPRU
NE+hWojIBmRfW6RSAu9a3jDkDJohY3hLXBwpRfQApp754/PaBKibDcZASBycz0i6RRGOmgv7Qsgq
Ex1wwo+RpMIzA/urfTzMdVfSYmO4YLSuOhfSx0ytN8X7RjnA+MMqdl1w+HBaP5MUE2l3FKSKX9+k
/XmW0U1JrKDVWnEKncaIMDgjUiBKzr1Z1tDQI5zw8fP9YmmChXzEoZj//PXIyWhU6kyKg0DmB1N+
GKOwz9xXHohclpV4IeGA2mv0jPuYX/2mu9evzAqdZBCLHhftGmJq2UTThQW1jGBUXUOBuwyO9hBn
OOQ56Bt26rBmJJ7V2pF4xk0gL0pKZC+WhEhoVoDSu+T+B7i4n4g0xPldTm7jrvVmGO9/zgkFNYxx
U9d5aYWUxWmzX7H0VkbWwo/ZOdiYvdRTlxDUkabQ10oL3zI0NtjPNsO+qEH6DOVtBDor6Ockd/it
A+R0EuHmKJC1gfYSYexE6jz/cra7EvDC43q/4f6SsAdNIFhJiOWOWdllhI6kyGwl6O9lwIlVyPKU
AcUitviui4Z3W5xM7FLd2ItGn2rFR8qPjL445xSSnwq0ZaiaFmPkYGMpEJbAP9QusVWsGGUlISDR
frz8KCElQ6XniQbGnvtvv4L02HiliTeoE9aiIK9AUc8xd+IaR70rqNB9Ch7wOzYsYb8oO8YxpIJ9
X6BXT4/AGzVfDc0+yqDL5T+koNon7tYECQPjBk8CaYS5lWl1tyFhhFwu1+/jlTDmdhHtGQXwud6h
hTmPSjgFZz/vpRJDkAUzRGZUHGvS3EjIoNYyABXBH1jCuXYFAbAHuvJRNeLko5sZHsGnqEOE6vA3
ATyZC+t1zoNjyWkJSIpkr11DCwdr7NoYAa+hRTZHNighPxEog7q/QBStHSnzaS+rM1ivuM4n+YPB
bpt28MPELKssxjINl/CceQdyL2H6tJG8qHJPe1Aov5QIfmGUYw9zi5A3Y7Rmh5qukRIJQlMe2iAm
SVic7cgrdkT35kI0tde3gPp8+zbVT8rTbG1H+2UqCJI46bkLsi3wbY92LRDt04Efm7vqptQiSHvz
hFOuGwbEuOitXpunS9ZfibpSx0S7+YeZ4JhPE6EZNLW0qTTlS9i3TeliwNNKG5nPa08Mi3vfu59v
rCQEAu9vv136c+i6OqHA0a3ap9hUz4ai3Q2Pnr9FGw5GbDJnC92/OBKsIhXfY76uFcsvuFxgQu75
G7eTFtsMLLrZbDESAwErCIT3gCPUq/Xhm+yg5tdrbs1CtDU8QuZbMQANlPPoMyO8/Asz8jMXNiP2
k9vHhY8cCd898fWlBKTPwv9UpY6N00ScrCUZmj8cRh2XUYF9wGfV8r4iiN5b+s+v+FYeNQodWu67
oSFssg2o72ZwjQww2hHo6ltHNPM0afMtTTt6iWmvGPxEeBt3jb5NeoMxvLGLImHjB2bkcM1v4wQ8
qUujptCgyb6x5/9/6q1hRTuxlhI24jf0krKyUuci8dZGD/BXztzqwS6sG4iW6l6NspGgGGouYpRt
7F4LgXFbk8LEGml/V7diNkFpdhnR3MJp8PfHkgPyodprJAkBylpDdtT0twval+nuhs8WLnfI6cuU
+2Gg9h9VDYjxK+N0x09fBYZxUMK52dU0UvBZ5BLFxhddrFA0UMddaxW7WuYzqvg15e2NOS7nOnAV
vh968+2YDtODld6snVTLUtc79QumC/v0kcMAqln629LRevMlG1gOsfkO8lGeZ/2hru4h6Vx9IX8n
vkn9GXxcZoQAwSmx0ZQh9bdYqgJyi7SqC9fx/JMpSXNyLJl/uQPIbCDh+MWi/g9MidVU8vFkncAW
KvWIMg8W8QJNO+SjAeBDkdCjZ7o2Z1Gy/U4EErBdG7NSr2mKIDCVMldqlk4iVWviF6Yp7OrOqw3C
wKasTfKnGjFgINbKJjWGZRhTJWzS9dJRgRPQi3puaMGNZQEaX/IrGZ6/gFYPjzzQU/a/CCm+ORAP
UrkScE5kxNseyZ560Yjvq4AzC4TfN0+u06LcjJ1TE9ewetAP63oTLV7UGae5WNJGtYjFSYxw3Lz+
LJNRY/AkqqdJWDIbxLaCMdoNVApiXhuWANjaiLY2O7u4W6pxAi7dzp856yDNKHLSkhcl1nyg4YoQ
xkqHBhZwDlRJt+Hf90c2VzhBhM3P9YUIpuW0rdAV9zKb70gq6AMXZ5f5QPwbm6zuUBSKRDTn+xRo
vH32yUmwiqtylFouLIU+I3ge5sbvM9Nx9xcq1RD8opJTyF6NDbauJ42oYPk7xQ3TaRjXQTBX4Mg7
HS+bkx6yjwlK6lNlQF9TXd/iBNFHUvuZco3eFOcWrMZ1ghmDyhv6KSpJIpDmODWv79bZ36FvLrhA
AfMFWO/vnxiy95iH/xdeJ6vGdCDTCh3j5YAE+F1MKePfygNWR8hf9HratUnBo1xIMzXluqOfwD1u
CbusaaBjEOzeF3kNBkYlGZT7qGH7fXICThmb7aUiQFgcNwk8wcqLS8rEGfmQNE3lZTAh89+4lTuE
r2BT2Lnd1jKqkdpFTyiWzuqKckLDa8yPWp4tkwQFIrxVnSepLxYbPnEjXEBjdIyc1y+BQNkxWaW6
dTKjDoNj8urMcN3xXWLrEWdfJ83K6La8G5hvXETibx1qVxoLG/LZtE1oJrfHqtMIKl+2TN0XmSy3
BiWiUPwFJH9KULhNg8owwR02U51N6mq9NCkHHETXivi8OVIM1vt9t67wxoWmN7/IBmz+cxFHAnFw
whleA+OfswJ97u8LC8PsoD7IXm/zWsY6O7EF8wgvRIh54DRGblcnrFTxuGOrpfdCGun/YBK0QLby
WzrcXxvoWm6J4Fa2jwSoRmmLjWjgvhhr2RuFEaggDakdf7nNPCrbOkO1a1h4CDMGTxOSGueql2Nl
IaK0vgFnMRNyK1FDAKBevoeFZl8kdZvdWEZjM52a2MNd/bWSoC0nRNLFqHMMoQ6XUSliX2eyiIIK
kvFYpF7F6zKCQx+Bd8UG1QGeDOTQ9+uhOMwHqS9/UTDxWBW2tdzKlWAspV128zSZ4zG9WFuePPXO
2UeQ8zX/Ok8fuQtgCYedn2QmbGHcZ4Y3NyuXPC1OQKPEMBeeVDJV/iWKHzfHZaa1T5hDgh2XnYP9
rNPWDVt9UDFKl4nzedv1jM1RzIqTYVz/GdKq8qsFWcHbRGR1R8X7WE9g4S9Fd7HZXYKHgwLNgbiS
tr2Uh2HXsm60wrvF33oKOcB/pAzmWJJK2NhFsTTvASuWz+Qs+Yx09la0+rwao68yX8RdW0mBJemz
OUQXzaqr/TP3lbzrfM9MjksXyDMAjfgbAHfmCJ7kJT7cl9l+Ma1HZRuoaLlW99+cV4nNT59Sht/u
VXA3alHxnt1gsIrkuVoWqY/KwOK4edklzH9BKYMatugA0k+FnvcK4dYxWu5c14euwrHI9SZ/24UC
/edEcZUz6z887JDlcW12fuYMhAXihIxA5yGETr9oiEpvzhY6MBIIpoacVhV5xRN2ipPb8eIwnK8l
LGJHOMNdg9EmGRsUfMdtoEdm3lgdcOagNUvYcZXS4x+IIRnwZptoFj4GtSLHL2bIbuuru5fZWZ2+
kXRPBQZg2ZjJXyizpk/hVZ8Uc+ydPCqFrNSBOxswm95o2v5JuLlntK9Pv9JNPT09ArkoyeVSJd33
PudxJOHYd0e1xgnaT7gsfWylIudNUr4zy0364x4bw9qKWK3l2QNWAos6RM4WjMTRnSidTESuSQt9
9b9wOMT1YYH86gAZMEyjYu6SWWyVbHrMZxeanAOcvWGxfX1GtZuwirVPlxlLNPFkHdyeGhUrOMrN
2L7XbXfELdfwAmSDQiKFqMQzr3AEIMAswXpvo/tEP75fjvLVVHco0BY0ta2oNuWZut2fyeniyTHS
4DNI7d6yHMBY3ORmVj3GTzq8NVswl+LGGqGQ6eGtb342GGjAAndTbP87vEL2iGPM2LT9cDYFDEAT
yYp6WfAz18/WbsyB5Xot7qZ6hMaYlpH2xnytiorCmSE8jrVhz2wKvNte1JV1n+YG8UFQiD5/NApd
lapsXsWXDpCsIImLpXkvjnqLhGyMkSezs+EDoQo1mWwLAmpI/1ShvpxDIGhqQWVmvxw3FY4LUldk
ZNQ0/O0BCiAEtIOoxLFZK0kWCsQ/mSUHDH1WyEpWsJTVmjJdcZi6TC4btp0uyqogHuaq+dNV1HjY
YUQlAyVGq691BncFIrJd5yQ9ferH1d6PTScajppC58ZUv5IAtT+02Bok7UhyRMT6kctJ0I+ufYrj
edxByusO87R4si87yLoGD7Z/W5toP7R5QEorbQrEq4rYecs3iEUP/6KKLzKLbbwmXjudHCtYUUQr
1EQMW3ytQL0fhxEtQrimzrqESJtBAA4K0PddDIxD/Hq4o+D2ruvR7VE0MeYItHRe7cbM8Up8AMsH
ZmHtWuBQyvsG0Z+tqpsWc8odfLqlcq66ud/NVq8htqqK9shJ6RkCkhiqzmzeQeSv9GA85hwGkxhO
EECzb5PTkIYbs0t0z6f6IAmL6ecBC5IBT3Xd8fiowvQ/F56uOITRp2XCoa5p1s2xSPK1Rz/JQAhX
9o5U58HpMRNNXySxHBaeWZuPMPYwfboUB+1zH57tv5iquh1MYer+p60Ze5+cMNwETkLRFbrYkJkv
WHGsOKYk+tD5ALgRuo9X8sP0HRDjGo+99YoVOHrCX5Og/K+CsSl7yzAMHNtBSUoM5+SpaocL/ymS
baoTOtT1k50HX2q52M6AdOipKvHuNz+y7idNRJMq3zQdDO04vPY87n7y1etpggpHQVctlqeE+na3
6DcAk8EODrxIcEz2/SDGAtADfJ5oMBGnHGjKYALYC4tSkWpJmqSSwyOlF2yRDyOwTH7hxE53W4wa
WJyom+40JynE7zcTGMQJPRpxwix/7icXBamKmQ/Uv/ai/L2jLooeqnfkCBvIH+/XTR2Sem3Ip2Yv
mF8osspk+vdFZKedRisKyl9djhKZiC/M/+3k5VpEWiSwCiLjaViRyWT/TSVSMKQO6osOBlgeb/mG
doXJg9NZLfVNPKAXynlYYP03TdlSQ9Q6oH4Wai18/qrACKPr7UfDYtv1Hc+XhHcOIWnPMjkE/exa
1iTAm5oUWJBTpGTDxIg375tnNJmUy67U70Xn4gXI9rROBMfTv770xvKJYvJ8ZWBzF+IBvrnOikiS
lyjQHE/8lNa+I20l4iDvEMjbSuJUM03JypGv0Fx9/vL5TT12DNcfuizeuvwfPcdQc10JLHf76/gW
KvVxM2WQSeEGU8uZi5iUm0h1v3puOFHwgbWG9fiQDcPDKXHD5xLNjQaSZ1ljd1JKi7mW3Du5UHXi
iCjlm7H3BqIL/iqUtPirpWV0C9pEmQS8I0wr45fTi2QynmLeZvENmGGYVAR3wtB6QyVVfhlhYpeI
ck1AXKYSUf4/zm07LEYkgIsZBp7ESOpMhp4f7s5ZF2WeYdJOZyhgSF+1HNctQrNqgjWugUyVoV4I
suskkFU6V4SKfHASzoWuM3uFh9Pjf1lDc9NmdxP9AmUvKLP/CKcKr61Vo46CORQXGaWVw1/DoZ/f
0Fc42BmKANn8TNEtBMaOixUGhlxjY4PClgoPCiHAx6tUJeMhYsBINmEiRyBr+woqPOO3BTc8VPk+
u7L3JZ4Ymn5BgjgJ1WTNt5dBmse2OPHPCw/miQDnWdRpdk0FizLum7TXpnBxnTJKhx7d+QZbVurJ
ULjJ3w6Ces1eVeCb632dnYGxlmoAW7S4sHxdFmKwr0ZYlkWIYAnbrtwLDl6tobRnwNQmIXYbS+Zk
IxmHxQz7nB5E6CTDLtw26eguKp2y04Z+wEOESkUcJim/j/YlTsRp99sbdE3dbgTZN89i2MB9IhUk
0b4PIFpqmlTF07o/LjmKODpujd7+m7wABnC/qBxlggklhRTSKJEEC+6LuQh0VdnCP6L3mHaYR5xU
TuA59XJ6cdApz2WTLXROIuKPwJtPLvPAMzvvMtlXBrLnRzo0/OQFzWqRpJR8F3i7uMlJnmJtsahP
7r3C+75UlCdOervgevIf+s1UPcIPZyxQpURmcXhsgQ1VwsThGdtczbvaPXR+hz2y1R22v8woLSI8
GjbcdaS4TS6RQXA4mCf99ZU7C4KxRjYgmdceygVrM4gNED9lciDcV9jxMp8N4gBLBjzaQ/jywaKz
YRbC626VfpHrA406+Z6ka+GIsSMNJ30lqWhgruagANVRWKeFL/8TbiyGck7WXB9jmYZAjNiQpaYD
tNYhBMSwD3BRvCYPfKtYEWmYY+QCGkLYXLT8c/BujG5Sx9sAlCKzZdWQqL4OcYuIrdxN9XF5+n3H
Z0VS0HVhscWpbZKXlOHPXHnbVzubmLeUxAlUqvR3WarWDDhRba/nKJIMM1OlY45K7EGc29gOl7iK
kcdzfXpX3BrxPfkOGrA9TduQa5bd0xWk4y1scw/lIRpTyFmyslG+Gos3KGOivFPrCvFTmcGMRPL2
9YV75h+fk0xT2JPNJQ+aZfeXtKCnJXe6bqC8ey0VOuye+6mK0JSKpHO1UwRe4y6QodGtxd1pKtUF
xMqjv6UmPQZop4Jfebe+Nvg4/Uex/RAqYuqphrSlRZY/wFl7q9hPvmnyAsAb2+ONJnSitGdBLeur
caTrXrsfDSQ/HNMF7aBHTicmmZ3ICwozHK7OZqnyKoNaMcffN3kgmCdA4p+KCnLozmsIbbC5Sw/W
4WAEspvwe5mAmglCLkwOo5vhxRxQmg5XPw9tuiid2xjWr7CxbvBLtzihPFbHPgDqiiTLITyRbViQ
KZriuC3M6r8DIPUbCUczHdN/8wEGco43bqPfwdYIhqbiKLpIqPe1S/qjijbOqudPcyMQBTFjoRX5
KfIEgWs05Cy+97zwc/YdNJ03luXbXZNhqHlPZIOvmIFJiEc4dX9slp6vodOVWVFQhX3a97FOqvSn
tQC2tc/kllbrFL+70Fmv76r7MJ4K9fOqER5VGWClDV5/c4MVJcegM740GzzmbYsPsDpYLll5j2Z5
AJq+z2HzI64Qyh574HbLrdkPxAUttGuIfz7Wi9XBNJsZmnCVPDxddTQ6qoqwR5xRvljpys1GyeU3
Vqsi8+rNQk6P4K7xsTuNy8AWsQiHS2gmuQnwvc5CvcauuTTVqCF2F0AUzlKN+bebSXE4/18tL+Gs
w/UTTkTSltsRQCWBtYL/DrNdaSY23e22oJjNu0KQ5jJrhyx4+2uu2dU8xY938IFP8E6/Lb4khm34
X2qkjznYFiSdUbTli2LWNSLegB5rIUAB1fImOT7E58Ew0SU7Ve1smr0ShW16uazRO/o5PCa8Inwa
O377eWf4Qc3AiZfFAbqc+QwIK5wtGNNYDBFyAXPMsw6vCzXxIW0U5LZYksMTgNnkK6ui7oGWigIi
Rh34fnXPogoSjWnQ9aYnQOlBbggmizl2MKGMoNYN2RWXyuroxIg2FUWQCCeuiu2DMQYAn7h5o4GV
jfYI/aVCduNaeV2TNiZAjC1gdYSvdbOQK8eSDtl8Ca8rm8IXzt11UyRru7d6PkLjRDVLUBCUx0or
vRvkaFs8rNci2H2UIP3MkckkGpi9+tRUdvItVyQMtuc5fq8xKu8wHNIzakJZ9PRzBzWcYztx+tGk
DcgY3L1WdyYW39Tgm2tROgxcI2/FWNTkbFA/AbwEeQtOXcTFrLJZIKKnjmh4hZOApQZBV5/hmVpD
XGEwPXBK16q6P+D948VrQ5uQRRt03qoMUTH10PBYN5Eagl3u53+jqjlq7iXJ4jYI+R2mfAqO57Gs
Qqq3INCGLxA8/P1iOIj8QswIcZuFG1iIgEt/FJECRFFdkp37prfz9UVxwGVJWcZXhegP8ifjp9wU
Ob05xYC30pSFwcO8mqi1RJdFs++esGLerDbiA12TlHYWjVqsujnSJ4dDIqu5Rk0aCPtpgNkXsLgM
kU2rzk4a5HDTZ8vqlGLYk0Mp26PVsOHTYk8HWkK7aTgZgQ4SyEzD822CAla/566zybjCjnvkd2xA
0Mh+o5qT6m1reDCgeJpLNxsbEnTmNMcnh/7bHZ2yBAQg6fQT9ZJlmkXznK1MLBHkxqJDImMkZ9cc
GW0qWoxjPhWqMc9YsKGTNELbfRsqaGURCtT0EMASfpG35trRgI5Ar/kDPRxtP7CFegCDJaAGeqbN
az1qKQsczIq5vP4jexLQ7B6IEP5E7uiPXt8k+XdwUm3nIhHTJzItjQFW8ep0mRQHTVnysbuy8qH0
3lZX5f+y89mfF2YJjPjDqHtSEsZWb7Vhqauba366580AEm7BUFYCQPs9laRiK38gKJAMcUOPwkg2
L+97W2cqW2QO6exGop06lyqxvU8euH7aXoyTWKJ98m7LwEqvgUwOht/MV4tw0O5vcVwxkJ81+G29
j9rGDlVt9n8V5xhyoDvyRBLP4kxn2qVsP7nBu65mTcv0QUYpVw9PfeeXymu9SgqunaytQluziYtW
XJWI+gyeXcGZtwOWiKDffg3lP6yO+JxIhGVj9YJ9JRj9/pQ/idNqpa8D7Z0vJ+uq0fiN2y89jS3M
BKqC64sf74IeqLhqh4cE4q4ehh2QjQ7uP3qbmBxorkTrp2ERZyJhGxcu6PBdmVGqHKT88rrNGP5k
xbcIUG1LZdghk7Av6Y/9ngq+Qg0cEy5r88PeCm+XCSJb7E7l/UlWOvmR5GuDqvB/L9iohpsM36f4
5H/w01YD5/JRcVkWt9Z5nNWXKyROC2JhrFE8RN9X1k8QWcRRPiJBUWpls7cuMZiu4ZVtEwAbgZEt
PXUXLE2TEF3/Pzy9JF50wPAcnEQbxVdOiHxAi0FiSRbNbUMNE6MDNM7m5FaFSfJWuJ2Z04Ijte52
y9rwE86EA9DrVifDqvOil64zX3WDyF2LSS43Gq13INOKcZk2cnSovrWIS0lWUBjhD8Hd2Ap59cNz
VD1QA2tJscGAYobMCOA9i1QhJHxgr4mjsujGZ7haxdlAsWi33q2ZxbwZsxUWRyvKd9IeG+2+oF83
XDd7/0QMorTrK4mkJXVX/p4b3zH2cGtQqfaCHnsadgT49eW0RzEyuGOHpr0tSb8VtazGvm2mKTaa
ZQ3k6qrXhtIEwpC+y6nPQefD2R6l/j9jQymB7LK8iK0QiOYIrz/D5yI7J5G0fQ3QZOxpJQ1ySuIL
dICRDYhNhp8w8cPXOqnTgq9PLjjZlJC8yNx3nP+a9rRYA0qDcrlCa+eTUh2335dKh5jo0i4Unk7l
5IIYQIVTFE9Ql01CPv6znJ9Wii3+bQBxNKc1r/EWMRS9crkw/nl8WZvbVDVNwRhB96DIozNyUZF1
zb8J+tMmO4T2h71IJX/ehgr0uGPVWlfLhZu3q1VkLaEAxmckqQw3zS4nOnfl3mAL6Y8RU8Iet1i1
kkqBhBoa77nZevp4EdZhSU2gCJV2SH5Akm3AhIVOYT1EcHVkh9nU3wF+4UCliy7PsvS7+QLmMG7h
loRUFx8QJYNe0iuXShRA87gdD6cMSdacPsHJ8txgZ3K2px9DygHY+lHhPgjX16WAeO9FxAXgzPBD
ClxYZ7ddeYEegMtnLxDG2VsN1O2qK/Xa/mLcDicsjiXYzxUh5Q58+7ppFg8dUPFsaVi+fOinCnsS
QGAlBOzwEIXphTALgGoFASJxQyOd3zzI61YDTrnGag1/ipSKZfuO6BnYwDbDiGIvMEla3p+p9wis
4H/Wn+OaTsA7efbj7upliWbJHce4YmLqRRW+Byi2VzKX+OK+YQFYnACI1bLPvu7fXqE0IO6fFB/W
420smMtvhhZUfWfwYNA7Ppb2BfEgeDgCusESHYkcgJUeGfmZeEhjBdaJ1Gsl0iG0A4kwOjP9jeQO
Ja1cLVKE40VRNi3iBBWYtSl41Yy0F4oP4dt4BTJ5/Sd4WCAFWOqL4aL3Q7xZkLk9wCtdFDX/0a1l
31m5SQyboMv3F1o/7q/ZYl0rmBwxJzWNlk5YLkMJtqB8dYdeBRsCA7doPEKzc5CrMRkeVrl/VFu+
AAFLk3oG4r0/f1aPVfmGNEalnljo9t7126NyP6AuwgsZx/msP9b1/V5djmbwVgfoHpcURmtdqHCM
htR5jNTSy96xGhmMJR74Q2OysG0SUXDlsYP3TbcytSHaeCwidNkbecoZehib0+Le4u0R6UwkLoQn
t5ZerY4z7/Y48l5zg69YPZs7qEBa9rZmFblo5FO21uPJjnQmf3MBEB4U6Mx4bUOVAQsLvlWCveWt
uS4d5blzaWh53hY0l+O3tdB23WoilxGUvRLg+z8/ptKk7vNmcuK8q8w7jOS4soMdB64Ys0rUlUQU
tOs2D9t4ueOmx5bGI/zJWscG7BAEUEWDTHInieJIsFbRK4StVPCQ2zDjOo0diLiIU1vi62akzi9l
DiFIg9EE2bktCcFL7dVX/wUWXMwT1Jy26BoY9kr2zcfzQxLwDdGGJ5MTuUY2Z7/S5kLFoJx4OFtp
YEPT/nzeXKN2kv99yEf/QMcfq5PJUfkQtK0gH2TUrBbtH4qs44qe35y7McNn153mwE7fLhcyvvXK
63KBAfsAxjMuAjJVxvPS66rhCUKZLJxVoGBKOHc+b+EWzMoZBGDxkWPFkHlzdE4RZuUqIGLRx3Se
0ccTg0MwsJ40+BKfOFGMGanymRUHXaQXuhspAJm9O0XDT/Y2iwWSL2dSYjDeg9Pf6WGbIZSJ5Hac
EZUTkqlVaNF4+swUykBIx3u8DVnwvtIrkgh474BhgvXImB5ocwJ3gStVlMwCljsphtsqWCZ21piO
jiMcoTd9Vw5cMiWTJPeHvTPLnxF7QjSNJq+UmRl1eT/pS9O5SVNihAgwHW6oILmbt2RddpaE7fLE
kwP6srHO1aS5oQ1YExdeYpLqgJTCj7Ah/SQHw6kOIdTIjsPY35WQTy++BbNkCLl1eZwwwnF8Wluz
BxjAQ1IAqsP+cEmQZ7YGVVcxT7GtrF6f9wKOsKJNClNVp+rVgE1ZvCaR1qd5F1dLSHEsKjKd69J9
sbebiVyEhmmSneQQ0RKVQb8UA7yaqiCPDPNUSXRk19fjQDY8B/Irm4d8H17IiX7xRKDE14R7e9Ss
AauRl85LkuJWrNT3n42vrDXD0U9qOK6k8SjIvuKRG3saTVwRn58/UOMyH/1N7Dl6543oTOUSejky
RyUdQ3o3IRrcG1kvAOUqcxdmcsIFZ8KSBPkacY/ox/mmg5qfNt40llGELc9BbJvGWfjN0MNPtUa5
SzSEJo3kFC1MG/hw0UsNaoJWxf9qbBrxT2/A/ECmKkiJbY+ZV9ciIDIChaiFmL36q7Y8xbir/JJV
PD9iqclPqSZr2S3C1XpuzSEZrHjzEvefc79EF7w6ymZkeC2kxCL4Fqrum5Hif/UFGCN947RdUtlb
YKjgkSiar5JyL9iWYpHhAENvwjTHlUcMyGPmDYF1Idt1zDVJaESIgnzGxyujzLLTG7mQcA2TkabG
5Ta7mWmkhdCSBE4iERzEDGyVnqKXCPMpUr8k5nTlHQj5TZKF96sJQh3Htwfg50T9bEFkYmgCIfmu
WYq9hoi7P3lEykuWhRj1fUhOlsDzDeeatWNT6AKw6leapyeSwJ3EAYTIKwFyDhpeiYbjAFXOs15a
CNI4Sq4A1xq//+pB/7rQirAL/yYDOHj3lz2uDBC0yrBY8a4M5KIpRx/XiUGpW2kGPbleNgw1OQ7E
xro97SAZleqpwM2yPb6qdO++8dqbcPn5KHFH0yYopkZa7oNYlhOBBRkBh5DyUQFj4CmAkvSFGEvR
6CV1B1pA+6Yo3tJGFVXo3xXJVG4Nw1EmuRbI9/Hd1Uc7w7C9wIqEmTcnLMfE6X8jT3tLSsuMmA0P
BH4WzoFxX14AU8GFdcPtppZayh8tfvtP05/A4KvsyhzGIRunlK05MO7JeJpPTvpP+qZLx0rkIHjH
VznYoPnzlO7HLlUMDr6Qt/0aI8k4GAnZ01qPqvx6s/kG/CalgzQgCTIyDXDdKytLs5ZtddN8xQK2
xFDPWKZBLgdSWLkihKZCmrX+sHtMLtUh/EyATzsxKyw1a22zZiHBCydxc2AolYiSGTJ9joF6+jwM
B907WvN9P3U+CJtIkfKrbh26Nz+9D9T4f6FKO4n0ZmaRRgJui3UmvtswgpxnUaDlCNVWmqGPAiNG
bdNNRsz7gunjOMLScb7W/zg1oL6AZDJ3ve3RFi+n4MGaU5aG1Qel36jhk6DWlnl4c+Sam7fr/5tR
z3Wwjlw5pWOlFjgRlOjBC3VhitnGuvuASYUiqAx69G9c0PwztWQTs9/1IMi7Q2fKlK0Q1GODY+zO
CgZYZBSJ057+Jiwbs7JAlOonRP0DsZ/l28SPNLkdCOftO7FqEhaEmEHJfUkh2MY4oAHFwUc9hIFs
0EY+tiKerydhYZulcb2OYfWwmEb+P4yw4ErFgKtxVJ5likVlP6SSl2r71R5EAy5WL8vOxdTbqs5O
N4vxIJ8H7uJZ5d1CI4U9jVs6doi66kZpWJ4eYL1DCZhM1wX+VfILwuIMEzoFiGOUYCaySqw6BH1O
86Dv9ViFKdu5G15L8ViPxDPCAtt2vc8qbaFh+IzM9tg+h6QMIwA7661PKHeXY3XN3v7tqQc+elfr
fqiSQ+0NyHI7TBN1L+3oxN8PriJwl1446z9Kozu/0t8qer4re3t6ofgErSFNNOiDGsgNrTohCqcN
0uRpRGORWcVDl1TRX+LDvs9YOe0kyUBosVCp5oSqc48F7Z48CYsDRghir+j5WxFOywRaTL9U+xij
TxOX31LIsJpV5pfGAklHxXYUjY/NX1iMABpR2hkX0C0XujfWwZvedSd7wmMuzsf0q2hdHKevULEn
eIH7iKPhO+Y3GD7v87vfZubMBsO81Z+VggeCmfMToZzmv0safLlSl0wruSd1QXAh8PcZUh7/fzo0
9hInW7WqRER7iUvOZiwDHRM7oI94f4TzcF61lSroyxMMub9mpciA7awh6FlAzY90d+mC5X4gtDvL
gwmCPgaQsfhvXK1aOr9Kx8q0X74R+V5t0GtJ8+5EAFtryyD0wIWjq2gfyz0TgT2MaSbTS5GxlKKg
Xpx/M44Vs6SHL7s/KrGiy3wes26yfDDAp0XcGzurFqFZuI0bpAFlixqLsC72QoFzwALn3s60B+77
hkPyGrTiRog09z9vc99EPYdEyHK02OqCmGlA+kt+uXgm/5ox0tGzOrF00i9Qr2vcu6dNjA2BCPE5
yoiS2VZVaZzdB30+FvUoeIP+1SuSi2x/hVzfBZTqmuh72Q7S1Ok5FIUHRbNvWvluiKBrKNL6DR9y
F8LxXgIdQaLkfJQrMdv+YCavmMBO+/UzWUSIpkUAs3pjkSSoZRwqzwxnfypxKz+tTosgwamgy3aG
+MmYdXH5LcrD9bYNZ88SBoqPGJhVxDMceJx9uF9NgFKUnqNfesuVlIvky4eF+rEGNUdBzO22m9RV
dvzMOyPqg31j/YktOdLGVcwsnoMn+L/PHXRpqJalEpcaXKKhYDWEPLbucqRbL5TiHk9ErzR/A4b1
bHyYYt/N0wM/0+yHArc6MzW7u0RLItUm7wLCCrzIxnnma9WT+z1m4/HfNTnK00U1VAZUsPjYkzJe
VInmIX3IXQYPjwEz6JWKeCsRXH3WCqhD0SukrIqvPYsDS27MsalOWkE8d2Jz+0MJfBWihjkhRnVW
lylfxF2O8qLlQRvQI5OjQlzy5Uv29vM5KvnrXKTfeBvlGHiZAtXSNAlsB0+13LL9KwRIe5VPqAE+
Ge+vQt/Xf0k2o6lI4aBcKfaQHsGwL+Bo4LINr+CV2dDmX0wLMqpBaxt4fbDAD9ndHqnZoV5vcmDS
dBNW6hBRwbqIn/dD5OpIY/slgg/K4zLGgtxtcdB8CZVQes3ZtyIWK9R0XQwExDTMQGTVuDtyrJ2+
9RTgVob6tsSbNhHMLMa6cJaQ/2xhvXl+W/dWOTX+aPLpWdSshiscXohDnWJmVezq6z8SEZ9EaYMC
0YBCVKczLdQLMnut2yWBh5j77uVaJIxzcEL/7sIQhctZTmzCpm5GZLlS+Jnex5l+qrisL8xcfhHS
E5KNXzDVL0kIwNIf12rbIXnB+22gkFiQVX3SIaiH30+deggN24D676ELi5Ox5agu1orAPdS6sM2V
RnLZ46IZDuTda/h8yMkQkMQNJ+AiVJw/DzD8I76OjkNbLe/vugrNWeY7eYDDIgGX4rv+t9VJveL1
9UTypbuxb89gqAni2vfk802IbzaaMo+/paAD+544rUazQ5taHDjpOdeqFC0HL4WOf2KVG4JqnrqP
vZdDojCDGXH3bNE1hITmDFk5YA08xVPxIHqO0lwa8pvo6/FUKK6PEOyiDBYKTH/89FNk9yfotBUl
1mwmd5cT6VpOpkMo6gVrT3aYfvAYD8FagU2ZgKbidviz84ayGG9Cdd+GqtMubJFPnIfU0J5espyV
J7ApYCPSBkEhsgOPaf/Wnwi0QjxPvb9Z18JicVd2LUXyVIvYmzurty7xDm72qmPsz1x168HNBowt
6ZPBfkTMe+dfJW6QWufKNPHiH6WLIBrCJu6ge1j0LBZPjSbCzPBHbIxShR4j1LabrOGRlQ1OWhJ5
/5waWxhFIGmaVGJdFU4LaAdob0yd1e2cKQiCYaC6nOqL/kiMqN9O7eEsdDo95o81vBpThCR6GKNa
0NMhwxlWZChEcQqkI/OpMcqQPD1Q3Jmj2SN3y+1Pt6WkVR5jFFDpDzIDquyJvb7a50UgPkacqyic
NWZc7+X+QeiTXtyvQgKqinGNvFndcUN5xlujdtbMVBtvuntZHNVphLJDAo+5RHf/hpZ3AHv9eEJq
trFS35U6meRdLnWiYeZdjSlwlZ3X71cqsIR1XVuyySgbe+t7qmvlciO16oQyjpAHjpQz7FwXB9Hk
8P0DlluovOjtervFADUfnd8ITUi6BamFoTKRk2wQXi03MX9dEAOvobtf//23I2Hus/YEv7UXfzsi
t+27rE7KzW/o+Rh8ubhgSbA9c8Sf7bEyFDJbHXiZKyaPv8jdSluL2burYuO+R5PYtazyUWC2y2m2
U9U36wdRKmsJJ+gCAQhQs6vgTdvpo3QEStuVE1xiwanoPQSSGFEZPpNtW9tOZXV34ZkHbsBhEnQQ
hNoiNIW7+iwEL/mBWWApfKlAk+NeDFBpkapR+ZbaR7tQdOb8HKLjNpEQ+LcfHILd4nWlNFZoJ7qz
vYiyaoxzoN9qb2V29yQa81icrfcsiAE66pA+8NSSjkN/zPTvrPubDUSRW0OqIU9IAmWz8QLm2EYT
ODMal/+IVeqNlXmeZG/YSYzcDWgbkENgJ92Y3p0O99ZMin7CM52l7gaYRGFTi2UkXUsBzrOhQMG0
E06UNFFxR0mJ2a3p55LTAbyjZq7sXnbe0Agxy9uVM3OMoCFkn22Z6uUj6NNikhQDeJX7Y+NyZKwy
1c4WV4BRUK4wI68nU/bNYoMTw/AN9j+7NzOMFUcgOeURu11S1GJ9PMNvsQOj/Xijqze0mDeIWIgc
57lAaX3isASHtYglomYtGvs1kWQmquRKeEVYWfgxLb7pyag9xtGRFzFO9AlOO2W8Yl6h5PlXN3Q4
3Aku4yDhhiIzDyyOKi8wxH2kPKvolx+skU6YV0cZ+7rTpvE+poFEmMuAZdHXgsDOPwKOkJoAVYtL
ZLyGqZRGbfKqjBdRlORwqlU03jCS+CbwWQfTYccbDjIsuoqz6ljGdh3V9lVR1iVNuoEgebYsZCrF
JsHXWmpkA2xEMhyUd1jycAu49pklayLIb+ZbHtDh/BmcT8lLJYHR0BP7fV9Qm7eiYfxjXFO6QRF9
J3/NGPlCXzTKFgXSqTUeavDjiznoFRTPioPqRyvx/bcP0n3nYqw6Ys8JDWcfU+G2+p1FieTxlR1r
n37a4WyGj6YJHpUa2X8VIY6Fr4QkT0PCvRonpuRlcmr4iRVzJlU7cAcdj0NPMWrxs8cwjH84c+XD
2dCd9+w0tK99do5b2YcSJ7IxKCRici7mVLmBWB4ErTpcJRVzRKAaYIZCHbVv/iu0O0MxwJwab45O
BBiVdxNyiFJg1K291Djp7chxL0AbWWC+aWN2D+2Ev5Mj33EZ7JL8ckju4168SvwK9HOhsdy5uMXy
mhQF19cMB10e/Yn+4GrSQp3GYIKp7YKfMsYzWTg5dswUxjc4svOsbJPEqU8O/Dw0zr3gHnSJV29J
oZ33ZjVlyuYLpFxbrnBnShZBm3oRywmTCBAAJOAk3y9xxaBDaKVmD05CXG/1IhpKRz3B2Hyymtq5
0wkD9bdyPf13Abt1Kz/0Udv38A7W9ugSdI05RYk7CC/d1Kl4z4qk2s6yS7mSfM3hpNkCEwdeFC/X
tFT+pWbcZyYjC/X334yYivraNiUHO9nrbjP3gjLISpJvKR1Ibj/qLSSox20Rd6PsAydMBSG9X2kD
OlpW220IGSG4Lm6hN8vrXk6L1SvBb5JxYQp2LeF5f+UIjNXq3Gf2GOVChyUlPR4ZA4g/7XoBksbx
oBVBZ4pLxIPPMJX2rjuQiKtVzEusxG5rEH/8AfHbht/MYyM4SPJFC9NiT5oIKf+LmWt+9P/KA8pL
sn+tCTR3JoZSZVkO7Ed1kSIWY2cpMGLmloBoVuxTNkWscvr+Me7i4nGKB0Ls0M6zj6F8j+ZaZIiC
jDhQJ8o28rmUx90iomHdtyvzerHgMZOpN2DMSbj6egfwdQ6ig3T0vN+uxSdjB1EYSA5OySgHWzHo
dTk0paQi9YbWsEZCf5srqlm+UBkbvXmxhlCdF+RYMSliCacXFOR6p9Q2cmbx1UrWVe0bDaRLgBW3
ZDnvEzusIrj7GDt07B2XweiMXec20UkPnnkFbc4fNAkNTBu60j2N+ffwrgMHvphXydgFDaPyuoMq
GKEhe9PYuLJeh52S6VVYFNeffn9uoQDxO/dNBRFViMRuHaPoNLQLszfZ5reAZY332Xp/5ZraTcGN
llpB/JSBdNYE+lsK76zAQrnYYmajOu9JB32kl1g1EKLKNTK/6n6RTzo9w3jGA9vq1hMkxWDBL+qH
8LAdbFyecCK46EL1Y2MovuoXf3HAQhBgNcjMDZH6+LgV+8xisbCS/kXNCKpCQGwnph++up3X9q+V
y00JEfdCAS3bfxQFOxS8lRCyeED2Y84AbHfD1fxNCSwhx8/NQoCpXZrPSUkBp/7Z4demD2OCwtzn
Dfe/bzbfhNnF7JoHAUwfQz7rR/GNPFAGK2keaDnD96CWwxJxMKmqZg9fSVkkCOTsLs+WN2+WFvtu
9Uk3tJVTKwyJBC7iuaVL+sso5rZQoLwuNoWBpAkyNrXQgjpKb8tPIl9o/+XOw0Ro8qK7mg6m1tGz
Wf2aqK56B4oHK/Bq5Fo7wG2HTj5i5LL0pFgGtDFaxTdXQbcxwHprb4HazmGpCJuMnQZAnXJRUd+x
ZpmHv9lL32jcy21IndBgvJNNxdPwyPDFc799hoPVbxd6hfcNfP2Bai8UIc/kGslxvLprSDLNSbwq
mXeyBYiQhu4y0UKXy+dnDKs1puQIMV72bpOZ5UzYLl2/LpOiS8eQcKkL6OQyj4hNhkmN9LgZRuUi
vk4DvqeNNJzxJ0w2SkDvdpkBgXzLBCfEBqps/z4sgmkGPNFycfKOlW8gQT1pfRaWo1fLMJivFbbv
/jmL8j9ltATBy40e07okHV5QIoma1789zBS7hmIJSqC6ci0ED/iY8ExvgKmZnUgKmprwEDEd6Jtu
a3dIVeyqz1ASvZoE0Oi3pJXFUv0dI3uF2eFijM0QssCyWJYGDJHTIjUhF5PAdor80tSthx9tOiVo
nyAOjYisH7lQ6ogHigr1jiz0Mw10diEE3ZIyc/R+owkje899/oqQRK34uVLCFIAW6OCfgXLPipsT
wvrAuJPEFTHHQM+7iDEDmvtIUsEhh4VgB7WCgcvgh7lwlttQftnOwTHDJyA0e4Bd9Oi94GijcBh9
f59nL1uho6qUaF2PRIv9ezJHlVM44/yKmafiuE5ragz1yzpQ51MCDseBJyISU0p4cHQghwR6h7jF
f/2AnKdE6sYwjPxwBVNU2odqgwhuP5dmXtXf+btFTZn6h00HgmV3hOl8orel+I8zkHLS0+dn779S
of6f8dC+9ndsP1SrRPr1eeDqUSXOI0wGUy2airRb0YKz//21aQQcFxxF2+z1k5dmVHNhQGznFT4H
xX718NpybMUpGg2jPkgT0GU45blthpqdKFrGE7WksVxFJJJiUxo9JuKN5d5MsO6Pbzn7hDAgQmA4
9dI8xaz1Fu7d31kUBKQS5BmScO0hKUL1I8Q8whwqtfTtFnz4f2zmkSLFvdXScarLvard+M5+kJ3p
9gbNkdip2RDyNmg+E1jIx4vyBgLqrBSD8P0ttnfuxR3L8hJ73UQFUoV+Z/u0Ftb+1D6rdTv/X8Jt
agTveIaEn5xBpGPd6SYUCyC5DRwQGq4sk44WGZ7c18myTw6SsnjUxixJSNIc/ThInL2FA3ICwgU5
caoaikxc/UCV4gT/9yPfZTuJHP2WaG3+M5eoIraB5NbuIEE136S6vFZ6lVXvcQThyGnOhdlueuPy
zC1m+bxqC56YNiMOLeKryVwJT1AV1htE3KEqcrgVg1stlQYv7a+x4QCDXRYIZFaQyuRilPfoCjTa
+j09VZr725YV+78QHnzBKVRR/4NC1SP4kykjx0pqV9cpnrFRDqEBzLvPlXTHotP/6Jt6QQ08sGfr
GnSOOgdAWBMpgEKtAFfuz9u9RolYJTLsvljryr8XqxyPH+GjUrvtuUa6APTRnMgA7GyTv0N6EUBm
xQ08NaxybFoMXBKf63iMf14ErNtubKJOw6zTeWAbaGBwWSOeYgFNUKT9HfbGCk/qzEXm6u+aja/B
ErRsnoeXzpSx5LWnviTOFx9I/rHSN9rV+As9zb/CJUDoGgTeqjVWwwucPsF1gx7iHtty40psjphW
4NEeQAUN91cpheackNR8I8ubVX40/b9jwJyJNnmWIu7dcaRwhVENCvWrhGqjO2pKOGdfW3jk7OG6
oW3QLzrpIS3LyL/hk8dkXmDEiNMUUF1ztJuzPXpPNod0bfCVGS6XblPMm9xODiThanquJRQXozQa
T9bY8DQBy4J99rRlRerffvEKXlivaPuIm1m8Dd4y1KTlfNmBM9jUdaCyVooqCLTys5/1P/fiQxlL
HTpFPcNO0WsJsz5jfiYhuvFw0TGlv/+0hOCmaaXpY2zz2hUqeazwaqo7UOJBQ+yR3vvKYEMR+3gN
yvgb7+dI7EulE3JUIOt2xLmi9X+gvvUrPEbH08buIGKPL7MXJgULzDBGwb2zFh75Jl2e8+6URNwv
7SJ2UgvYOjuCSsby9R+1jcY05oM0aIOvlpZ4x0RbuqJVegb8YRnsX+WnPWOqmeCW0i7XNKZPIxBN
kr3pzUWLjy7BwaO8KLloSZuUBrvmniE0DkVO55E6El7EssT1JBHxmUb2xPskPnYBFcN9EpaYxjma
m0erQ2mvuN7VrsT3t96PBYs19YgHjNtHHPAGy/sBg8QfnJQCpUuk1aQFlxftMYjDfqGbQWmGXCb3
xgsJbgLvEi5H43d17GNudKal5YHHQXaZ1Rl73XVrZ6O9xH4lIODNEJgalYzas69ygGnPrpT76d41
OtBVziNB7SCQwvWf6HyTsGb8Wv1UP1VOVisH+cMc8zgLvwFBTlPmBJceFVL1kll0wK+hmss1NLYd
mnHGB/KGgiFVMs7MCXNJvPfKgg8Zy+/OHo1ZeLd99pVLp5bQHcMHRPr1Tm9xyfBDjunrOD5H0R5J
i4dRBTyRz3JNri1fzt9K+NDZR6fo2wW2NRV8eI9e2j8HJPd2kLSPBkRsVymxJaLaMRCY8zhBxkTG
AVTq0LGGBVDrZg0x4Vd3uhZJz0HHehqtkQm8S1K4ZGVj2ZOqg22tj+o54Pelzfsrkw7oDXTVFDjC
E5ALpSO2UCKbx0ujBySsiCjDdGUM/UXychmip6VEcT/KurxEJxrWneeFx4UZw9Sa/1OzhxNbkpJX
VSNINFhOMiF2vUDsev/BeSHaH6Amu5ptUwc0GLG6I50k0GGsHk2/TaKbzq6C46s/9wNSnmgsuUdl
C4tJzRiYWS52hzC311cn6lX24k+dWfJQFHEqZFJU4ISMrMmCLw9tTc/1hUTBMs4bN+oHmaESy3Mc
LR5IiHQRc2EEQ2e4Z5lt8dhg1a1EALHCHje+ypXbn8YZ7uBzLkbD1l/lLWXF6p98gUKwzCWQ3g88
ju0Hjs2CJCTNsiXpsA89jOngLMB9b0pQjmWzhXZ9PxHQxlYzmPGpQL2KDa4CAke/8Wq6WaH9aV22
FMMCFQqMtMgANQkLrGPaqEvFZW0Z7fZwfK+Vf9s/KiXhIyO9nWyII2yuLtNnM6so/bU/yt7UyuJs
AF6r1n83Z3W2dCKMVjv4Yt3bFWATalxIK5CSvLmO82KionKuQxok3tBd1rUzGhpVv8YnUTvEF/qr
EmBHD4oONLYE8R1YAJ1W6PJkvipsIqipClKGBzoieIElPJVIJm9PjSi5ujcJR6AKGANcDWa1a4TT
/cNkv5mHGxk3xrmUffsnr+q71u1gFXBq3gtUD5KGLYtI8nd1EeJLmlyu/SF/kR/2VyKUxGyvRzG/
VQmMf4ExuHcZEWULcUxwpzPYVoi/6VadrnS8eKqVxVw0WXwq8DkkOJklC7HkK2Ov7FfCNP44b4Rq
Pe2Y11WFyXPmc2IP6H6xExtOZPD2B0IWJiS8lyFb1ZpnBo5rqcF+0XjtsEBkwB0pgvrFr3XwDZYf
k4Fs1X7DN11y12o6gZAd3+YWc44gAE2B9DDEh6smNigQHUqOZObdn3dPWkWv9A07MAdj+Wu++P9s
FLH7bHo0wUeA387Gsxn5ppMufBdWDJc/BWqJ4C5lSjcED2TzZic34r/BBPonuDGiW4K0glfZT5i8
QWlDG1L/rZO1izoGQGdVCo82GeZQHJ4WltPm0XWzcQ3VCqD32MaNtizSo4FhSoq4cgym8eayaYNu
GIlImwoess9hwZz1lV26KdQLfJhKJfk26/PYH17zcTE9viW4F9p3nbo65Y/eB/GmIDni2qXiXvGB
wYGYpX8vRSMOq/4Po4XLEKf1T/qrcTfPJLBnCqDOhMRDlzfCJsWtfn71F4ojjjbCRV+aks7WnhUQ
8Kr7PuizjOhSpJu10acgqAp1HFzSDRzpLo+r5hQ9vX51IgU5w0GoR17cIV4KKJXR5qtXaPUoNeaa
S5QUTT+1AZfirNmGL9QexS6whgED17UEoGKHLDz3a2HxEtQXrUkO9pVSNGNiOQVb7TcSeJmcoDLK
pbQMa45RmR26toPJQIEqphu44BMO8dmxKzmTdqpGaqSzklmgZDixy1Dz7hRQd/hsfz9Zv5rSuFv3
mjhGdS82VU34Y9lwHXgXy1+CnN/bnQ3CNs+Z/NqanMw3LjyRPyGNjnC2p5GKdV4X9snO2bhA2r4Q
M8kdTHTFi91HNSIUL4yhnNFF/JriKBkrAB2mSuNBLzcULK+Wm2nD5I3kU5laGwdWFZgh9qydnVaI
MG51GKUMuzgBHWGrIOeMd5squNeIoM1Bf2nV6LTNhpJf+EyPa6ewaRBQWcTfuKoWPWkU3ZPrrEby
1Al7VJT3cHZ81N+BsJsHCYhm+FhR1oPeKMN2v5pR8qZWJH3DDJXY3hb/RxyY693gCVYMWXUZvjce
wwjZ8BYNAMZCRzFfRM1qzWmwekstuEhq/T1eigKeh4iTdV8D8MlTMgbtvfCgoRByT/O3T6S0A6sr
nMxmCRiyBycKNxxz5Cwb6xOZ3LKEsDHbauHRDw4jIryxHiTuB1ufdXgA2bUS5hwPduriu3LbKxw9
83ywscJJJ39BNCELDOgF+WMmazRvw4Sd2OyywgW8m1Fy9YT18MCmzfqz5jzC0ITHE5Tev5by3auY
j1cWSrvOyrIUx9aZZbHmLBXoZFo/ptImQdTUzllYXLmb4iyDustMgO0YwfcyQXsmiy96eSFY0jlr
UGwpi+Zv22A16cQzpTpyN4KxYzI6wDVWgsuSACflCXVG+dtPpEDwmMwe/DdqLs8fmMZiQlqM6jwW
aDveJGlrAWDmkSvEPB9ufkdzLlbsDy72LaFJTZj+BUX4QjSjXtJzrqbCGCj9qSEPwnpekZT6UnFU
tbG/7VyYK0VYIR0WQdgj0xKw8lxqG6sd6UtP+aB1bYHECSsdlBmBakNe56i+yuJ4BD6/UbMtOB7N
1FjpZW3nYcZ+3GVIOA1/7t/ft/FS3PX2Wn3YKRWkiKEsxwEmOifUg8oQns8RDxKLW05oFeS9gDe5
VyfvDuB6CTax08gh8UUBdSsQOYS3qZLyRS0ip+1qvPb15/UWkVUxEJvp15ayTvsKr7uO7Rx1IVn/
/xwYOknXbXRjGGQClLkdhWeeI5gnk/pjFTpwFJQoErU2+VnNi4WgeiOO1MBgh9+0qe2mYBtt1lWd
hY9la2zIbOYbYqXxJ97pZZjyu+sIWB88DqzTMdNAKGkEaBEAtP68w9iIUOZ5pO7v8g5Sfxqp6ycZ
hO2rBZ9ixH+JwaD/G1WR5d06xydKNfrrnYH9SEei+rsjegUZY71b3wuDJ4qnOnkm8SAaiuZi1xnF
/MPWchvbwzvLvYKbyHT1pdmWZY80Svha7WUakrUPB3nfumqNF4tSbYRH7T/dhLiecTlpCJ4lrfwO
QSP3uJ7jeFhUgz0HqbUNn2Oz0K50t0E5uwKwa4o8jUpUWogIc2bvt9Zz5VEd7kgtKcUZ76+3m99l
PLgesjLYrxfAbp1cqu1J6INlywMySVV2x9j5Ff/i5ewsazo/jTgT8EV7xc1Yv19dDUIEolgNYmhW
d3oMmGPP3q4edPoir0X+kZ+9j3pDq7Z6o+ZYPeAbheJx2BfcgVeuHbYHt4R6/vo/7/zmspeqBen/
QSSpHbHUmNyMEtJtywDpGM4ZEhvqizHVvZT1NUo5EHtz4HYzZKVy/DQMWWiS2yitTqmJ6VYfQEyQ
lPsrkNntBHIjkgfZmM3rSmKl+1m5oqZBpZyaXwuDHuaY0Dcj1JOnCoCve0GCFMb/BXMbuSpvcGzi
VCkgl+U4qlVUXb/4XrN+fHlriS+V2rZEspXzHcnuwdvPwkiQdqQxeh8FiJ6MaR6agdawjxceahtt
UaqWKX1GCEhjVpWUZSANMdZReHQKDRrfDh5kgWsqRVTK4ghA84BnVeO5ahGBdyejftJNarzxunqP
X84v0eKfsALCkGOvqviXBfCJJ5+s6D+8yXuzvfnETQHFZJ5gA1n4c9WvkpkmwyfTo3Ha4Y0K2Xfc
MKP19U33AaEjLGcG5E1vxzXYqfidO6OIo2Kf+oE5xggELgogZv47XdK30RA3crQf+/VlPCzytl7k
wz7wzV9m8DkaPBqDb2pvQZ+HytXY++ZYVB9bfniifxgfSmYJZvBoGYs0KKTMErWRWbRvnxbpZpDq
R03x4pizlLYL3ugrmAhDGa8Hzma8hleNwAD1OKxV8P0YuKEWpVzZnpDEUPX5ZVE/CGW1Q6tKnHw7
nCthq13sOcftBTRefmnPF29Ff+lxMIdt8ng1+VQurpBeNotUkpeo2lGQsEGrPmV4j5rU1BcIk51k
DqkB1zA1NI3Qjq15EcfvKlKDK+Cag/4Md3zKmEnO6dG/8MndKBi+BnfwEmWJUoaZM9+JdCzgPQeO
Z++0FtAErsLlKQiypYEFXmoq0jnjDFSALnmRMbR7h7CNKne7iTrDBCEjYgXSuc63N0+LvnO/p0Nt
QdhYPJiaph+6V0W6VoobL22uAe9O+fpDqIPk7vIDthDQxh0nmDtFcgw0U2ucm4nURT7C5Te4c+oA
n+aYQxVWHd8NbEdyuCkHVWIWv6m8xlysEPjKqPXv+8Fx2xEgxesRoB2s4zj2+UtyH4E2YRLsrVqE
jGLDQChcWIoM96eh5x3CFbdCW5NWYiJqjC+DOtCq60zvkrtr8vA1FImuqtrwKRJBf34t7UjUJPsD
9TNZpwWAGGjL4skP9TxZj7Leb4kpp6u/e4RJpzyN2l3yp8LwUpHyOmi6IBWfSz2Ghe/lLnWaRBD3
nhuXG7IIXJeHAhs/zMtSrVE8zkkOqCiaI14EtO09/dA41MfixqTUhJNCMPJaoR8+kfA1kjHYCb0/
helv8BSgpI/xZwf8bTUk1x0ibqDsKqSP1MySUR1ZkauBbpcqOqfK6VAmUF/hZN6VXo8mgWq+o+s0
XrasIiNWIuF+bk4W0K+ny/4vIgqcxPoVJhJhvIuxaeWtPZfO9/2bja066v4/O/0d8xje9UU0NVxJ
DD2K60vj7xUoNNy9HhqUo2GDDAFae22yDhLGdfp1sKB9kJcohctxVzu0CYGkwMxw8Siz9Qi9ynWR
KmMS4nz+R1PfRDMFIQhnHdCVNpHqjlARN8S/Slu89HBxm33bZYkV+vV1/45NYv76/W8YfuWltEBb
ZLVeTmwANyEeQJYN3OwHFqESwqDmRWC/TQIM1aHS1CZPaML33WclTEeWz8jLB8YYCutluHDCcXqq
nsXC5ilSd43tA9PuoaaJJfNU2vkDdlMVzvQNNolaOieu8LJZ4R4Xeg2fF+bNY48/keOQM33R9VUK
JJMsBpEToJjqevE9L3GVOg/pv1uqqLuR4xSvfrsEP700iQUrUdbtqIN8Xn1IfSUrQucKeABJ/WSK
f+Kz/OrZ2sYzKNGWRoIGMBbqlS7fdLPF2d6GDdQ5At+bxLXBxWPyX4UpUKSh6Ji4vru6th66HE5m
8y923E6AfwlYjDfF1Bcz5Qogx8/jlKdzt6BtnDS1lmFA3ucoNErQGa6ZF+uonsExMSUsJLgkA+Nq
G1KpTJ9Ti40TPs9dUF/9S6cPmOjKKwn0zs07JF7rdgZuklIT7eftSBL0e8pTKO//euE2YlPWRaE7
3kqMNQbaxSVadRa6PBJuKPUw0DS8LiSLSFfcvFYHkfd/7qJPa6a42h2Rwp06661oRVAJZ+2sOBEJ
6UxPeOlerDMuvfuBzI+PSylJxBN4XDPw/LGd1VtimxcgvKnhrj8Jm2zBvnyqsc9OTQO4RJ8vjNoA
Cqa6/09cN129IHnKfVWvmGLX2PJmdy1NJiFkNL3yTKBoqan9HQs37h4naYjYjgY5yA43+2YG+b09
wIkkkYoA0ilOUyyqkwVTfNf4YNJN+tMiEgeF0kA7RgIF6BxppZUdOjrtLuMdbDdR5Crf8UXDp4CA
ejOAaA4eIulovGPK6RpOxIznXkd6O12vlYeNvdw/zuw7JvD6FdUBVVNZ0nZ3BIKWpTkszfYSOcWB
j3Bi7f7QSxIHpqExGQDqRGS/MqSRT6+giH32r3nLggRKrHFEYIBNHpjE/VmJPLCvr8thTfWwSA8p
R/eA9oZluDihbfQakNXtyGNChJAAXwtmxQpMBblFadhtCWKESa51+hls0OOyTByomoK0xiExqGPH
i6Om6NxxALJEoSxibZMg5eHDNIrgyFeNet0D2KwLZArgBFgoBhtE7P9wY6GEmU4VE1RXypZnzxo3
kqX1okPWyEJ+lSZAbxA4IhMiUQN4CW4DCu3iG9Kv1rDEEeVQBOOKpfUmkb3bZvpXMP8jIqkoVOk0
4/H/hnPBCwOVfIASYDisM646iWmqBUCBgT/nDHu2GAWREImDZ4aEdQfakIHXyP7QEBLOYPz8Fu3u
PyXNRMFY8L5YewWP7GNZB6SdL0mp49efI0a8njWo8jWc7yW5SIew1MRdRTrhBVuJXRRPIt1x6YGr
SVnpyLrZMfKCYl4VuGe0Uxxkn8CUzbpQEn07iOeXHOBCB/J8XPOTFEpeKCSiRWnSYUjFoJsQzsFf
DitiQ2B3xN5N14aaCLrSvMj7lniw4D60botJ+T/RWEGSPLu1H/EMsi+LtBusBWx/gYWsYdip+rH4
THjp8iL30SYvg5Z1TLwoCMnIh3F1ChHUbFjebpE/iR8Qk3BUjMVKYQTvQNbDOeJ71xfCWz4w2T2m
f3fWuuQnhG2P4JOGK+bJnQsYE+CLLXTFhUz2AKrqRm+kebl2UoMFcziDxSmTx0zIqAAduLp856Ki
TRxpW99C5i4UlHGm6HQYF1T+BeANBaZdnrbXHhbczVrpO9T75l7RGBhQVpihKqw1Lbgl7Acw/UR3
A6zPRKHcrMmvz5HDul+3TF1J5kpLImUE7XyJGCsNGzVloNEOpOE0CqbBaEBaVOiJZOJ1oqiy1i3s
Pq6Kwz51P3q1hxoVKnjbEZEJuvwoDZMSVah0JJMvz/KgYYGJhMvjberGo0p/cRfFTuH4H25NJza3
B+o/btweHI3fv+5OAL5UwRuim1T8Pa3r0i/SJYiTxzujQRuBFyirEDE3U9jPW7I35laKaSXjiBtP
sK3bFlf67KTw/0BPEey0GbWk+4GHXM7kNDoSOPrTI6hWeSQjLj4UajmRZJmROIXko2+HDJ8SydIi
mXWOW0vvOMUzLuB9eA72SXNbo7MbjjpoGv+car9yA5YegFrwKOgF65V85NvNqitdqAkop09sSdgG
HWor3mdpl7+Wa1yoXhZoI17P9iId6SmmtSQNuWMQa3/G1dW210StX6T4C6euT2IhnoY4i//1A42u
bYIxpHVYIMkEtg9pu+3/qO1PkyBIrDOZ3dYehFvHGc1v7edGiphizKc8UoO/k6dCFMllf2vZoDqA
1jv2el2jMc7P7gnK/gk7kt1LaWKhuMKqMu6AvY8uCR7GI+1/ymwWuScgQ5ToK5KkJPcXp6bUAnvn
X3qm3TGyLZaQvhDtfDq8MCuEc4WF6qN6trTrxQXDYtuceEVbLumG/DiOqrvpBQjm1vdlu5Rt72nM
QmxElstNRWq77DV82vuYdz02vr9bekWQ1g5yWaBmA/lVC/L/jY0DjBqq9JIpl3TQ1DkWrOW8RZ9N
o/SqcHWa4nMtD5gewertbqzOwwodsk6c07lxoyrrERdsp0UU8+F9mgh9BQe0TzzeXNfaJCeM8EJu
YRbbie7qXGoBmVEjkXXvHVyHk1G5e7oGPnjru2rNtcd/FLcuEcu2UEKyGCaFrVG5C7LlEiGChQw1
fnnM3OmM3w0b0TSw37MZsPnpK8H3sdYQZqG6CZsSnYBjLcy1MHFCDJVIIsnl1rnAUCmX7LGipnm2
KNUy+MefxKSslbqvYtJnbU0CNBd4sLwXN3VrLiMc2h+dt5uSm+LajBPEHHoTcWLMbSAxBYH0smpE
mWDGwITZcKpFphuU2mx+TGzaAAvdE/kV5z+t66A1YSWZU5KkCjG63NoeRm5Z/bTk7zUQPicn0kZn
P07jGPhi4Rk7N6uclfvvlsCMUUAFtM7mYlS8JOoeQkaW81xpBuokWoLEYFIwzlHsg5pDP0CP/oaL
y620Ikfshe476UcUTsKpE58cSGfwadPUUPyrP2eO0OZalbW7UdAQsEKjrxrmJQ9VxPR5csz2PAmp
aHY6au/B9cKjfkJdnLlGQMEvhkXbrCgNVM6/k9pSuY+WZsNHmKLaygTL0WeP+PO3Oddk1n8vW11f
HeQe9KQQHLtwEKteQQK8YOYusFL+0CzaSm650xMJ9/lKDQio/mk9EaytCFcj39WxTAeojNZ8gsHi
j4b9H844MA3l9cOs44D9jX8AT5d8EeYgPP+H+W+VbCdZSOHz4QwM6rjfOGFdwHQlATZVW2mpX1KR
cUirghuCEGC3jTS507p/U26yGzNU4SxsM946fZaaCdn9We7evNfhQS9eJiXOr8w4yuXpWNRkU2Ji
w46fYAYiyKfGZ2ARp67BZZ1RGh8wCsT35Oo+HL4rzRqyDGUiHFp1mocIdII5HKv1cCqMCY8XwaVl
bfSvs2Nfil8HkDTUWPMTNlnrVbVVvFwCDnhpwoWKYxpqAEF6ar1azq6BfE3xj028nl2AY01AjQMM
XSfqbz2UWToxXhmZ1rFF3gQBzn66XiPNbUiy8m9RBb7ILMjNMpw/V5/9i6oBpvNPfoOogZE6oDOV
2P/WmqzuSueClUvW04x0FoQJTJ7bh/8LmDxmiG+6Z8xVeHQicZFaZ01DGt3mvuBD34Jy2hWA/0hv
OUKXMbGZ9qYlshltxqrJi+HsVMkuah+uRIuOBg65KQh9aOvAPuryRqX4mkp4eVSSkNjuxF6Vgc7O
+aHWH1rguOnoF5P9oXa8hJr41qlerZus+hQv6UHMNeT7n1dlxLWw2Q80IwM/thIxcpzwcuEJvhaZ
wxwXW7waOlqFC/SweB7KVbs6TxN8f0qemKpZRSXIBtY6+VHA7d/WZfGR8nfdG3/N8rbqLR/xwQla
9oVCHg34VObLC3jyFzdHv81oA6zBv8uP1lsDmXb7Ejy5J2qWQYJHnT84yBOf8G00X6FDv+R0KUl5
GfqZ3J+O3DffI3OI5nRxmr+kSeScMHOnCTDAV9UclakdB/6+kCww/Zs+wGViVFuf+cbz5MFqagKe
Zngrs2jGQc4tV7FGAO2s05m4Y0ZolpbjVsGDdwW4L5N5emrRCnNQpW5/Zj8LxzbjfmiEN/RUtx6h
oGI5F+UIrBsuhzvzKFM21c+ny6YFW2F9Zz+s8aiGhtwZyVeWPRdwoDaD/q/fj/yHdaCvSWceqm1c
KVWWx/PcjY3b6OKLw1MBlAgYN5SPs8/DLtb4smnDjQlv1Pzb5ggOpQFdl2zZa2CwPE03OE8davkP
tHrnZNu8+p2CfK89b+Wuj8tcohMwUMJwsETjVdR1YXdjPfBNKUncq96v+ramXVxhsXP0M4zlbI0c
yratq3cssfh/jhZEOBngdKHC46/UjW5McvexKF3p1kU+u/5pjLGToVGgFqpL4uPhNz/8xIJQ0LME
u8HMeJm9+kSpMw1TDyYAnduBsHu6ZP2kE/raAo+UcpTDajz7+o6TwXab4wAC3Pu+0CmB9L8AAsYi
638fZWoTvcXM8GFm690TD06T4INMVeFsZCNHsmUjh4QKnb8qszY6OmrvI9BdcYQquRp8h0qMOG0N
fXnqy+vaQIIQ9cdV6QP80Y2Uedj4gozWGcStcebo83Qczp4gzNxvl+dHQ6LxHFhcakEr/yyqprXX
hYv32/BdzaOBJK30Pey6GrwT1UGXCDMMY1g+DeFVJQXs51yaP84HyV095bSJWDMPbdQtPdVZ/K0Z
oUqyzhfc6qoqUET7zsnkAfW4/lqAtsqOabetI2h+cNZkbNDXqWWnKSOSxzxxBLkBlsDXYvoWQ6q6
gIy8QwfDjVg2Jck26smUjiHgG9z1I5e0iIhxXLLN6pxA5FKQ9wTKzuHwlv5Z0FFHNMZgT9yYiopQ
kC9uu4uFRkk48daqcwJ64FT9A71pJfrStHj/Aff0r17gNc6uibO9OIg7xH+B/nFfVX6RDiqbi522
gTZ6qdGLA6xWz4wmN9fGfaox3NKEAXSDfE9kJ0C0IUckSmxJDmAqbUo5vZxSD/dUsCX8dLF2j64V
QZmhfnCauyvmsFOkaWr6OOkDKuVQ5qfWqR+WV+nfGfQ1ITlEpP4GJWvhg1VhCDf94EWwA3NE1ne+
se0ClqMqLE67DkadevWPbDkZcLEkWErB1eLhohzuo9ldAbHyBNQS5W5uQ4Q+/CikpApSjrJo9Waf
YxIbYuCB/BJgk0M6UPEhJKZOCDCzZgoDvB/44LJhyn++HoaZacDkCFevVopjQ1g+TVnADZyhVguK
EGcIGg2CLpz4qezUyk8EHENU18ZoHRg5bp6mp/vw34eNLK8VU6EZm+RfcPQMyhUuFtMujymxjLdq
zGS8yZslEe507a9a7T/aFFqUWU6QWYgKT6Ud/jl6VSfRppnlU+slJTh/cJVXG05QuwIwxVUAlTkr
drEvNpv88yWFCbOQhm7maMgsoe7QbssrrwK8WOUJsF/hVHhtLbdC9OtRqf6wwamdQ2/z36PKD1uJ
sc6wv6det/PCfwmd/xGFYnUBu1vGRPVF72pVbQU0Fpg43VsS14XOBkvztxQPsQZpcgsLzGb4MNs4
XT5IDq+j3UT1pMkYJPQl8wvHjhE8muoSYSpF3NOoVINrmyWF2Drcpu2CGzqedDsypl64CpnegcS5
YraMukeHEGMVZ2Ew7thKruOAmakNAswMvYGZpmQe+Q1wu4+qfwX8rQ53/j2EVFgwMLF77SaiywcK
muWpQhSPK0rJMPT0g00Gdd2p8RiM1yNGymycmyCzL8x1rfyif5jzC0Zt44UnkX9AZa21yOSjfhWW
NDzuwWeRpEl5RXObPmf627pRVWw2m90J3a2NzCVIPYkiS2ZcqKzhzcTRryF31HZ6FhyKkdqnawHP
OvlGeaH9SYqEnANIefO9jluj3n+LtwZfP/4aEPMsucYSbSTRfREjImYiK5AnWioiwRerywICRqHf
31SJJnijT2SzHVSqg4JEylksxk58I9u2Y9OkFsM6H5TLb4IOKkUHYofmrT3EV8zQVk50DkiaFniA
7x52zivQTawkTZd155eOJ6T3+oMLsRw3vBgJowqJGHvfw40B1MtkjMyUIXt5ZQeTMYylFFcb2At8
kBD5rPbeW59PVnKedNKT/+hDpJuZ3NKLh619WXfDbXlVRn+i825oFhnRjoGvNDeFIJPLB77ef5Jd
RFcPWdFPC84OXYFySRtEOGoM3fDwsooSkMQIsozKi8nIguEH2DLjl77STupTZfvc6/vJBuRvklyt
VVVtgg8gSS8z7J0jiWFeS06tz7N6B9vq4STC5tNq8wSBvzYy7RCULbX//5P4e1OvAUyhKSlo7w3g
F7QxlJl+elqK6kI+mcdK50ZWb2JJ3ZQEfeOxW6Cdz87CC4sQZVevlAis1vIn4kufHj00EYulutNH
1qPLnTdFvoiVZt7Nnws8tffPEyoM1JJS1Iyjhclkhc7LUc2URElZoW7R5ELPVOiwj3tN5ZHS5E0n
Z2C1eH/cgBf1j2gclWCIhzo6n7ifRRsS9QS7a5zMy2cmPHLNKT8tGrpmKiNjwDSb8lgklq8v6v/W
2YMT3eS8aJsubqTQMgPoZIVGuhtoImiduPOiFbTHk5QhJnfAv5lRJi6ptJ9vJ0wRivbszc2WgzLO
wgxcHYzgVquHD+WqZSeXHhe+QtotyADg/B+qrKcCPtlXNb2Llc94bh17dBV/ImK2zo4pw9/oej/v
kpNcOXkYr8qL6SpYIV6/CmyTCCDKZGKp6yF/+wb70uO+FtIt8ZgtG5+alVaaokiiXNY39o69OA8g
8mTW01OroSq/qWv7IA1Iuhs1lXzHD7FB5Wt5v1B6PAQaY5rhOVMX/rsnbLtqMKEJcp23KEZBlnkn
wpa8/7zQfnlyv/3JHgZ0gBoSA80Rs2FcGfWhxddiAtzfrYCNW7c5tZnqJuDvMKJbzuMMTfU2dCM8
EhhDMO2jhwVRqPsiTcCpdZuZw7SXQyZN0I4/eucQsX4o+PXKVTcE4cbcimm4oC/Gor3wiVGU6EQG
CwWxyN7iJQBu74Gn+AK4m+CBZGdCxmk30l/dDwZN6CNxGCAhttxg91hKirXndCRl2QAuXI+LXvax
IjZlvIUZCVt/3cTnYY+6AHgTxEwT7wNIzMFmaGbDMNxgOeSiyJiRs2ix3aQ3hsOobM6f5/pDNVYL
cEH/TWY7rVnt7IcIOpWvZPF5lGBXbOZIe4Ka2JDUZsVPO/AY3YTGiJxE5A5w3QNAnvET6XWH910V
+Lh5FRpJtfWTkc0MC5RwWHgJzTtbmUd4qMSj1oKAZKiWgD5t2pKs0mEtP5Zf2IptgVUfkKkO1H8X
J7J/7cwLqYLF2czo8QseQ8trsx6BC3cIrkTT3vV4E3Q/DYkLUjD7sc4LYfl/iRfmmQBKXq7o9xmp
rP4zQSxIQttNxSLTV6teafiPLZ5jAbZlwyCgq8SvDBCTXfqKWf6wfTk+kaO2ugtG7uFIkyECqyJF
qEeJZt+i1NvRYXzIV/gEtimbvfnTJcr72Ct7fIDkKVUY6yno4BYEkwA0ej8mk190bCtJ4HGoST43
WFWdEgAcFFqZ+XvYvbCCRQgws4M3LKk1KNWqXg7pTxczhJkUyXRK5iJby1EDiDImRbuck3vIarj4
lQXljhr4uF/QeMb4WqqkNBgoIs7/2T/3L9MDkZlf1QD9W991lNf581CXUlqgXRGKajEoh3Afo/MF
GNw90dvYo02oVqmrrK4sXNO9FIWI3wCMw73pGQFR+QF8SS96XrbhlobgTCHfjfetcD42+WNL4eEm
VQkmqLuf6Ty6dnv/Ryxi+/ERyaWBJyR5lvqtkIERW4465SCdrDTRTpVKb83HmY33qY2uuDj3V0J8
53i9vCpLNL03KQ2AERUyfTZmsc036Hw2h1uVwlqGSE02eyKowkw2OU7XZQJe0HXYaxD1STml8QUw
Qk69JIm6RgCAfqS2KyuWRvReTIiM58HjdA5AY1JH4awj3QJnE2TVVr99QRBpMwLiylL/7Qq0lFxG
KtA5Pv2EYcbDjjGXMfLAiMX0mtQd5RNWEnvRRmIT4/OoKIOaOB3EUFrG+hsjTq1hw5J9Rl/MYcvU
xmH51fJI6hBxHsblNfPCvBoxSfUzRX/reiXqOEg1RuQMvPBdBiV6+WdhM/83yDVGQSIje5+qK4rH
iljcGho5qa4Lhw+0FwB80EA/dob3xPojEKkfxInIIcOr88eo3kj/V7nOSZLdsx6KmUt4jFc1wg/R
8NPB5APJMNMZYuiRAiNBC3memxDcnKTkjid0WwWcR01lYq7tc7VmJf8MyX4qQr3bote7bfsMCqPa
wlyeB9qDlQRAMbZyw2zIz8jZuwbtiYMWIu9/hvN/DYvh747EoUI9K0jr6DdQX9JfcKxamm52fqGc
jCkbGZ5aF28UKKj3FsdCVjCJ9rw2FZZY7uGoUhKxDjQhrj3Sis4OEVMANiAwLhNWPl4MyRzqoWII
jZi9fcvK4vS7BWE9P1aQPOnk92ZngLh7bhQjxGmMghjpqXi0wfvPrn/YZJIWcyCJmuMgPUscuCwk
VQXHEfaZlbjrEbg2WStQkCtXaFGvp3ba43Hiz25ndMPRPam7jDcxJps6CuWtw12BTFZOswSM1oIx
5k7YQ1E1+aZqVjtBxXH/ltm8U1tdek9TELDnxGS546afETI2irZf9dG4VM63guUvGOQPUMuzoeED
flpfeeaumbNPZM8Cj++BnQKN+TNiAU5iFvSElCcBhzmwblRyDSERRR31hO2O/OWHH4kJzU2U3m18
+FVr5OgaADsxzmqZcoI/YZ3vukAxOQLYKnVCCuK5gMdFBgADEdHYIXhzxT6SflBkfJzjc23ehkOY
6/nkbQucbzeqDgq2LSm8LWUhgo/rvMBM1ZDWgTFGjq8gmaqNMlXDVlnSkA6ngrN8r4bbi462K5u7
t8dGHw8dE+5J3HA6BSdIWja0uv3OEfryFSrV1/fUyxcap56fCJ8NSeX48MP8mNzEfMc7F6KarLE9
mDg4AKOlwdw0AkA6qedy0NzUT3XFRA0ZYntHEkgLhxVzaMwZAmFCQ/9E9v+BXfqNlw2D6IhsIlfB
3QoyhE75+e1dxezywhEau3/mFcgPDzkIU+RWIhdjqeHqD+NHqeYQTSeGcZHqQreSI1bP7MYiADQS
CD0FMuzOsZf7u78/QPphOGwPyyQGZHhdt6WYJeU6KgvnTBttumgEBtGOdkdzHOsJUdFZNaCNqoEh
yOVqTTAXP8f9HjkfdY3XHkX5rYqRhPiHVtv0BHI36g/H7YG6b3eqjvP7jcV6yo/aUi+TEAd79j9G
z3UsDAmqp6rkna3RbmfXomGIQhsPTMBOtlFTRk0xCd+mOOdJdwo/T927TPlCuTq50Z227sdFeYoa
nI0omZQIOvTYLBR6MUwaKVLaI/Rc/CGgbi18tY3ke5NAqjzs3dpMSHoHa/ww6TvoGTTf/J6/rYiX
ErB6yS5lfLxsPYDuB8MUNZpwhXyTZvoHXQ5YVY5uDxXlNeRgG3BX0ffJHqa+WDbW+YKp0sNKQily
kwZ2hREGyXdf3Z+J/obBzy6qE3+bCcym04QTKY80Ceow8F5JQf8PIQ0IlehKPvo9v0d5BS89P/I6
5YH82XkCDBqUT5veW7AV6hqkxUKa1xPnovUv0zrnDTP017D0GCMgPBnT1YUqLKnxch97+OWK3cbu
vBPLUQ4y5FKdWTRFcX+bMOQQDJJ8XvJVdfIXxHEoHTL3X6eiMsaVyAJTcKrAPg8wxuLw4PxlW3MS
NbfV3rHd9HT6+gXNOX9TgWHEZ257QbNZ37JC7IEzZNtmzca09EsRRVniBGYX84JI5qzz8WXpbTnW
5f3OUokwGPgB/fQ0A7YOnmN5rfB4JAW7i/8rvOZFnq3S9MDSu/fiqgpESOaPBmsj67YmTcsitVlG
6QTGTvsA8F+leJjEdv1jwqiEzNI7yJYb7GkZwpg7eTqFQ6aix80/kSofHoCEgmYUNIjdlJSKr3qa
T3xWXWebWloJtY8TuTLNmaRFOF8xdNY+Da1FO9Qs5xbed9X8Vk2cvPorU8CQp87fLnCkNWVj5cvT
NCL2boE0EpIjLSNndobkdIbWTiiGVMXVE3tegngPoTWtophbfBfF1FhZYSuLEu7Ka3id0/o22Uf0
4pkf3p4/2U5XY9gcHu9sdtc9ovrUkOWVj4ReJCxDe17jAekMhhZ8EKbmWiBgLJ/fZMyk0L6Ekk2D
4pWyakocDXguP06XZyqdOmF7Xfl4yMRLdEpvhb9l/7J3PTK4kEqGxdFv7oobDkN/GSnt1Lo/JGA3
gFBmNZqp2flqgxAvZ7zdyFDAYpfHfutaWvHj9JOmlilu4/gZRGIVnOJU4QBOYybBfZrdaJioTyoY
SK8i1Dq8ciH3R+EsufdSb5WM425MmXwkcutK0qGR8Xw0S9odMv/kYVw+H++vImS9lj5sBj9ZDMfC
e0Sowng2kRI3dDyPtAzKmJl7raR8n/FhCrQ/kY1tiJkVSlOl+MtG9loOjFyuW9NMbVw5SYTXTHa3
5U6eZ3aGaTEfkmRGdbHHuSskqohm59THJYW/2rUSH9w9W2PnlJxN0d1h6Ma7f+w81s+iPcwiRRcZ
KDDGhus4u0Yc6w/B7I3PAy7AaQY+ReLLYPUsmA9veWM1Fk5bteHfBCYN0U8X0TrbvsiHwGubxwof
Md8sYmFDgonTe1ehfHFiupb9P4Gz/fIsCsAXzC5RoBndZZQX2sn37sGHaXi1+VNOxkQoC+FsMUkR
V81vk8tUyCf5LNRKEZ2IKUOz4f05w4c8Quta0EYqlAX2yku1tOQGGFEJacsiXxEt1hIKhq2he0dI
jRmSWymzQco/UVmvdjt7/v/NoXjqe9CgD/NQrlYGHPNweXm6nOI3X0Gtg+sH71PQ1JEOdN0FS7rb
KbT0V/ZWlYdfXOSYbV1dC/6B3fNDQHqlwOEsmtvwSwDkc03UIUU/1uBAqZeh50+VmmCqcjZ0ZD/y
sqdnZDDuRHR+mQrHKrdvX/xjqlG5mSQI0c1pxV8gxnUumaFTBgFOjvi0dtkg/sTo5+JpOz9xqyY0
FmQNhC4hF1WTrQxoIWwHNe+UVgaBs54ILmskRW1nmwHzaPUw01x2EVogEcRfRsFJU7o7HsKJq/iT
90B6TrBBZjyseR2Z9LyCboXNfeKQUDP8i5Za4VYkoEYMhQJPeTcUfr83PlTP7xhSvVlMdRtmHkTk
aNczCSqAj+AGi6fTFjAuiZPjKTsYZtbimqeFXXGCfUkjT6oPZqA5NfLJxvLoSNDeoSAVElSmtxCq
o6VwTpZDIITI9qAjNsjaEC5GjDq3ES2dtKkGekUMD0sjrrMzNgL9eI5pg92E0acItA4Kn02mcyBZ
uor3dgQuKulUv0surL46MNS8PXCkUNTESPy8L8yKLnsfr8vC99cUu+HFZQb2ufOwTSubP0+xaag8
CgHcC6HyvEYrM0jsfpnl+GHQRHN1/4mgHvRNkHfAL4G3PlMhkU+svgYXC2pT5wwsQorNfF2kvfcC
s7sK4uyQStabyf64dTmrT6YXGqQtAy0pzI52sGT58h4oHa1Yc/TEFFOx+U74tVWEkfrxeAUy81PK
rGHhUEb34pCFqEnsVnWMfCnrT8k0ET6OyW9U3t4ilmzdyif/fm/rWj5nfWtWBP0Fs5j7liee9/Cf
KwGOidCkwgtnQnP8Fy7fqsD1MLyk1oCo2CWGwkyuRY4HtPwmL8aMS7EVUTPtcUNHH78gpNeBkVcg
/3d+asQK2OdXTZIpaX7CBmpMHqroyNdLyFCxGP7ZcEpSj0yqRbkIRm5WBL5T7ofk5+MKGvYxMlAA
CwvinKgYfFNoMCYLwQ4nEWC1NV+BZ+by1v38DUAqs8OQx4SBePLUZYnUBmVVxEJ6q+SivxD5Cpq0
4HzaqUlrzyErfyCLV4F9t43Asg23vrE3j0tc/EiBGZXYq6ClfDC1npFYmZWTCwi0YcdTlvm89cqY
mG+3UmYClfUTMMBzUBfJcDF4VRXu4EaUphuojD86MW+z7VJ2FcrgDFEpKChKLrHlUDR1BX+n/vwH
uiaPxZWg/79iM7T1FBA6y0vzjeVUbFOezUiOjqbWIe8V/I9zXOUTkjaMV5XAnoaL66scIw7GHch0
IU1cCSwQ1qrHC+e95cGROT6GSaQKwDtmJVN1EjBzicS1bR3WE752s+BJw9rppnlJLEil8r4R5XkR
8JvoTw39LRdVY6GrskDB8tPVuO/sDfi6+8UgV4og5rttFhs8jh8QtHH+55JbSiTsrzzbCwwo1Fnz
ySYJroWKM8V7ws6GKR9ZWEKXeCeNsWtC8GNWpHmXIIeik88bEeXIIKmTe/CQaSW2JDfHVTdFYuWM
i2fYuC3zYdihRgBqkR8UIjpcRp+dk2Kd+ETcJWLz8IUnPrPzur/1WwGBwPwqF0+FAvQusW60dHeI
jRb75y3wXTtlpwK60N0h71q0ORDD//e77VKrb/dQcgYdiWasqb4C++8nM/XQsYqDZUu6CxZghpZv
wWGao3X5/JCIh/EF6UvvVt6nOtHjwdxjTzBvdzkLys4sNaMwNwIzxRJb8ZWjLC5JGU5CtY2tQUhQ
JTDlyQBkEAPChuIiRkeR3nBsc5sopB97Do/xHCP6794vQWJFWOWB1dlB5e9ZNXMyUFuldZQh+uAs
gLxqmgcrbymOBh6ONcnSSAibU1gwUK0wNvkJoyQFwbsMallCFBdxtH/Lp/bN55npiGj/VgORyZ/z
JYovjhD2pwAHxZ4vpljfcwqs03EjBFJuYXCOUwnr6LAi7/cDyeMCrVCABHnZHeYn+4g+oAUQp2tj
r0hyyL/0hnUmHMrGNXftMrJCV5Loh2hJsEtaSMdOwxneZffiRMC4n0GeA6CyhBhRN5JJ+gW+11mM
dT3WocaiUsZgEx79D/2Lrfg7s7v0MCYf75FnSZ6/Edf+ZDKeH7js1VDnWVIx0yJj5znNmyl52VUj
NKzfFcYzWkeXdsj7ExYr7ivoQjy60ykNwB4hMpbJ4lZFIQddtkuJ/XKAKG8ibrg7fRQHIOssrluf
79B5UL8liqeCwa0zqIYdhXfvOjac7P3kq/zFUoJJFmsxXERg8u0h4O/Sg6BL4CoWWNHRrQ9yyMAf
OY0QLYWl4Ineu96R6NrP4ZFVV5nZUiRcpjq/+3jTbskKFyh2ZteuqvIzZhYiTgzV3gByF6jATzlM
nk0QW22IJiINk0nLohd+W211YKSSijezQQHXUMvUfAYLVASc7sM+ATb8en0Jn85uA26jaJMu3upS
2wi6TJfLrjaTehM3C9ti8mYILCVWPBYxOoGqc+mtxo92sQFrLhFB49UdsUZ6j2pSr5y5N/7aZs3J
ItzQniaH4BnZTm+0HMrCLPJzgjNJMwetAZpLRRljt8SQ2evXZ8/9fHRYG86lVPVzr9lukhr+PEG6
06GigHgohCrHdkxM+2UTB+jTZWNCSQkFbFUS1SEY6T0p83TGcVmLohNhSlijgRECGKw6ixVxJ36k
W8snXq+wqDXZZENr1Bvct7bUIRG5YFwPaoP1UMLw2+b73xbMyJuO7BtBVU/uy+rI9DygJaJ1324o
XXXsMzN/izNd8dccwU8HBWrZgFGg0B0Kxb2hPQv/k9NCfBIvj4JmcdzqibWnmOM9cKTFch0U/Kk7
CP4zszAIcqXzfUdgfDae9TQey+6NGDcow4+E1a4ndAeSZan3k9AwWKA4O2eIgsKh7QHucJmJLVEn
qXK8hoaSx/S3e76vLLyZ03r6IRBeafcECEfWEVrfDlZcU7x3H329Heb3zdaEKL7YJavuij+GvNBa
EeEjCocWTJPPZpdXL22Ckcmm1L0g+gpJMzcrsjXK27kGiAO+GBUm9UeQwvM6R8FLcO5/CewtgTgE
6FbHvz4oo+LFO5zb6t/YXDgJlWnMI0ldsCYrBvFjN6mQSGodn4W8SUtf663rtf+dh9uL0hey+9KL
iCbn3pYWeYwr5KULHLIg4Fs9HwwavJj7TkkMPWBjn+jL/p9Bs6ia6xdFVjQ2RDv3nsxtEug8wpKe
l3i2l3VXgiCIqcWgOnI3Yc//GAfMSUiN1rOUgzHHLoKVjB8qtFwsXYPvnXIhvaSITR3KGK7WnWqX
2toK7+KAacbJXNEdBAexkazI5yh4Fzp/1DnWsTn9ATJ/bmoHm6Yp2juLOVdMZjgwTe0DMvWBexmh
/XW1gEluG2dgKmnWhcsRV4m+YyQqj/I4BwkWeG+YnNo5jqo8cDA7ABBg8QjePqCY6hskF/RSDdTW
Rb7XpQjJb6GlSIWJasDQu3J6rThloyio1Gg3nqmrgwrJ5fnIdJdcSXYdzjRukXYZflppoXooSzpG
T3KifWq37U7ivQo356wQ7X9qbVSsfnjHi0VnzlrY3NDteu0x+rZR5MiBVm0TpKCfmw06xZLxmzJ6
nc/7wWspyPBpDPz6oMwd1I0Lh3Kkh8tAaH9/SO2DciwQutX+yQXLEIn3XABUpGO4+yrkP25PAlj1
OdM80k4gya6WdUcnpEuJFq4DEKM239mG9Dbj1z1cPaaWCnIySLr5jGK/TWweCM3Ck3lMFAHV7GCG
KXaJNs+ygcaIJtDWA1xK8P5NxwXBj9NeHPg8KaguF58Trwk/1N5cGAn6/0ERmJBgV7zmfIJ32Fs6
AFIFdRhebul6ihyZWyCiA4b12WNVwZSaoMyG6kEk7ZHKK8eWdi+JjrFYO45O7FQxS1jkh/Q/PGxm
Tbi00wTGggMWLX5xEGbeqnyvXwM+zXsdJfdrbJb6tYuFDrPxUPaSiAmu7VbJv8VY1LFqhTBT3lLz
s6a6g+kesrNv+v+eaKHQmgMhri2JOs+69Zegggf6v5nX9bLHW7d7r6+plcC9cMRBQUYiHYlVY1L8
YS7yRGtVm6HC8LjH6gFDm7qcFRMcjMn9JbxSMVOHkA5cuc/cl0pvVXhpIbJWia6+8p1HMnxr3IXW
xKfIRtEpDWrM0/HSP+lv524Ge0scYoEn8S68NULmnCyfypsUicXN059/j/ar5Nzc4DJboDwJE8qm
1m9PZfjKZWFPXjy2OZFyUXI0KPr+4MfZxMJJaVzmAg4e+IyvPlBFlZWWrEcqVLYs4UDMalAtehKF
mlCYXa4Tcqb9855fYNg/hWjd2zyx1uAC1/4ah6dKXbsa/NsqylGvEZwXanCw10TyDKp80gimkcIj
3jcENHAX1pIPsa8q/WFeQo+75CFFsZY8U8u0fS558vWg21O7d7eLOtn2mp43UK35uNgRE1vFh9Mc
2joAO8xorJMTBShzYmf7DHPXy5CVJzcjRnTAc85onTRPL/FOwDH7HBwuGlEkhtxWXlWnatnWz9Vx
lwJFKURaVf+xjUAnWhXs8+efvqBfeXOHTP2ZqrLLLpFTcInXN3BtX+2iYIqpeqqzeqUzpNr4yZu5
cQlG2gw9KkT3u3rLBD8TVzyuRo856m82fedpRdhywljWWxygQN3YFb08R3/NHdwS6G3Vu2Hmc3wN
pC5eTdhKc5jDSx2jzosTo7PAnQFKAr1BjuVZNDO69NiLV2EhkEowtQNyEsDrFdT09d2pkrbLuqk7
9jxyo2lE0zhd2bkdjRAU8UqIF+uSPMTUc5GRzbFrUeZPLkvGexWIPdgwFDrhMz9nPL0/AtY80KER
7iVXXz2mthpiBxHqC2nZiJ6mAC4LbgrTZ8D+rI2rq9lRcDRTp7wTddsZ3hOermwkrubtpameIRuY
4tdCbLjIzUROpCHjkM/4iEcPUdugy4Cy9V5LAsU7S/+tyEWcVvzH5WNUbmsD4uKqyrUgqIwzYfnu
XQDXkjFgKcI006BpI9opbCj8phqWuAQIWppGMVUYF1tmMeWh90w4mxwOyRN6wrEnCnLCPDiLVLXl
X0V7v8ifhv+PKm35zVsCn3TzF90KmOOLoOI33/NBg3SZAuiO2tNHslV4IAwON70t/cz9TKsTT7UN
3nHMkfA2OFMgin4XE4WuVf2FPq7KfQnWpUWB25M+YNpj6GDacScTIixSThDDR9vx3HHJMYf81cDc
HblHJFMJW6eBNHVJlO8tIl3FAf74vRBRjIfyrHrL6Im7agXuTlnY5kpRx4KbqeOXuq+SfIsQjt7v
vgRtpfFZZcsjNy7oA4598CLwAqSRMdRJg5PazoQCkGzOBZVyQq8jXFHFPVUzwpOzak0CXNJBViVt
kFDUnJY7aEODqy0c3mIle0GLKFyoqII8ULuldId4h14NEQeyb6p8o6Y3hDBxojjeD3Nr0UR5kd9S
o8DM2sxMfY0lbmqoe+eKKjpzbcvIzf6r/iA9C9syb+obfWFhAonzBJkDBQuYE3Dj4F1Vb/VCgOG6
RUUktmc5zzw/o9sFVCS32Fkud9ORaFwp7fGK4Hye28tCHdYaIQHfJii9fFRO9BTloNcT0vVXJXvB
oqr6dX3m3O490CZb6aP7OlnxPyUhaiHytViV3qNRxIAzS2F/bh6MozTRo8id8sSxe153hJ6RXAfa
8/1Gg4bvONhune7HysS7P8LGqr+w1E+Hhbf88p4hL04f91xYlh+lz6aL1IwNC5/gyEoSsvzXU3MS
JGVvyYxG/+LX52GD4MidQkhD9BPP/zo9QFDPOHEkicX+E6X/sdVXdYaG8MCdsTwK5yA4NVazxMy2
ut1LssxTUSjgWN+rpICdAyRF8pHu06BN5R7gKDF9Y2GBjNNDZyEKIfFTPLdnwSKR6G4iugy/5uzb
2hmiwGQaANdGRFFzhG/MyoNoI9/n/5vfohqAE11R+2eJ7biG7G+eoVrxwq5oPolWJdxWdsZJgoaK
xH2f6hB7sZlGi6IiSLIjL4gEcChGe/vYhgYO7urLq+WY/1DajuOJysV+2xDY/2ZZ/Ymx3YLktWI6
ME2JqTXwF56JQhwUfW9xmE2Q9OAr+U8b4UW0RXhTUtH+FyxwWeoaPQ6ftewwAfQvWOA7HPwNVTp1
WJj/KOqqRLtrPyXM5LBrmX4pagTIFP1aLAwfYHiMfnJUwnuY4HIh4IfLGSAQuD6S3kDpfBfehF5G
8yS+VTCaG2GSBToOiOc+LI0oQgOZ+5o2Pqd8+wVHNbNsvhPw3tU0SkbOq336yiGc3nWgLcPE3Jrj
rm7ltVWsKPEX8t0US6rkFCCDV8qIXWJ+ZK1MqXn+xLogQr9zhUOpT72qc3/dlY1wfin7CYEIQ3ai
m6ZYcAEuF/rfjbopH5rSB4jHgf8jDqWbn6PcmTCrcn9CY86KtJJHEbe8Uv85KEczCS3AhV6sLMsQ
vHYZNWkgPCvL7o0/5kiwgQI19L7Ec4sZMYJpYXI2YV+54DUXV4N9Hvu6phHOr6yY527IJBTZF9VL
wWJROPCjN6eWamn1hsUsBq6lD28XZzds/dBu4ErijV0reNJliJqYwztReOF1VbFCP/uAWtAjb0ue
2M2tFaPwbi2r0BOmPFg74/yrAdVttuLUWi+VO/lX2Ch7HB6vkzyhKJejWivnYCrbn2dVoWMBXbDm
2Pc2cwu+uFpO9UjfBVxuswgMpOwyNMsvuDrl7WPA/GIO5rTF/EvvYSWEViRGxizc3hts90WOuncX
JyT0ois8z59AsHyDPopSLZ/XGJawTzeGiXs+ZOsyOrsGq8bq+kmE61mj9mnAkUZ6R1EdctDeqrBM
lUIEjoTFDGH5lCagPjyQgf/cHqdCfAqj06PNXeaBqnAbf/MlDXAHxg9p4rWb/K0qXVXp5dBTiLnM
GSzEcXA1xwfVXnzcbexEHse6Fs74lKOEmlqKtydpOzqm8pzcFP6Iu78H5VSnouN506cD0U03Q7vU
l/7NgzWKBCDB++hi5Dbk+kgFqB1trJXq92bdSkP89x6Np2dJxlTdLanuTiD2x3l2w+pelaBI+Tl/
wJ2o+I0bepDtkJ1lu8+3hwtTidEYZA6eCl7qspnqlGmz8dumHdx+51fncbmWnwp1v592qi6RNJot
O6no5CVQcW3vQPo8+/TVlR8swvd1Meh12OwOs2C2xowVksBghH2SRzoZLn36xmDrhxzrDCHlgAOY
K4ZVlsJXwblO9pER79hpwlMCrraZr1HYbL6Wmkn+FTzdkfRMutPytQ8vu8tLgEfSa/C3Wl6AIKFJ
qT9EMFRqOODn02BUljksJDIHfOibGfMnEzPssYBhPVe79Lg5l8LX3Li1VwC4OqsAi6JYVvBqb1vX
hB/hhCIZiFzmfncSJwKVKA8cNmZEc3NGq+92bRzYuf6uAArIsNFPkeHiAlTWbATlydFZYbHnQ9uS
3RXuCsMh6svxmwQPmXygiNvdM0nwfLmFvLtKTqYt4GPWJoBm4GC8JSPUpYoZH0K8PuznwPzmpVbx
Y5nykUS8vbuMj6Du9Mhbz4FAZOpA37cJcVi/j/GEhq6nQSniVcXu3YueLvqAFsG0Gc4DC/DH3Xb1
X2FrF7qFMYdNw226M+fpDUSJ8TW+Y1YmQ9VDla/34sZWjzIswo15Zv5ElWr5Zg/ur1puOoAosJLF
rIAIHwQ1+/SnDG6scrryaV6+K2mqKRO0YvzPttpoY2fiiKe9VjhiHJ9u3bM70NX8OpKrE7JHKn9a
DArnOBADzVGItcTEeH2Mh3T7JZ4xkq8Q/vX+8qJClLLRHuWYcPNzAlkZMECw8Fj0uk8MFJdsAE1a
fnPQ+XE5HmxpDtkAhGac+bGvu1vLpRxTQrv//2ugnLu4BkPpjl1gyDAgeGfqiqYB+i8YLjkgPjGH
q24UbS7SKvLqqv3MxH7fUXQzYWdh/L+ZJJGSs57gqxEYKeYz9kNvnsbtUKXCT8FXuMg9JmJ8bmtf
uMv+pLuMPRl3OsGUnvCBVuqAqe+UsFt4tiogiUGzNtAZHYZ66he0okThBbVM3JixlTuK7x+R193T
/9iJnDLmJhhXzihwzKnt5WCV/AOkWDU8Ipjdk8cFAGMSDsLhfzObwHjTQ86qQJRJFZSQ0n2TXOD2
kYIJePf4SJqOcasDlt4JwST7FbVnoRYi4YqU9cYCU0xUTnN3Vj+WymlJ/zanfdIWLdBrQjlmwKw2
cMU80CrmRbftMA1liRE43vtYWZtkH/9Xa0SobYemKeZpYy4fQGU9w1N0WTVT556iLeTmjHPIMZhK
wuN4dQv68DHDH+ubqd84bVaPiQSIOo0HT3B/EID7i5gmTMnknk+2LSDWf1sgBDddOV1Ffk3teWY8
Q/koMQ/TVbJ7h3gd6CJzFVbaU/w2xPY1WMj8BmXJPzoQNgL/zdoWJAq6WQcoaboZenO8X4xpL/ei
ATwG2QYAHkxnT3uq1lrRvKWQOf4rC11BgEOVCvGcPXR3STJu3sUGYfGdMjLIdGPrgvDc+TMHLPIn
uI8L5P7t99/255PG/hBBXX8kz38kLvpqaIdFlQXnff6EY3vM7qf2FV7fOITwVOUx3yYIwzYD8/WJ
sidM0SOvgSWXnptDEsspBFqpqQXz4YOkeV8w3K6QfQppt2v76QI5JeUR4nQVHyCTfDBb2uVAbIED
5gQguZuX5Zjas6mME7edOnjJt8ISXRyI3GaaGeEbQ2SbPz1HrA43S8KHpVGp0TpJvi87inMMEdhw
FN4lApZgF3f/g850hV4YhQDCpl1x8mLwbCZZD/O/nocjdbh0dxf49ARAwJhJz6yLoOzclWhrdAdx
eL9+mTU216Hs3IRWWVZ4VzhTqq0jeO9vmMDFKFNr2O4jLKo0bASpIu6gRPsd/ke2/kaOoJsjzzzm
iX0E/E5ypxSEJFdpZTYJKdoxJAEvLql+uCoE+uJovrO5PyUC2/duSgrSO8T7I66hqgMOfw5FTche
oBl8ZNqZVjQGNEBw9hbYHQkrur/VyuTL34eK/k3HwCxNCsQnSYDg1LnQSPlzPftXKc/INzYmZcTV
zQfjPjnqa7ADd7v8IAZAj8xqaL3hwjD8ofW9fbnpQX+hlBylfbccFOzegPpNzRtnpY5gWrMvpKoD
xqX03I5qGeRvxbsrJx9nNDk8Wl/APoZ4Frq0+7mX/TrsW0qAuy+xGX/J/WHrhuDurehHSl8Vom4d
uWWFsThSe90rK8EhBZq0DZezF4PcQhz8NORjY+aMsFSb7DuhOGeONTDF8hqqMpuMrDJC3zrK/+fQ
k4CzuZE1GdQMX2SCSoY7TQWg8CgHHmV9HWP7uu2r4oEDFLNzeo8NEJ71BNOKnmEub+x96fDljJw1
LneIi5zlEQzh/dCM7H3YQYZ+1z1pc0cUWtHRMlIAQmI0hGlmEie87ebkJdQ9ijF7neor4REmYWys
ve02LE+T18Ob9FPSkjDNIfNTPCnWnQYOIamdaXMGnKq4MVSOVX7L4+B+vB2gLqtqZoZgpgFTKJts
Ro0dJQ1b9mHL8zN230qLgMTAwJVTv+GMJi2B3IgAV1Z46ky2/erW3Cacs+g34JSQ8AhMusDhl0em
g5WVrVe68x6p7SJQvfmWOFvPNkPsf61n09mYPeyc/sQF+CvyOEzwZfjV7dI6RuxhYbBHqtEv1WYL
mn8LTD1PhFOcvX3HahgpHIjOwmtL8whbTt3Ak0nii9+w2qshm4JfsJ2S1SFe//T479GeXIoN8O89
V8ypozSoQ7tfjHh1obQJ7vFBdTcXCZ1sNxwvue+tPN9Uta38wfxEZ0OB2jYk4wfedcGBQAHOiKyY
bFkmAtH0tRc3A3wPEC0mDOSem5PaIKqv5pehU/GFjERf9vcprDuti2c5TowQmgKTHnS0BB6ZtKm/
6GxvfQlVXTbh4qDxxQzw2NXTbbdvY8d44gfwKdt8Hiy1pyKV/fUeVBcaZQ3F12BegzjZ+l768+qA
Ff41957L0P+CE/DEcyIfd/9FMYahToyh97MZ2EhO0iocTYbYmYR0TetysCKZdi68H1JVuzUcmG43
ldrJ4zg/EkmIIO+jWTV5/V874j6bAKIrdC0EK21LZeVFdPQdPpGw+ePCSX20pHFbpoSzRAGMoAh1
IAtCfP1Eh0xFa43CcSDRGfNBlEXGF6Qyl4ix+DF76fxzzThlWW0leEBP35rHJW4X73PGRB/7FcIt
orejyhhVytukJiHhLU2VRBXtrnm6l6IqGaoWtNO9V/UY8CSGDhEK5T2aQitK6fwnXgZkPzh5IdNw
6yA5fmosatRvhEMMnqUR4bF2EKiKfJHLhpd+g2ALy/J2ZZFvuyz5Tm3/IXq8gxSogvNY8Gh6M2ys
Wyz7fwg9p8P+fam8N+UhzHYSOsaD6GRNGL/D365mc/GYkaNmxwA38hure7qKjGHuwGpUVgJMAUl8
97p/VdNOwnXZrGN2+nHyj5QZ31I6Ic2QEQskJlnN6iAU5eT6AonLJR8mLjUaqyb0BBxWHc0mJOS2
1Htk/yz4An9h47CnZAcm7qeS6uby5mZYAZJN8UkmrNDO2TifYCEORbHYdBRUOX7jPDTrTNKjigWI
JVKSkGbGkimWaRKPgRS5NASXYkT34UJRAiPuQedXop2LDtiFSDkKmtdBQBuHOWFTTWcsLAgBDBf+
D57ieMx9X9Rw3hwxrORhAMWB4c7HeQNYarUW/Ib+5cOA4i3YTEhlTEfdr/C7e0tmuF8P2QCPOYdQ
FdnB+qUXk6YCsGe7WxOy3MDUu3V+af0yVZf//ugDmpYMiTOh3tmVQ9yhTjkyyUbASQ5VE1YjToXI
IJdbxkNQM9OFWoDrTZijnLuNwQozKEeLQFhHzIdULahIUZIf7leJgYuUOrIHh9Yc1rAZKl+2UHeF
ui5tMttAoun8UvyeJ+40b3yXX/oGBdtv8MrGg2iUcxKS+vieMyxaZdMeYYjjM71R6DJtW888SK04
VvhvFzNtt7oo1Byd1GGRK1XGp0CMikwBLlUCLSKek6GvXJ5I6H7KmXZ3kfm45EOCO5D7ahx6ebZc
HSQFZsBVKYBe8Iof/5VjMbRufgzQIDK1pECCnq53CGSNQkPji2KkKp0Ylte9Wps0KMzOBjb4htKa
mFS6/edxfpKGrQyEdTiLe2ZTwoJOiRuMgYzl/HLoViHF57osqB8n20Uj68IwYdmK+SGPgZm66e1q
VqoRKruPUOoqN7viOkK2LIUBEGlmdJiKT83ftGmSlq+gvS38brPEnlGsWS26IHKxvOobrVSLQ1LF
NjfeFNwStdjfhgxfNEyJelVSuHAZ0OfZXew2wCkL1AEAw0DqYiMmvBiezw0c5SjoY0YL3jKxPsaI
FXtdASg5C0EzHNGz/u9Aeyo0dpw+qEPmKl6CwPdRF7FHHIwuW+AM9aQT3Ws58Vn0RGqxu24VA5Tx
mumBnqdD8q8iTOXAQLCIolCrhMvLVpf1mPGQ0NNEuSwcagoFtv3m61qtXdIN1HzAA2V+PqMgkEL0
9Eg7rGN9a4p2jdAq1aOxW79vQzWK3DpUrYog/xCPouCzOWpzq7NZ/tFX/uvUngZGQY2BzCfD3mmH
2ZtrhYoCZEeXNh5/RtHOEY2Hq3TC9HIQO144GI035IZlPm4nTaTGhb2ImbFHiF3PUhJukmFAnQI5
am8B8ypi5G2H8Qrpg8Le0pyKKvyz3vpllqmxwNc/YevC2oPbSMpb/PrWWYJ1joc54bWEMnQWau1b
UcZwse7I9yWHyVkk31DZT9CIs7Ii6NG/UYALlWxIvCO1lI+5Yt7tj2YbaJA0yTcgO3bqIrmUo9mF
V0GYpXumLcTz9iZ/BOcIXz4iEyFen2OTANgfRAS5b5WJm2Yu17DfQ4EWuIHagXHscENQdD7J74VY
ZeJ17uqj9aNZ41La3L6OJ3NlrO5ueHLJMk7bdAtQGCc9wQg6YkWHButh5XrM2oRd1mOZjvIVD07j
8R8UO4n+iw1xUxukWrRe12fWg8R6b39VHpdns11I+3XH4GA1Gxr+H+o1PNdZ7GIM7C/e/8VSMPXM
kO0kXjXTtUWKfPE6gvKRe3yCZZtIhXfKDXTU1ErnShGAiL5mHQHxDf1z+NAMwHhV5E8BgAv5QetS
LtB/q+n7Q0/ZjCVFoTHTe33EfVEXiIetP3pdYTgR4pPRw87YK7XqvMMOd4zc7rJT3dUBGguo2wor
b0fsOAmenOfS/7ceLwos4Bgi6qGCTxf6OXPGmnkuSMsQzVGP45C6phXv5OMel6SvLCNYDcOQss8+
rlYjdDfCR8G9v3lyS4uO5GtPv06zmB0SZt5DBcrMq6gmowj3wfMSliBD+I+ezPU/yRulDaZEotbW
DO4YJD8vfmQTaksC5DgVqY+bGOwg+V1r8hLKn6gP9tiQ40meoPyCEJtMwTDDzikRfXTUEX6+Cgam
g/DyxBco087+BoosYr7spy2ae2ztBNv8ZOH+srQUEWCQP5pJM8OEedidVQifR8wQb3lOsgSkownA
OYtCicTAuZNjIxMtSgI6sT7eXIVCmOHugscUdqltqGXdcpQwmgTDV6ZRFHDkWt96deZeltJOaEpO
Vyua1+bS9p0yeXCIW4H/oZf1ypOz6rczgh+vQW706o33wU4D4SyTV2952OZejZG4igm/sAnIH/J2
DyE4ziIzbcVb1lfTFHerb5nETF7M2xyIAD3Hn2au50WeRw6j8ZgHTYeKrQ90AYcNagbQnIRi95Ua
hmikk/Blo54P3LvZpWrlbmhs/ym2rOE+8z3H3huj2AOxP7c3X6LtVcSS+Jvt84C4aW77xnSS+9uR
o0RUK2E9SW/ErQpH5t2DfZf5MyIPK/lhBxw3Yc23SNQQwqLUN1UGdj8ig/F8icKJ7Awe23w73HVa
bwCfupboKZLFrQ1wcUu0BzgNgH6sPUcQu7IrPmcjmj1pMjTzTAr51VPAN4yGrqBAKoCROp6iy2Ut
TUgRtbck8HvsTnx5Bg0W769ziLYrRioMsu3jscOY9eRE21rkV8XZP2O8xek2IiUNigwFdMbTSYJv
hw/SbFVMifX6GP0m3NgYn1zWDdk1ZaFzfa0E2o1Px4p1C7G3UGaWhr/ZPQC7c++gA1LgfDy6pAra
jUU/Giz6B6HeM0dYALuc8dHX4J3q9GohPTZRpQs5k75EvqZq+M+FYvMTXOLCfohthiBv1fIaQxwy
X3Va7lEe6RPQ+tuD1n4vOnDVuusGdissHiRXTyMP1SRGl8tSWy/H/HtzWrSw4CPrtbMLT6T+Bx2W
FoK5KDnGdfZ3GtazlYQKyIst3/yh/kDsKb7Bch2qvgL2ykbAF12U5WqAEkbGQ7U7m0kAuYVqFksr
Dc4/OzOHj9hsXkIVOOlAOYPtr1P1LbdWXw716qJXIqab6Tht29Qcoc02Awk1QRGEvrCmgEZ5HNhu
AKPMbh1xj5c5t7n7k7Xh5BBnycJhCLZttfqRIvpT9DxNFESQiBREXX/AFHm8rE0s84uBvvgR9z2R
MxAg/eYNwRvlFm5/5ORR1gc0BN5Hnln3k1M/Hyga2ypR1E6qg6v06uKjCBC8Qg1SzIUuUr6GIdrL
1r6qodfFQ4FSl7N7T1M2cbt+X+i0ii5r2FqTQ6u/9LleImM3CIYXJWG82OKQuNxdEeIa+p4XkAS8
lk4KqP8fuLN0JvYUCBB2LMCqha1viI9zqy58VLQXHbwDIp+SDx0Qq89DZt0ZcJmTdIxvsMmH7p+M
eYelhvuPQ6TPUTmsrfpIU2KmgCahRDzj+IKt4Eo/0gf1xLdypZDgbCJrXsI+3C94NdKGGfF/Wq0T
/hCINRSmnFicud6vqGekKx0yrRQEusTzqiy9ZJNoYF/RUwuGGviKPFXJQaoH2NErkIbvRhZqLlGy
a9mNWbsffXa5U5iRUTT48M05djXlQ7eOCpkIxMs4d+sVz4l3XeA6gEo++Mx3R5OCbJBoqJOI2Pzc
767LOCRWt+SF0Lb3+rQ3STGebFYHR/eduaJk29JV/a3NB7cVg2xdczEFXXl9RmTyZ0lVlDeDehTs
CzPXU9BAX416xvwPQ0ym0aYEZ+ZYSlkhPDKcjBWNvRSYlrN9cKzYAfniNgXzBNd/G+FxwFbzIzul
tGcBGZyRF6zyrt0GeFAxwIjAyIqHCLUilgYewFbIlTFQcVvB+gbkK5Rf721dNoB/0OsjHzoDeXXd
G91kcwQ0ED8KwQ64hcgtlQWdvpHBRiddXuCmM4YsqlL5WgY3lejn6O82mVEyRHoSWNl7ptk1ttzW
N1MaKDwmO8MwTo04GHDxcIqc8w68z0F4yvYnP/iypl3iSO0PUznEBhRsqhvxd1pDU53X9er7Gatm
4811mCqeumbHJE9rDmzUgfm2wEMhrOQZ9t1Obn27yP7nGDFOeGK9xS7jJnpbUslN0L06rYeZWs4b
npDueeMvEiGCVKq+ICwXhG23McPlHE/Sy9QZ57AjWAUMfdr2AkZBUPYBbXWRi8xBA1hFo4s7ce0m
3zPlVmqoyl/G71CC1U+17UqP0V9q/yxqLTC6h8TISNpJs3QBVFS7Z/yAekNt3AjskO/bx95VOqeE
AJnCXW5RKo6VHC7gvLQyZaoH0CwMEIdjq6D8aSDzH9O2jL7RTLjWcYd1qpZ+IRhZhWGtY/JZa7Ds
LsCAtIYhQJ3E+1HoKcDp/G3q1jCrt55oke2Q1X9+XLH6zDJEyDJTv6vmoAbBxMU4O37gRUhH/ISx
r2BoEup537YkwehTGBaXaJ3Sur17uFeU94vthuspDlNXx4fTmwN6xyKomWJTN1Y1MvZw5lKrmE9b
yFhlFjU1NYQ6Wl+nDpYEvfL3XvKn5UE0irz0UK2hGhGZXA+ZmH+bFD2uj5UZIYuLk+Z7uG9ifHvd
lW9wKGP2/le+so59SDpBDyUtgl9jG8WTiRmFbog8NNmLZLe18IhpyN/b8H9G5oOYcYyKBU+M3IpF
cCrmlQQYvcyH6B2US6Fr/9Bol/VZcaVNKor20NY8T+32xOg/vaLVNt7BB84IokgsMVqHy1q9Phaa
b6QvfUTTr56mas5NBztrKrE8P1NKZP/8UmL/6AE5SPAYADNekYROsgX6Izcs1DXY9ZJVzg/YgdNm
MZ94hCzcHo0uCXU535hprab63X4fAj2B59+GN4VMWaV9B+04i7rqq///33O4fxsZrd6aGz7rQh3z
cYkBIJ1e+UPZAeO1vDCwy2LaHEvm2+1Bgin/UCDcdsgzf+9Eauj+SbvnpV/2FlrogR0qdFmOgM0e
rGwzCTdt6636bEGIMWPWvGZIsX06ojBMGD/S0oD6OMlYl2FKm/Vy8EM0KY175k4EPFcPIpw5rEmq
VUULoVy7dd/C6Om9bpbfevvetOFyh7j4GdUEwRkTJyrtLSEpyjA6BQsn+P1lC49L+0Gy/kBM8hsC
jv80YTfifrktZTfQIGEu/LmNW5UYipXQ+QwY2ngrRTeXf4gMGmZ0ndzu4MbJ+LD9G0jaCwmCIBAk
rGWcNfRaaHTHjCQQVCN2M+3OIdU14VP4kpk2RWfKHHbPN6jzZw6+lwjsE7t7HWxQsMfVvDYVOqBp
5cv9gqxk6mMR+VbCuVPMJSLGqmwywzhTHnd/gw7nLoCpYKP/Qdnbg4VsDosJsQbsCFTA8yMmIOVF
W/P75hG3p2Z80G/JP59uySqvE18sMlMlI66WK4QXd4RK+/xm0C0I3oBE6rzf6jAtIjFBEi2NKGIc
l1cHNDE2Y2updVbdhWnVF+R3qtfV0llDcLFTd1F49ROj1qhXke3sIqSmCUvqDuzWgmHgV9I+gt6B
O5ZXLL6lImam4DfkLQUVwyQlUA53qH191s6hzGu+34CizAJcYslry3ndy6RPooBPhW6rc63dRqMq
GqrzjFDkHMoyaF4SSqWasY5TGj39tTiFCADK/iGax+UjIqZ8CpcbID1t9Efb9ht9BjYY5Ch2d4oC
PGF02tsWKslMcO7W3LOkJ+1B1naHNfwdF7DlMfUikIoNRCLWjaRsA7lBRgxhqdYdUFNCxmFCuVzh
hAhdH5ss7A5keeTn7seTRgMsXex0j6GyB9Cu6z1jh9vg60tQnwc2jxIqC5bd+hVY3ZG07nQbXsI3
fhYY/4PCfBb1duKlFYr6DMIrjt8V1qKiOxSx7PzzZyqXgz7AirtdjlKBN9D/eJqMDNRBt1z2B7xL
o7RavBlkfUdRIHRF36slqMw1s871TyO5JkUjoacqiJwjishQGr2OJJ0A7qP58FbS7nblrE+PWbbs
R/i4vE6H6IR6xYr/Gm4JZV6d1ycRchmkmVpdLNCpsz+VpBYbiRKI3gjMN2+iwxaAgShA7Yxw0/ei
E3F0VjRsJA0csO0hYNABb0wtA3+k4c+3BB3oRoFaX+/VGBBzZ92Jz5HCThhZWSLQrGpMYReOoyev
hpJ6t6F/2EtpOtznNLEk23Xbn6HRY/nxkApN5NhynUcYEF1Ukb++C70KgapkVXb8uuccCamkHtP2
RjVEK0uCWS7e50DsWBPDyCGVtdx9GyrSWlLnMqMjgWeJYvsQv8pyoXPIJEvpIRlkuZQ6jOP/t7Zl
GF1oHWvFmVA159CGbEKdeBZ65EBJ2YuS5HqsGrfA54QJJDEkLikVF+hm8BLKl5s007sMxw9iinjy
eZUp11oQsAMlDbWxV6D0NLxmpMvfsGThT/0nx2K1Kp/CSdg1TjIBIMm4Bh27mV+x3jOnUECbt/qi
bHQlmLXisrfTnRuZUtpgufa/D5BSjtZJ8OYNAk/RLkQE/hB5OH7TbLPVDzotV+AMlouDrsW1qqWC
9JtfO2rfEuf+8RYV3cVSYXqCOmN/3lHkB2GSsK60CdTq65y7e6nesh4QEX4tTr3pu9Jc9g/I0DaI
9md8vrw0u2QxD4oqeU9bS7V1hPJZHIQE7/zVZASUC7UY0kHqaY5CnnYPnk+fTG+NKYurZToPncp7
h7lR5T8JK+Jg6PnwHNphsIxV/qdSm2IXWfMra/Y8QSvid2CuVRxdd6G/2KRsKrPwbkiKfpkb1fx7
t+spxo9uR40EvZfqtdwW87YCgKexmimioXxBwo7FIeLRGXkH9cQ8WqC7VHR9YhIgKMvgzeMmCT9j
WXdnKFSjY5xl6ch4MnVdmzNopFU7B5bRK1kaud1Yewd4GTZZ/KOPW5J+FuseTe2gDCfpnBK64glB
pFG4XTlwYSMtXX3+rGj/HqmK/SYm1VMt194EhoHENIoi614m/yWgbvZBrU6qnLav4q5Vp8zuEpVC
qpvFjGm4ZioAUeNtFNHkThVESjfz1eRVpySQUjyWeWU46C8nKWaqi8dfWigCxhs4uFBCLQw5QXvM
xywH55jgHubv/bvMzqX8DdrrApHFHH8fhOG7g+DdckUv/3pAJ9ODx/KTIkOoKENmJkwyGy4oYwxT
UhOMYHSUa/ZeL6vyBwwJTe4KYPrhbnxBHrfnTrWlw1ab/p5bNq6dS5ExjPAC12Pfm0X3spT3Mh2K
9LUJ1W3oZJoCIVzhmyQIbWY1Xf3iy5WFdeka291Fhb+ESm3nbFS1tmOMUYJk81HnBQZ1pgNXTHMu
Uxzs2PZpihpuRcyHcLYIrjWNafQAqPCJuBtJTQzGUXMQ3vZY76Y8GjnpxhYuVxI8pygtLGW09j/E
vL9fsAAFgsm9aVolLnBUm6+IXXF1OrybWX5IfIuPJUNTEXVFzEtPUdUrPuhw15Wuxck0REZGrWFY
wtetA7e47hHIX3V6JOhholMpqHC1OI2qbF1RNrOLu2UhhuVbLX/CVcqhF9g42gYelWZ/3JHWFQyT
L6lUdzW6f5/B6a3ijvJ2TU5LYX2EdM25HawkrrScnrV/uWDYhAXqm1pp8i1w8lMzlNOQbjU3rF4V
rkk49wawmcK91XuM9+L2hCYUjtqC/U5UHQ8m1Zr8NWOqd1eb75URLsdww3BzBGFLvRGs4BlSZYQf
A/F27ph8LrBd0mQoRjW6gYJ6XNm6cWYSZkY7oNRoTT8STYz+MYoHA+1i4YMNaH2S85s5wbarLVNc
VFHeoUu9yt8LkwSTkuV4kjSY8H6hq4ZfGCNAgUCNU3c9a/AnHDgjKMLdXvK1NBtXAYj97Nuw/X8B
444owTtYfO8U7XHMnRF3gOGw0Qn9qmrh5EtxMuRSaNK8B6WdlrBw/UFWsEku/pOR8Xqv679z28/E
x8rgarOAhDP5JPfo+D6kzd0jyN0mi4byfd8gNonJNYsv7VA7NBJ0t+5hrwRlYvrXf1WMGLZdclGJ
JuWBYzQ2xSTajmffTyKjM2SyIvO86XDXhduPRTYrwQpkmtFXnrOt66lW+vIDczlvd1ZMWTi2MHSI
2Bu0JhCUfImILpCnYsZMwC9rZyvQ3dhzZUcCdadlazfRjiMCVqYPmBoH53DbEsL8KvLCj06zL+NJ
nUxmXMHXn7qHjoDFmwOg7GsNb18+GF829YDHPew7SjQ6VycsFwCuQ+5kXcFIxS1DZYTRMuX/wuLd
+hsg/AMx68fWNYxa/GeFZtEEcoWgH7uzrreeALtotbN70vtWckIQvmmH1GaiMkDsVp/f5xHtgUTk
X6d8qnlFB4mZ0Vshpv5cmDxv3pfY55aveRFhO9DDb5tNIgolO2TD3QhILYBiqD4QBz88ZZtLwEHY
I7yrrtMwv0rxJWrOSyipVlKoI3XOHe/Wjay4K+Jpr5sSFJaSPGb6GwRhsqfex31XBkbkppnPxt09
3JDudz9BasNXA8QCeIgPTV23msk6w0J2oaB4KRvW1QZNNlwoqw/QsxKFePf56COLz2RiCsND3vsC
mcKtT419WhRfXKkU9GylKGQ9btuVhnODqszSv6zj+YpqB+d7sQKM+PWq9AZOwMvOSkjPXqksjR6A
J7r4Kmw2GZ54SNq1YgSzRCssenACC3P1w2+OKqkMiv7mSKtQnSV8R+gQd80Ekr6E9BxkcK5T0d3R
rfrYph1Qp0JIbmMiGUsjYstlSSfz/OEzDIg2a30Db0h3ug0/tSgBss7FZzntUvvlu2oa2vkjQRZB
9aSW4Tgb0mb89G9dc19CyhZJ/1vjSYB6G7mvoLOWXVMz+xCdMewRZjtYZSUq0Lh3f0uukUahmno7
5A1VZjiISPiC1p73uOSBgHNQoGNvIbCI5b4JyCYpUGm1CdtITeWbUwuduOryzjps18iJPQ/jLTlP
4rhzheJVPFBlvU5vST9onqZ3kQaQUHzVr/93O24LwtDtt7vcIYDTg4FvYpHmzV48WtVOPIVOeYKR
n3Rq2GU2yhKSmPxLa+Yqamo2iVpVS8nVSSCJW8pssWlkrg/aKgB2CaQV2q6awljGU++gFDQlkWNy
HtgIQF1/69D526CW9ZYKk1wV6YBnV+aetM/UpbtAYJ6N5pn4YRSFUHTXj3kBmb/5KTVsy7bFyFia
ZsfPKEzjBVK0INT55oUSmeH2DtfoU+qDfIzSmX7hNrzDrtmeYiRFE2LvD6s9qwSF2xsF7zhUDnC2
oZ+zS82UI7MOl5EclYbS28EWhselgxMt37D8J56Eupni8WkKGCb9mD8pkzUIQuqY0qNwo6zeJeHM
7u0dkiJhSngFy53kJ8/nkjeV6bIg4p5G4MVsweRwMqGr/snPIx6+PAw/AMwRR2zbxow+xxL93yFj
HALw9lJST6Pp6/UMOF5jzQfsNy9e1mD6qFMYMpyNlCPbpFK3VZfK17bJIfZV8MSDrYrOrdUs/ACr
dHLY55AhWGPaXJ7w6UwTzt/lNIbDD4kAzOLrHwnC1MYkWB8mD5FMKVyca3gAyqMeMiJ6GreFLUBx
E/gSYS/zjJKupfLOQTBObz4Csh7AascZ3r7e+z6IRAt63pHlYmKQrIakYilyp1+WZLJkWAcODhWa
MDod/AzifrepDXg8Py3VFb+UcPs4/jE2F+JRhC+euN5wetDbYi3HrbahBhUnSjAYNY3ZrhIHn9je
61/ZR+I3gDbPmY4ynDlf7YERtXcILirK59ayNo/LIpYD7bIzFrv+u73uvrPfEpJqmsDSXmiIJ4u7
UfC1620dPsmKcmDUWtFQceigxnP94aGR7Ojc2D8sltt5dHg0nWruafG5ctxBj2XiXq7ZcP/0reVV
dnQg0iy+/IhMlaYEYePRZQYh12XlGvOCmw0qJHa+5uRF9dXvBmxJerhDVXSGKR5xfJijLuHDxKGG
gopSj0QkbgnkjGepsQASOK0WCjnuXPm5ts+0tahuA0Gm0H3mWUZ72Fxp+hhNMfw9bSSPIq5SeKaD
1JHhkQmZBFCEP1GV+z0SDenEst9q51RwomJBwbqENneUkw+6N3EiMt+MECudQdjedPxLDJRD1Ver
Rc5KP1J1sCv4eFH7rn8oLG9jKVlNaoWYMa5A+kYD4S5SiyBJsW2HMK9I009ZPaTboOC5IffjKIKQ
A8NtAzfzKCymheFendZIt/dm5bqKaVGEZd/TKH9rwvUGbOwJn7JbpX1Ue/c2Pewh7kJmyJztnl8t
fEwRpo3O5cv8Hus/huuI0tzNXE418XNVKbraKcGboYCWL5TAKSi+ZxC/iAVcG+S2IhHHIU49IVE5
zYoLln8ggJChe6cdDlzpIN+FW2Odxcgpw7931kmztnAqrSjPR94uuywl9uSL9ZB6vug1oFhIF3J6
GY0sa2Qj7mOF0KN+q82HBpHSAT4s7Heg1dHPlCNJKJ/RPAFzAXKm0N9Wmez8nFKiwVukzqx5zHys
1u79zwK/NEtYxahieL1f+kxTfD3nON3Eve82BUaOJum9xP8OzgmEuOKF3Fl8GkESFpTQX9LvLuJP
3ns7e+5mBIVnE2hVqHPBzpgL0hy/sT0xrsDUNkAJA1D2KoAfI0awNQaIwYq4kVBWpfoBOXyruv0I
XWLyAYKdzgX0DEROLYZcYfCG27QubebLinUu4RO0+E3sgiNhU9CYzWJWthuvtLs7nWDfX+I1g33R
zajzG1HE8GJGKe87DBMCMW+Hre0U28lzaHX6xnNwK9bjRTTb+hARkjdpuqKKIf70idojkxdbMM4Y
jtNW/xzi4sbvdnd34qo9HW4f6C4Z/xi+rFz7FzJcgAsNLMb6W3/FbPQeBeV+P13jne/k2X4OtiJI
W7Liw2Y4yQgWr12HU0WziyMFizK43fJh/vg5/t7EGm72N7JsXdAffQcuIKvwRXsE3GlYofjWJqck
71RqM05BUDl7dbIYxppW+wEbBg8rSqKIrocuTNc0iX+vEkEFIcnrBx+e3Am6mv9L4ibGGttiftb4
gOiXX5vVynCFyDH9yUJWMmN05nby2e69YunWjtYIUEq9cPNGPesXR2sSrnAuDzN6HBZN3KQVs5Gt
4OmnGH9XMTm2MbHOb1z0+LlxcftsNWqzFMdhPbs0gnd+VGDYcAA26yKqaM5oUzPj3CpRBW1MA2nc
VVT/E//OvSiA35E/BMtiwccQ8S7Vd6/CLkpDMrRPooxD+B/EYAahYTM0Cd1Eot3zbfHAmpqsswAf
X6aWJ3c7oHqe/BF1t8Nj1T9M92AL79DVI5G13cWZq833igjdg9Cn2i0RbdDTTFVoSbawU8ikdP9J
DYGmZhZl4B0Zd3Is8pYu8alM8tof/XWnCTsW0jl+fEbdxx82NRRW4NNJNzbqf/yb9WmdRoOONDJD
8yVzs5lYCQM0aWwxVTKalRdT1ht6m7hAohc0IGjgSLHk6cK7D3zsgxPBe6LCrJ/gwFlDc1cXiq4z
Qy3cVFsor+d6O/al406v6ql2kgwsLMJ3cY+5Fsc73zBOEGilf+4hWMJDquolS5MYSOq7kijq/nT0
WUhhsHqMTjKQGynodteUi2ZsvAf3qeoPBsIkL1lidj4sdz+ferMKFfypwsbHSKs4yIv5Elpoalb2
NBYDfwztV8V7F9tP/KXzhhaohVPDY+qcQIZpexbKYM/OTxfFxsjy0odRX6p71gYMTv0O/+Bd+/e2
sF+l7j01DwMkT7WKNJdCb7Vq7tPuapWBIAHB4Ic3fW84v3feiRpLI7/itoET0+RSp9dek8i2qqaM
uOHsuVbArHvpoa1LhZG3qiurMHukSWamedGaHGXd6dHEs2o42yG3fKZ1BvFcqGjMd39BVBl2zjwB
W5WxvMCKm8KQJjV1FzGtmoOXSquDugdsyACUX4VjA3oIIKLRfxeeysqu6vRYHZ7hcff22qRbiFWk
u1fSxKufbH+d+vRfYFkQtZAY4RME6RJ7h5DS3yv4447oowopNNGUEBvxmFvltIIJDXvBPPzNDcaQ
JtlTP5bq+hCiN3rldlNl65CZqG3EBWlrEyhNFP4MU34iQLiacRAowT0JHrs6wBzJFizllzF4M2Uq
Lmfy98NOL2WBF7Vv/7SUTSFeEMmikar6iC64kkrvhH8Pl7YEdsM6P1PI4cSiicpKGhz+NFFfQreJ
bYyDE1v135nrjfFF5X8bQiCX/GHk6Pwn6sdhS6vhM/tm9vp1Vet+kNC5T/eZEh6HfuTgYV+R0lvj
oBa7pQ0wsERjBpgnDXTXIAqQHkiEa4OCvQVjDkYofmbqLTXJFeDwHF36L/KAgf/ndMOK+4GV0hcP
5hIeK3AM5woURnfxmWrrw85nyd62SwZ5QU3fO698bVSdJ7k+pHNeAdMwUkWpt1kKIOAJzydastT2
xGc6wzC9K28D4ebXJGI1pzBeTH+kq18QJuYd41zYTtP6bKMV9XcCeovHJjkle39xk02QY5YD7KMX
ahKR/R7yBb6Oavt7YzBqhcsckTIEtpmVHf8sx/UOceNp/ZpVMMys2DTGYUxgvbWLKWygcaEdLNaZ
R9hF85ZS/PNyOzM0+MO7dFLitAHJnI6qpc/ClvYYuEwoAlcyQCaAJ/Mmr/CJ/Sb5LqJzkeDxYhFI
m+wAg4tKgbgWVaPlGCRMTaNjBvzcObsC1+g/MkYryf/pces8MKNEBWtwuI84SOSH+b63I7cBnjoY
WL406EZzMcDhx7u1WFT3l4WWeTsN8bq/ITL4ouK0pGjqGpy6ukYqYh6OndntCWRRE4qqCLklBg3Y
+6PP++vnExkYyXTxe44KOQqpfZqFkWUTnnOe9n/zTtZ7k7yyz/xALdKhAEc4fVCsdloqiesrutSp
DX0WG4wYKscqc8YTYdIv1WMkqXy7QkNL+KJLmuH7W/teI09oCxHlX5CldqF7X0dVzVhtekAZU72L
BsB2tlvHOehmcW5BCes53nutYPKrRYKB1cQ3OWx0QFTQjZda48FRfm+kzyGXglVG95Qkl40PrWsM
01bjOwXoySpNKZN+W+W+3rzo/AmUQr2xEGXy7VngDCgf2er76rl4SsQTu+atl4Kw/xIxUXI0CCDv
JXB89z+4gcdusHW0rRzLHbQzlW5ihbu4kS0anwdGkcGHsBFWAY5f6NmxE377Wfl+96yPovg0E5Pa
+IrJL9UFjeaqbG9d+6Fo8Gx0zyoAgLhyfJNa9lWvqo7fj8HCrTStb1OB3WFlybGBajAuumsgCLNY
FxchVWqL6M5J3j+lgkn8TiStjkPVcNiF6WljRhxJbPeTuRcRAgQvHY2ZOoS+TP0uTW0moLcPc+H9
rFhFbn8rYU8NT0o0b4dUX2h2Y2ICOHKqHsNdXkPT0xxw/6APyHo0Up5vmvr34VuC2oIjDbYnHWPv
pkYPG/ieTLc+Q7GkTsTdtbT4RG3UM9JIgf9uS2fw4OjA8n8m5sQdcDAmxWDCc6EKlavgjamvJpGw
Xwo/VFcS3hlN0NwKVvwx8ddSMo5w3WU4zFXG1A+/JEjF78rLqZp5czm9+WOQ6F8Kxy7KiEFbcb/5
0++7aPBbMkLETfLRhOHLrN2kbrqSU3y5DfXc2gBN8iwzgZTxHHvvMeUcPCEIJNSXNqn0il1IEK1M
CfkgD+7GY6E38AKh/prq6kT4+Ujat/Y8drLippChQK1kyWvny+LqOB3tsNwGQayasscxDExdJjNj
YlbWP8bK8UaBT+gNHC1VooPulZlIQ5tU292LPw7f4GpbNU95pAVZF1ljtulelSRr7iDXdWrt3hIH
o3Y1jo+ilyeBmsvyNubTHCCuJhi/vNeXFEJ2Etf1WqX1yNTjBqjL9KzdSurBD7mOsdihQSsUKh36
X3ZFhVB40CidGLWoSdN3qb89+ASjCh+dSR8AqnJiG61cH2pFmwD1fZU0dMtC74+qHLJnaPzeFohw
RPMKKrm5X+tevLoEoRhB/9WjC7AuwH7uUjrZ1lJibD8g3i2DkKdmUa4YliyPNdgFDfB6SRFrujhk
p1deqJHjoHi+Mah227pmMHpv/sbgHMuU9guaadH4MRM5zR1IOKqz4arStijmaYKO9qcbBaifu7qJ
k/HISkUgQb5QSuDJ3c2kTFGnWa9DSQ5qCcrs8al1HRkUpZ3Lh7aKkMqY3ASokqpxzhCNUfcEPTqj
PRk7fVJ9mQOkExgTAgWbjLrEXnfN8+x3i3X8zGWqkRzjGxxFdPslWSlyh7v0zWADCUcedQIVv/XG
tubWrAjNrXU6qXX0opoIMijKtHBQ93nJZwYnFJTTg2Icl+n6ToDSZUHfW5LnG3aYOFHjpwdl1yJO
KQ349m7unXZ/Ov3UyvnPjAH2tToJ4Q/1nMF0eZT6yc2SApLuyXu42nV129FDLqpYQLqVNreZ2WxR
Q1Srfst3AuOzGitavHmV+JR2FXXtd/Fk86Xzoys2J52DMM1ssqHBokwqdPrka0ARpAenwoGv/V1D
3nIbzslH+WFw52GBLZJzAvEq03pYv1AY+hW01M3q2w8jQO5roggtrtpvGIwtIls17AIF7XNNOC2X
XugncycgM8VKV18xbZQC2sjDOvRFe/Qxr/zK9aiS7xB5PxX9nCPgEFXkLsU0KfH28A/5SKMxzbze
8SrBC41bCFuEBKERcZ+FOL0JqYfwH51g60Nb7fFSf00PU6gupGZBOdEN9rREtaGubVW8dnYWa+I+
8n771tgseAx0djgUBspxO8NvPRDs/B3Gqxpu+NkBEeTh+Sn+JqzVmiwpBEjE5OqJRTXGsVWOjowa
1/WAoLGK3mir2xc6lOL8XIlk83kPQ/SBEzj0dpBf6aFJHz6i5808RutmqYjhPMO2Tv08AlAJwM18
RZvSJDvy5G7X8z2Zdag1vBqaiimPGa1r1nhgCS4lomzrL/WpahS5+Bv65B1Yf5PGbK+QWo8m2Ibf
7qzD/w0+SWqFG5MjJHMSi1UbFA1KHG6VVFul3offhLgt5Ru/m7gdHbYCGSWii+7W0R/OIPn6IZ0V
erxf/fl40a3gw9USIrMVunogLVp/XG/wQIZh3G5v9TJXnfl2FJar2LvI/rEloXCl9N9Q+OamstlV
QwXV+hCt9ikw4Xr5iw4qsR4vI5R5i4lQON2xIugEvsztGkMosZtWiGaoZKTYi25GInvqu2Z+2FHY
dliUqHDFYLSp9firx6I2G/A269+CrQnau8hPQXmcAmHsEREhWcbRymJRpi1GWOn7H/8+9+oV2/Xt
StmteC6mFXgCq7vPvCx3OUV+U97/n++N7lso+hD+l48orQw47xgMGt3+eY3HHx1IhAjGscSWq1Ng
n7YPii1CSU2Mp4pq2lWBOe8P67FQC9lJk6l7/UgoQg+zBtPHUUPC3JlxR0f5gaLFhx7ZZg/hxPE/
AOfoVmpeFOt2fFM+J+5mlojGziNCYEuUhz7B9SZsevIKjEOD1SA828/AL0ul+uRsfpmHohXcnL2g
7a9mgqMd14ezlIoKriuoRv+KfM9xtYIdBnleX5gBaOyti/GfCVL6EYs+1HstrFXnadWGUSe/fQoI
QmOmAVQmj2L9xK3qc3nlLdlv0q6OH5QIB75l/5FYrTMgn+NBhyg1hbAlQGr9IjrfNIAncEaCLD1C
bTNzJ6xaCaAguM0JBtUR4t3bB3RqvmOoy6+zObXXEa0oq3+oh+Ip1OAT4Ft+kxwlZjcGlyVezj7b
fNLMk5LxsqM9RSvCYz+OudGbkSuIdpkZcF5tQqFa9I3wUcZe2eLWyzEB+HI9V7zhueNuWnhtqEHf
FCjOa3pCzjFfjuqbFTy9UUX7XhKegsbh2DtRMozzjUkKlhLJWumi+c+l1GI4Rh7tzAkHVghVpYlk
HPuYl+xA+cws37IVj7RVFZBWUiPHvDQiCqjAcEDwYI0h+1nk/dRZ9Pm5gMT2hq5BFGFr5uEG9EZ9
0wkoYFWhiI5pX4C+bPocLj7HvZvcg1OXXoJfZWlop+Bw9kaBLfxO7n/8DoLUwGz6SNfPlqTgVgt8
tdDJNsBuT1ZnHPnw48dZ5TJ7SjXczA0QLaDcdfTNl4ZZlw/OMDHJtPtYSnr+2BYZ2oM+T4Ert69r
Zhfq5Z+6HyrWBCQ/4yJv7+MdI6PMjWcpv2NfUtq+7oLuEl2hfOKBtq79yT+OTrqAf/TK82ruEvCB
MLWJbjD6ss8XHaa/V+V11uC/WV2uj9m46pSa+0s+6Ht4t/H0kF+8hkbTn6yUfE/ZmHitTJuxZ5l8
5p3AAqDxPKi/uSrxj0EobbFihS043FhGqndUUlxx3ytEvbQWyTh+jv3DMS+mYrXogti0rsSBn1Up
VhKbMUyVVy/DCia3l6RLf3MCTPMBfG9kme6+QIXG2WpFNdkqlkNarUcUEwMc6KePVDTBy99wJH4C
DKOLqpATrG8gw6BPw5bNwNTevadMXMK5g5NZof0eY4ASgVjdUj0GmlmPhk+W1GYB4GTwvooYwZ5c
3v8ze1pNgUO/rRbY7gt8LTO9+v8C2IMxWYQXplEwtTGelGk8GRtqw3DWfztNkd54Er7mCAHzBdI/
ttiXh4hHhKaoGruTIIfOI6TqCCZaSztbvtjgP0K4FxiVShLs1O94Zwg0Jtb/d9hGZHoBwN1QOY3w
k2BM4j+NqJ8ZMHuBiaaHPdtjl9PytiSqVtbJ8BF+oxwp5Vd03934FOmxQGBx6syV2kAQSayJP5bK
JrAkqNuhxWKl31AQVjuTPLZgboJ5lFvLXct8TMouh6UKxo1ZU7i0X1FsDJLqZ5LMoqGQkVVwYc8A
v/R3aloPfMvT3lPh20CA9QjyflrJwE8jj4JlBhCKCZNZ8HGMMhLGqkup6ryIdA7S7aZoW1rkhAUI
eIHIlEUrGsnO2CKXwAiQYzV4I+azKim8OZ4vtJyxvSRXxqI6bpXdxDwbbc9jNVRPW80G+lGV3FvR
UzD7DHHuc7oND4t+qMBhULF9b06ROIFRyPVVQWMOpapzL6PVFdWKnFFta6z96E8iryraGULpRgOB
r05Bv4mBiCZlfcQoKQ7SVdDjoYwOcRWaBiEGpoicN7HJVNKPYnMXMnQfLXlFH+T+dySiWQMRnKMs
CbT7MFgZV7B4+kyyhRH6lWvqzVHDvsLK4pxJeHhZEswGM+6GX8BIpIgKxyyxO3lr86PhnnA3f3c3
9NbJoZPBG5/zs29TAm9ioZPbLvlNwkDE9CuPL45QlWuchlJS1P6WiKnCD/ovZcdUkXS5VwIIiRRK
GsCuiAyIZjCsfym4JTuifVGWc/zIWgCHqx3uJsftx1frkBZ8A8Y1/Waptl4DnL6NoWaVz0amgTEs
UZ/+yUqzYHxzLRM48kcg5cftM0Vl4qcCrNUbiQh3O7QVpVQSr0tbruY0yj2DW9eR2JS6zFw3yGP9
OFNFavbFVshnbCLjFlPASTiMG5ovMg1UCBO8SbdffJiGBA2PJGCNYTH/3bSiNBEPcp90/SQgzmOj
mGoJdajuDYTcyekkt8pBCzWE7vNSFzmrsDLAhWFQVhRQnSULwHJ720OiNK+6lxz46ieYkEFTHCSC
NYwGFegC/uvNeJwe41ZWusbp7H/GWTC4WQzr42Qv5GCLUwHJKkZnvZe5Za4z6g+6nKsrfzHyqX1H
9i36jZtA3GU1tIfMmQkHGNbJ7TUM7haSwpnM2DVcdPXkz9I3R/vXA6bxylSKC1Z1ol4IHxqLlLI8
R12rfqoWepwH7MWAASriGeIS8DVssPf8i07eGTXVj22XkS4EyhoSfAipHS3yofCNcRHc5ymufDXS
w4cxJGEKs+h9aqhsLE4cJ2Qzuc7uZaf3DyqCvKtqQtcrE0SrU3wEd5es3FoWhebRbYwg6+DmZhrJ
aQuC7o15eYdAFrsjc9P7EQ8dzAPG7t6VOoVg8R5n2pU7IVQajA9A0ddsjKGU5yGiDbhye8edWHD7
dsmw1JeqbFx3YokkMxjcZnCwkIEQqRcCK2VmnkeNVlPQvcA468C1vjVjo3KnI9DaW59Zv6VxEfH/
GEiJ+mdD6wtGwq8FiRZakwAOSjqPd7awnM7PxQhz38/UiQJMWXyqtU+1VRw4reZB9pBr2OoR5NkM
tOVG1dpjgYoVK8FLBq7ydkh4PHW5RQPmPsj78UDBY91vVhOD/txun3Gm1AAT2PgZ2zm+F6m2+Kr8
mWTvu9pwltW5VQ5hf6coaxBdp7pAVLEGIOCdZv8gKnwqbsRJSnvFJ/MFZ5P6x786q7vJJnlAysPc
isd/WvCpkVzPN9OpVuClugOB/wlx4rwLhx8P/xdRyA+/mLv9SJl9mO/HlDQbX72kl/fY4qAeLKJN
7xPyEcZVD3dd2Dh31P5yG/K3sBM7udUHTkj+nNdnST7IZORlbdd9sWZXmk+neU/3ufWlADOh1t57
KOWGTZn9O3L6iw1n8F/sDC+Sw7tceKvclSdIua6j6FLcSYq8ibGPBDw7qNOjEOjpy8Xv7Wf6bHeQ
G3NrHEMe8RPIWduI28cu5AwC+ajDPJWLLVw5hdfJ1I9ow0RTabBTmJIToo51ebNxgbqdaCb9W65T
yCFOvlsfrjC+WtBM0WZzVr9cuYhx4oo3UTGSRWt9RdDwa8Y7lwn6jaZOOKnBg0obL9JkVrleayMj
83d+Fhyweqi61J4yuJgneNEmaK0ZdDDKCxRcGneGmI/+/+Z1PYHfPB0+1PjjtDhLGTk2vTx5yPhX
y8+DhB7afm0K+kcGN2fRK/VACD5b1tD4U7Z0+aYW0QPGp3jZkXCjIaBjRbRPS7detajMuu7XlCsZ
09ZVk3bK1epK6cTO2h4jXFd77xyxo7gc3SRbMM7wrobNSHfHdYp+75/bAMX+Oy9B9G5xbc3YgJ2U
ohaz1Sd1Q6x+DZoPkjG3S9QAKQ4YwoeMoj6PTyvU8NRtShYEj9eRlXGiYs/wndtUtCdIuZL41d0O
geL6pu7pPzHrAUSA+X6u2GsZufAJUMzE1ARs/DFNpGqfibL5KwsP8FacxAen8mG+W2HwLXHY6yUk
behBgWqLSCqrVVeATM45rA9fbO1be8IAZaN7oJOG3I1Mx6m+Xao1vK1wV7SsJj19NxsG3SLwxxVH
tsNnEhJC4OKz1KwR8pI1jQ1m6zEtsq0pLB9kfv9GZqqiwV4kvIB4b9taXXjZPIB4OKqXqsoU9YNU
0mSZvEymC2f5uybCnZnNYclsp8bYZ1JK0FYxpDlzXCfnJJ0+NXXJHwQ+XkYt0l21kZeMIVMJBaei
wXG0iXwDn5r6EBYi5duMWzopdt/2xG20IpfHGJBL+sTbeSePfo5E6C/sPxD/CG9ogXDPfA0Ri9i1
1lceHVOxIW8pSr1klKLfrfQVTjHP1LKuRdQcdK3GX29AGSFELpWYm6BUZvlkUz8P2a966TSskqvg
PPDL+lj76rRputMALCfil269bmf5MtL4zHI1cW4Xsoo2fbSMOZrEeccm92AI7coqx15iVxALHRK2
JLseQ73DMNMgwmIgTFRdkZI7x5qu161rv6skLFydaF8uaaUBA/f4wRvburWFiEKAy88K0sCYKOzC
aOGfZQTLCAyXLH2uzjK++PYFNd677JhI1mHr53qs1cvP874hPKPJffgtS2mQ/SmPGdRD6bgADJSc
D/M2mze//g/lp+jvPEWNFzqYX/3H2HgcTETDUSh4xSuvsAU0HKjA3Pf9objcrJWj15K1i62CHtff
DTVhVZfEHNNe3/7VGUvUzaNaSshC/Nw1RKXFERPP1za1AhrxzcUURq+UbYuqIzKLA0tbzNIw4/oG
S6meWO8TROk+/4ENjjeGJqNb5BCKMRXVzD2usMUaDGvmUB7C+TApB3iWdD8Mg+CUld6/W1ijmTY0
LY8J6ACwaUhYvQYkVkYwkfkBzjSYW9CbBOf6sryb/nlXOpKim/FdOoe1y4xiDJJ2DB/oKP1+eOWo
S08PTHk2wG61anR9RFOAxZDUiAiHAFAMfVal2KXfvhmHXsuLbneIqWNrtW2kr+sfh9y3HaliUk/9
uuBXHraq6LV5R65zylUGnU9Cuse+AMFW5ZYNs9Wm7pLay7wg1w17IPF0W8nhdInNyFVGo7cuI0A6
MYtpLT8DwQbCN+K3riVmQ9JuqispkE0Or4GYlEScVgqEAM3kgq5qlK3fftruyWeKIDGrD5vi2/QP
6ludGTGAbrYRgJZ78h3BpgAkEo28AYe9kpQMNh5iT+0I62SZGHYFr9x4vKCGVKsXOTgkCOGbYjrB
x8dYcn13zbDDbJST/jd+yGP5NfM1sJY0BoIlQooMH4Dy9XchlVUs6JRsBB9jftk1nCANaQyuv3/W
LQES3SFwjv33rJPtPIG81H0BuYMZyNMhgnGIIpQSzX6ZUwvgD8tnbD9u0gs4lsyvmCNFUdtkCbXf
rKct4eGhKBfviG5W9KB5QUTrg87nwCIZY+mOiTaa3Brh/cMSbuNl/N+OkKBd2/VCQ32ABQNaFxdz
N1oPrcLm2DD7BBh/ktJTKSBkKhCbSl0pX2cNRfr5iTNclYlOp8GyPooxz38LtCPIJCWlep0nXO2I
T7d5epy7VUr9D3nr39D1fZXyTbPxo7AmvS1f86BdD7kz2+e1njdFVNC3Y7yfipPMxmU7tVRBiQlX
Fva706hBluL5dsz34mj//RcdPcWYlNzEl7z2cLU3xyAfXupwJXI3ThaSFJaroxmv22TVGMBfjAmk
G3OlbgiQAiBFNj/hkxkmZfxTPiJoMfbNRLndig6A9ozBqGjsQQm9hl2duYCQ+zC3uYLksWWYodjH
ZkK5ZoJKz7jAeGR6MdsjEByPJnyFlIMqIMuP+qD6Q8z/IElDDu0WyCSaNc7PTOjm5C8/1ZHDGKQr
JZUn83aIxcXSIKAEAezyBARKSRFN6MXnfp3du0OIDJLuMyWnrgAo7cjVIE/5BL3dT9tIKJSUw/gj
Gk9sco37xID/wKAgqUW5YwfqbVPfnMq9NBXrKbxGKJ11k092BCxfJheaOYMTDrdyT1BpVwaNH1+Q
FSpInW5bltvayGwwKxtkpymWzMpqnpUDOaI7cZIJZHR6YyPxSVLyPnPVK044HU0Q61acHibaiQXq
SIJmPPgtIN16yT/WnAgA9PaDgrHW75Krj4+ObniKKrDI1/AV3e3InEP7hTrschS8e86J7ANQ/d1y
dotPvnycVINc+LPI+B5BAXkKdpJHW/L9ySDeLlnanMWG34hjZDRtQtSPi/8m4SsTnWOhgs9YrIgk
99cIFaTpBBzBjXOvTMqvIrkt/NQ7j90NLocNqEfobERrRqxYqyJEeyInXKjYvcbEbacjqrAaTH3r
5WhnnDRNHhfcujz6+ZiDvjhgykMpLVo37sQHrmxGQyW4XSqoByNVsj2mli0CPkCB/hnjA5abRn/y
T5RALGQiLuhmgEGNkYIwAbTlkpDUzaZr3PuPxLUE700Vafxd3uqdHhA82aG1+/ef9f6dRXB+lL7Y
ErGaxYZEA1gLo7DuNGOYsXl/EUJQ639ZOc9o3tEU+SNYrmVNhfCGjyVKtwHbxXpVp36x66pd7cO/
6dKclpFjkh+ajGvBO3hipqEk7ywCPbGu3jMiJwWa5RXDDzIKw3ZaJ2Apxg4DH57WTEdD7Wy5JDxL
FBngjP0g9ZXoM0LGZCRhAb2ItuWvSpMeQadjy5AyitAv68BP3izlKbklK3wxgG/Fmvdl6Z6lpYuR
5efjR36aARIvylucrnoUWg4f+c/Zcggtsb9dLv3uETJHol+gi9PUx4g1Nreq9PozPV5RAl3Q6IlC
Fg/lJSEdYj9jGMpDhBiNsX+u4AafXGcIfkIHX/7TfTg6XpqJxtEemN/t0SlQDIE4/yAl5dhNQoOr
3ngUuIYfyfDvlD5DrV/d3wwwRUaLh8NwdkXVACjWu0ohmuAnrWW+NoX+AeEXCofMmVmKpNylzLOc
Sz4CUP80192iXoLCdnbzf4gyH2Qk8ZatwzQEG65T+npvr5EA+EDxtL20IKsIz+cO31THGt+Pz57y
TqBnmc7Q0eDLkiIcMynZuJPzZ2zmsIusk/l5mKkZLK5ii8nsWBKrc3FPfIJDa18qFf8L2DqyZJRF
GTlYg7hRgSJSHSywDo0Bh98TCK61m44HNZSY+EfZNPQJLOYpiGNxJ/zljEe/9AEtHctSbONRrAq/
3U80qiQGRVI0iQz7+voe44VGMs8bb3jebQWequEgiBnSSFl0CtGpKsZRinNAqUPUUTaeYBgKWhV6
sm9d3NiDBjEsy7WabeSOOtRUotXSzfCd4oAtbzngMny1QkZMgpsMa5ipEywoFlZf67ebDYXn4qz/
lnZWx9p556MG5s9u8lwlLIMdSWtpBBr7mXXEf7aa8Ly47lkvvgRX+La0oqO9N8f1QOGYQFhwdXJC
zUl3nyj+ptjK3TtRZQEjWctEdabwZ8QgaLX70jaIKXf2sbVkR7Mm9u0LXunCVxEQQnRqkNDEOypC
wlZHxLaPSqDbswbKQDZIHaKn8eR4vhGn6Pm+aO8z0z7D1x3ukRdfca9+CeZUHC/ThLP9JHmLA12E
tQ+PeZR7RoaSVfFXP5MUiEeFlna0E0MU8qq1QhFH7SLqeWDBbp8Snz7xbFi1bP748krui4nwnxtc
bfa6EqHrnXNesatEY4kaBxxp2N6vDDw13z6sKQ0GqRDu5+4apd75xOU6ZIHuWuuL6yE/i7fYrubs
HpFHeot+azByUPUjXItVmb+VK6Vs+l3SgN4boGYQhI+SCfnOBaKBU71HeSqFXFKT6Glz/Y7pG+en
lfV+bA96MUwfkdTyvHi09TE8LKL/qRKVitTPz6Gyb7V2nEXQ8GR8DvCr1f46rIHCBUeszR/r4kT2
Ixmsm5lIRQbmbdwL+frjiFkQmLMX3Bm1qVVI5wtm3XkhvEjTPAWguxoCVanhQYW4iAEfWUm5khvt
WzjH3UXDr0vSIjVERBkPlw65avtxFxX9vSb5X3sW7LsmSx7ywkH8bnAnzJrJS1AkohmaLJreQmdO
Gb+v8mcC3u46iMGekke9lbKmd0/DvCelJI3ywnXCARdAUPfsik2qLW31k7ZsLnoBXP1UISZTmdlu
ATNp+tBe9IyYb440HlZwkseDTGRY0GC+DBGg63PS0b/3U9o+x1QKuzFTGSkvddwN9mS11yPBAVhO
7HOVvuKX1Xj88+yJcYl2uF409GjkIxULCzfn5SUvyuaxRxlDpGfJWVPMWwY+bOZc1HlG3xCKqI0O
IiW+4bL9FDN65UGqn8MNi09zflEN1cIJRN4pmbA9fjlNVR+7GK0JspfL3pf0NMf7CUjcVKP0G3pU
10J4D/V317hn1UExAGHZpOuEAwe7qE9XmxmIWQeLuQFBXGlqGzZJK09UlEcFCeEoJq6lZTtnCpiK
I5eqZWdSx1MYwc24iLMRhv11S43kEAyTWUGMl8c8nSExYyIz7qJZOHAn+TSHPCzvJ24x+D1fnI6c
sIePPGecoMg8JzsQOR2WIv4IPiWLsJ33L90X03i6gRaZkKVRLsG8SmVRmJA2oucgzLgR9/5Swiav
Yk0/VBIqEgr1DLeZqpfvc0uqCLpMJN6NOmfFEYmmwH5KVqTe7Hjpb0ZYsmP9Kqf3x9ouq+/zAOED
Uf2KlICMYY+Vlh0beoF1uB6azK2f8FQUBF9n0O2CubijVuOtBHyM7XopnZZ+JKptdAaM8T0Ca4HJ
56VBq5AOYd7LihaVzypV909vJESICCumoh0d3e7v58gbyE5JPvdQ6Ogjor91KWESCBYwVqDlP4Au
Tc9p+ukqXhId65DbqsI1N7DVe5IccMDnYzJECdHRXDy2GUYwkdXp4DjDRLEt7rUy4ZatrIrWMkTK
EL4uzuIBlQ63yu1CO3Ww6StOfKPSdINDYtpB9qxOaZ9FSQJ+BKautB9mJ+2yVswJndvpPp7IWXI8
+blj4jCdR29M+UiyJMju3+Z2SFr8WUkHu0j6f55TKfpx9poQmbrpGGZeClLdpGHh6X6eYdf4AZ+q
c7/168qyG0XRevqYzOLDxRxlGOyEI7wOsOLPskCXzn7B42Y3XELGviNVtLxNyWRp4LhbgspG1BYU
4CE8meRjRQc0a9CFJ0sSP7TRJWW6oZDjfdwX7mXwFQHobSXFa8C45wJfGaKKUrFQqF2ZeUwGO8Y5
h73l3PJVFINqNHP9yTs87ukahJtfNGf9cB1MwWj30ICOsRz+LD3zw9uy2sxJCZvOfXm6CQe8Ss8j
CURl3s5Tx53w7kzpgasJBc/v07/LnI6FTl4b9+X1ucmt6XSDaDE5eOXAdEfmHOeYC917g/UdejSV
AfoecRwFKx/RRq4UYwwP2Epdm7L/UERcPd1zNf1Q1JTCfl5E3HMhGtuMPvaDZNkyyK54k9HK+FYZ
LEsF2pjpQ4C7VfbNTWeAQteTxReArJFFHpj+Upb4SV4RVMQKM8hQAsLg5y/AUPYS0q+nB12mjP3d
7pS7bTRoo2iSzXNrB3qn6LxaXZ10oQp4ay2yNzh43Wuayos4F3ONa7IyQtD3RXYNlvgisvE+efJh
Z6kaJoNOUEP6P5B+PVgHgCR0kUAsUZrkSKG459Wx7sU53IK5aV8vVwMDIeQStrjbvp6bBagU6CbW
DpW9eXo2jKXLjA8AXVzTFbofNBUNfuFzbEs/z94XG5vzRjCLH8tzPQdjsVqhmdPRO0Dd7zJvWHZj
qPXvaEOQDemQZD2vhZXZboC5dfuJ5LwLOBY1AtMnJldiJe9FYJZVoOA43pTE2WeunT7MEpCsCigA
XglNm3F6r/pwhyfDQw4Cz7QQEVJPwJV63xabnYItgFk2YMVdhBwth5naXKtLvvSigHVygTP0LXMH
bpVcnzjLTt5OP62mSQV+dggy5jfGXmBGFqRSleBCf0NyegU5FUYCfDXQLTFrrIfZrEf6rIUgSWhq
bNGvblsrA88LTQ1q3aYXfGDSLhJPdeKGEUTn7FKmHRrGnjgg8btQX7XS8yBJJPfAPjbJZiLLEMh9
iBP2FjqgoUNCh38kilzpKYTylld+EHFOLtygUGNxurDik88R6sjF0zsOnfaHzqGjK0meJwb8UVQd
koKVkUHwOK1DOImBvxVYL7Ee169bsHhnN4WfLsGy0FmKJuxS++QOxXIV0JhbJqruoDBLM8Vkl1z8
MCh18JXhn8eOEuavNdnK18fpHBqvCjlG2JtNAVlv10L5daTVKfEIH3TyfZIqSszj8KMjbV04Iubo
yBAzt324tw3xKb94pmqHyHo5Wb0LpIw4gLYcJc7/7IdpvJbB+Whtt6xnK8hyX1I95McprJKleFku
Y3Qj8YUKxNmfxngqLq4c60lKMsjOd13TZh566ja0EnE4dFFTJ4mFgz83P7EiXY4ykKn9VTtIqkXg
7sdxifbxKnLyWR7tDAYt7HPLUIFpPvAzgRgSjEnTpYNIOtodJWsjxFl9vIhmpx/5zyVmBWwKjfhG
/fmQ5iFWuwMhZ+RdlD2fFBLnrZAiNoHdIfu5+bEtivlU+JjG4UsDyHcF8KGBdr9qAKvBPQJYVLDG
39u+e/WFCBTccViF+4zOfOcw39lUjbKfkb30fe8f5/dhpGmmN6cu5l+Q41yz+eIAtI2/Jaxyt6eT
YoFRgdKDPGlioxbv+5Dkd1fOPsJ8Ot9O4BDN1lX66D3XF5rJdg56iDjdw4D2KDFwgEdLZ48xhyBy
53iubOhxSS3IrIahXImeez/ltcczGRzlCwEr1VgHL7dDAV9AjmKmHz5rBmSv72qbERhNkBCCIR4Q
6rfdXh3sM6OU58CJhG7yaJWXSQq/1h4PXusMIafztxKQ1FY/1wov3a4/eJn4Pmo6oBBFKys4eNnZ
JaIWarNIzSMBP15X1T+1eUKLjquMBtc3SuDeWNQ609/g9Fz+HjqF5XidcXukZfK0AV1UfeDxp/gT
VLZ5fNrWzREEMfx3G0jYNv8eRPO8I+mjD6ctwXxPBU+oDkOQ/syGfBb7fMMmGjnH6Ljw+FZGs7j4
1jzIsgCPgA4LmLqbR7LkGN9CfIvdrmsK4d+SmpJBQLZtRqx/M+G00jVXZYt2O5dhnQWldlTfnyyV
SE0btECyBcn0ZldL3IzefE853GbaKxymzclTqH+eGxewQBSGmhOsxEJkOskdY850POMxeyne5s1W
Z7dkuKYmIeIOn9l+Iu5+R7bFeS6sWDqo2uozoHwqkpSLHCA3cYBeeBoHh3DRQ7eQ1b5Y/rqRUFFu
8+doSoqG0Meb4jjPWlLsfk8wpG+dEhW+KK2o1tBbbY6X7R8/nUoV3gDI2lJi0PhWngiFJxQKqb1t
Vb7VztypVzx3E/QxCjCbQSG3Q5old4ibvcOX9B4Ki/dOqSz0v3RfBbWjK/HWehGbSihN+hxSsxac
1B7JLjlZrDa0QtQmCFhoa31qcrx1zUe0EI5smIshXUSOCiQexGat1oZ5/+GfLgu0Lzs/ks8uT9ST
kSJ6dmHt1OgT8J6tvtIsGaWXbFXNkHtU1pZvMNhZVB+iXOowAQPnSwxhu1bmysTRWCO017EVbUcv
DkMcZnAh9dMmqv6T/rk0Qmc0MYpyIzm7QP7BZyKkaboeUzHGnljbJfRZOWrjFkiBH5HBki5oHI4i
rr+hAHG+LQLo+qwUqtf8Zj0HV2Bq44ePGvZGtzkCNH6XvNcMIK3b/sgoTKAIbJwOBlvBuXxrWSaH
c2G3XwQR/5j9Qy28By6NavRsu+wEK95n/gluR5dXVRk+XYKSfram+Wby0z5ECzIN5byw4bLogzWG
uWEr+C/JdaZXlE/0UdfK2dG+y+YVYCiuxMk71xfxmagQezf60bT68EgE0eAOnf9+Za0TjAXsGGyt
+LIXawBPWo+Ygn6Mn4/1m/HUY3Sw3UyaC+bGRo9j0/VSUX5wHjLEZmouP5fDz7Q/fkQqkNPd7ZkT
o1FYHExKoJstGxwxNGxZdzsfR/21V2scmoRcSeQluarFK52TLYEj48fHp0f1yeYevny8Y4BpvltQ
yNjknrcu7elm6QLNakPApHTyqgefNFl3N+Sq2vR5ML5lu8ODBTkLikcVGDp55mxTsfJF+/BEpfT3
4NGDykeYth01da5nE8YfyxJmisaiMXMyrd500AfI87TNVpHY8IUM/p6GWTk8AqAlYrGbhwpFMU+8
TpCOklunJ2UapFVe9phQFFdl/KOjuNMA09ICyzXesEz6GyvkNwgSf3Sbu1hf1xUNt6P/QkuEcokT
d/nXuEluAOhlqjzGF6um0WpqS08lcbgYkisIaJxgkpZWtFPPk90bQRfvkvMmkocZWoFM9lA/Moxf
OjmHKNDgM5h59RP/4DMvokEmrSfiqJ653QPlWLxX2tmUt2cOkmHyiT+VZHUGkOHIltf6X2l4Mu2I
37nNDMfto8VAzTSGbmoHjpFzApXL8E8O3vYXnX/4tSApsADHkeZWve49b7n99WIGqQLVlkIRb5rG
XPudgC92qqNdUypZ0B/9jIBcLuvPyPlUjMVDJcxk4gontIb4uMNxWQkK/zhMlDfRtjUj7lF7q0iQ
FIoD1XYIeIETrw7GusyXqhJ4o+pdG5HydllVgYuD0oJEg34RrnETWW1cpGYp9slx+GFBcntcbsN/
yK9TMZCLBnAhyPmWK62VBtjaGrXPjj888Shgmik4vS1S+cgMzqqQUx3zN0RHE87VenCKHpxmOi46
7edlsJ6h/EdOV+06npJbOOlYexj0JCIUnvS9HMwTiGUDo81o8T2SKpCkAmjrYaZtCBnakF6jhqAi
D5bObYp3Dn+ImhGBIqF5KJrBy2mfeU90turYwd2tUgK7wEd+buJ4VFE6WvaqDkkGXppjmszYOEhG
lneAK8vh5rbOgC6c8crQ3F6jEUYHwig42qnXcaL/JwpXxpOrQuPmG+jo+VWN9W7ek6Pm1GgssK7N
X0UWn2iDOJFSJFAP1pvA3QMXTIrb9ff2/I/yHlQtoE66bRnG1FZil2KyPYiLI/oCr+nIE7Kr2Rct
42POX4iyA2xWpN0cj5c49NadxD2DnyS6EApvtA+G9M/vT+YB0bUGeDNzK3+8+WqBmlwSvFHTF4UB
JQxBjFFxXljalOqinFhEcVl0o2bw+zSYHcFs3hNx83xOm87/OjsrBev8o295PKoiUwPFip22RmYK
PGi8bpi3oDrXOg8QprdKKHB5CPEhJdGStq4g8AU2Bs9ykT/uv5t5eYimOk7nHm8bXh+sXFmu5FXL
zJOqwWIauI2CeKNWfLyKnXeEYbbOX0O/UdqqwbsbtiHcqrM3dfR9SDVZbpJ0XUJCP4vyxQ1CTY4A
vnVaI1N0KosMETjzzayiLWzq+/z73fl21gjHKuwyH7ARnpaL60eE2aNcAX4djA3ZZVxzivztfSnF
PPbK6IZTw0isEdHeM8q26VgIc30bYHV4ev96wduKJnSK63fQN2l94yCyUMKm5xvxMDktyEWVsNoG
sDmRR9er1knJhzxinF2nk8icvTfbqdQY7FR9MixxXCbOaGD6qLP2a7jQwWxwl/CAE/XkygQWSU7B
DRrfDemapUDroSjby7TFu2stTrdXrlzJAub1U4Ke9+8ZcySG7JtABt0BYK+rxInFyKTtgFKu3Jul
7JiGUiP1psfM/FeqeMlHEvMphw0H8qRK+8qes7l2l/ucmgA2ENaRpKOLmrYBclAymx+Wn5jtdMR4
7WdpsEs+272tE1sdSUigz02EccXFmouTu3YAG6aPnCOxv6xa79ooh2AxkhVqtb6ljyTDpFyMsxwD
Jh91l3kktVPz8TQ/DhSUCQTIvpmD9UKjz/k70/8Kt73y+b/w9QSp/Bk2jB7N/+INnom6FzMyDFg8
rI3C3iVF1/s/b7TTw2YM7QVzv4T4fUV5l8Yv1QTBnBxWav4JIiYF/UJcmx/JLPB+wmdU0+jPCmXE
CaWOagW5dmnXpGk7fCpV5IYxxqWMVDf3eGFd3bkgnLXkA4Pyen1jdmbCtGiRgo9vKwdxniCtSLph
7LQFNjSd5AHzpVOK2gxh8Na+UlatQZ09S/+wRk/ohcm1MQ1cAQht3/Oe+Euo2CmGIAIopDBbHsnr
9WVyqOaFz3SCChgyoVGY1TxXDRPEyw3GUxWBYiCHr/Mvz3kcx7McvSe8alIlxWf4bpW9W3JxdIxD
erl3nqGBxo66KFRL5rKUe12EcDleYMuhWLncT4b5fTwzb6a9LZ3nlnusmlss+socHyje59FD2NnU
lqbmAMC4KnZcpzyGe8nMACtVSsuOji30qlKR0hXmaeb0gIl0lTPmytVNsytbVIXGOw89HcHGQ1yr
yAW/sqZ0BxVUTsUN7/eTIDLq4A6b7ffD1mhYBR7mGxsxSyiC6yHlXDqyZkg7NSAB5XsViju0ICPE
J9SUGsvQGuBz/RoAHCiPH4kOCKtgIDgOL2iQTL4kwaPGoCOpM0cgNOuWAwYIrVuO8BFti0nSkhLz
F0oWy7EQtL07Y6rnlEaPldKWiMVTWY/UMo4Nvu1kkYMMsE1tvvjM6ALKY8V7Qbh/NHLa0vKneqMK
hyyn9uTpIIutt1zCSTljdIv64DXmm9N4pIza28aQQbWiQV9t1sJZ0wnZ0NjZt9Oh8ADyh6FLreh8
+JuVn/s8eL9t7Tmavi4OoRaU52KY/m5HXzdQpf5Sn3IDtexdW0sj9ivofXMGk5yEuud8OneKiHby
wSiNOuLdn8Y15FzJ9h6vWoXZgDoJ7iCRhIxLfcEFtDmIuQFYETMOQm6z29e+/hWDSe1IOtrTkvqL
ygUEtkC1eyiF7b4ZKj7MYbm5hOfKUepZodgGxQ7+Yf0SKaifZU9llBR3tAh+Pabi9LlPq25n2Fc2
stehpPKOZvmI0MBfl2aU1T4b5qoUNPI813Ar0Ocjt6IPdTABzXhONK7TdLbJrcG1yV+0jHj6A175
eQzV2mOto6KpQCrY8MfydwZX+KsCklU96OpvRgmxQ20ugi3Yowo3yOJpSxAXE3U4+14VDC+BgSaf
nnvgKEUZeYfe/wPLNGPjfcXeg9S6d9IFGSh7+5CV8BNmANfdtj8JOKESztZVStDDM+BwEdHSKidJ
oBrIzfrofjsXG9zk4zHjfKceTnhXKNkJP0Oq2dmDUNO5qoJAThEsLaTOW2S4F3KydZC9kj435oG3
c3Oq13D3piVTe5R89q0Bp3/uo+aoIQcXHnVtIhsUYYJtjlHU1Ezjly7wBGVrMbm+EbqT9iNGkzeU
ForPWda5EhPsItSJMlOEnE2bXF7FnhwOnZsUEz19UoAOq25I0gjQGiOJypM7K1wPh4YQo6sFsH5W
e+t1pRSX/uO8MayCvC6lSb8C9HX5+JtYlQFAZB6IRWpjbmTKnMF7xEqOh0v49pKp17HqnQuvMI+M
Jk72rDcLbm5LfWhFCp/SNZLMPdv9MEuA3U85r28oBV6WHTt5uVoqpDne+fjHKJyunPDK60LoB+ZL
SExNNmJJHoNS0FPd1XcgWSmj11czEXw2fSJb4ZQxASzT+qtFYmfbQ/af4SKF+fvCx4UfLj9nxbbK
E0Lfc02O38Pgh04drGzjDR0yuLfOqE9d4h9uFHE0O/WV2ZhT1IaEVzu2/IqKO3O3CfqQ8PgHvAG/
BTNgK03XpsWG0Yowh+fSXF9F9LIRPPFqp6pMwZuPbC78svsdbKwuHAmzMG6VZoIg7UvLlg/MrQU7
U0FWOO7v6xDHjWozCEbvErIlKWgzOXBq20+TRstTRgQY1btN3sJJLufmZn6dcn0LRZW+gTBgtDMG
tXotn72fIxzmn5isSbHvucNvOkhH+NXu/LdZTnhp20TgFQ9ZhvzsiSRLkD+CMkW2NCXdPnC8C9q3
aC/w/Wm42z/L9b6ZbFKIB7dZGafSp9Iv9kdIPfHl5ivubJJzjfuscZ8ea7VMO95RZf+sUirX3pem
sqVlDN1ByEXHEu3Rgu3s1/ZFfamz5B7CFHhPvspRwah4p3IRieChZ7BJ1bqq2ixwqte2dQzA0RgO
VG1fbd967kIzVdoofx0o1SeQ5tg/KODqaShfXBH8eiuRzbuSmkgfBPCEvp2URNFZVzbaRfYFaAJC
hdONSrQBJVQIwytpn03/b5JLvIjKaPfWPA0mTi5WjTEoVaPjK+TsV5t8/vfeLx2GQ6+AkTYWk8sf
3qK+myEOQeQDRpjHiQqsTFWblVgkNQ2OtEqKAXSlQ33xXF3q7WKFab6MC4blFKfdx3byE+Wwumnf
7hUBAsBtzXPJarzZBDQOMWLU6hNz8BU0WsIyozSPKSnl3Fve0kLgdTYE/TNY+ZzawuLpitQdANXz
i+FcVHig6YMYsMzOv7U5BRgv+WyFfQu9jZ6zTYFHuddMNTcSVWbnnHsf+JB9tGeWSzB6GBBcHcZi
Kh2wTkNkNAyGn3AMBCENBP6B7QZVYp5sEBurV2CkcLrWDoONcJUN9b8mUevolCSyswcjN5R2u0VK
zMVCIqdWt0LtS20RPSWv28pHxQQzPxrebnbCSbAMBjqGBnwg/UU8CBKxoYRbcmSUkzRbkEt76QH4
xTgx80+wqhz4RDUV4Mu2xvK4Zxx0Eb9yPn5pXQbnE28w6MvSPss1A4RVWee9FNj0ZbooVfrJOO8n
QkzgR5432CuOyVNjhiEhk/dpHsGM5Aij/WmOWLikfemUowuz7Acu6YKolnLRHjcVp2msGt1ddabg
bn7jtnBYwD77whQE9QiLKlVSal/iuxpcaHg/SVnppp/mapHiHfoOa8dmph+W0xMJpWYSklXpQBFw
jdideSjNzG1JNrorAxUmtr3rRgO1CoALGw0QAnroR0f8wuGRE3RdHp7ePe8In+rKbfYXmrXNY4UV
OnrKRRe2/LnjcVgSWErgcYqJV88RQgVvn9W4dQQ9p+os1j+LTvkO0q/GuMKZ7HNAiM7fXTqkuWJv
zB54lx4ub9O11QgEFq3pAYZafhAf6n30jcl1qo9F7fS2iEhlaVzKvUMt+hidkdnqy1m41lyPekkO
WcQY8ffamKZCXsJAgcDxFZ1x9pejdatnoA+6JVXh8i0JyB2iEOZPgEglzQtmAhJijcRLcI4T5bw2
GUnjTqHVTCC2Xe9SitS9MmUbQw2idXjoERv0PPzN06Y1nffS7eVRKr8/cH3H7Tt2nJKaUFzG6vvV
VHPekButbRbsb39KGURE5VIJiX+SWMscs0NxUl/Sk2Kv6Fp3hduQ5E0HveUSKvMGS6kq/lUiTpch
up8V41BrrdlVLwwPc9UzMfFYoeH78HauGPKXPcsCjGC7V+bTSpCGwWDnJPpvMjIvo8furVGd5Boz
FEyOsF+aXi4M121qwN2oZN3MVjeKJ//Ai1PLxE/mdw8rCMi84B6T2nxiRMtIGXyj0GndxZxnlnSb
daMAayErnOTYxcJS41XQGxUwDgEM9IlAJI6ojncgw/jBaATUoN/d63nSdo7lF56En+i4CGgGrZIV
UEDg9fXmNoZqTsU+yXSQJPif1rKDTTuLj1vTYvQ8uVJgoZFY9TgYM8juN+dwyPNHsB9zojSjfKiH
ZCQ7oRg/NwKhD7Jhwm+HkZUFoR22A7bOYYTodwIuxpsqNae/BcaJSl4Mst6cTxa0Ob+1bRjpdZBR
kxWQbgxmd5tNBXN+3ZTKOBYPRiMeoIxBkGM9dBMELHOtOlL9KhOslEm6sbwm96c+Emx4G5Gnxd3F
dNed0Oc2U9eg+qHsW2Q2Zu2VJ2vJHYeBctQ0G3sEvtmTyR1UdCYWtFbqlUrePsBczKuviivOZ75c
ZClHLdTqBBvmc0drm9XaAHAmF5V7awoQ3bcSW9Z9yeccj8ni0mNYyoF9C1VlUB+6ISJJ5eEEMHGO
Hjv3mOVbImuqTbDw8qK5Fxiwaon0voYeAj7SVc/DkYzveDvZ0vMdZLZCJI8Jl4WI0zY+3Ar+wnQA
Q9eueTAxnn69JadL04np3y3zdMuwWZna3XFHT+hlC5IZQTXrBEkMlzl8TxbeXxPlkynqHxpWY/xe
OvsYRnH3M8li4qLyzLtvep2U/LIkSmNw6fNTl+kDQHyHwg0Q6FJfF3m3pqA6YfdBu3mfPVJiEKp7
0NpJE6L9ydD2J6a/TDtT9WWQaEzDGlNYXmjYYIovQx5pw977U5eDgBMJt8zN68WTY9nC5sszUVXy
nH2UxSgGXkBhP9vnKC25RxEpEq0TGVDN6tbr6N9o5R8SiZu31xYlafga3giFsAVAh9XmBoay8UgE
NVRCUcL+c/ZIHcI83Gczkn7dFPLXRCzJafSTTpsu8pT8tXZMufhLKcVg+HBFiGp0r2OzkLSbLm+g
CFv3pneOOf53OgQHhcNGwUph1YkTEz00z1i1UVvGw0UFQvuE+cw76BqNDh6MWFHVf3DMavLLwoE7
XpV+tOmpPmzm9PZVvwxC0hjOMXQz7HW+ejySr3J58q65SkjJNa2NWSBjfGZIiTSr208OhdR5JvMt
4ZkdsoFvGuJyyjkCxwfLrWkSEq6EcHp9AJUmL6t9wxSKodWNbYvs+whRh6T3SZz2kzlsSjjpQ9YP
C8oDoT/MYTHqQ6vNon2ubyTX/sDIH7srjK9VJYWSIoqP5fL7XnNNCP3SkHXbf+osDXqYyGdTn5v7
XN0gK49ru2uRdH2sIzOnD68j69XxgXCzl0er5oVfU7M54QLG/Ukh1RmNzkul/ZM+fh5LlrwV8rVk
6B3hNhMugg3yallDoThQwnpfgoH/lCIPHLRaAp2kKWm3foxlwrfV8xhWveM6/5KSX3hjVFpU3UK+
ZNNI4FICOQn9eyu+JiOHqZGLzqbvlqfP8ADQgc8fujuNrBVG/fbp7VcTrA6pD6+EDmBMZVCDEm9m
9MnpwKX+ms7c8GKfz9xpRQPe2AjR6t06kBJGaG7GQp2lP/KOKO6hayOgZHKGNo3rC7PA1Q5HA2wh
B0iWYQnV0Gbj479oMn63jaSmh5GPjwkD00/W5yCCjnOzn69r2KzF5SJYD1c/AuvP/O53cAmVAN60
bxfjo0Y/sd0rFDVwlEtKmGp2NVPCPGvQtLLARNmRmx534pkt92ZqDS0w6gJ4CO6PlpW/dHQkZCZK
HhR5AhTHQ+fnpUftygq5P/9Aez5u3cnf6UUCkpsO14zfR4pukXI4jtjhq8/cMM7HlC6+awLBTIfY
HKZolkqJY/j6nWdxnnTUzUD6f8szf7fKRY/Ew9EyWcIcheX6rJbKS7YduoAEAtMmmG3Un0chD+ZS
3pSQNzcgcB+57CDzwTvei+lefsABmcN71XYlQ4L/3ZHk74Ps1y9xMQvqHoYJXcBVhB8tD+NMVM52
Nw/UOrqaPYOU5YL7TOldvbw/uMcuEGNa8ENzk2PmdK40sQDgblDqsJCUNhEFr2trHrjeojP0yjzw
QNeW4bBtFfYPZM0qb3IvurkXD6OBovlEzEo3WK4lBs580AVC3rZqm7jmxe3OCuAytWS14oBcyCnL
oh86YaGbkPl2iohgO/VpcgkBJbZNGwGUJhnegMkwemXt+REB7xq/C+oH2IRGIsxVc2j5GfGi5EfS
+rxj5b55pcIwfFrij8RUX7FySOzHmfJ5d+ejiHcuvhPu5K8mlCjO8y5eVCCJplkrkMYW+V0mX0uy
VLM0uJIbx/ZvtFtQ/t6ezVk+UlnVCCqtwYdmBwlpYKf3kXdAjxsyVSLTcg4vsYILbP8XRlMOABxy
U1UK3lv+3gwrwinZjVs6yqQKOCWwxqoDJHsGOZPuLt/StuhdAgy0jpwVPqqemj+keJAZ1wSsXKw+
UKmWqvfTnDiyoVVszaGDEydPpLrsadHAzbID1fg4s65kcU2kKybf/lOgroPyE4e+ImQfhdiNXOZO
uAPbIqE2h3ji/LZ5iF+wJ/6dFDUeVRaRcVHMcqZ3iOG3DT3xS3vpBi2jiBlxiZPP8GnyL5CT1CLi
l/VcPjW2n80dz5RetUXtIyJJWuIdSt36EtFhK0+UQqwT+cKBhbFUZlDYX6Q9io4qxmxp48mIO6WY
5J72hVC/ovp1GKB39DYnbpzAiUvBaims0cMSEed7kKObFLs0SarThzj6pU6qdbqmMvueVk0g1vB4
w8Poeb4sz2BFxzLkdmFr9Kpq7xmimFrF4KsUUwE9CGqMQJSv2zTB1mg9/paISLRmOXkZzkQJa669
44hEkLEk9PQu4RubFyMiRpNIIg1ELwPh8jQRonuQGrpsBIZd/YfhmkLbvkhyLsgh6zYG0ipu9vX8
yVDkF7f7Teq/iXGHLCeg6RMxqTgR7aUK4Ocm77PuC1+yntZosist5a/VuF8O1dkJ5EMwe0a7nkgI
1cZAr0v5Jxx+TCs+zBXPN7Bz2SrVuQ9LDIXQU7NWyXH6JSkq6K0I+R82FRvAdae60WvhPQkbY/f7
TEDMSrOhN35s9e/KxPkCEz4oMizv4eoAIuUikAF9tPKWGbOgKUO/rrXmpKZy7H+lJ0TTvZKJkJ3O
MvcrRkn6XIMOCgP+InT6ujElZ2WPSDAPr1uoC6TNbPTsiGfn1kh/YjGgP76rM2XRx//toFLo4BTM
A3e+FL7N2zDTrbgR1ZOx2A3heTnpaXNYDaPpK/HTdk4hyz0yIXvxXW3n09i/HkoMpMvbpQ28Ao9z
6Kmio4CSFRQa1Q4pVkH1zC3QpHbofEip1va6JdybkGlgJB2EcDxm3ttmPxMp7rSqRum3mes6Y1yi
kOSIEan/gAYHKZcPv+yO0fd88v8DMbyZb+7hB0ejXu+q+6sHmq1MwiCDIlqx4Wcqff/90C4OIgEa
1MPZLEwhDnhAISgzvfs19di+LzWEltbARAw2sr00S4las6dABFhMBQKMMLFGVSzffm2D6zaJjBxQ
jW6idE2uHBj+Of0JeM3SNntiloORyx1q7gzfWF49R970o0sQUwJpXjXaVSluJYjMSHTGnBdtQpq2
ORs2ZsMcdGqTaUEfzpUUmAhoItLApUNjzw6TL/ZKWSqUU9epoRNKaR7MmvJaH+1QjF42vM/JRjA2
0feJaIOBCOiocU/WfPHcpr/I4dvf+HlbY54P7BHRejLbAATm9i+8Gy6L0I7l0cVEMZTGJkRS+NGO
EPcXIDL98IRZwKdn67GkJeIe38J4APysjKb8AXw+AuOnnrHovSkKRdxejTzAihLinr8OVHlMn4ra
hXWTLA51cngPtnet31aSUgYp4XUG/V4C8bQQycRvn6JN431wCz09Y8JiwROSVmSGeEvIZEjKCSOx
iYsx7Xifzy1/4Hf7oZQNpDxgi5gacHGzYpFtWVpPLn0cBGfBTIiTbrJw7GObflbjiyNxsRgAGar0
7rHB0HZX1HFRwRTKwP+O8QIO+NTWizZNQRaTMiAkM4NwfRfYa79OR330p22U0A5nIex6NCZTR9Mi
wZlWdvCMU5jRLvDgb3QRW+ohE4TtrqVA4x6r/Gulfat0dOhEHAGC9QCnf8rm7P/HN3nMqGmcGwUv
kLhxVJogVKwfdbxlnDUZCwu91jGBMyobPx4H4erqiJZ/OXto6gi7zRHHHZHZNgnetTHXZoAwmh/X
ljMUrVlUSg6Axl5uzIAiIeb40V8+R9lqDK90LLYWGHxGP15MxO8gRydsqLiFnzP0QRi1WUdQuLaV
EySDp3FTF9n5dKYHzcGDGviyZghpseLpy9q8A2+qQg0IqrmWyMhITnYT67ix7ynpM6W1w88inUTo
j30HYfIYR+zDdw/MzKPoNgKigxVAgTNqw99vBd+WYYen7oXoovtdLTfk3cael8ocRzxsEez1C1It
LEM9SQc898cBfmDUY9xRVodCNRNJsW65P/KzRRk8ZGXYyJfgXANjWXU5uIgqPQbU1Sxjt792ZSUh
OnV220sS+K339QHmIMn+kTRzaV1xqwwzRMwVKq9IPsTkJNv3ChZDmevlXrDw73gbhn+R9tMgF18X
eAPZ1DC0MOaTQyrHlKhD8toAHdmiiFoJYY3aJIExVEXHhZLykuA+Z79GyHm4h/50/JKtWwEezsdJ
7u3pkblR3E/lmXv14YP+g00zH4M1DsbKXMX5AM/jJbOgm6PFsh1hs/JeT/Ia6BpsUCffHZzRHX4S
RqLaxzov0LkqVcs1scfnw6QQthoGOmNQfZhILP6j2lHU7+8h9tfi/PYBhNCObLezkLT5xyFzsEox
6x9I+TDyOLD4LrPOahDwynKXPMnp4sBJ5/FZdTRZa/kiBebQx7EHvQrIJwV7er7EEk2MPBBVEtNz
fyp9v8wkQWAWJRjZqzTl2qEG71Jozv5+MP6jYH5PGGbQ5JBvwTxASHUUfyeXvXuNS66MVubmI22Q
vs35wRZD3OprQFhPrEKcKylFjWhHAa0kXSWjOhlCaf6THmhIN7DyowK638zVpaWUYZ8BKbdLmz6h
LG4VBukKUAp0fU43eynGIo9/f29CZwUBu5R98lJQaNBn6nByA8MoipyDLMtLxQZyxd+spyaf1gG0
0vZOWLRD2EStEniTrzTPsyTOJzmHdbPZ71VpT4aaTi+aOcuTJ7eZbRe7BtIG6f0K4soDwO3En2vd
BmrlPI/iC0UOYEUvewPf4V0jSS08b2sYbAr3sb0XYF44ENeHKiS5WMDSeKYFb73MuTXtY6DhT6AU
HwNWuAhD+n5hBzlzvM4Ir7rv4IcqqEmUSlgqtC0YyA5wtzKwkHkbtEZ5un+e48zprl7nCeaDJIYL
PmO1Dmk/kp64jXwDMOOpL6uEr9dg7YpbYCi2OxvAHYz9ZtQ1pwoxpjuCWluUqLJGg6ux957ggCWq
pBA5mBNBI9LLbBSJnRpag2I5HWd6bMpmQ1ddgs8hGgNhaus/kVU3UQyrONQHjUGn8M2bNT5DDl/W
U8FXjhhr9XEgxZHPQ4xrGr1Qg6k7LCancgmCw5wdMSPo9sRbECOkz5BgXH06KAvdhdoChJk7FAH+
ajKrIJzYB9UdbV8Na6aszCa6u1W8wnUAVHnlNuhx7CxnZlucLR6fLMH2RFpqtTimZtHVjO+hiVJ2
ao2dkgYTmNc+gmHjDY0v/a+QMaKhn6zIze1TRxZ0UUanOE9/qC7WTV417/2m0LbO+WRe2TeEbpM8
dS9ibuimKoZUpPVWrmDfmF/PDxVSYV0xxFi8pyuzMEhHD6wnTQkAXTeGyKT4TpOiq1AhD6n/9MNy
noxvh0O56Cx96TEB0MTGQL1lIW8JuvVlYICHSuFwUuMYYKcr9vBPcu3wGFxRV1LIBrv83wzNpk+R
65AWn+qI4Cm5H44VyK21WMOGXUMn4HHzSOHzHwA0BBSt57hfX9WY+ISet7sqpklRtiC9V2Zvl+m2
/Go5iULIRLWLmYeTw+RDufnSMgDxey0a4OHXxFNPX59U6HXDONyXQaGbv8Lc7O7GB7XSD+z3JTBU
SPvUJWzuUua8x2ZssG3+Pi4F4Or1pr/zC69mwct67TL9W4rxRrpDUc76KDYL9OmOVDT41gigJHym
ycMQL4TD9OwUMaI995hfVWf+G7FuFCMW3FEORMyH/GIZiOSHalV02FBE/1E5GJcW72DFQylMXjvt
+lsSPcIxZ1I58T3ht0JSUnGo2OiubOlDyfPdKPT8xCIC5pBxnM64VgzurYJf5mB0o82+ji8naG9g
WUaiakN4b1bkag6SUTp0ffkGtCIVmgFoY63ynvspcL6gZ3ZertyqLXp8DFpfjZe7aG8y061Hg7/z
mW8MiWTcNdDakywAAKsgMIZAVORJtXULNtE2IXWfXe0ks7PdYd7rfoxn9nCS1g+YvRShZPVBNXgL
Dmt254vBcNFRpQSlRT0r/g+XyWDR8Sc1hzmC9Dk+RwHh/BddTYrnmGgKVaRAmN0BbenNr8g+ra/j
C2tPDBjMrIpw7XpUW3dyaDYTXdS6c5hAMKWcPelwkJQ2u1nNW+/3zojJCBx1N7M1RYbcFg7b4Bag
s3bVtyPOo0LiQfg2vTnQibr4uqdWulFr2+pEzLwssMPA3jeDXURjk4LHDPOQsN1l8vAPhifBqdvm
wpzT9NmYbu/jLbb0hyRrIAnRrt2ufCBpemvcIA4LhqFSl0mT/jqwLSG8Jg04tF3M3Eeewec5UEx9
hONmjXWXj9P9IFgnZXDmMX2PFCs+8es84aiZEvmfurjeL0MYbYTrhd1uXMTHP15QtqIMqe9qPKqx
40Kxji0wPm9RFPoEWe16WQbR20d58rg7z6O3KAqscAVo2A6Ybd/adKHi0KzZHa6uv7QNOFfgTiF6
6m/cOLI8JIx/S7jC+mX9f8OLwE2AZFOI4Dn0LPZfKMS43DYlD3M7QQnekFHCuKFsMdeegWH9KtLW
Brsb6loylDdfo7TQi/iKe3KqyjI2CF20quXus+ao9tA4Jpg3zOLRwb0+P9caVSdb+WmtXIkC+vAE
/pVp8u2bJj9vnpy2pgdR4oQNUuLqLCAwwtbpYYGRHayWM5NAkPRaVgOnAymOzt9+6DWjDl1Jtg8W
q0z84oWwvzbLKdIrgJBT8Y1HPMbMRYon3dzhXnCz4bEQY/pIENRbZK+AmzqvSEYtGDCEOlzM57as
E9MDhtZLGSas3byLT7ayWpOH0ogXBo64APynX3nPjSKGTGPoMIeTp45jPVxg8wSSZfsuvP2lqmfn
lTBnQNSZwXlGOG5XDU7Npv9qi2nsWqG406ErCmfFdiWc82Kn2mglnyPP/47ArPxraoMPZqHPo5fA
XJDFJLk3DfsUrIonZj8NUPDu5lE1GGnHdWSNmAEqNTO88j7yKVxuyyw98XBIZwmfeh8C7UcGXDV2
MJeVIsnOGD05SQwHbquZbAXB5GmfvcZHhPHrxT6tyU6pfDXcPgDDre7Uo1rAJwEgH0FFWJYVvdmO
v4w2EFhPXRjC2JOJLIqZb1hXmXWySKlhwOErGypsiZST+xyqfgYAlnKTXe6WRcUYfpE5WtNx20In
8BEnxUKfOxdOKzoqrWieH8qDvKV3v+bhD/g6RjFB6Lz90T94V9tl/wmDRRulTv4zJLiZvoWucE3x
CIn7dtz3xonT3wGbYwpoDJDWa3Omk7C+esEQNMwBmaQvSBrZamodHTsVdfofhHC9N4o49N7GIwEw
Shekfmbl4XpJLHGFV2OBs2O0viR0x/2x2K+DUhB8oQk0YMkThwpoPq4Duc65ZueFQqKtMyGqT4Rh
3qj9jozCa+ZD8zTwuB7pOFfoeCzczYqr7AUjlr8lgpepowIlMmmQoxOAMAP7NkeSBnZ5zVGc15RL
iD2AuPWP5wjQdqjazSbKaYwSfJMy5d9ZJQ2grHn/YUwOlBvhIdYmxHzhjBzArHc+1rPkhSdhf7PQ
E/W9Ifyj6FVVFDuQIQGtExW9z44UWlaZGKfQv8sq0J9zXQzEbqRJW2m70wtW+M5vnCBqtKsfHlbz
2NFB98pZdnPCx8vFoDyqzqgI0Nqo/b7xm6+ZH3YUjuI1nV3azf42EcsXddElCxccUUXzuAexxM4z
1slJbEafN9b7/yqDzCnm7wqE9lzI4I0z7Empd91wkHUgnEdvO5N4icSPCjnzaMW7DqZW3qOXjxFH
JziTSDHLZj2plC0JxX7ydVnsCmEQwMo2MgHbmor+uW7kNOfhMOTDjeuk8EbtBtUE+X/QB11x0GoW
g0PO2gnscyi1STH0M5rkPbAiUbEu0yD+DjOb/rOU6hjB9Gr04A3qmCxCiTIYCXb6qHAMCfbj0nIf
l0loeniBh03ZgQFQslEMAEPPA4SM3hZvpYUix1Z3MeHmHGlHepKVQl4DHjFXFCzts7IMV/TzmTER
4zSmQHrmgsB0Igk/guTCra5qc6aEzZ+P8IY6INRKX8WCqpX6LoqbtP72KPe8Ss3yl+JdumSJcefs
qm/S1w0Q4ZzlN4sWLWU1lEr3hVoGr7FdZPOA9TsZeC2PVIYYrz6mmIjgrJjUUxyVZdpIGq2ZufwC
2avMKE65Q4B81q7V//wO47mFWRlmcWAH/H/O1J205uqyrANdvN6ia4hCMnFaCw8L7Zf93rzvd9Wc
dSRlVy7HV8eM0IODd/kp/nVwFFv9Y8GTkhd5JrmOby8bORRxe4Ow6uo3H8udJiKAN7ipE2xpXUwN
NGIERwpHmaUs0/fwZGU3uFQEJuwy5n3Dw2qaM3uqxiNH4E/aazRw5ZG0og9N8qPGKb8PN9Pk8zbn
veJMBOT/ZLL/81DRhp8Boz2hw5ctcOkJTvKCajODJFthQ8tP42dcYpd39hWTPzKKV+/Fy/s3ffnX
/6WTCDQljVXHYFKXHbGO5RVzJY8g1RrixfasHLiU0ckQ23xLEowImdny6yCIISuQm2JtEMfpuuAz
jFXj9L7M8iiu8Ytuol3zIjVZTVM7xImVtdzU5u840xk7XtoTCsEC7Fo1/MdPX+4u2qDqfhUhtPuG
/N5bdPH7lTJ6KlIEFPHxZ42zkqG63UKvvt4UQ+EAChaGSwP/B5DC0b2JdYqknQ2j6XnfMtmqZRkL
tYeej5R194HIP7OLHjbdeoOCw9TNlgiO6/6tqAxRVgb0/13Y36j9ezIfrzoSv/+JD0hNbzZlacno
cG60F0MiW0T0AWWSeI/ECH8Xf0jpYu+RCuxMjBLRECBh8DGiIVXns1t0KvcgxvXQYhrUF8zDdXU3
FXaLy3XrQdISBrnqUsGohDIMYo1h6SoVSaHeoGE4QAYCKww340SgYONMWDbvvtbxQgWAE4DpMagT
LlLh3cvJ6IAC9Ss5HeU2B8jEEit48HpKaiIpccLb/rbEZRJNL5QVx6fjb0dkn7Alas5KZVRs3pn5
YIDmq2pvrqcX1HNTxDSqefVI2/BU6anAJbHS/acVB1vkEgqgSucMksNooCIvqkX0EKZAwUYblA53
hvIsyuWbxyeMKkEr0AlOQhiYnkYdKI5Xlw2k+Dy7NXezHQBV7sEae+Ttxy3yf1D1KzBGH/v1fJNb
nIL6ReeWnYjlFkNQVtCgyvM3vwWcgdAp/o3uYCaKE5tMAfYTOVqH6BPkBxK1mtlbvi8s8KyfiNnI
A0engt/Vo+38+1R94Py4se+P/4+DtkanFLKOZI7yd8Y26JyPGqFOoIGGNWcuYpYdhLjjq91eb3He
5Vk0z5e1gmQLpuGqXO8MhTzkxHwQJWqS9aLLaYKuYLqJz9La9K+ChSsptPC1Nysy+s+iEvR//uQV
+rb0LuUmw3PESmvbZeEEVYKGmQf9L5P45g8gyRvxKl5Xew4vDDaA9nU9ZQ2Lox/mufgRttTLRuMD
Pi84Mux4Lemxhkfk3Jaq6nVwOBk3e1U01aBSeX/heyFqAp7V8RRwaUkCTr63iaSNWaJcg9252nq6
LCr6sqap5quOXHURROyDXVObWiRyX7wjS5fQho6Doz9821eNzcB236ep2s6MV2+IXXQM1Mx8p5Zq
QqEaIO6esp/CgE135eaQ26tLG0xbtFZwwA6lhldVG7f7I2T+R+4m4ngpoxzD9LENVMB98p5VdkEG
SFAS6dKvATmzPAGz7naUc8/U5HhIcbMr0Bb8DYIlb7r55XtPgXtTXq9gIq/ofGx5s+e7HB7FUOCg
QW3wwIBM1+l94hiyujnyFgQGNB4RJsvcH4aXD0dfQ5STqONii8z1dvkUB7mhIAqNPnLefRvyRMyb
q8nik3iDL5j1X7aL70b8BBLq2Rxsxa/c+L624L00opF5frNL6QQZ7oQrwqOwsaCB5qp+CxJg4Fa3
G8JBLmvluSztwFB+9YceS6rCXw83YhR7xhEYA8fHO+lBv8zQIaClsl9+TLkWY7Wt86z8ytYoqsWu
G1oBJegjrE17PC1spk8DaaMNyXykQpaQvdy2/1FIkFy9JRpSmoAw9LJcZdvUk4S5TwSJOMRiBH91
umPPw6g7W8Z5uJehZSSa4UnCZLQ5K9HDESjgox333Wj/nduW10SH1HXt2fupda8LUunxyIMmQ7/+
tDuXunag3ykgpP4IrEzJfH2PODfM8VMn3Yv3bNzfojahGARWOPodkE2JAYWtgaIBRxld+NJJYrr+
wTscLgymOaHlQG8UIws5e1pZxPHudSXZed+4x/O0Ov8FVQl85nyWZhw4Im2n6wlMYx7YM3NeZY+7
7hy3At7cyrZe6g85tmKx0cY+ogGICOPIUkVYmYf39JWUOdYKoDrQpOsO5er63w/96amuPSxwCHMG
nMIAmurfOnjCnWCDMqbYVB6xXrkuieLFWTHxrAN6hgqo8ez4Tx4ogju2pFjfIATFP0vB4M9vCGvZ
t4Vp8VkvzK57CkdfG7ssiXJvIoy4TK5CiBs/Igz3SfMK1eJlhoRRDvdGgFOG4nuFZFi2yP5IBzTf
GRFvJi7i8wIitgqnvAO4DjE5fS8UlIfdZ768Y9h6bRWT5/qBLnHATSKGmV/ZSaPd68tKjsG0W4Dw
D3jyRZfcmOIIGHa1Lea6eMKIarg0GfAeY4Gom8GWvdYdmNe9YOEUtwyOiubT+uqIdDSOs1Hth/N2
3nZswittzbKMu+359HT6dHe3ZksZHUPaYX7IXRb9N22/MgoUZRo0m+DeYU98sjhGEOIa66Ag7FgW
GbLCLJ+7oluq6QOGR+9Vp/39f0tf4RQGbs3R2IKw0Pbyb1zFdD+ZceBt2bOcmWZauqYpIaRt/xX8
1JpRR5ghyq6bKcl0QaYQCEX5a+f6uiZzYMpIIaAlzKUM7Hu6h84fLefMEtS6oh9UNGW/cqm/FVBP
gvl3Yg8ZQcKt+6G9kCj54sBKUKYdRsI1Q6Isi+fjoWBNBlg70sP8icegYnxRZjTBn3QoJQ89lW/r
X/2xCC3x7VaNEkEs5vCYopWo0kaYy5tnTcT43NLAs000eGzVQS9dAd1/NoZDcVlQqw68Bf7VwY4e
87vDlcXQIfrGAm/Lt1CoTJKUvraa8dxfPtIXGw7R2lZ8ryzgaxw8uvHifjtnM4UBNcQ/at//o3zs
eSuolV+DWC0W+A05VBQ4lXeynMV3kY2EvTfPtaadBZ6KA/HFUuIk6y7T79dfzGtwOVxOzJaNsXUu
3rRf/b5yg/lFBkYPCzke5ebmb8AlSCQZU1+oODJSvv5B1YT8xPssXduzwYMBYeBxQRnfnTglCVGX
pUahwc5xIyQnZL3qv8otLKZOjHaBFz2N6Lo/OEmeOT4JUcE8w3OTOYE4a35wyGJ1M9zayftfqSAF
2F9ivIz6KBuEgaa+6mU8HIyk7UNOwlAV2E8d7f7J99YVnsyLLgO1KOe/GIO9h2s6IckYaA+YMY9M
IVYafDt/wq7tmRQ6YihJUR8dPFYrng57YnLgUKugbbvOM1TZ2B9gtvAP4tO9LQ8z8oVAB9MPsU0b
72YIL7OHO+NfSVXcPLoPx6IWHwe8RRdJGETKSxirSheR+MtzzNho+XvpTyJ3/9hEMb+9jtAm0L22
/bAO1zGk4E0+1+KF7fqxzWR+Hrn6znAvuztkPVCJAJXP4AS8ifd+wHpOWkE0SoDWWBuzcyXtfAKk
391Euj2WeSLImkkt+eaMzvOdGQdjjYHBHHpq5H0UFfShKJXajGOxQFwG4lFyc0ad38Ij9axbZidp
qfxFokec2gqV9WbT1dVIKo0Vlepl+HK2JpsfTdhcwT7NLMkw3zMBw4DdKPf8E0ya1rLgIua7Ey9W
RPpyGVvrsynwb28IJ6JFMhEQY1a5XZpE2cPTRzXmj+GH2BwI28kUsGhReESfnV3N2QMReIcTArwD
3dxrICNfutuE5V8IrNobZa2KtoYQobqrxMmITriXvNhqBlk1pQrH+rlqKhxvYYoJxELU+hDfZ2Ik
zCcDElYndcyXUAMtXVsnTxXSG7gtb7SILgaoZU1AnED1WJA8MWM6nai+DeCTRjf1QO1q3yHX5iU+
DV1tAfqX3LaCQNL5fNLoldHBQRNsrML4+cmQtYNfbPZYYPu5Yrae8KHzxQI/cdfEoFFx50ANs2cP
TGaU3KFgdD8T6djVib39z/VLd+E2k4TeWy7PuCAl2Iki8Vi50PzQkF8KNv/DNKl4U9R9VgpacC9n
aWaErfnpqHU9hKdmK1ik/MT8H5Pfb6PG32VKKX8bSHdnWy+wN6Wn4L9K6xg6Ze4e26BJ0jI/tq3X
BKsN52GQy0GycWXiPy+fUqDJ6iOpkkoluEZnd3TSlWUVz9vfV/VHPbDQcv8XpNVPiIny+qdtQrZ9
IQ0QMmrdbotsWg0D0Agi2S0H9xN5ytvjdfBtgl3xH9h3HwWKUF+rz3Vt+V7oPXWtUBOOIhmn5xOB
FLYbnuIrMek4AqUBmeyS4rk7FRv/zUJhqb/AunlcIZvGV8xTqOTAypeIqh9ghCuBDgEW5mQgbFXS
OBgvl556V943hENwUYxFiIwSRRqycOD0W8DM7X9b+lFRKLKoFaCKhrWNR1k+UQZ+iNds8KjM0Wrv
cLRo9TN5k3QPmlWY2UX7tupFUmfaqb8PLtaFBMs7uz2uuKdIZ69643sAoBLE2GX+MmAUk+/EH9JW
VjzwgqKyx3Lglmq47m3IBxt4ZlpRLnBgdZnyVv1BGQjg6t1328Fm8WndDg9HzdXmIuIukLpHxjM2
uJ+CY8jhoUMEM8Ua0rFz629kJfOqvpy4e8d41hM3UyHiMC3xh80AvReUKkOHKEcNL7YIFGT2uJ14
YgP5Dr5r8P30SusZrYvW+L1CE6iyfg8opMCTuYI05mKZ/uvp4VYpMBAlf0JwW4FdbpBCCNkpzTny
LAhHFyy3Z428SNF5dqLQguWAeq2ThtAOTRW2bEnlzdbsD3XqzEADPIEVHkmZ4RxeU7dlfmYwPde7
Ym8BNJaeFKAOinX86CnTOqjnjR1ODR3tPD5miDT0lNN++htHgmTsmABNbt6JA8GOi45BRU8xAS/f
Fh1CcB+irE0q3jlJ5tU5sSGj2NJ9NEImOV4BEEDEMwem09Ft/hBJ682OGTx6oCb/q5xoOr1hSL4r
qPqoH88Fwv6RlcQt6jaC6iLJCgTVNw64cenjMNBH8QU9tA+xcXtd2Z02Zi4fFQEJAAKc/scdhbtu
M42u3Q1DyJWZPVSHEnidpuYyIPp3m8Ie99eMxERbxs2R8ksHwCmT0nrkJWvdOLhYjpi9dAoikuhh
T9JeBSEaj4h1Bv9oJT6WK5MJeKG4MbiP6XpW2zFhTgV81yr6X4Zw8zyYNSvt2zLnwl8e/3EGxgvr
kvMf05CUWhZ9YbED06sOBdLsmQlscCu0dcoVa5sYQtKjndkCL0Gj9UvdQxZjj/vBUij32M4sJvtH
c8GIuLFxPyTccEwX5FTqIPfS1dmgbL0WJzeUyQlmORoPPCC8tAh8GVzNnzzvy/+SzDl88sYiImBl
23tDJP/EDPPrfNdjHxVOBVlZDQ+8TL5p7XUL4YCrALr+V51cCzJjMnxt914IbBeVRpi1iyzm6y64
TQ7D7RXmFrD9p7DWAjeH4+hZVP2Gy37Aj4L2W7+DyRBaKNW6SGCBAoFK5LhTgSl1WLiXQAWVHVVV
AjkTCa2c5RHAXOThDuasrQZl0RtnaGToYwN+Xxw09QHN+8V+Vl+8SLypYVLz6h/uejLh/UK9isYf
zxGy+emNce2SLv+w3NDH8w7iZlU4J4H+M644inmPNTB5TO3vstH/Y3cTv5KyntdYUEYD3XQs4KDq
z1xifu1jePxQPHh126dRVAwRwswyFJgvp+SXD81+rETamzzbrl70eFTW+pGsnRXbyq+snKax7+sN
kCyI7GcKSZ1Kxmv6gizQg9ceERaaZYbt6vQDY3v3NgNO+9z65hWPRVsQup3ukaab/JPQpCKXbWzN
/LzLulskqv1QfSDgIXhDqwJkCfjuejRcy+9ZNUJqpZmaf5Eno26PpyPnJ7UH7O/NKwAUKPTXMubO
TGoScE2799B07oIXIzzICMjKG2LqfRR/rPtsMMbu21kNveC43AFBGWtUty8f2Al8ocHkreR9Kdj5
9kj+rteKyqLXEuzCqQSHganLgEhoYlY20DFUbWoMqFK84SYV8E74RqhHcaVCbdEbOs0TiyTw/Xdd
r5rul441jNR/z7oTSWlh0o4/lTxHNZZCZKtJ4jOzcNNGHBYGszHVmlBSWUc4fHqIN3/zYQ2MJn6+
fqbJOzMpQOXA4BW7czrCcEX2E2Kv2cVn6bZWChGNy9hhOebiU4tanRxo3fO8+7ypck9sEBrYgUFv
KADP8TbMeNNN748qZSSYSB8sEpd8/MeBW6006TPq2H1iywVxz4Dtt8nvfWF2g3ACwU9fFawvM5O5
U9g9AZIywtDBpP58BP0GTIOJ5vjG6Q2Z+SSKj6+85n5tqGvI5SagPZcF68RNliKzAamct+Cag8H6
l/sGjmeIr+O9FDT9sMxxBnUsBh8EVOaOl83ttoxnw2PCa8t1Sqja7mm1UxiKoY3BB3NGoRqU9H4y
tNKqOBhE0ZJyNrG9RalAT64zGuwIv39ooS/NuaAiqdJroNDuiCrF9KYBuo6bT6LreuJcOlzp4LOT
W6kYBh7CbKH85r1b4UXf8aTx1uiWISHTTEt5IfDJr45Ma/IOAYzU7Vd3epVYR/OH6Y5VeWbRprWc
0A4/9ExUni6WhXJsT/dhXp39tsMwbyCYzRqyNMxmbT3w8sUMDvFoxs/MYKrGhfEFeuSpqAg14Ril
hytzZmFxnZ3I45MbP7u8Quf7FRhM8moKBtC/6HfNLmj7cqvjTHTT6zkPDzMgzExXQyD9H2TT85+p
w+MQtH0TUFDtJ4sx8rkTDjdrdZcCrmBElpyPK2wAwyxErFNxMerwzPLH++FFkLek1lSPZpu1wQS5
TVxSAohDAjb3l7GRMKKwE1teriLv5mXhs69AEXB/yg0NrDdz5GQYtVewMPVQBAVCdDF5BfvzESZL
/m6JfCV8yWJdE1JMEqpUjyWqD9J1k+mc17iftTuQz0s1Vt3AfP2EBU3Qf5yGQxFBMCDPj1lIOFTr
fre6qhuKYt1SzwwSGw6weoch97xE6klfIuAbaV5TM+227G+tYAD25onWm86q8zJEPGKiIdT68EYl
ifHvDdEJXb9beBgH37htBwJn55dk5M9pCSX8i8nlda94rHSVmIdkGoS6H+RpA52jLFmssa/CdN/o
OhSZLT/bZk7XjHHP4aA0nqLjPJP/DO28YL0hGnEIXBZpib11w07Q8UGVJxc4eahJLB0BSMYP9R/H
NgJk+XLOzYvh1OmXAhmtMjqhKCebM/xd84hR7z4gTWxjT9npCyQiQx9AYxYiMIE9odNi7zrYulMp
+N2fbez+2f3Qva01vPCN6L2OOL72PJc6XsaJxoydYbw8RzZBVPU50PWaWUkFmAZICxW4P9hVzjWW
zoovhA3oOpIySMVcNvXuH+gUdO7fD98qtAeKIwltx2/YI+t7zKOL0pFDglJND8Rnjc8HWoWgUSUh
YWxHzImKzjydaVZpFZksTJ7wZR9w8fYwjAA+qkO+gibopaPMkw+GAdqErydjJgR1OFhZsFypD+qV
c0BfdqnAWqdcbJkY2huPcXCy0BpfpLd4DDWha93deVgIjdQyqZbnduCGehj3Ig+r5NZ7ChNoiDFl
B/a6uYIp3aPr7PezfYFaLHQ/rLUwBrMqKsgnHIWhbje4raPcxkxrC7R3ulcn+94XIdHtrnffG19D
0MqpmJxwU12rMBpWRRbavyF3FeaeDozfjcez9UI2DoT02LW/R7PRzghQ9mPLhzx0apkeKgWQ33bk
nRul2dw2vFjM9f4GaEIBlGq5sIEItx5ZE2sQvg6OfLoFkjfBTYyEAuWybffe5oij2LqNn+tVH2si
hZtIaWqjH8U5UuNfSMxwE7ICPCIdt2V99/L+0exLhzmdA7l4FClrohJP4++mugHVHFV4KbSWHlXr
T1j4FUeAy2q0KbVe0PTNUREml9GuOxm458vXRvvKoGLDFBsU7Mw6yAowy9SSbVubnYa/msayAKik
PVeqxsOnvQcQ6o0vYw/i/209XtDWZzeGODer4cMrDSN5IJecHHFCdlLi2ivgmcoOkHN+3TvfXaO1
Jdge+MbCuzpB3w4gRT5K9IGCtPygvvD755zQh22EDPKwwPhwQ+F9uniSKn0HmdrD5ljDzeCXDUuJ
XQlXyzB/hVmAeZSeIIFRasV1DTHFb7F09c5WjUeC85JpFg8RcqDzRY5UdABfT4eQZlJC6KaE4Ni+
OSd0JcGpsa2CMmSDcjdVK31NP2OJSjEMpACXp1Oq/UK8rTc6Q0gOqGueK9beswpgvIot16hDwaPG
lLNZdmU6nLmdzDWjcRUXAKfBMK4cpE+99uCRmVoSvByAHa03cmxXrHpekWmQrNOM4Hze2YankzWX
1qUKt8xPit3APfvLby8ltTomTjLgW7TsL8q5LXw5DH9LcF9uxsu2wTdpGUe3On7bNO7M6vN2JlU4
Lgc4MDJgtEAgxPx8rhSlqhAGeiJXYmcJpYS7/cHGmI99JFsIIbSUezoQylZ6/J1n4vaH90Og9tGc
PEnCUWP55P8A3+fhc4lNvX1Ercxb0CLFnzNs7OTzW+hYk7lFEZffZgXYNdd37W5hHXGSYx1wUYNP
hLE1dWX0TTb4+nVp7RA4BIapJJfkpsoIxi5ASXxmvOrzerhF9ZGXPY293KYg5etkFVTNBz9lg0Xb
gHbWHomDK/qZoJD+gr8NHLxSZYqwYlihrvqDnFx9eLKyzCUuJvDnWcEYXnGcTdAq39rf/Mdg/Scp
DSGdxSWTYY+k/g8hSPlZp+JRmD0XNk1VYV5ylcvniH0Ifjd61yRXZEnLKJsLToHhqa8rrD2+KR5O
dKr2G51Cpk4tzqqLG/rLq3ZhYioSs0seNZhRzvfuM+lv5+e3nWOc+6ewP6LWOjPv1UOVrYDwAql1
BhttcKckl1rs4mcinBYpnxUQfKj8XfNVbTgXfmPBoW6E4WY1bX2GqVcdBeu1pgUizUd5bI34oON5
ytYvEEEqhBAtHXwwaIJdJnJjB/Pn7pwsJ6Lfg+H0496RG35lnRGc7ABZBRDNXxjA8lw2mBsDyQpw
Mi20GIaLpFqbmDpiBt2bpUCTqfA5J23T/jbU1WULkWHpPHIA5+FXhdL6YT0/7PDnyNHfHbHaQOuB
V1mEYG/pDQEeOIw0srVQVVHZv89ioALMqvaRpFurPPt6s20Utky4oq6MJGs0N794p+VffJ8DXev8
IrOpxsvWpjvr5BQiwfaYr+UYWjM7T/hxrUSk8x85waOUUFtlaxKeZAdlG4jdo6N46dM0Bc1Gd1QG
0tMir7ogfT2YR5VTvlGg82TE0dXUKsA19QzF8UjzTLW4EtV9zXGj4RBLB9PSwGoC5MCaV1y8zkbi
pcXvGAhJLu4JZSSze+RTy2tFznqtQ1hCPIi3nl3mocTbIzwWzz9UNHixOTMAm2g5JmtP8Vpw0mTD
27wNJlvK9UsNBmsT1/7O0EwTA4g1MDJhizY2zywOqL2kPLVeolNwIexH0OBFpTTegfZ28FW1uOnV
FJJIge/VfHY6mWkatjPZsBCmPaq9f8mxcokds7yVQWg1ginn61+QR2MDTGJ42GdFQrCHmFN/yDyh
NpSJZf/R4TmyJaeTXFQcz9WB/2UqxG6KKLIziyCdI8DP5g+YJuq54rz2VgPId77XchaMePDUH3Ma
wNXQ0H37CAoHPjbnnauOzzhCPtj4vLPm7x2hPktelmt46vaguv5dOWBpqGYsK00TpglEpIwSyQMi
4JJwvheYD3ssKCLfFLNBO0xvKCNUZ1wew3AivY+JX95fA3Bw0yUL69TQvp25Az7njR/Itp0vGbRi
kc7piLdldH/ZOpyj122G/x4fGnMDrWGl9Z1hti4yM2lXerKczGmYzDkvGnt2rTZRaMawWm52F6QG
toZQaqnfQ8NZ/fLahOjYK/oPCiK0gmLEHIV3UM/sxktEp5Qqmuq6xr5S7U4YUXSO4kik9s9Ekl0s
VEDnaNt9YnvHxV0WQbRj/YW8cZHxqWdTBKbptqZGt0yKUztu7T9YQyQNM5t/cmk1mO6w3cuzXnzE
0ClgWXcGLRmUqfbnf6Bb3l1LL/S9XeEmQCPhL2x684uZkPL+RXYrC3LoDMyH6zOgHr4PLZJg31H1
iulQRr1I4WT6SH2GAijdxR5SiJvzxzZpNdynyvx/Zg9Kk7LnC/ws5mdyInzqz3mDiPgfeV3atX6g
CVa/lJaLF+xjn3xEKWutt6YzcXdJm0o70GQSNlLhMp71w8BwYqkg5TwDC4wYuRsInZuyl23zeJr5
TKSg9MW6yL/GvSA2gIx8lZ4p6eWjlgk4tLGu+4nGeJlN3fDwLGpFMxNsTw6dZEp2bZYxAX7zAteF
it66C7mx2mxS5FjO8QrnBkIk4zVd/AbcHNnrQCWV60Mc1vjEpUtSPNXDpt55al5aPblhvDvbV4Jy
63U0Jp2T+rG23UN0CirEwjG4+ns0TRdi778HwJ/Uv1o5zw5hm4OaKViH1UQR/O8gmdQFNEI8kujI
iWnBBjJ5ObsBbMYI+RdFIxI9d662FE0e5kunvRYe01DuL5whsnY5oQEhCtV/CJKBUO8tqGy0yN4Q
aaavCE0p7eJxqYY7R3t5kviLzNVK7g6CqzVQPLFNZ7Q99By0mu+zId3Rm84BkDvn5i+4zYZ+v90u
3yGko9w/qFdyQDZxe9XdWpE4gGn+i5lm4c85wMkS5pV2ITYSbbw+X9os0JGGX0tTmfmmjq292dYH
R5WnZGmIVu4DpSwjZmqGuhAXCNu2t5HS3HmhgUNqB7Pi6yaYSNeG8Ibtqs2/YOx1w/X3D0Fcfl1g
FTcofWnpFpCgeHvSwicpigXRMhW+k8nr0aH1qatjbaewDM+Awh6m4hVPCIncsINnL5xONothSM5n
ZwHTJGfzpy3J3BGfhrED+5AHtR2rq7f3rzm+pVXn2NlWV72S6dAKuo4rD5BbTrlFNAuBZUl4WVNy
rVVR6CBN/5FgDm0Buz0ThSXAVV7Tm5qM6b/uB4VyMM5rGEL9OBsXrt2dDrFIak7buzqD8f2Icrvi
6MS2T+mzKraw61IvCO/kHJgIDcxx+8YywGBLNRHyySZiWI+Jm5pnU8Cvsf/yHVeriUB7HHzeYsKl
vLFgY3Rt5U8igulXkxYEiqtH7rJ2Euzlgt02xPZeg5ghal04IBon+JUtyMREMWOzeLByItjWuTTO
064bfbyKAs9VFOMuntUHaqkLCEphwBnbSQI0fhrHSb0yxB2YSTprTIx2atOThrGXGai3jp90W9G9
OKE7VxNdSXhG4ielNu8P1PdQrIfzNnqqVYSuMop9spCkWExB1YLGE9JcQpC7RHb35EPBulT46a99
FA2PrdjedFfutKJFlcpQPf5rWITRVvxmmumwLlEa9ApGa8EAuVaPBsa/K7aDzKPHD80jt3YjcDFE
EGHOvzozHySN+6loXjaP/znnUfjwlWfZ5rlEEhRlcspAqYE7AYooNUvznZ7g83dqvosDQ0QOgnkK
6F5MmpgHKBqnLEYJbSVrWELIRKQFbnvG58H1ccSVFFOLZjfYQeq/mZTZUqmmaLQSNA0qi9oPx3gG
aNAD2RjJCSTLedjVnlXfIGIne6QUtEjOLx+6kOjpaVcW4xy0pNzsOw5ue4aW3B9V/jWRjAp7GtMK
kTvFkQlvF0iWvrE/9iPkPioTbaJgTLVkzxzSytk/Z+rJKviO7o97nWbyDXzYLlE0YL8utc8mjsqC
lEx/h2qNY9bKYtQn1GSyXaKdldG9+O2479T2yRsrY9Ib0NZhBmUm9mr2V3+BCUTA7gqZEDeZFnEA
DeIMaecvGms/Z0kp5FA+7Q7Iyq6Y8kQOX4y3dc/spQQvyGkgeuG7UcmDqdM8RlJC17N+E5AjySrY
vc5DuXcsFhSSLvlecPidZUPOnVqWJ7lfKtrgk6sTygVTKoL/uR0uBWuk4neXB5KfP7HJpNm9VQXj
1AFUKf8Qyxu8CibzNGLH+ImZvej4aHS13/NqPn23eeZqesp4n3lxw8BFu1+++bI1ii0SJiMzQ4FM
zuFyWzdHJijvRsAOEs/pbpj4o59mX/o59wVO1PBlgHaL10FeiP3yUBBYLc/ySZl2yLeO06m6Ocql
s11yJvK6Eijdwpd3ZK2vTUxdttLRCOtjmnRC2dt5JG8iDTj13h90JJF5qblCeDnbbmUPxTKKSAz5
W36g3/FHTUIjDMCnBydbosThq7h7IE94qCmLDNu0825vZ6VwW8r/ZHu5e5629EqRVr4kX41Ap1qe
+R5qhH3iiIysY5JURjZxtiBieFCl9EytyVl0jBQJXY3+J2xPyZip321Rh4pDQG+7EQHe1NrznX3k
Bvl4E4b748LDZvCjvcKAny3fIM8no9YwsMVqVEDYTiJOJdLDTI/mmcUo9HQXas4gUhl88TMkFtXB
vacoVuZFUQ0V2Zr832xhLQGNze4gTt7dp8Ehlg94I7v/kBnTBQecnWNp80bA6xx2J0ZkHYHgp3Xf
1aL4PFkpwZUauRsBIjKON3c20U3ZGXMtkkDRscgNNfuzyytxduE5i5f6WyAnd8FQSm6vv7MNLa75
t8Rf35SsGzSHqNSMLuVLCJvH9ZAii32zmfSXNxtdFSRQ7PcbNU4y98zZXWA5Rx7qgjjODLtHsT+F
Lr/fnXiU4aB5B6QmqUchrEXHNdKBlO8wf8EiayyazobVQNEX77Uh010IKbgq47YZ1ni5qcdc83qi
vrUQm9Pt9CnCFQjVk62ipoD2rbLXfZW3pxLur027s3OAZpA7rRYI5WoDvmM2xrrP/Umu2Bgtj5mz
+z9Mzix7AAfDbqE8QBZaITIUzKRf3nJchmHNEB/elSdOoPf/2swKP7AcN6cqstdDyMnV/BF2fMkU
jxyomzwjbUxY+3n16V8WmgSRPQwxhlkM2JcfNAQzLT3rZFg1jLld0hxX7wxHv7OD01DPMwl69Tpy
7qJzoxTb8l9gBHWLZvchLCkH3uoUDUhfsF8QmD4K6ZS0UHDKXPrWioFF30WX2rtv47RNPltkwls2
yYBf1cHupAx9ttNLTdi7uytDGLoXIdRI+w3hDS/JwHs08IjRKQa/jJFzWgdFJeqsgIbb/Gt7KApU
3MboMIswQnT6Jzw1kNyk7y0j6xEIiiHEbFssguYypl8Y39HLx33K5BBPJFocpy9NZd2JGLC7KoOI
7m6sZ8zr0ANXWRPPJVndPluEzzCh8wwNHgDDv4oaaGRuDzR3+ZyVhekhSdDREznAjVgCpI/ii9h6
aXHS4GoI2Lo+mL78p8XmnF4A4NBdZJO4OtUS6iBoIpKw0+/CF3UTYkqBDz7nMpPHsOgVJGHRBSui
cPEFzCWINIu/ZN3HtQTcfTbmOEjgCdWt3rtl2ojlC82Qr2EUK8oIABQpbnscu0cR915oJBgWSlZc
rCxm3u33wefmfSkXLkifOZnLZQqNcULB1mNW8xn/M2SYLRgF8/PHbdrmjVJyUrVsaNrbQn6a7Vg2
HSCOr35pKnnN1+a8KmKVn+oJMNEPVYkmYV62OoV8HR4SyFBK9AIA5mEVFj6MBga65V2y8LQBI/fd
f3ctB+K0o7PrTlUjwA8iAE2mii08Mc0dRqk21jUGtAobOrUq/1ig4Huv8gkginQtpS6VqrFy2zRQ
JTF7D4pQvPp31+oinzjhFqRgSYO3k/gV5CIr5WynviCfdOZlcwMcgc0cmD+06+O4iPomns0bprAI
YkPOcjN8GQTpA3GHv7+CTEc3zE7LTVqplEsE8B3PXXH6ako9ZwTZqoXqvvMN9cIyqNXVkPHxmZC4
NtYa8G4XibPzhz/zkzHSJoezIILNTvS2ZbK27wZt6BX2obaR1Czup3Z2lNjnmTRC7jRbAEQNGUdY
po4eno52oZwbliF18spmg1KWkScOgDQFnvn4Y9RUwhhYWu9oXhP2TbusGP8taazwlsfrOWi3HrmX
6RUfwK5ov1p4erYUxzUie3VCpTSCBfmiSCGgCDfI3Y0wPE8HrsabJ3nWZzFKUZD6Y3Hvl1Rjopk6
QiDlQ7ub7TWcIn2jVRUhaCZ0FOiUN3FT624wJOUH884Bp+8v9DKyA7OAFNvQKjNQ5ThQ7xGH9u/H
0x44mMGfEaEUkvSWZ9qhmSwcCGrqwvir3tubh9qtIBZf9GtbtUJBT39VNB6ululkqhKGFZurwFRz
EP76I5S8bT9SqM7ewY8VcSj0WYhLMwQJ9CiAre9ygST6bC/YZhXZoRc9RUGLMrKrslJ2eJgWgTGE
GXRjGXLYE9fQLpjAN5ZnRt1FrF+yva6YcOJjMbKRnXnL1RAjO19/cjy8A04gYpTJcX0SY4yNZ5ql
SaV+nfPt/04yzRdnL7Vb5IHkH6JOvbxA5/BXfiq49JijTuKrozJcFnYhma2H+ulYr1dBpYhBm0FX
AT5XJH32eBMbsvDa04Jp9LTeQ++sQXWVnthoau3U1uJt+2OxPOwEziSdw4XUAsiCpN/ykz6YJoJp
AWoGm3qarWXLu/l2x5ZTda7KraI7dehli+TOC58widGs4F2jtDCbaJkrCs4k42eVUY50iv451TPy
EAsjIDqsrwcN+02USxpv1migiT7BN8+Mxvx2ehwaEiU0sQrZ/PpsBU6QDs93v7OCTmoe8Xk4PMsz
xZAEgcSLJVXuDVNS64xAKLWEQhwVRGMozPJvEGqpALZA6U5aabS6eC1qK5Az4rLpCc3DFS84GYb4
hfFTntZTHs3wLoDTDTCl59uau1BTGFNKGwl/aTf+jM7vkl46CohKMdUhinBOSMY5s1HcyNGxUj2G
5NOZnK3/UaG5bSEdgml/Xcq3iEyJ+pV/qmojyBP++nRtWI2VMI14MW8gXGBFeV8foMwfwsKy4raZ
6im7t57gmUVUTI0F5TF/20q72GrLXG0CW8qEjRvewtTC5FrSYe/SUPJ4SOU1uVh/DyYtUTJ0/3vN
gM+mCe3GZUAvJ0Cd09PA608N89NQPwXO/24/2R7hpyE75IIhrsqzptMeNj5dBh783eA3QY9ntvAQ
4ecq2nCpjjzeKMffcIqnFmQS2m2TOcrG4seqB2CAICysvvgxeQ+4Xl5cxOgZmBreQjiSroy27buM
nWNp/1TOgbFo7gZyYbIjVjguie9bh7TbiGUfY/M3N2aCoJQ+KEocVMKZGAmxe6nod+2VdY9xudO9
P0u70u5zkOUIJj3gu32YF0/f3dBYf23+S53c0ABd6xM6+sxDCZ30ThuItrTQvz9G0BTfeiYILz61
pey+BINCokhIIKNzqQGDGZ9cYwsRXU9YgG0GyAnDBLBA0I6xMuGMPwtNPoE8+tmEl9jLpZh3WbOT
kDRedsNtUdmNWLsykDYq+JjkULXiyQUWY6/MqK3azxyDhII7xHdv1xCn7TizaeggokDIrWrlEOWU
OCy7jrNHT34q/zuQYTxwLPe9AT3V5JwOy0tZIFj2Q74jz7UQqjm1rQoPWTYbyvDoF6mR8PfdmMyw
x8V95ZZHZr2qK3A/peuVhMeHO8nwuTCbdE6CwMICeLAwRvHkNNxlVJl0pmOLyzDYyr5yomdvK65w
3S+tS3Xi1wZkcRIbQoO2nCuw6c2uf2T0VBp/TVsQa6X9xKr/xV1Z1tWcHQFI0lvd7Dc+SK/nTL80
BIysAhb9kgnc5fqTa1cK5cCFmG/TPe1jN+yqbiyT+UhgGOnJ00zs2zjTrvXLox05xu+41xtdKi5o
sEAs8xRQfaK+wdaVJQ0Ejz02ULfHq1k5Qob08cs4hIz7FkMRob0tjz3/THRmNR/UcsbPPneiBpg9
T+RzNQdW5VFI2Y1rLwaj7bJOOFuTQb8PqTF6Y+TTDtNoHo3nHetrto3F/oeRCMEmZERgTtbLt9at
hCdOOcKUulajGcRFMR0goVFKZ6UerKkbC5eOvtMSrNTvV5oJUI5kXNsZhH0+b2NH+WRtoBVayg+k
Zkmt8gecWAWAM0motmPIZyQy7z8tLnWHB8wlytrLKo6tcSA4cVyxqh4eDGXvdjhen804Bu0f2bkP
AbD3VHGahwHiyB7Lad1+s/3sK78ofNvoGMz+ST49AgXWIX8pBXqmK8pQ6hPxDL653yaQE5Ioi4WW
Zkwh40eq/eeTlLQBDIHVP81Nl4LPUP7nlJStCZ9eEBay7DWeFM2n/u1t2U/Q6QxGOfwsQZGlgDdQ
H4fAy3L3jX5UrkHRxpmPxXe0zFHBB1vG0/qIAPNjxrYVGaOJzSSLtENyL14rG4CBoFGdRMMEXRV3
z4B3FaCTkRrp5K6JgS4eLKU9rZfDpljo1p/4cOx7IZLVw16YPBgnQXA3oMKztsCYVk7cY/bYXBgX
K2Q7e5nDhZqO2NiGMIdJonqTgWrfOaMYvM1qNuBJ4QKUQ1rmLCqB+VM2I81ZcOtHaWRw+JR1IPFV
fw+pGngPGj4HjKzUaO8lB1YucDSKWlRQLqyVhIFZy8JgKO11fqfCSV3vG3h+GbIBIQbQgyRSUhKo
FNqjE4LCTdxWmBfFmhoLGt/khauGy8CVEPrV2EARI853wZSlxQmCuqrQvsG5laI2zWSLRrE302ZT
w1NGwJPCKDdcEW234TYRd9A9++xJNVap5E+2zmiVsIDEkdeGGeJ5wWMs+81uZHUqU9sMx9+cQ3JQ
ccbK+WmfdUuH+mJn7ni0VtU7ZaNUKFW0E6ctFPXDvQZ4oNLCIhv30HAEhW8JGwA/rk6EQw29v+CM
C6l3cQda2gUZNBEg1ZtxCuq3lNlNHc2l62vu5pIbvktNIzwsnwxqYlq+fHTwIMAnEo3B6HghtGeL
ZVkw6/xkI6wBBcLqNYioUiT0ZFnPLC5gl+epqoTck4mrZxmWpSZsiQI080noOikD+eyfIuQjkjAW
72gIkE5eldJoNPqvGw8W59MFf9y+a/QA0F6aKjKA3m4i+l8XPvlX/UYaAts3c9bnpQJJcgX5H1QN
n1G4O/Aicsb+kSYPxloeWgcTkk+kIqjtHu8YVbyi/PFMKo4gh6CGYAPQVJBwl2qCiu7G/0iXwVwz
pspz+1DDrJCee8+5eBIbS4jj12MGr4wIhQVX5tF7JyHgVDkZlbGZlkHnCwdH2MfidbfVs6gYLuy/
7DpR9heNWn00NlI7b+LCD+jdvBzJwpj9Ht0chsUFRDurWkmVcclOGS5i9IV8w3yitG5KJsN8ujwW
rKsKWMqAX8LU1wcLV/siXY8HmHhYiAdKKYCVvIEXOtwm3vBSJKQt7uqO5gwZnghqJ8JMChCuQc0x
k4YZcW9xeEqIOdfixCVkUptwrLrwmpCZYxRf3g+c7VwsFkBg+q58AxUdoMGxR3wLwdjXQbhq/yYi
UUe1GMgEq24mN/Fi5iBR30m+urqAkpHeLWmBdLmW/q73Xf4S6tc8ACvBAhHmjrVHsjMcD6P7U8+P
Paq1ysLaUGo5rnDWLx7sceb0q3fW1AxbD5+eF03+xrCfCUba/N+GYxzy1Yv4UYXeFLNdtRDup7LQ
fO32UxPAShaZA6O6rEGGuvwmjwSXgVpsdx7zqmh+9HHLed3E80XA2QrF3IoDnwMv746IhCurER8J
Ec8E9BC60icb2AzNATuuTvyIYZsnJ1+ldUyj4dnsBrL5Dl5XiPNrqAzVmXWTg36RbxDk83qzRMlv
W2Jc8U2XMcjUiAbXthdurMCDNUEhi16wS9+t9tR7bcmN6dQOeUQ0go2dBxs3cI8o830PHu92SVoA
vNGmT1WxHZ76U83XgdFLRY8stwwUmiKoGLf98kBnfi6IFmAxm1VtGaYgedvjwtfGx1gZJLPYC3Tx
YcIfvHG5fH1y4o7EpiCyOt0NMwxcU4Nx8i1e5D3DKiGLmRMfDqOMFnCR2WeD/s+sTpPEYXkKCj33
CjioeX8Mot6NKZ7kCV/p88V0I9w8yoi+PTN9d2o7nMiQXk6sh7DeOI++YtkWbdJklWCUl/mZW6D7
fZbKbsDAOOJIfrkhqkW94upxebZmwozjx1b4saXAIaIGyn1991ZThzcnT9CFf+T9KM9fUHTKf7Q8
NdNsnIkwtOpqvJtYb1nyPpQSPgQMPW5TNp+4SmrSrV6biCatA2i4KJMLtcqWaosBGI6FYrg0v1Vr
WAtu1/x/b7LWu1eXWVmxDRozqpFjiUO5mQxXJoW/WWYUdbhHjSQjIfPgbczjAt1QKwuZsbYhk9XK
oPnpLUiOqrLRj40IGlTGFua/m+C/VT4IirY/F7/ZExFqG+PXkmBf3PGYAWe6EydsWX/vp8zpjReF
VDfbXZKbMhHsN5DEDuhGOLruqt6spTeebyNjOet893SFzqcPS5eREHDas72wWWW31spyGzT4XnSE
Ze10k4QJ4rN0zedGgwJ6NmdMcjGsFRSZW3UplIEM7S8Ihcen85HXUZ98VD7PDRuKOOoN19Pg62f/
2NJnGj8AkzVTRnNZ5hzKtb2gqG4ukYLWdaVr+9UcmHNbFHmDuBt8OTubom0XQTFKiqTSjM0ucTeQ
07CJy6veoewYBbHV9oBZOWERnwR8ptk8h19Sn89eLafzqwKwK1RYFgHOi+/PK7fZXAcjpuCCT+kP
81LGsd7Tye6CldKIk4RrURBq4Ud7Ydo1uw3y6qyEAbI/fRjYhi1BgqyX9miQeN7btTgJeExA+xwS
2youllTcKfxdGgXCoWJyQyDFSMdKRvmJ1LMX1o70aTIJaBHYwVc+yp9Oj+zWHe4anVtmFhX1Arm0
6SjAv2xIfw2yIelaBjPsjgiTD7cgZRYDzf4hBTU0nPrQrOkDryedwE81709Rk1KBKC9HT8J5OaAQ
+D3FZmf3SPm3rJRk5BPz0kkpdJdgW6u8v8dPW9tLeH0UhsDeoBaiZahh8QmKK5GKcMxEVPC70WRn
O+2pAVgJpEvLPKy9N+XixiDqjjcbAaqI04WKkHEe+Gl1udk6VCsTeNn2FI+FJ4c9lY0KbsUob/9w
qtMHwLJBeaFjgu8dYGOi2a4u07rdu9G4FCgFa42yPsYEC905+eoxRQCzdpkaYgWrNe0IGbFr/I2y
R08vyejFoJpEJATKb5KtElL79Z6fH/TACTz4756D+3YrTa7K1m3XBP2SgO8m86F7mOoDbf9q4Uyr
yFQXl5P8RzUe0lxKcDFsHcO1tmG8A/Tt81w16ScvJlFcfDySmE+i3a9LOSDgOPiR8OosY/VS5yfe
UIJHs5b9hbcygekezEIOgDXndcXol5XjmEVkEA906k9qKZXTg9tz+uIw1Xod0sqZinuVZ4oFakHG
figb51IwgTdNQ64IKHC54tK/3iuLFdrU/n2ct66Oc+ADj0zXkU9Bp3Uab+7B3zwH4ROCWPm6UFWR
ZR9H59OYkPceiGMJpovC+agJ+Dk74TJUx1X/afztSdC5uKBqBqnsUkvjcsh2VeLGTYJx7/omR4sM
+ka71AdBxFgBr/0MAHjjlEhWRTep+1+kKlLoBmw+rANu8ZTkOFGSFe0kE7UAezNtaoSvW04n8OAU
ix2oSDYQWI4cDka/YhXEhxojkevpZF+mZOUKzST8/Mov6OQ6bzsy3o1JVZ+Thb2EQzeUecJsk8Fa
yKJyo9pIhelQ6LTG2VIGmnOJpeMsTjhWiSaxtwRurFRLdmCzy917UkhPdSjeGbQa3wy5gUIiYYAD
Eqq/ajwQdZ+MgmDF3jFyaKMNMo3urxLQSbbtjhcg3AxldjVXFhDr2Zpg2k2ZjWk5GpL3DcUN+57B
ysxrd+Tfmgd6ht41EoWiFl73fn7zO0cudbJ4CarvS24cEmpSquTo4Yn54ThjrtydyX9t1SYvkru5
7sJ2ZqTMZBWcNPRaJxTqHdkDa74xi2H1nNtC6ipo7pCZbPC6w/Mvq4TF2xcC/V6NpFfu6LhcP/km
brEhdKyO/l/N3EKhmqNyDtsemr6Nrd/dH2btu5fmfU1DambzuJJP5okOmI1PA+AOWhjQGq7mnfCv
f1hL7wTDvJioiQXu/M15LQZScg20ODjVXkE5VGd14YrQOvJZDMHFB4aVzsXnPOs1Za6HnpwkNXxP
Q/xQ+FbQS1mkA7mH+xutj7FslGTfoAQYYbkUblIabJlv47z3qVA1OFemOSCbScoa+do+8FSWVP02
5PCv6mHf2m1h0T7UIinu4AHKCwnlVzGOoD1Zxn9k2F887qT1332OW3i68+n0bZVYwHkbtmrK8FsH
rYK8ZU3N+Z7OG7kp4n7c/Y8EtGoBXNzxKsblwfXt/VW/LFjhAwGrZiLo1MgC7FSnmlC1lgHFtWU2
UbKeVDug0uP9nn90QzsPZJf3PCyQB/S+FiPsrca4CCYrwTto7TTs2WNpa6d7OdvQB31MAOdYVBsd
869N5nf0DfuPRSv9jSNtPOoTAKAHlJdBzGRhT9/PayvQlWcGu4h2J9+vs1MKqIvxPPNsngcH4GnY
AhBCh469all0ktw/kwKN8ra0AVxHSS5r8G31C09lCyc5M6DLNQF0eLb02wCqAzAuBOO9B84B46zd
mfG5LmHJ337Gh68p+odc8K3nrY6KPkb7QpBgc61QXjRYrlrth/iJhBWR3drO+/Gu2R3QRPG/4uE9
hA8vda/aXg+17Lh7gPbscagk67lScCoP8d9vXeUxtQ6dos2Q4Z7Vl1maOtrHO48521GQ71Vwx5nt
VBpESCcvwPnN5u0h1Aaea9gL4OUMK/8WW9LWxqpS9ZNbv7O6X/tiNNOFdy7WUEw1D00xSeVJoKaC
as/4bH24YPnfomqMxqmY8X+vZqvH/Xi2RSi4L3fpxDmHYsAtR73ZL2c97xG94JnRwe5YoGY5WG3I
U7M6Bg4+TrA1x8vlyE9GSyJSY0IWtm3MP0cVL/csfMnJR9f9koBiyDfFmjJKK5bRspmlxTcqQg1N
3Or5TXhstBKvTKJeYFLR+oryU1HpJ44QN4g91aRy4qS+9qlzcbeKQUhi2c3hjY712S9G74EWn1G5
Xq9E/Jy/plWBzwVm1LeYCCUm85movGA6T+KUjmkEbcuaygv4zpDDBu8FhMUX8u8l3X8G8s33Kgi+
nAa3U3rues8hdGeOmtOMVqgCgYybuZFN/FNuimbMz+HwpST6nmPYqSiVqE3QUIQTZ68n++3L/w2m
zCoGJOsOuNBCpMuub5cCoNdTV2aV9pgavKqLEfK2l/2xcwhFsrDr03v/qfegeg4hykOFTM5Rwocf
95UlOUn83QruYVXLvFmQKSFquGdHaezmLLNDGuNpigfTk/5rOnSfFNAcPP3r4cdSM0ZIB12i5pkG
SWbb4LO33S7HLskmiigStCL0ueZ+xwn6Q9876d0gW1WXGUJ6BtJnILdWC9/Qk3rKMpV8dOcWe33P
2JGMLDgwv/q5C35wbCYLMjmmPYgLx8Xy5OnbivAL6XClz9ynJlrX1iQaQ91NOrz9Gf/2ApRZlPsz
rNGaGQbH1F++yd5UhSdOjjz0DiZ+44n4dwu19LIVCgYxf3VOrAsbuk5MTQW3UfOfXgAB2T7KQV7j
7u5cFuKmXn70WYyGRSJPSj9sKvGoovoK8Lt/rs4tpmhva2i9KNSo1AZTicg90WiMrhWXPnVkkoZL
lG6cbE0tHgMaZKIr8X2az8ly2UCl/BymtA1PXX/VlEw18UAr4rZxZgNwkIRe67zPCt8Ygi9FjZw4
6NTCNowmN5HY2SWjm5wVQyuP21RWuQ9M+MhnJnuFK6iprq2goNLyE38/qoYj+OORbPLy+Bu5F9F5
PnHp27+IE4hLx4yMLWPWkPsVBYR4Cxo+pKSXo4/jrAW9RezY+Oq3aeE3PsXGW5FbDSaBUnJtNOGI
724JKtvBXmJfv55i7Xf1mTP4UXTAo2RJwhdDULOGaxf7LYYt+3nbNAC6RrnhZOhQboSpM9D6PvLO
HuDP8R6DJTSaW9IpUqEENR6YeMSNeaR5FnGSUVSotKkZ+nbM4xGvunG7UoE5fuzt3EoWIano6kl8
aLS9jAG340hkM8hSpJ2/NjU9WsKuWP1FmUq0vI8p6s6yPMnjLMSuBBOJaJLs1OfnpCtW9wTFLMzK
wf6DMUVgp6o2kCkp1/muh0EcomzZ2jy15XqWSWG4PXuDDx1iz4J7EEKbtwuPEqeb8iJFNCiu3el+
q/LZ5o0fvQVV3e76CjtjlZwMEAoyh1MbaR90DW5iArQcMJT0JO6bB6z0M/Ry6ZhD9TpSGKq+cKcr
kvNkpzZ0gNgcTRpcJTiMDcl7bb3mW3iXEGDwlhad+IsCB7k1eVgIWB5NFTMRWcbh6HpLvVE7xFKw
m3DpsqRJxgDg5VSmbc17A3qCBdytJmsqHbDroeinrZf3vCoScuVI3Su7A2L5YCgA45zKQZxHkTKB
MrRu5nbKgncmRO738mxbJd8dQirf8BQ0z7mLV0vlTa84mc0x4NsXCOeyxPn1YgN29NqJ4sYHyDMr
cZTwQWDlcBlVk2mdSEL6Rna5PT/WYMt0Ub4dZZVfavkyQLImDLxVjO2885tSFHOjw33IO1ejMh13
yEBRPGk63UvVQJPwdvdoSmr5fCePFUDePWLVU1zPLCpBDAMQyTjRFsnJBvJBRXRZJWIz94Kx5kBt
aanLXc2xX4LtJByaJ2Eubb2u4SEFnjVzFbNBMsxzxTffwocLPv6XnTSVl4sk6F/N0ri8Mb+FOmxt
IM70HBy4B4mc3kndXPAcLcG5Daazt9QM/S7qztALeGtEwfwMrduU08JyMj0R3+9mfQMte4uM0JQq
Nz7y8OfFtHS7WZuh6krnq47fgNtlf8jz8UiLVNcQIo8ZwaZMs6WsbRdvLtG0QJx973rG5n9UOwfl
8rIPMJ3KMxuNcbPjfZ+HCbRq6lHr5b5red88ic0/c91R0LnFxusmLYr/nxUIlHAf9uNZSmdQ4fox
5KMfwaoAye6QXqvI8YvqlEqdxL0U59sc84VdMr88i45TplgzPcrgvkJf+cmty1J/s/CA06lBxcCq
+sX8pxUZuXChFUnRquUu1grWZqtNW0uTrrB6rHDWuy2p5HrQt1Fg5k5O9qiOpNT85MJUdS/XhIUg
F+Mwp145e1Tkeh2AAFNQ+bXaMN0wkAHTEWY9zWNYqEVkzGxtiveSIhQH3YnM9I7jCc/skohiyzAs
uCE2JoP69cu2lLcB7dhvWdeGm95OYNxxzlluuQTFiN1GBoAkKoOZyKeCXQZaFZqMHmziqO0eSKa9
Qk7OyWY0G9uyyWVnEF0LYpOAPu3/SqpZUWUav6UpTwJx3tSpd7bYn/DIzr95hS+JH/Gn8NqlnfYT
dDjsPID7B00DdpOT3rlW9kVu2/d8hBYeeydX0J6zIqk8QOv+MykhNtcWH7bYa3yzMPwPM2Hg0z4y
3stzqICPdvY1dipUY2zOKkmk9kdF52xA2ZhdfYf1xVCDSk7E9wAodhgmZGwuUjJ54JgHIL8Na9f+
0sM8r7ZkgCMEavz/dNgGIGUg4EMWRhDopa7PWfD9fK1OjjWC0x6VZQgnJMuiEHJZzRVa7anr8MxE
JJpyJ2YuxBNWt6prMU3c5rAOBqht3Y8CJge3A33bG5mWChIUCQOQf8Hdu0aY14CduJWonrSMeN/X
uou8605FVZPfAdzirogNTqGyPMfKkYwDUgTqqfbe3RDiIzhH9UY7DiV+63/2OY51mfpMyDAsihiI
ktY7UKbJrcbnianTL9EXtm7f5HRkX81ACU6ZXthvA4krpeD+GtlI9WnHflxCya9x+nKqRzQQR05M
WV+/rtY0+wW4a0FWBxqLKjZWPhSNnwT3Ur+6u59h7+N5kDTE9mJSkpGlW/afoLViECFtB0jvelLG
D5W9a9daJvJ19omo9QF11FB/PvUqXiC5DwDdxY+1JdyB+NPgrseP7EERF4y2Yd0M2A40hEmGoXvB
jqDIOGC2Yh7SLCM6nDYZSVgxuATGCG8GnT2JCP/A46sTNnjofYI/TCYDfbRPl94mn9dXi3iaEmdg
JNUzKrJdWGHiTo255XElmWiLbDwGHWTzSh/QcNGLgzIpiMWm3YptZpB0n/C4xD1UutfNcn0ej66u
dyihLTDNY7EBXfVLejAViEwnM9WQd5MyjrhaqPY2ZFsGEwi/VzGNrZun83gibkQjym+cZf7Rmo+M
1GVEFKF4WD99XoTmZgKeDhR8hQMEOmZfmhArCRxXthT0vRy9ezAEFuWShCyhtU5Y27xBHi3+qVRT
n638jc6GZHH6DiduchvRpj4xJmPSFttexzRO9C0TTkJnNlweK+WYuM07yGFIqUrcMFeKdIEoyI6e
r9UINBjUb8wawHeAuxGfkeSRMUfDn3X316LCfOhpA8KF6OoXDhzC7IAKVh9wKcDTOPqroIrRo4BY
I7OeaMdxG22gP2Ik43RrM/CsxRKcgqRSX8KX4mzz3b2FfoFMcdYCwPUV8XpJyRUPF5y+tIo2ymxB
4JOnNAo8eppluwhw25fNGHfHLa26SRcZLr0mTN4dBOkMGqJpTlApUvscG6zls5vhQLfaLIUvVYAG
BhVuyO3Qx6Ay2cEmKqG10Lem1botzHcoobStmh75H3wzRL9nn3ylbW1fMxFwXbZ5jvXFcsSvjFe3
WJVH8yhWLLmhM/ojfULdL3RVtn6mYZlqafYV8t8opAHTU2EwLLUmMmEzz2XB/E9xM/U8Ot4rQNS5
PAYyuoE//PCyjAe+XT7EFF5enghZSFPXMTJawBDXgRWpbMEiAHLeOky0SYDDc2/zlUaymSFRtIxO
G4x7LM20noUxDYxn/fSVgGkYcfoEeFYK1Us08ZW+3LqM7xYy6vOcqESSVNxe9QsJHF3B8aqC7As0
RidKLmgnaLte43AwymPhbeqasCDLRJTgtNFOCZR6NUrRlHEDr/NAud2MiinLw+0YwvB6bnJ6lH2J
tkbMKovxGhTQlxR8/z+MdYqjmt7P/K/00jZIr7AMD1jDuWHS5XKJPIk5RuMKGjUJmTjvIyDGxXpG
TlOhneTSDc4OPrnXOLWlJQhQWJBgPF03O7aB5JUEMl1LxGs26PulhqyC+geARMINv/kjO+ZpqqAC
FiF+8hkjlq1hwAhyyKdclDVOpvvNUlSS/TV7G11vI3a4+ZzaDvhUcwM2levw5HJqbnVWBo32P5ao
6u7YUheDc4LaiQcUwEGUzQPhVFKNmQ7MkpKzwDspLCChOTYxQlg/x9LKAA17UJTl+EHSABw9TGX6
SxF9uAHJzSZzvweDBfU0ih/ZJD9fHAF8R+2ixHkUIYVmwdbP41Mf1I6xaw1FZ1Ox35BuYYJsfC8K
njNrZQsBHEHXblYnx+mK5LZzcwo2azFDpgwJ8Ux7SPwXpBUcupBsJw49VhuG7ZuHteYleu8AmVHo
eW89g5ib/OC4Kig9wF8iBACnJz63JwtTiOQIlzUuBqDf8CMxhFW6vs/Q3uJcU5NZ4KsvJc62Xdfl
xtfPHwqvXThFkZrHksI0iKcz/p93fRCh4byTPohsmCivPcnr4FLN/yMt9nQnvEP8b5yCsNLIWxVs
WQtwLW/5NuVs/AMDJbfgwL0Ypk8321kO5AAN9fAu18shhpdmhHJhAuaGDPQ7mL59Egu0LYKw0C6w
14Ukjl1Q83w3jZuTHrHDc/xxtnM7ws4wd765Vqh/Gv6Q4llVxnHIx3t0WUds2LpU0DuRL5ZiIH9M
x519SHYh+0rbeSTLhaPezgU0/AizWlIbX+guiqYf3RzEdfHs+DnJJecuTuhP1FDrn6adj2CYcLu5
LgvMZis8nfZORctfOBcTZNpB/c5eOriSt6rzJslTH/Yw7kaWvRemuwDq0tVqTMH38IbaMOZxBznC
W6GPYuIlaJf5235jPNgiFWWEbc3fz8jPyRVfMAEplln26i7Okn1T/WfR28EjYKVKQQMgk4rsW9KC
vijdgJUdAcDGJ/poQiSJY+LT3fEbfcLpbQ/t5dDCJrJaeJ0sEBiC2BLjFBMpgz0doiRK5QbMpqAl
MQni6HlPNUuqVLeZmyFdXvpf6g5is4mKvzpht9FTkPXoGBdIBEJMypzmNDzo9fG3DqGXnMYXaYpE
3LjkxvcJBVIGeVWg/Ka6MewEyOhQRtzUDehItIixtgPC5Dl+ILdH11A00x44yVN271eq95DKGMQj
PYvJX9AOtYoJ8BTykagV+6YMtKC/eEo7a2ZkaRD7x9ITMRtdrfmVIBMVZqIkxiVr/am0NZUNhZvK
KujN7811KXm2cse1wnwTEEtM9TncouIEWgf49gZLMUJKO9FjGvfMGBGldNiLE5qWm+7Z663OBJVo
CE+mRKfkjYAWGFkFJO526UKMlsaVCmhHA0o583yh+Pz0afynspxafqGh6xqulFJ2h2DT+2ThnEWu
U0hpPhChJWhCps7t+kyPxfGciikXAjScsiB+DTwG8Z3nVl3w3Bcy7xeYUDSZ7Fv+KHTGYVbhRzUv
LLEO1yaeq1cUIl0OHYOrsahOSD+MIDau4+fZsfcX8dzygaxtTIC4Vlcldr6HRTvdFd5baFh+xgUK
mabc+yKLiJcyNjbJJjliMcHX3YQaiNHP9E8igrjNrOa46cctTGnw6R/a2VrBqDDvkVLfGzeQ/ZeO
YvgUucD+nxVcrjNNZYDFEV7ciMfMfSOiXGe2DVwv7UtX6zAaKmYW3qwCwIVbbkiKrdelrILMqIco
EnVpsWLUvR+b/cLTnurI2JUq/fzcJ/tVmeNJQJ1sgPJKmQtiKWtqQTMpBybGtW9R5Jv2J8PQ8C79
eZqTRFRLdf+iXobn07My+GFLknwO7kUEU+oK04mjH9m3B1j1xWPSA35nVHdB1cL3xbcD81+AEk/Z
sXQR/e5ytetswJ+VLRpn34mapSqDjVutHMiOVruFnEJN7sv+QfX+EC0V6HcFpaFd4IP8+0uAqMDy
9QxZdz19jGeivTkgbbZEX445h7866ZFuhZC+oTm1kF57XIPwYt/mksvYTIsujPZZt1pgCOTawI1S
tsewji8tXti43x25M7fRfoC+21LIcmLcujv2cLJkurYQAubPC12MVemweyuRA5EQgxtOtaxcx0Bn
xFoXECIsm2qpLSmQ5kppkLNEzMBfZxATfUtC9bwyzSZpcQ+tDTdcauKOJjlwIJuPNSLJJLZpxuaS
Lb6HClWmNYq61VKyiA33zfNIy5MyrM0s7yzcxTCHYuDUF6TPnJgztq9Vsw8XvRwWvU8zi0mGyTBV
izco3toTSNpHut4tUDj0mm5/5X5AOTXrLNGnnSBYoD1yKiNvg5tv+uSZ44dpw4W07ruy+VRZnIHq
8/8xU9XDXxmeVN0uL3MMLL3TzwkqnZKR5d+ImNywI8VxDT6KJ6tNjrtGQRivPSQpelzW7CCXPjUo
STNYM6zZ2FB+seC3vNNdW8Hk6lIVxFDafmYCVj+M8vbwEzbEIsUNDl9Im/PoJvXq5BLNLJyw4m04
OcAe7v/oVcV9Zzn3dz5Wwid10GHUFhNDySg/riKUGNRYC/tzsIrDhZC3iT2CK60tQ4w8UNKkK/4l
hgk3AjaFLyhUv5vpBG4sKDZPbM/CCez2IU7Ffv1fIEaZVwCjdWB8zYqR2n7VrSK2DAfwPKvK3Og0
2AMM8aI56EXEgAKASVLSYCdgWZV9oXa9hoDTNo9J58MDrnpFYQJhCtmo2HujLExaQp3VCI7qmVsw
J6pgAWACpMNdJAU0Mn2s7YAarFoDvm6V+uOdYhY0HTHtCyOJMYS1I5tV+8XshK9x6fttXSjzgXmP
bHR00qYfAX7/uLRalsZ2G1Qehvv/ziZFp3iw82ngtxNDBUsblxdyyFPqtBCJW1nZAjrA50ntK7QF
XCjbU4ttKgsDhXmEGykwugGJx6I40IWYbM3L7tpH1b18czfhfHVNw1wWgsR8I1Bv5JDzOW49I9wU
J7Kj7dbG/NtoP0Q8zJ5QX27q5+sRDyu86asKjUiBCTPaswSPDubld2k5S1KI/5mXN1ZouMcyasr9
+iPcHB2jYZnU+M8h0RwjPwQfmurYyQL3X4nVCPpYpa/T69/O/DlJsCV4aDKbTdpNyI1z7WaYMJTR
0DXIaXCgJZz29dcs59PT58y6rUL9gBa3n762p4WT5dOJH7UMYiFZ8FAwxPuZGqB6OKaEXMT/NoyN
PPG6idM+vUf8Dtnf87TNwYxNspqVH9LavJypqH5bdus2WnNAaj7FBKG9sc8DSIUMTpXt8J6hBXyr
2gpVS2tRFqUzRsGgz8LJRR9QN8IaEsf918/kVMN1t4Owdxz/mytovro/LLQ8WM2tcDiyziGnJSHe
+twiiDt41CwgxaeOrOL2FQs0j3INpcE6D3yuymO7raSeQiBNRAe6XPcMbbBFLH0tnYppR5iSoTfe
GLiiJFv9DbqF6VLSnfSY2VXhEBe/oB9trqDKEdOd45fP54Udbn0p5ocDJdeHdtNIKWSmUaHlK8Af
MhFtIo6DCTvUHxcwaJ8JG2ySsDOIgUFmuZURLmQduq0H4AM5xBTb5guWeLwaKjtq4oqUM5F9iXd3
8Nd5//Q8IW9r6HVB+fDcFCJw78iQBxZqJ5B3lNaLU8xwggDHQ1Epac6LB5EmLwT3R+bF9QktiYQR
Afy5tph+UJHZEH+WkK04s1dVB4yDk2FikRakj//n6djNbgLRZ89WmQOZqx/xZ1ZCsUvX2w6YmOux
paEJ3YZp5t6EvZ3efK0GN/nACUqMsTU7u+6Mg2trfelrTPgsixDIf+bWJ4c/GU+8frwRpreDDOhc
VNH7HsIcEuZ3Z6lC4DCKbWjpjCg+UprRfuWM/mFfCoEjetaqe/iVCzoiiygBYH7Vu4gQSEc0Bavh
HdfXgdwOpYNskkqZTzCpRqAN0hga5VeKaRg5R9vAKBoeeJ+N37dYC/lYWMSMxpTY63+vJ8Bg12/r
Kn6t4lIwL5OWHa274/uFLQUTp5FtFVXs5cPah/8mFhlVGUnhn2ubjenj13oAEhYjjPLPLLg9bbNA
SpuZ/IgvCZfskAyxiafOaVO7Y80MwyEqz5G4XwVxfXdiOMKOaTWAedOGaNaYLRpwGVqQkImOpqwG
3Iod0npwhew27vVaFVRVeirPR1OVY+Cz8iVtNk64wusSBJr0iY7gwBBM2iuzPlfSE90UiEfmYRKb
IQzaM9od5vbysC2nxhHQ+YEt8Lhw0yh3qW8++AIELJUjGuTOWlIewKefWRBFFrEejUz/z5x7LejY
CBl71aBFIwD6Tor0gIq2hiUE5rujcYtD+e09iEcgWPahjwhmcDyHqEE+JCcsmixn6wAO8PUNm9ZE
yM1nFLP00Q+EkPHiUkv8N6uyD+w8vf2XVPiZ/fV5n6X4XSogm10fkKBU/FMZ7Ey8LfO+nl1FQ8BT
ZpFMJxRDCXs21tXXAurdxuFT/2chg6YLZKfkGgkbCHKlguUnXQvahzeg2vgDAMvda+smgyZ1tIPI
giaWL8y8dhBpsYIPMiirK9sBOiU6pAoQdAeCdJoRGoQLLm15sbC5aBeDJD/p9mcuewgcJuAi+cY4
D4LexgFp6BUIgAEKDMogAnUo93ad7v34i6jXBBjgBdilfNz5tUCli0HzA59SKQRQruD3ZHzEphoT
UppFWzP2p/ndfIobTwKckW1HJwn/ZxcnO+R2OiHKqvIE1m7WLa6D9cFjIGQdxlK75qWmaYYhPqUF
p9rR+ZzagFQhokqDFXo4cVPSKawLqSuQ7FSR9vkqbciWU+a8O4G4oe3C9jqo7zwO+mc3z6hGpZvI
ClvshgnZA+eUWpzDi0+RkBRvQGhUzNtAJqgaIfHIlFZ3U7VJxc8xSar6AWajCqWfTDcHV5vqjsS5
47sD0WBC1Asv3NABkHuF5HMI2IVO6T5gGuuGcvMo5Pxm5MFB0GYUjaqPccyMuUS5KQBnvSQBeK0N
3+reh4vtwsTTc+CWQPcbXyMYbGI+WiPEmvA5B04/g8kb4Ltia+x0+wFYYoRvXYcfmfdq274zFEi5
wudtkUpcMikHtiUc+TEhDIvTyAGUM2xGiS7ZVgCr9RWhbcDgH6Vy9hCFcqffbKUFDXe0laPZjQv6
OsakU0hCpdPMPY/6SfFxd/uVdc5Qybf8mCA7OT3GitQ6+Cta4oEG0D21Y+/jD0qA4t8g2Bj1okCL
S+hN1pkEpr4OvRNYp3kmdbgR0NITUSWQAVmrjfwEBPBl8FsgnJ5jFuTBocQyrU1Ws8Pu0p4GuwTz
yC05JviWraOBQKI4dZsnArK4Gh7ckF6usoyPDcsZ/KJT79kMqT8uVBc8WRky8Zr9Tly2sN1rBeAH
fDLF/G5I6lSiyFz4FqsNaJTsy3PUUku9QwnS3ZRgoM8K0H9rjM+3AX083ExPKaDOzRz67q+iLY36
qEKNMc6VmiYTILCmQxmNYHQznbWLoBs8zQShIAE++zcsQwFIMx0NOscHCahg/tPXQJ4CUHayp/wq
VXVouM91Q9ODdCxISPsbESjw/IoM/LnLNwCk9D+HUjXMlOW2jMxpfSPh7oYAZ5cR3c8WQclzUepH
oObeqHqHK4shHk5PdOpZW9BxiOi5jz3VKU3+L+kMSHCM+dHP/V4nOqe97CVOHF4LDhCuEkddYs6o
ViFAGl3RfR7c4aXztDI0+PwaNvYSMaWJO9NRCZWgTOhK1iU/xl5bX7mjcwmy93CJxaMthj6Grt6A
uTe0kIF7lP73KEEAwoQX9TfhfTgWm4H7ioWjMEFbNnMiPLxR2wbRFG04aLFgsaTo+sM2wR4JOQcd
waEqD9VYu/1b2n2PXu4W3NmYN1A8OiDerlY+ykzo0rbAkOI6rN5jh8+JxEM+Rl2ckW26BE38TlVw
3i2iAjMEmIkM9YoLJPhkjo5DTGrjKZXd027BBwzrMLUdJ8FrwAii3XA9IrRWqPFIGCVwEzBzd28v
/pIkTK1azCmPEuGGRaXtzW00os5f84W1zqpUTh2zmhiDSitFRNJqm2h7M6QvFsnr/uGcT1koWlOc
42VOhVBj8hAWHnok2azszH5B6ZsBImni1bt2BZQ48RaXQnYrgSIp5/qvYPrtjmYRFgvf4rlMq4i8
KlJVeNjYfsxsVo2wg8ZhQ8z+hNz26lttTa31R2rx6qt9i639NQZjJz5c1RLTM/8Il/R04zxjURq9
WJWhUNsOcIXGyuTazwYeYTLJ0BxW1aUJYHdUqH2mNDBxV5KIJ8ciliEK3LJTIhOMWEhvFPMSMYF+
O92F6pEdtdSyvg+CIDwoiKhw1+L8Knhnqjxb6tRIJ4P0h+roXfaVjr4Nmc73eKRq+bicG5Is90wT
SkLo2dO2Dzd/TS1AUrESVAp+NbzoWog9PvpgPErwKJ7TvfXm+INXCO5hzghytGucJ36N7AX7ReTp
5mG1wmiiPfXLVeJ0dZguqxeahKJP0mVwj6qVkE8hWWUMV1B0gxqSEo/HzldHQzd5F0lixrIPYhBO
dN9HACXCusdB5uPt3YSegT7Fz1fKAc6BNjGGJopgSkg0FltjZgfXXbFORJGW0fs4UjQxJfYJXgy3
3ZVuJJFYjmuLsi753C0hwF8PJKHPyQA7ILbDF36BEEaNIdd/pqLanc9nTV44V3vFWHofj65TdC+v
hejaaW6RWJowzdjco/M3v2WVz7ZzxkyqGIKY0ivUiim/eM/k6955/GGhU0TUDeM1iJJJwvZ4MyRK
TD1OvUsxGNCCr2RnGeyozvC/vO5nNzV1/S7XejRY1irNEjx7Z9RqhqdHNHKiDQJdYlvuOeFKBoFh
ALS5KwMWyUG2E8PkdlOSN3WY/cB9yinSKIyYlHKxPccHDkR/0wdZeHavib38653dWxCEmlZLaM6T
qwkCAuSey+QPxnLBH5ylYxRtGALjQPGd7XqJpXs/hx8EeVZdwoBhjDFbs92sL4ySsSipLvvBzgZU
KHbP/LGfXwrXkUk7ZvyhrPlYx0KHh38BBq9klVT1LGVlqbEsRZvu2USji8X49QraI+96jQkR9ZW2
CRtcilzEJKnEIn0JW9jRvyncRROwTVlDRyOUb+amWLnQdI+21zW3vqwKmuJVH4iRVg/UT9O7qnn0
Sm5EC9233D6WDjLUtdrfV2DoDM4M8ATJ7QqDhDcPvdnkMc59SrQ6rs25lEAOAnGe/VwT9TZ13Lw7
3+LeDnU+h5Rq/1b5TWRYzFG3VRKgHm+vxsbSwge8rsCz/0W2zH5NKH76zGmr0GDw3C4NOANh31bY
MGJG9hOzpodIw0IlL/WEKa7TtYjdG+b+4eopMATlfXPy1au3GOLr0RNaVxY3kH+o294CR4oioPMY
MuSp5PLW9lgMBvZ8wO/4LDDNDJSHUDNQOhUmprtwegEbJtlg5b0lbpW+/lN7W0Em51WWs0cPbUht
Rp1vDcvm7oF2lY741cH470gaUTnhiA1IAJ6XQ2cqTEgiZyReFmSgdQkXGPTHtOcAcTuuMHaAQgJY
LmVCgIGTtcfCXMOyFrUDWCqWf3Fli6eX3WPY6/Wg/l0TxG8iSeSZdizVGRpeiOcNCVy1GYUOV7q2
pqnmMry305i94xmeb2XbXbq87YmBI/YghbtY3gg2b8loSuMBg/GUhYRCsvP3TuJKiaQKI3fqf2sX
aoJT88E8Ux0jl0qIkxJtvye8r0N6E5BI7ehtDO+uZPm43xonvB8bnxk+6Unvx+m1EJgkGOD+H5oY
OJRd2h+Q904TCV6DRBh8N9tm+m9IzkDXZtv40rO9Cd9K6t23Cd74qV8jApDMnWp2SEQCfPOoxwjZ
/POlbM5CGwutqeJk0q3U5Pt5UE52lIX2wbJLLvE+2icG26/LCIAkrAFSHA9+YvgOu12A6hbxJrvC
8kh6lP2X7UW+1t9g0Axc0aeYzfK4Ic/spd0KC4qTEvcLJQkaHW3mMTKD61kDfiFMZJY9NN5N76vJ
qnr9CCxYg6ggU9qW9qcDkuBWEgJVBnSshSTRy05hOTicAm45rULheMeRqqMiW5/PYvddlzTU/jCE
UW5fRUV2cvH/ANt7gOP1PcnVR9B4ArfP0gKk9AFeq5X+V3Mcgb8VvXEHuq1dGJkr7QHm1D5y8nry
x38lx2Ct2xCX3BxscoS7/WtxuADyXUqZNa9FY9a/WOuk0ZWZZfOr08RkOZvWp5lDhMAGHmL1HchB
CEA6WKB8VmfE67x3t1U7N1hlptygLW2BZKEgiHjAJlSQPNo1xR1wXP8ov3ozJNDfEYfLOC7hfpNt
4BkmMuOxeNWR4LIOPPgfsBYv3o182rJYiCCdm2lYESF/uSea9MvgxNck4ZmWRLu6s5rWmGJ9goQu
cTyuiF2HCPsMvu08s7gvYNoMy2QYpzf4f+8u4/cfGACu64F2UP7xEvRecHhudLbsmiwBihnCUZ99
gUFx9qgLM5Hkw6TLy3VZiS4pVXZqOpF8hQun/4743U7G02vCtulEwyi5k6ez+nD+iAcuDhfW8n8a
u6shq6egpU2Z9OoEZI+6PzxXl3Arjd7YXbkfLtAFe6AgmNpc2cpn7AHL3k8wxLqz8k7UqerBcUJx
maJns7nBFGmJR8UqaPGG7MYwdbQ1GhBcBP3xnKVYzlOZhrmVwxakud/FDqQzeIu8zDE4zc2jy9g9
s3x23PA64AdYakuLkqVQOI4PN07IN4MeUJC91bXAP7hXn/P1BapvHYD0V05waTP6EaA0eCFMahPS
KtMi/6TzGF50TsxnD70KQu0fnkBkAjMEasTdpn1foVI1v17D5Lex904ySNgyBi+Exk5J762h0xpU
j7MNlx3vhk4dO3mOV7JOhtcOv7sS0mdkeKqr/jgmJ11zONmE+Tv/gyBL6POp7E1yWZbvdxjaKDWs
I4uufgXrqidCbyuqKfhZVntbHu5sOX11PbkgUr63KYZNU6cMlgCA/7t3pVqhErjNyDbQ+K7jcp0l
iBHPvHUu3fIU/EJGd+HvRCvUJQjNfrooxTlq7W/MWM5w2NIh5cVXAoRIn6an6C23mFWp2StMDNKR
fTC5AelSznUoBkQbqUW/P+E7JXpzGfae2VoF2HWys+tx5zB8eaF5s9+0B7CxvpZ2UxJGe2Fef7vw
EwRJ+edc7GuUdcDVtkjYf5Lq4Ayz6R4uZ307CNdcqrsluVuxR+1HvPSrb1EbLfOSMbRR+mGUk+pL
OZ+RACIZvfxKQRsVhPdrvpPjKbSQSJ5MN799JtlUmrlWxg3u8cZWageaafzDi+1elk0drfhLNRqe
3l+sYTn8Z9Lc0Js9nC+/Brtt7BSf//sM1onN7eFc2oMe6QRw7j3sQSNTvZ8NYEF+ogSSBHUbhY3B
wUcGbldf9IEdsit9ZQ/HmpohNk8AFw331SIK226KQI21YTIWHtMvE+7MDOx5m83cdGUAAzYwkKCz
MhA1b8IxfYjw4gyqJV7fZ23NLy84uXHoGvwLW5zvflPsPG0X9yKPMtm5pa1k4r2oXCVSNdT3pKah
mQzILKN8XlynBinxfcjY3JY/iNgi3f23Syjf24E9n5af3XYw3iJdOXlkPp1OfJWDAChP2O1CV8ib
hvnZCbUqPvcC0CsfL1qvMnyLR7JrfGCpUKsZBbftou2IuFsR1Cli/6wgXcCqI5qAebI8zdCUyzcz
wL+72JTNyzn78e+UpRCyEx0jXKtedvKpiMcOeUbOxazYKJZq41wKXtDv+EIJTeMXHH47/Z1X6ljU
KwSYOpF7YYN2vqgrhEYjuW+CzoOYcXs2WcqWk1oRXpULOxcsUBAg1qaUAKtmkgOCqr4KLMiiEA6i
W64CCtF02phdazeQHHvFr4XBW+tNLD1zY/MyAXcL5R63FJdRm/prdu44711DjsC+ghRlAwD19Ysb
IsBzfu2hLet5M6JAiLCxjWeMD37JCylR8KQuykkzosGV/CuwcBBUMIEIb1im9nnUO0EEhDkkXiXD
cmO5xSk/+ZWpvoP6ghPXFB9uK4D1MLnRpycXaKXRHa0E3xqEmJPBUHGO3JfScWZIXKWUo8A0jgWW
Dym83rGhF2F8UaIvo03oAI8C+MFEorJjxkOoORg/v4XpKT6GCFaFXZsQGN/2hAsuQvieHTPI/mge
iPpCY+raTuyDVMfj0oOLH3ahRxwg9FUpfhWZJMYkWkjGwHwUelXPFzXiFgUmXBd8DklpoTa1qNmf
Xukm6YpV65PExvHjk4F8VQHY277aXZVfMyrTfTXxq31u/Wcdwt+uvPhOQWmEB85Y6ktEZuE2VPaa
QBcPDW/B69hZV1XLz/1jlioZIXLqFqeYutrzlSg010MVUEo6PyQRFNWq/8MF2SauutGaHBoVCZAa
vkmNmVdG+8hECzm2Svg9WhqHii87gSDJ15ocAzReorbI/z86mpvFKjlKw5eOTWmARFYTgVGPae/U
l1h6BfaAzN9qXuC8ioy2McxcLID/W44Ug9GsNbREeA8Cb6sE1cA0xio436iXa5XRRp1WeSmuJ7+t
xjbJ0ow+20J5ApozC9vXqlEq7UOl2dqXSb54/3g8QXrR2TEBMlWT7i8qqgsZxvhG+UGVZAJr4eI0
wapOSL7ig7at1dPFJcB0Eo6kPhoBEsyLD/gNUAzOKcUtTgAF2lLG0b26W2/vVMqUq9TRpMTCSl9J
AQ0btcEdFLnNBWOCG2mGrvWb8RaxbKfsT3b3T7R9FJgBKuTyomvIECanUyb7xzm3Oi/Kkic5Fk3K
d6F55QdEkUAyjWt/xLS7DNtWh/2mEs1fQ7w3hrMb//Hf45XhLcLL4oAw2Yw2/pUkl96oof8Rtkss
pynT0n5/sm/9yxPqtd/wyxYFhcWqyfmxBopb66zmD2nRsJe82qnSAV8lBSRySr3IvDWdNyQA6CWg
XlFRI4pljQ8DjpYwiecQSmL4uCWOCCMw0L9U0B/zbOBf36puIp5ZoF76EqZ8PhKRbX04wuYViuU2
8/N5R6pkUG41a/EsiIOo+x2SN/5fDLqFR6gxpgqMW5p0zzBYYOfA4glGFoV5uMiuzPgp2+dAaNBm
XSRf6vy1IZSkZ6bxe4dY4yaz5ariycOEegUkVQnOejAvueT3FEU6BC3yYRJ3X1YDcjzgzksWsVF8
2wacTrWz7J/yjI4hTN0hMtryUHHWpJayghzOBADsJ5yd5vwmpxR1ZErruttFNPTUNIjLDCg0kLST
i4CLZ9PURuS62NmBSXnnF8MDTIFuxC9gaOVZbAWuqcAOAyuwgYznRwv/Ala14CR0FwKQkwWn46ky
+HzotvSdCUg1hVxv5g45bFiwzZgX2Z5T/96C5xyupsiS3LDv6DfS4jIj8wnvYJtn3F4F30tXhhNq
qS0YxXui5KArvKax176Q9vA/+mZRGX2ndkn2+z/Iu+jIUNyHCesjx1bqiAArsYaGdl/oJKL7K09I
PLwADkL3d2yBJo/3o9FpQ68+qOEFegIO3wGxn+0klOmhojbEVBbpjH+5Nos5PeKKxORIBo6gAvyN
+CxEWnxJIYiEI1zQRLtzAchHbG+TuN5dy2rb5DnfYqCmmP7dJhTO3BIdDMrPnn7czNcZf8J+vdDj
eJcTfvIheYHFR9iI/Nh77xaP3EQwndCSo4yvnpQ/iRTPqAt7Ll8/WPZWtX34rOb0/k/DABkt+WCi
SVC670nHR1lsO+qWFVicY7PWsX51NAHA+irMVdkrN3BCtq6magxyi0AAs9IhI2HBfnRwZe/6vbb1
UILYhGgiclASpi/76yXKfDpi+K9Fsrlp1MyFYDpOw//2TqjpV9iur8TKH9BxZaVMR1CvDALlH/rl
ZMhhJ6YjW/LzFxi602+IHCzb0T2vQykpgmN7MhOduEvoRqvcS77Bzup2ogvC/pcMkSQLzxM1OoVg
VkZytTV+rJAWjsfP39xftO2qbh3IIF82RzXEfAGuHqRVMxHkRE7Qr+OUKw3lwxZHcFXsIA2TOqOH
rJJpO2u+P8h1fNDw/WYNXSM++bQWlq30xFV+T4qAuFiVlOxSSv3WDdX6jQuTJmQ8EeEM2wob9Hki
n4kI/tRvVTA/SKjDyRm5PConWes0gduqA4EYk1h/f96wndDfxIMWA3q08tfcyl6X9dTRcjN4j5ov
nsBI8qmsC3sVQjqJxJbbu5Xgsov1W4Pi3rh6uf4mUTcgcCQHXmQH46oRWzCWrufcI5xP10E1u19b
jAUnOQWZJeHE3RroCXWRq3qmxKkqkhQXTe7iOCCVHf/jCaPMp7x5evtBlb+CGnez4kH6PL2x8Gje
dVfy7X84kn+NuP/J4/6Xdml8y8a2qnzPzxb9aBgxyoLsej7BkeIEeccj+XqAGRzJ4y0ftwFGMHIa
YX9eZiLkoG6UwbAYCrvlaVGYdteLVGmA0i1bhpmF56G8yDDuPAxvgX9hD10Tv+dETC8ft2eU0uMM
qYshsiCp3hb019Ee0451BYxQDnVAS7IH6PX+fQdixymKJ0iSzyIt4DoFAE/+4oZj26jYMS+2jTBR
h3O2gtqMQ/e8Eym3HS4jJwVhv2u84y3zl9z4CtT6XluQL/ykMW80oUTVfKmSgubkywrvaOmrZilg
BGdo1ykrAyMr3kjgu95pnf5+4ffqVCKpdghazhmBXhrq9zYOJbFIrleVJfHn7VQVwmz9hVe2kkEJ
z9G23K5sWSNdgFaMcyxpOUaMxb3Q5aKcYB3bogkNZnS1alXUmIfKkDXwz5EzVzMKFcaTmgEkNSE2
vZpzXFgZlcAWwZqbwP14xvRG79FKo32EMGY7KZLL8tovNSJksQ0SKqDgaQRore2Ty7YShUpVnCDV
KktbWOT3xLSHsbfhP8MfOWn357C5fbqIGISpR3kvGX+fZ1RXhslipSml3RTml0sNYulJLxfA4P0C
tCPJ7gUKGirCWo5oZShoY+Gyq8LqtGhklGlkfXia+iHxKCHJDmDqx0ZgeoAnoloQeQXALyUfnsme
bfmFu/cFIsUBFJVEKPl83FtIx3Y/IFYTQilIKP7pr/mHe+qyEnRtbujzpQ9KNo1fGtl37EsoRRNJ
X9s8yYAGF/JgvPWO3YLH0//RVJjdreovvyyEXlEy5GVmkof/+iCBsCbcFpTtH8A88wCvUKja8y6p
GHMf6IxuX9YUgXEJhtPNLauxdzTCy50m51bR+g5mceeOG89Bjx2VxosCUoOvM4cxyKMy2bmhQUFV
5rXrzlST3YSIH1m38tj5gf6yFFy13/l/ZajITQ7p6YOmczTMgDJjs012dk4urarWrICBMpVahCxZ
Z2LkYToQpJyU9GsukBBoI86AbdGN7LEVW4pfqXZkIBhnLLTAcy/scRCX8lexFOwLHC8OpdZq4Of0
l1LlfyJB6Q8GV8d6Vp4ovVAxl+UGbU6TMwa1w9cw1LAs5ONZtnPnevKgLL/ZMscGlGE3vtOdVzFS
NbR/ybW6K1jRTwpy3poaWYECBH2GX8xClHbelvGyYjuD7LqtM7qzG/jEIUVbyt+UoGil/MJqOtCB
8rPbp0jwzkyS3AqcKqey/M+xhBcyaA6+OQhnIeWuQryHbdE1RMjxQN+BzwIm7Z/6DBOWVD32Qu+W
FLq61IlzrRXA7caPrCTKxVR4TdIs9YyJxE+ggUyK4nbbby98rOnFJt7pD2zDjBsxoT2AFGjgbqBr
y+TplBl7nzyfhKPlEWEFv4h5wnVYNE484BIhBRRbzzawean3P4NNpUu8Oz7At195mp/IpqDCZMvI
b2K/5b9xyVyEEeZLixBWW+paUMXMarkycFXAIFrSKTLQzNvGw5/kE8KnKHe1C+ODs83nRKG/u9AG
r+jDJeF/Ad/KqSvs0HQAk7Fak8Q1GyjZr9GphmDmXCvAfktzeg4j8nQQbbSvTvnXVDkBx1h3Ff2q
7DLxVBzsiQylxUz4EFV6S3lbWTfAIJfBmDvcxbhFcepX6po534yPbEQw3TWqhiiFeviAoG3WkMn5
rGQYR9xQVgjR4d2GLEVCMyKUgt/BUYmbZgpM1JAcP5f6iPFNAM5a30Me/P872vT3be5grKK0eamq
F0smdpK2kb6qO/+M6w0CXHtEi4CwBqEXh9WxLVYtnzkZYv3oJnTumBaZLaVfI8dBD4DsVuBlQFlU
pbs6fcPiU+YxrXuPrv2nneIUSXIjZMz3F1A2wH6z9bnl6/zVfQWc9ubFg5Sma1fcLTLdoAfqqdFd
gyTCcJX2yXWzYkn9n9X5M4bLVvbiJsF1enCkvpHhcYjTxQS9/GWsID8uaTJx4HAh8JBmF4qOldfV
5ay/0BODTxsio4qlBb5XSATxs9GdTwp45wFLlBP6XBuYfP3jl76mwoi8ZcrTD0NMXgGSDLzmdBro
S3FlvQlhvX4C7P/7RNS2MoL8fZl+F/fzB6Df5YUd0LI5KFO1PjihjILI9LQMxndYGLEbvn+WAbap
capC4Msjc20+ZFDU+f9anhodLkWP/eU3JNYHcochZgyWJrK5gZjoGr8/9g2X6mp1MkUdb5c1fJ7o
5ddUp9grRl40+H2JRpc+KZqN9E15nCEJ2TtkPP6A8p24aXQuafwhx48P5jyCPFpFlf2jAqbAs+6v
TpZuidJGMtQ1xxfhP7BvmahGG3Qzco/luVTjDw253bWSM66IaUocdoeXLLPx0PjU9Q+JTnQvTozt
eN7vZALNcsNLf8HgeEnC+LdfPdMqOuD6KeUrXNm6ZkbjzlD8IUComf5Pxpz7vLYLE5vCDJhse+uk
DPvqyvP8mnBRIW9Z3fW9GebtnPjaIn1U1dpec9oMo2v2WQYL5c9YHMUPLbwU8BwBzo0JazN+ub+h
AEHjpRE3EJ0pYNKwN+Ab3YREKDWx227SojfPosUxoBsW+a80Ca/7HkQDD24jyZSwkPAIcRbLgzCe
HTcindrKCZGL84/c9fDbPOo9nMacZbJC3zGH8ZNamZx9ig/9GTC1gCdocplY25jLY3cZG363TbXh
ltcR9MtuIEO0kEkd23cLjHkfhhV8ZRSexLTjXUnxtrx9JCfoC8mncwal60FO/gBEma7gTV4c9aJk
mYrvNULTJBPHSMwxaq1OJ2NMh8f0j7cxbLhVhR2fR5JhmS1NOWuy6zfR6Y26DIa0Pa6TBBC4mVla
jg9Tz99Nsv+NGhFqC9JnjTDu2B3HMD3d1MTN4TZPyNdpUdznFBYIJj7k0fK1MSkpntlgP8bgoqaa
3DSn1JNqX4mEovJ2BunYTdZYVULsdUrcEPjsuu9vdxRI7YL897fp3a6QG+ensw8A0oFM+F/cgJQH
wmLHPCZeOlK6sVh2qnFjnjCsEJMGoAMujtVZcuHBfLmUFMDyIG90zNVpfXeKvZ/sNvAlrRTHhfUs
WNtHqklwZpdvVkfpJYxaRsgVwTl3Kc2LCVPNckXnusfIOcubnKR5H7lAEXw4iZeOKYMQpVUdWduT
yTfrCU07geuqWBMftyDWZXPKiT9t4AT8GS4P6R4PfIPZzSwT7eBmqfZPoauQhTokpgQRdgxD2gG1
C/T4ZKCP3TI+iFigtV49xLVvkqcGf0fGn1qcDRTCC5oBmevOSjqrF7Ov6ZcaZvjvUDzMbWe1zp1v
xwNmOboWbwbyYUqUtBarTzSqOZD2opS4/Yp/weJhA6FhWb5lkfgVgTxcDYL5Au4HoKHpSdpqUexZ
GQSaE8XQhvcmJZEorJxio424TOtesgaZfhAfRBBxPRsqgFUBPthFR5Xf16kjsCma6IlTsgtlHf5J
EtRKPbVkiTlqw/ZDeYMPPFL3ztYS7DWBll9k+L56hIe14/OCoGX5CdVLAcgENuQmbJIHo60a+lin
6AU2URd01T9+drnjQ53Ue+ifOj77O+XYsIgOu1tPd4IKv12wu4tWhZX/U6RZlaY0EthuVIPNgITJ
CJdnKRQyl/gSu77wqsT68m5iZonFXKRzEUO88fhiB45EWSky3MDWORQshZkr/4YtcEBRfVevG5Du
BC7koRfxHfbXdD/XIpguh1vjOLe1xWtFRFD5UBsc3NMwX/LeLQc6wr/FOubsX5BvjkkpnAChDQf7
F7hlCtXJdik48aK6wb37VkTJ6IMsIPVvByWK9uoG4/u9x1YUR1btP1Fq4OWhZCJDIxS+FL+mQOAS
yWyCdQnp2DMhiSEavMiDF7C2YahC4JKRkkUGkvmLZNkNzaeVAi+EEA56DvVPqqXwV9k/gMQnq0D1
RTa6KzkTalKxIkQztp5VPIMGlnsa63ENUNP+6tgZ6C1cc/P46E2gtjr6zevRA71R8GLYB/DyxM1/
6jmpS5whsXKVozWOL04cQfc/jsEiJfrV7lUbZMsfwNFD1Ld96ty/hmueGmsvFj8qV80NkXTc8RyV
sFGKGY3sbaZJkurUavxY9oBttp1rGgzXfC60H88WZNzQbaIuzHU90Rn8Kw+BZLBmatTN2wkcuV9m
RzXrVVFm8z8QPGmOSpGtlkLfhZUNdOIQ0BCTNyXYjQ9T0buisP5inGZGclRZH60zQ8+PXo+5UyOv
LdD7FudfBBrVSlO80wOBxNIHV3f/Enmz/ECzMrJfyDsLrfX7berY32eJDuawWJbbqwgorl9CwxkL
mX366nXs3AtXertd3szMQ8Y6gJFtyPcXAckdBFRG+3HLv0nAe4SIrfp0S8lcq8BjaFh5bRrjweo5
NOTfVqPeEBgI7QQz/SNOVIOVYjrZvJepKe/I8YC4rsy6Wqu3uj68nlwNyZPTAbGLDRaPLjT+Adby
TtL3QReikVwOkxACOb7eXkuzKcV7fMB/xiWzdo/Y/s6gbWk/gm8QghN5mMME9w0GmQ0ILP2E9eHv
jAzm9phHTF7tP7BwQ3RNwL7FO8D/jN4L0W98IJH/31a6jD1Z7x4X/MRsSVPakQuB+Cgt6tO+7irJ
Vk+XWcGwNVjkFDLnrtJGcm8LWeTMgQv2gT4OTfwNsFSQZfevgKG+3eKkd31Tloyug3fbMFnTQTy2
QEM2rQ31BixmmBcmUyC0PgeKbettPCQQXpPt0Z32RSCXEMEy7iRuCEbj2HtTfIQGbgXW321Wz5EJ
t2spRzidZNMrNq5DekrPU/lF/xZGEolnkxi785GXJkUpa49P9ykKOiHjwdGGJRF9rVVgHJmbAaAv
0GUW3+3+LZRYbb/SHM9KFiBfMo5AuqmGPOxojGIeWnD9WSLRXdjdGr2Q6AEFeKlaofn2IFMT+4aw
QsY1cNvwN1+yNpDquEzVEcjS67VeQa1nLH5/Vy/kyicfQ61tdKGfw8LIfUqR8rUcbAZxH4zudfAc
QiT7Fg9KPXcR55gbzIf9ZPNaTLDpWmYpz0cq0cW5IuSsU9+nGvflwkAvQKzJs9oL9wzmvBIXkBuX
6SRmZhklDzB5rVnc9yKSEQNh81HSSZpwRjZdUc4ein66o2R4V/0Puwt4M7N5jH6is6Ahpfk7Ie9j
8CtUX3aNGtNYlTHe6IBEX+zxo0hKi3GQqin+xcSKmofaIRaQziB+norbwO/1EPn223UzOdhdPf9N
0K39rQfgnwpiACpo/yDfIHH1CVfwariY/BeFgPQcF0QDMUtC3VomNycDrh7JU8acfYotUjiITVRu
DoC9IGP4odI74zr3eCLx+zAc6ZWdpe3UZw6R5enV/6h8yCGDfzSAMMDPUrH9J5pij6sCrMKDnL0A
RbcFeKBGzXtF6jc5Wgz82o0TIXvBz6hQq32auJNNvhfSXnpaSOWG+XgY5FFcJdE2ajYtqE+XMZiA
jIkwkXRpExONi2GxbPha+LMEaEn5CtCrlWOqeWiT4+VjQE2akmHWIwhkqZMZR81/TomLi5mRJUv+
aoaqF19wcggBJrsrfhx7HdZKgSxQgDXlzQhtTpk9sOB/ysniyjDw89ZUlRa7ah/OJq1jYL0Q8UFh
LS1kZfmhVpm4CpukjAW7uwMaDN/he8OX6vbo/JZ9tDZAu+UFU+56Gujm6h7WsHI22mm6V1aAuaNV
9LdikMp6T2BJXBQieclSFf3bw6+hGSFXI73Pq93/MZbxFmdpql4v9i5zcAtJu6EEqc3f0VS0BjEb
2ka97M0yLBjNvkPCtHYSqjppPcjb69rA3tUaiyiF4HuSOigWqewtvlDxlAvzUsGitzcPq2noSgas
DLK3RJD+kDKS+J6TwOHnpkkzJ/sULso36SMxijAgvzQv5soVWkeughvc70MpR6m7ScD4R4w0drCj
U8kcZc2qlkZWyec6yhJRG6MxMZXTZZdhxq0ltZbFsSwCto/9WcOAP41eKc92aQSt6ykrMpwXzwXE
RfEehyvPh1fzwgClI04s79fQYJxjbvipUrIlkal6sOunmzLsiMNyPA1oZ1QkAhIVetOyMqD5rA4Q
KB4Fp1jo+6elRzPjfSUXqHzozM8Kqps9BEe1rOK2cM8uoiGFC6U+H4OxlCjglgvzpmXT0ND0AiEm
6xsGlDi4APiH+6aRI3OZbugb8VzDeYEkxXBKGh0AquuybAKJyN5PyMVtYiT71O9+oNdDxZkSYap9
sbBpscA3V8GtxqQSSSGeyz5bQ8MHwu/ROLR5QQ+IwNVsLNfHDYXAFRkU2SgvPu9GknE4Bmp01yw6
wTo7UJ9+mRu3Gwp7V4w0dOaDWGApM5pa7hP7HI7kVp+JPXElbX5ct2jYrPFcK62YYkrRUX6cEp+H
qeNljrNJBjtS9GOVOhyWrMkSAhZvZOxrPOcAZMCOw7HlHig4vRAp9/aNnpLW4anTlavdxgNM3a/m
4KaqnnRXGOom0gSjpxh0xJFAr9DoNcMfvbJ+182UqEJkmbhEhrT6myyFV0TQXzJ+5j346GLGwXz7
tGb2eDzQ4X+PI5HDZlel1S/4jVz7nep40rfMO2HITl2oBXJ9qbJ4tPIEp5EZKajZzbd377mDOvG8
bes3zPo1NlQhBY0H9N6VrIN1T5jHn9odKFbcJ8ZLa9iT0BJj2KHZdkKr5H0mJuB8uwdNWRqqzcjD
exyAbyQjCB1rpogFKvnoaxzJMN9VVa2X1AHCp7nR2fv+djWcR8++/8JZHKB0VW/S0jI3Y3c2x6lx
5QEyIbyPKsj0V1yguImrZsQpqA5pOnhBpOBYcbZ3P39Eo++XeV34tjJ0NZRFAQ5i4ibLJ1dPOyim
Z1tIjkQaQelLZunjGyCli4UrQjDHniM0f1LWhEOFHxUh/yyfnWTInrFqeZEZ6E66PGG38Ygf6iVM
aGyBV/62mZcSQZytdcXYiV1UkZknpDpg6VvnqeFAKN/XBQYuzjckMf6WMpZ9Au1FdNsezGzz3qcb
0R99CLva3DSDlOwdwY81TG/IiTmLALnXmw8lEj+W8oc+daBagT3pUUj7xFcnzvyStElyljePwVDj
wRHfZrJen+K2Wgkqeym3yTM4UUkR7U/gjdcY+izKR4mx5tdATDYcF1UgI6tOllFzBxWRWyOG2g03
nbJNk5quLq/7iSrj5CIJRiAnQMWQV/CAX1ALnoQSEiKaWYjrqA+gorhz3UvqQ5Yr6erJ4LnXWxhq
FvS0etcP8lN0WQtdqU4zi/mtjSUlxTR3a3zzhSe4wKnXhL9rpypBlVDso46DaHPNgDaoShwKOD8q
kQNYNLOCsepejG3KLL/+64wO4rPRmdMPUiTxY1sztUfvofeNOUdtfih0ue93y3Rc3ksUK9FSKGPV
i/+xuCIRQUfcmg/FCYkU2TjN8q34AOMYUAu6uvq3ht5Kqc05AeAda99qu1ObcK103vWUt5tf6yLK
1kBDoeGsIRcE8h99UuybQV307klP9J819+60xAEZ8GV70doGvKs++FwCmaAXWvM8OUrmIPmo40O2
oLM8rRqSfJuSizAnZgwJyCLpyf0Lr1hxdRkGpGtam7QbesvjONRnW/KpqHPFDzo0C95I53o4xDPs
WtvTMoGmlk7YRoYqX+zy3vf7EFBn7kO1n19b/HC+jF9CKhxVoqudYBNKDUH4Yfx2cDneuHxHK/Bo
DXZQF7++Gb4/mEPx+xukwplfntn38+7D1GujfC9NYL0GVSaespo3z6gnash9I/9fHd7vFM3m0M3Z
hSavyhCmClkSFeh8usOGyBSgK1iT/SbK9v98z2Rxzd6Cz8v/0E45V9OyUR7BfUXRKV+3glZPfuO2
683hHimZppgOLyAooQ5btSj+Nodz4S/y0965KhbwazkRknSYHVaW+2Z68EO/AZWO+qjvzrsAxXgH
OtTBSQyTGrLEi/U37JwkyYAbTiRe+b4i4nGFYDBxQZbgvS4LFypYnifFvoRdxJLRX5ucywGDCV4t
YZko7i5yuQLpvp5Vw088Fmx7acFNqoFYYnnjbbkEmzdpgTYvK29JLtpLVJlD06DvikioBY6j7qOT
EFsHPqeolo+Kn833qZdI975ssTdg2XDmrQdNorXPa8Rs4xTYqAFrPFFYRe6xiYakP8X1PryvmxO5
Y7eQIq2bt94H/C0tiYzvTXUnMlb3sUCuvFsYJ8Fh6Nai4Tpy5Kj9MuCB3XkxqkPSYxaCqfBD3Mpt
leWQ49kcSezuAj8RZd3KczmLZiHff2KeY25HEd4HQfCcDuvF65N9nurCIkHhETMWw3V7HLF3w9jB
1op/ECZRbQNAHRVtB30GXRI0R1zTMNRAxaXA8FD5ZA7vwJ3BmgxbercCQRC25vKj5e32OmHfev2+
zL6tYrpeB+KBHRf2GTkSl4Se2PkbO3Xvim2+R5Pwi7DXUkTufNum8sbQINCTBFmngF2qo8FxlF9+
FBUw3kIXJZLK69QOoRiZo1gXbRL46pBu163s8qab77dyv/TPE3gvgJadka2hvvvDYniRj5zf+hQ3
/c/hSKelEt3cNyekjk1+TgVF88RCVYQ55ctJkw146usx+bdUyHlE3EsixAsq0wfa3103W77XirrM
talDkonNa6a34toU/0g/X3kVevmH1KXsrQ/wV8etii0bkdEpP3hS9nSNwvAxu5J/buyMiQCVyIA3
9ee40wYyjlGcOhEmRvMl+omHkan8A8qXx4DFfx0Pbihbbj5ktB4Ybe3j7KPln/efBEjKbD33rPOd
9dnaCu8PN784CbsqbYOfKFRJ5XsKh7N4M5eHO5ZkVqAGI3oKmsa5fwsPxc2d4tvP+fN1tDoEB3Eq
YspFGN4NSXw64eluX5BWF2/sWgrn33Sl+Kf//y1N/RSCtgF6Pxa4NiDUGxx43Iiry6YoB6atteuz
6wkHQLX3BdHlS6XP9/DmSxp5BDu+kNdAwc9O1LmnN0FPx9zYOW05XtGcQ4PmtWfYJTx0+AMJF6vE
2PVHPzh42sod1f6fti8VhohBLLFswpxJvwqchUrSP4O8jvKY101kMZAWim4jKOpV6fPWbGT17MPm
xyVREie5Th2kK7h1+78vp3ALywQ8gv4BozjmB4ze5bkwivEt6PyfV30qrceTGCBD5ERQFqOHqwWd
nesbVHUvqQRJq45FyV+//wE/vRaT6+aqlvougSevKS5O6yPLvDLUdgFFj6lvgjntdZO+CEolmTsb
uo7xqWpzeIV5/wU47cd5UeqadsjrbjXVrnSyCMx23qtUSXnFqqFjS43QcVm5/1srg/Wc0ibnqhWc
iDo1ZsJHpm1dznskImHrM1G1aRFLNosUYWW8YqK7t2tIHyvK9TEAuBn9ezZh5lTcu758UPLlfX/5
WXQ9MSSpiNo3tlrEhTMTYrkiYpl1iQ/bE3g9bsJNL/Yd023x/zjMqYFYPatt2V7fuVEUKDAdi8xZ
vRdnUGTBcs9FED2uOz0nqjO8MzRcbuAs9WpwLJOQHcM30J90i0hC8EcD0B94J5KwAP5QsVV4ajS3
u2y7yyJVbQbUVwsW1XHOU9gpNX7ATh9awAsVP76uqDmBnnQyIEpxEZPbvp6XR+mWBYzIPhra2p/q
fCJE6z9QMpqjSmG5AlEI3l/78MYsDi9BrBCnMlncKQyxZrBEdtEA0urmF1GeaNPmrWVu+SZzekqS
eoraAw1aaf2EeycNbNkxKlKV/bhEwl8Znh0TAkNNGTDTwozU0xpyeiE2KTixovfw/C+KeqkwRAzI
cDjgPAQi/CPvljwWg5KZtpx6y9U6h+jPUaDs1tPdPBaBf7rUWdysxUkM0rWvAQH+S0Rih2S2SFme
NpUBXHGj4+Rc76Z//e7nhUzdrlB9as+DVvPUI+0Vd4GEpmrVFRJ1KwBj1t66hBkmuR5DClTsrPGK
4SNXOuhXKRr5Ut3X49eKUv8vjXT+/XbzHn4nxOW68EziC4pxtGCCaOP/4ofNhrjw/GxReHL5b2wo
XlS5i34ZDkf/KSrMmVmEjCYqxr9FDQSz2XL7ALlNBV3fE05GIXhBY3begpDOH/4MxTgh2obfD5aX
Vzjr48tT4haT8/i+7aRwL0falp9X8ov+p7Nrms7U1nMWMOGYmYROjSklAaUm9RIHEMH5hl4GruzV
1XgP1cOD8OsEJnU5y6Yafyj7vCsbnZfoAxWhVYX5wZUIkK5HqVh/E7MlYDMln8cuvdyibABus9SF
EbwAfdzH02ELBUIdQu/tIRdNOaVzsPTmYsATX+eTzgOGxkZ3Y7w3O+Je0sDlj6reGhp59ltHK/uA
4En2lpT2JrJIb9hfDC8dp/WCsCodGXQlD+Kes/QzVabFA4o76xxbAosAmEo/tS+37cIRPiy8wVEI
krXDFtoSE/Hvv3IdXzVud0h1TLIoHE8WY5RCIVAHXxxYZLHygc49/bbJ7eB4mh9OxYDWFzYz7C+7
+3hYlaaSAeTVHYc4CGmKScrcCPwpltRi0S3Px39vHxDn4qZTMlJrCYoF3wokPzxEzT7PM2QeVBwZ
t3mtG9TVCC2PZxrAyDSvCsMBAqF4I/ldTQ0vzrGGsJah1MtgLvuFuUGGxGZiosaM5+4x4/Nv3eTU
xWW+gzr6BOL+gGexafduguEvMWMV9Mag6nVnhnC/7WpxWPcqOUtiuMTom223kfbkDCoKfb2NPBwz
TTxKoeVCrpdG0fplaAwPdYfSGUnBUaEfw+z+p0Hat3/YHnmd5tN5vYIuuZG5P184BZVjxz3P3PGY
U58f3ZQ0qpFvmKiqultTgAuETb1FvMdNi4o9wX0dyycoZUHY+pqSMJN6LC80+/4FeP+yI51XnwBP
CE4EBRLKnaM7EhiDmEx4mXkvDiSqkVCOdFxdqHEB04Ir9z8WaTYK6KxJrzjGBnRMsX6EhavEtzuI
aozuGroDUZZ68RTClcYaym4g8mvE5cSpcDmLMDMLdjm9K3ymxzShAKzUkKJ1rHaT2nMFZUePW8OU
H/tqw6aI1exQPz92q5xlwG+dnEZ+9ih9AqSzJ93cHXngSU9Y0YM08IYnOid0O/vr/35LTj4p2RfC
3SC2vgmquMmwGXOvUA6UAIHONEpQIXddOQ0QExUbXTXL16kuZbdWbYSGFUOR9TcAbF6Q5TRNbyVf
U/jrkxSQWMuX2sGmmLyL0YeTd7v7S1FJs1U9y88E0De8eV7bcqTK9WBOqv+p+mdLiaRzwmo2WrE0
XcbNnXyay/pGKfzKnpBtAxSvll7iolbEzmjSku2/dHRXGzyDpJ1p11UdTc0+ZM7w26L1AJ3x9INF
3FT6qs6cgpcqE0ExHw7eeAEwho4zZ0C3unoFYLAnDbTzP9Si3GSY1u4tdBapUrRF4wfuhAE+ECOS
kcS7F+gYfV3Suz3lyrAdZXtVBLN0wt9MjrioMwDa2aizgAC3oVnjAqPnSa8UkqEjse6441hj6U+V
36MSp5672wREmMzDE2h8nwvAgYMEkodQxCggm6mpSX5u7jBLOp2QUvLi3nSBjS32l6SiIukZP30Q
wMSFya2qgsJUrCtl5Otba1+RNvfU2AuS7gxEAyvul+jLHdpF1bqQRJA9aD/lTthBWJ/qCnL2yn1P
OD5pt/qefeQZ8HvAgdRutX8sQEAJm5B9gVYL8jwljOeqWHfkkp54mU7ZaTpHPuVu8f6Blgcc2wKW
8nAFDEWVyBFP4QRC1JwtQemsZjRiIpWQO2D7D3V3w2NN+48Jl3qv5M6YAoXZI9Wn/7pHwfQwNpWV
r9vsf4E2sFAK3LLY1eZDlIipokz3+KSl9qWaoH7jeWZjIsfaXYh7bUwGW051C8cclft2r6yYK2cv
o0oQT+Sx/UYCgKxxkJ9pU1D4PdldxaEAwWkIcv2odhIwthJY3qjqlhzzfKug+SS/N1u991yqjYrZ
tt7pC2aSsCgE2n2y5x9YlKTRTRkQ7npxNYgdzHNQqNwdldwLugOlfU5/uBYcJYujCUZ/aY0faJkq
rfmw7tUPyQbg8HuNiQVpGuqplDfHhyUa4e+nboCQYWqEHg02eSmdwshAal+ep4Hftb/s0ZnrdHyK
1WnaDMSYcBrQ7H4b2ua1AfN5Wrym+lOD9at0EPihqqIJxlGrPR5T+jTvAU4l/XGI4PJct9YbhfHe
Bz5Tfe3LXaTGU4hfKHWwZ55FOQmfmUJjkrPb/ZuBnc0TMJhqM9+n1ho+D11Wjzvq2WMOYm9qlIJO
GUBrNCl+qywbOJvaeFbWjouWLToZ+2x0RIBPIfjFGa+skvPXAGEOWS2BCfDZi8sFphj22ppgK2F7
7LL+lH5HsfiVR/jdHSdArPyqeMXChgrwVRn6RvQ/JabdajqFpR2+B+iCzKmsCgRdIZYHHNuo3OhJ
CcFtBOdf4m7qsYWusChb0TbjxNKaFjwrzZsBZGRT6MYQ7yr0SUfmAf/AYWFkmJKvpkwQWhnSH24a
nF6ruezxAeG4FD0YeEq95tqeQqJdmPEvG8nKkIii0fmqFG37mpw77JFaEAePtk3wYW2AF1vL4WYt
pqUYG+7Q6nn5OYtZYP5X0ywRXKboDKAP9g2iTyxpBJCxCPIGGCj+0FPyvHPG8AQsCLfF3XkOyxtq
YgfSCo8XOpVsW2DKO2NGZuTljKnR1OmTXHwTG1RK5R+4fWvUISEdIkCa7uzrOGkFjVp+AIHjbf2D
wkWSKf7imbaDtPzni5ISaQIgCgmEo8JinNSU9zt5DhEzCpfEJ4kV56Ai9VRBuAd4a+WwhF7hXzT8
sDhM6udx9XbWjvE0Ci31BYkfzleBIf/mdABglwdibfH/2/ifQyUde1iyQbObfw+b6TM5fGm0OOzQ
bzpUijq2nOl0YAljdcTn9ZNV1yXwaH1DpvWv/n9dVbi51ME+E/qosaABvVL1E9GBk443859bRiHb
+zx73PyDueYW79Z33l1/4JY85tmIO+VtUJhxK6dH/sgWLNbDfWOakmqx6K46j8zyQJwa8ngFQ4J1
MrfPWSt83wJq5xlHfqqkXdLuhkdtTnNDt8u4g5vRF4LjLygtt4nFVo7x+Y5Xg7z0H62BPTfQ+lKv
7N3Xh9DB4WhYwe0/B7g6+Qq//Ia5opdB+YUg99QGTn+0+5b6XQ4MEY2LEDLAJ92XmIMSCnuAHZRq
Ec48iR5nnEAnhjvJXTwdN9de+BKWS5uYr9yyGx9w/iJ8GtJpwz5D+ibQRLtPEFHMJIFKyp5qJSaa
C9LUUCHgDeKEqNG5iY5XcV9AsIkRCDsdrxvubAcA+Ign92VLk3HIheG2U7imQnTQDV6Q0WUFjcw0
8dfod6zjf21gk1W06W+CRFtYU3WcBQHx0rr4ucqLu7kddfAOJdW2PWCyheSnQYgzlYS3aW3L1R0z
vi/3qtj8bCUlTdsLbbmU5+TWS+ZtFUpbNLvbn8SL4Ct0LeRKrClqvvULO34P4daGW0qpeULUsixB
he0I0q6TC5Uwto+Xylgb0WS3B0O6vR2SsiRdpwDvXmWla7C2H78rdFQ6gwflUeDDwkOVkUITYatG
Os3EoppBfly4r5qr4AQn8UhKmA7PDI60A+KK3Arwx8GUdrCZhC2QiaDCyipI0BdirPn7AvBKsqO0
PdsHkMJD1J+3OGGfpRL09xHEbs/V+yhuhqrxvrVn/22sK0vrNxYdplm33GnA03TmdZIf06vQdErf
jI2MRpzvlJI2dyDQhfqVdRs+IZq0nRH0WRHRtMo7lcW9PI9TyIknCViH1rTVQfc+IeD8khNhePGN
kqmC59iGiRuxVaCF0EZPSffnDoW2cuZ5FKWD7GBpe/K0azqE9Z8XWNmiSe3e1zGCMBHRTBQJawsJ
BVB2x6zPXLM69voFDByOM0h8g2YJkx1dRic186h/fdbGdorBjQqp3+MUvwB+6RJYYgHEO0MuINGG
dWmsdHwjRZFpnNJJKV2SAVE7b1HVwDv/lphSOg8qT6mKisWA9FYwXNzjCvbzwTNp8KZCZtcWNbtM
TxT2b+Z6Ucc81rm4PRoBtP26DzpKoKCsj2qzh4tjCksYFiHfGzOF8jjfADM+52BobACsQ4F4LsHn
UTNBFdeoJ5vnB9UVui1IgBU8duye0WLsg9nhBeHSCOZpJrR2DG+tIC7h5ej9zyf0Fc9RA8jKKxvH
J0dJh5yE+vHtM4DQzRx0CQllipBJVwoZe7gru+EgJo0APW4L5M0rib+n66PAhPvrxIf1wSMmMewt
bPWVRvGR1/K7+HU92nUwRpMK2V5J7LILk89HfER77ghx1pf5SPLeEzHzl+rv9ONNkrkzrKpKHHEZ
mcNAQ9fbaGU/5TV+HGwDE3jbHVzjaR0pdOsYWt87XjpyyshRsC3kSR6NA7bLTsDTiX8+d1qhPZBD
I7u3PgOLltuXIHvHs0CZGdUxz3CsXWJ/bU9nSj31/MnCQtMLmZI00GQR2JE7NvucFWuzuMvlBOWw
Qc60LN3AnGM0v+Udk9SmcPecb4TXAUZgfyohT8kJi8Mbi4GxpXdFrHeQ7WVkL0Ql/AdU2jVnyEqq
JdoHhy4tGkoL6UypsgsYnMs8xPeEcAc+xvK0FXZDOkD4BCjfT9n6hkYIdhOaju2jIWO82c7Mt7LE
L36p8mDRLaOoeFHetrrjbcoUgHM1fNfi5k6xDphNKyd67WUvn5K1Eex/Trr5wC3B9ZL7wpCVFgjK
E7LiOvPFWe4bNQZPbI3PgY7sVzHg/bv/9WJBfqhtH+wjNq1d7DqYD0vAE7xIhznPS/dXQiDCJyNk
xB7bPe8MlKqK/hvZJeJXzc5AVnxQl4X2EbPUlkdGkQ2/XmHlLs8+x37/SexzEuJZYiYvtvLmxooy
Nnip1z1uFbBXwGcS+hYq8jNSfOc4gbLDXu93Gw9t420Bxb59yQ/+xt8KlbUQUN5vsr05iK5NgZLG
7wh8ToVJXYQCdbILDlLw1DoOxzurvQmpxUsyob8ghrWaM/mg7ogiGPvSfiQBTnofAkKNB4sBhLKx
DTpB29Qnp5JNY3n8SGnxBUkOyMIiQXK7zHugTdbslcNpKjq4nyLFWuj0YROmZkDVf3mJhpSsJXmY
4vOZRV0q1DxEHstuehboeBcUKCYedH86kcY1ViOoN5wNddqcv5Nu8EB3cEs1YuwqvjucxySiUtGb
wLWja3cH6k7BK8O1KmJ0y+OzyBSWIz8v2CnLAOMvIcxNVNMuvypmj16JnQice7yUEUv9O+QW+coE
+CPZ5yJQvzDwhWEehWR3gXs1sTeXAAzu5EY+VcLVghA1OQBinjhedoGJs4nYqxVmIjp6at0Svpsy
+SZhlgGWmmDRXe6QJtrv76S537C9jHaGTU9tIjiAjfJM9QB7h4qIfWPyGpsMsKuLkntpTKB9ybaQ
SdWdpQT2s4ZSp9wq7qUkvxh5N035p8J4Y6yTrO179JsNhfWIryod/5guW8tQHJgGkUFN6CmxfEpO
jGzVep30LGVBgrmQ42kUcKFFo7udrgYxf8y+nC5LdQPuJiWkuYwD0ndS2+Na4WepWu+5EKLxUDqs
Mj8enaYcoRBdiO6JO8Od5pQ8to+qeqtki1JJnYj2hgbHYDJHSp4TJX0go/wIwI881y3FpW0aBwId
4Y+mlus2C2BYu/H+f1hQf5PdUVARWdOJl+o3g1VF0LhebnIjZJ3I0LCGhIH+Juvlqan79QBPxFge
WawCbOVI8O4P/wZ7+0xHpva156oDA8vUPPS1cUs4iOlI7TgaC+h4G8wIeN0CQkkIPVvQIm6HjaiK
3xsF2AzZ/o/5o+D4BJzNgLss97v0sbInSuPrRafypqGLdegB3lNg5oHj04AnHA+1eDzLTmeOhNlH
uFbBZ0j2ITqaUmpZnhUlzEAzPpQ7YYNJSxa7J5HZDIG4zu4wZB3nKelJ9GUb61k9IqN8BXj7FLFK
AI2cQkpxUxmS6SoGom4lN6QNWQGbd0rPIAVfQUgYyQ8COKwonKZVHj7fBbND1XZADFHsYUGoFgFJ
OGy2ACnLXuRliOQ+Xvfp3zQi1ObF46bK5RZJm49gbtzf5cfQppjFlY0np/ZMrQE1DBgOcdGkoR9V
t1NzgPQXj2QXjilYgPkFyDk5qu5c+aU+hOuiZyBiEnJY0o2CQNamjj695almqdhFWPzOLxgcqnI0
D6hbjX+aj2adC+pmM5owQT3BdwPSbIewBq7uFmry6oQ4T3+/9OfSi267aRyKD2hMN4jN5QZKsIoH
Gq2afUBqkT6kN0sfnXjcVHIOapbSuaBlMU7C6URZT7i2e/mrAwxnXv7qy7LpHhhb6wZ/kF/jD1qj
PJdFnGwzLq7fldRvqbDtnQ2A1nVgJszsl4orLPnrGPdEzZzqaYWdPJt/7Hs4vdADgs3Zk6l2YDbX
QMEw9hK/OH5eMADo1+WjyFikK4SkGCj1V6zXC2k4Hc0IEh/O5m2/jn0zAjhdwtH7m4g93xZkbsgt
d7JotCsnStqnR3obH84mPGZHk4AD5CVMRtqYj/vTFaebT3QMu7EOPE4QMFxUaXRxelr9Z+fIsFDq
A5NlODe9oB9u6cOO15keutn7c/Dyaauo3Yt180D2I7KOPg/DR2qetZxwBoE6cAJViNuKtZvSs2LM
mjqOjX3eozbkZ+zHSGNFsHNdTmtxj2SnOLYmVVbiL3Mybmag/67Jdx7+x/f/JC8DEM0DqibkuyPV
nlo4yEMD7yZ5XA4eFpCUvg/MeB2fszGqkPmK8QGHMp/5q4Fl5u/C2h3iDD5lugV6cdwS7zt55Due
Q5/x+iW/Wsxt27wLeFVT7dtdcaOc3OzAiuzIShHSJGvnGUass2DwMCnPCdOD1R6npPG1abnEbU/w
5zIcnJyHG5yZsXlEw6krDl3iTjzAJca0E22M5O5zYASOBnliYh+bEbWvNJ3DYpmj78SavcJge7Tn
rugw9JssJZGfyd8AHQcDwcNCgWrsqaGPcUEntlN7tBIttVdiikUlTRFWoxvbhQqqBz2aTKj/evZo
ZjuYmwqNCYruY0tRBBxbagEqi9AnByoTZhNM75DpDhkB+hUZeAvaX1DKyYF7QiRRT5qkJIcwT98d
/o8zOo22JrChTx6wOx+CZH8Fd7MrfmqgK/Ugn8d41el0RNnQmXn22m6YyNjb8ZnKNzrElEzRjOzW
VwrIEvcF1eXBWRc9dG7x8hD02Yd4OMOYnO1mbP1hFemUnWVcPO9unH8dJyA96eNwddAEuKWnHl9/
l6CNwyH8IAs5UFO2jwOgaD3OJdthxmpXx9FKJ6Jf1a904nkr0aX/KPiCzodjRZt2+tHfiVkhGFrT
ICpY462Hth7DvNllNBoMI63BnBjPbm6nZkPCay7emOFaJfKzGYRElcksqzEvVlvjlsGmfDGir3Wb
KPGPDWfhlbfpl1EX47/m6pTS/mmxF1sRP9NxYerx+qR7aaPBi5ISLqi0YWSRXVhQbd7vy0jwk9wh
e2MYbI5lTUvlF3QPzO/COjJ4ODR/Ur4132IJv2e5azZrmzkTXV3Nnpzy4L/VDh65Ky4lZPmGAsV2
NdqeXjH3U7vYbrLPP3aAJxrvRfX0H4XlBMXq192xTm8hrOA9/VP7rCvla9AKqECKtoCHILK4g6tY
vyUtN1sktsnNLSPFQz824ijGwkkXhIDsu6KQEj1uR+lxyOygHrLpfNuTxIBPi9sNDqXCLNsmRoym
H3rPh88oLdpPOAd0NorRdP+aL4PnXXaB0YSYNcClVN1NKsEoTGzxs++9fRMpqs3Zqis5vKM+rIdh
ocBM/jj6aXIFwvUkVCUzMvAYxYGuGDf8aVq6MCHXvF1YHspJGlggkwS8bD9b0dLUysJVIizjb9pR
l8PTFOthADsX4TlSs5MQ1eE/fgSIMBGLf77fa+bTAcGTk8/duZHWvaIBFUWXJzkaV6WnaSm8jZ3U
SolX7VZ5Ozj1r7DEKxV9F8kjikuZBs86rCPc+e3OGoV+96rrFdXruY2ZBQf55ULEmT9iyQH/KYQP
Njz6p0GSDkJje2WbGRLftnGwe8p6x84AebA4ovSj025tMx2DaKXVAPkyTTFVpZx/v6C5kR4iEDee
XUtPoflsT+U6/nLD3XjQY8PzqLIu1iIue5B05uxKiWN6V9fdp9BiIpFIQ/kcueg1A8b7pNOZElz/
P02bgiUkR+qdmg/A4060G+kPpdXG7eo90J/KXQ/sdEYbiFEq9ebRH8nfgQCF5kPTxNsMaVvTpOFN
9ereIZxBllDKBc4h0J+PDhFSdxB31EQQTjfeoBF5cTp5onzk0NJD3gO04exTQU/jMpXqGRxQpc9H
2J4pAXvctXs22lCMJBd8pga1LyLO5G8CFCddT00K5M4JzPWPcYgarxBQklQdfrpwJnTsfVsulJ3R
G/d/84iSOOGtMsmd9lsOGe3sduwuU+NOrQgGsezl3nWsEo7WENXT6CJsz8d6Ndi/xbk9YJ4isem7
rJ04GyC14Ya72EtucsCskheova3/uiZoGg65dXm9ndC2GPmhD58yUofaPCNWaOt5PTJtCaVdCYwO
xPnwNbO6z6WiduDplEKQbxDO4oxEuRU/J2Zabf6F8ux5EJYr0y1hXtYowc3eres2g63v2u6Yyhlj
fDsslnvDAEKZGM2J8QDmWlBdYPo+0n9qZvmrTZ72jhRAZ4yyE9dNdgd169cRcgheptwujIj+VMlr
GIBcB+mElo41pbslp3X4+hkMAUTgz+aP7OyWbH4P4IwKsndEt8eEjBt20K6xX6MPBdWC1jtTK2kr
mtQBi99/xd/nD6D4ARUcqHQdEdhamo4ceYFwZ1NIjnfrrpUNv4ttuTCfAoR+YugitoZo33ITzqk8
OEnzD/ac/r6gBn6ohTj2oDXrKg8bNz3we0SdqEamYSQceDjUaYRCS37TYDqXn1XsnSo3Ld8SYPnq
rg3zh77VsmKLVo261zMehoVsHLLMt7Mv7ypCTKncnjT6dqEbA0/xkLWqW3e7sRBbIpb187Qo7eqn
hvYBQVx5FAFbETC7qhkZSwkg+qRY4IysyFdPGEqoEngzU3mcvVxoAzDnkN7g3Jiq7tSxqy7TUkZK
P2UnITz6NF3TqxJgaqf27a0Ri9syj5mmUCuru2Kt6N7lEFurJk/8CV8ovDl1hAbfZVOih7ZhhmII
BBHm5pS1K7IVNEqanm4rzlL1HWxj8YutmbdP0xpTu6tCRqDg1SySeOhQ6iDOcfuIpRARMT/faq93
kgA4BsoDHRK1PYhQ7HsX2fRAlXgmCixBAUKME3FQFsDet4NdxS4QYqKFZx9YP+7C/pnO0N6HpUPS
Dk3L2LR9EJdHUwR7cbkRFw9jAhtjNZCpTVyqHWYervGYHwSPv6f/DxDoFLjz2OpawjBKt24Hnv4U
VVhIxjtF4lai5rGanElIs/aZhbuCnVQO95ku4s2pTU2RfdcnlcHUx8w1aSsWVHp/FpS1DtXsd2Wc
XM3QnL2Oy+aY7SY0DjnDgjpgMPJpmOJ+ml7AmJUur0SyADBwMmuIlL/GZ7/Zk4enFayGQ5n3Ql7t
MuSRAvaKzEmjjSeziiclxgqjCk6e6YIwXHwy0oJVQJsloXNtrUB2OAueTzdaju9fKJxC65D/p1ke
DhoH5FySA4iyl2kdmoxbM5JQyfYAYy6eDvYV2KLDGqGIHrMFgfPvk3Zu5Ys/i1H5YBUBul+7KpRo
jXA2R0T3Sw1AINO4aaEfoSOQwRlpSUOf5usebxpR9sf/uq8HHJLukbMnT7bEt1KQ3B/h5ZKnbmdO
wtG7AO+pWNU34WdQJ/o/HYltSgtPv7mx9u0/+gzSM6JR/A0McBwzxN26ry71pwI25FoXrohIdh5l
VMuA6qTzZxikjzMqAxdlZbQ9mpoCkQIIB9RsxZrgBRz1a65WhnRi3yIRAppePaoubFboF0zjmD6+
69g9DcrBcffkATC3foAbORNY9nz+rG/5SWJcbWlxgED2lEXzJ/n4aC5toSWYx2SDYhAfpNcHYPTT
wm88dbkESNBSGADOCY+cqvkH1lTuL2pMFCWsx1nW1CA+vhd2KeQ/LJLcNjJ3F4IGfMc2UEvv4Xa/
xGxv9lSMCHp6GPPaKWAOPmSnyWe/lk7kvvApOlwbRnt12mx2BM397AXZ9bFsE5/QvbdWhWojom+i
ImJbGlX0YyGlIquVztTZSIlyUA+icnz9JnN1TLwdO0cfRI/izlL32uC778wOPaL5leV6qxlVa7M/
Mu/hzpw/wKkqVZ1oLiQ6NFVqEn/Fw/cGBOZzxEJ5ToWmKtOUK3GAA3924eNjEg6qcQPsdsuKS2SU
xkHY3Xvo2aRs1IXRFe4ni+9JQnKmpcXAZktJboHVKljOUJ7Juiiw9DbdkZKvTTfoW8FPvRvPrJRx
tq3hN+Fml003u08c/csa8wQY2oIoUYRAHDTh71Nt/oFXU0SNVj9mR7xHT20UDY/pUnu4ZU+cYw/Y
NaM64VEGwTKeIUgb79H/dWkfhUDx6WeeMGibjRLryhZ8tuWNxq9s9ysvaYrRV0fxaTi7RC5Aqbar
9bO4Ow3PDhkWYyYdHkwEzLUzRNtllNYMpvwa9P2kJMogs8QPsD5yUaq9jgW4FiK2GoW5ATRFiNpS
RqbPVBHKsFdfOBWqG7FsjuzXpqhnfOwVhCGK0+qyq6cRYhVk3Mq6mVkvBga2q/kl0KvFgN5pKfUY
fO3x/odtz2xIsiP7vh3Aud9koFNcdcndxZQB8/GuP7yylS9LoNtkwoa075f2Co4gd0NGbPHLq6A4
av9noehgVEt0tKka1kNQ2hsdyc5z0l6Buu7VkW9yjp7zNRUuYdULKettIAGb6GSkI9EbBZQ0mf6v
vy9n04Yu2bTL/X5TsB3CEMZtuAxyMiEokubrjW5+aNddcslxXLWOqqCnZtL+isBqyAZU0U5o+E7x
4+aLAO7GWLv2hiZ1rr93ji7E0doLztOq8Ffwx4PWy1v4MS6MJABaJqFYq3vN0N1n6Og/rFvC39FY
URe6h7+jw5GYYsePg2vwO4htgS3Znmvp8CCM8IknNxzPgWSHTFH3KqFA88akGh/pEorSBYjpCdlK
+CrcmBDLaFl8yjjyHr5yOC17xV5r/oMwyjsBcx443k8KtunCv56wNefZLu6xw82tPUv4E0dni+SA
H6eOsm4tmTGztZdiJkQDY+iv3ugwzwy7OTwccu4nFvUGE5aDErwdx6oAsgfT2ZS5khuRDvE04N0/
+D+h3RuO9i3vkO7eSLdNckPtPLMJ9K4kQiaciAycFRkm2NLmUWGMCJCBaekS76iGMr5fntoqh+lb
gJrD/904fjK0vWAp6mQcnExfbnZ1SnZXyN38Zv54Gf5UAxRBYESQmOnUn+RrM93jL42/rpv3GgmD
nejJac/fwz6BCt14b27ZvejiDBGFq1yvKOxdMtkGmmrJjf/RFHMT9je7r31b6PMdL94dLwjKNWbj
zhVKNkdt9JYRsahUaHHkL8fn7KmUD7D6I5ItttDHqMxPXI3vklFn85aYwqY6OlvZp9o3Wf7K2uWA
FrG4rNDViY3j3GgCvDho54kjm+ThQ4xiMKiHaJhEf9O8Blc9nsqSI6W3nFpugAvVT80D/diLPaUj
Fut6HyC4fdZcL+2+xT36c03fe6kIZiHgpRtKDxMUuPfpHtspL2r2ZBT9U4GL9K58ooTbb9xSNn+s
HMybk/h4a7G+Ph73+ztCsS3o77RP0VjXyy+wF4q72xqLFptuQNctMho18Ihe57x9KBIP52QjGaYK
oYAqtSWkBLa6WZohETaYpaOh0kZQlsFjsfPIQZSEhWWpj8LkrJBEXGvP6Y7F8VBUdWMmIZ9fSrmA
rOwYaTfvnNxRCy5mmQU/mIQNotr1MI7foAuXaB5unifKZB+wvi7dwnhn5FoWiZkETqJYBOGo5MJn
QVu5TvZ6cunTyD4B69+yftzYQxmx7+oqMrVS+fLa7BY/nPMyo1kJ+GjLRMx1HpKsr/ZA6Cact14d
CuEYIeB+/32B1y7h2Rla9Aku9StQLE4V13X9GNB9EtfyKgrZiYCecGXtpZUqbzZZaV/ApN+Y/f0m
BFPP/eie3QGjdpHKmB4DSN2RQ/8R3Lo2ih7ek5G8RkXrzHfC+XT6h8frevOVZxfWpRbCc5XWivDW
j4te2F7yTv4VSPtqmpMf9NEJ/DBaM73RAMJR6GBVKniUynW/QRpyIqA57aChHvRQA5/cBpTenScI
0O1yYWOVyRkhSEWHJYN1JVbZ8p3fTMTgIykIn6j+j7t8CJctnUeB8nq0mS/iOG/EAV0rMTTTkm9h
56IoPUrF6rrbS/w+7ENMgF3Y8ccypD0nFTBHdTI4exZr2N0sa6Oi1E78vqLkn0LgwcJO5fIh3pp7
cblnqwjIATNQfpA+3lvZHKe28H9XZQNQwLQipKB9cgSrsPQn1x9gtGDln/GjweXZDHV1cA/rsLbV
ep98ux4JbfIj7OXktBC10fv/Vtb04uhYHZk6XB8zpnFfIXBIGNvTwRSY/AkrapTONZkayqIxZXmb
kBFP32oeHfVC04mtsjQhWqKN/8anm6FjrG20HQ0vdzD5MWrysc36SXrCKzpYZy+XXwzOnoVM7Nq1
uwVDeQkmDbjDpclkUfigSgQ+6U5q1Ez0vmwcmOTE80FkQXBp9xFuyfVBLlrzn0k2hU6vDTBeHQbp
hgVJxUpA+VztcY4IqKglBlrEpluGGfbmK3ecnqsUfqXE8y68Ioz0NQ/cRU7sYYl6vjR9d+sTtWG2
XeDUq8kRrBJpHy2KtqhRF6MdN2RX0JrvAm74tckTHBBkWjv/hNHnyZs5f2uBJoQHEU6PFsCE+tc6
ScUkL11P1dUzxNu0fQ85q068Ec8MwuzjaWNey/EgfLV/VFNwsZ6FLxzZsOmX6bKZybDACYpM1mhB
qnT8KokSDyr/XYM2hcZxNkwv0KzMB54s31CbMz81QX5EkGxvrLYcEY6DZ9DDahM2aIKoyrZEkCgQ
o5+lWnjGXkTHF4fK09lwxkBxKTVBvwgWrRw2KJR9FpfIph9vh57UTVz2rswM4DmSIqmQlue18N5B
tQWjTQCsb08mGOeNCyRxALxPO7YAwgVpsWzSZT69q/C2ppUxibgSnrFFgL2i4qKsAadREmMr780s
86KM8L1wzBxWfufknpm9bxKPbI374cS6A6AFGR3L14bkTnLJbe+69lWhHETBYeKEWNt6mNX/bcxJ
ConBX3HRy7ScJX+d0+dVwLcKJX0EVZFaok6l71u7n8ypqqL9QFYpxjb3wtA84d4XkPWErG19OFsD
toLoSsMBFZ5Owl2OznX7/QGo5De1A27KrxSb0hiXextrjEJzviY8odAYafLVtIz0GwUVhrbSQyvQ
JV2df0NuASVy81+2GUiNLxBnSB8o2nANCFFJzzhlFQli8uWtfkWbXfX0TRjz3lkd0wJAUM3vaZVH
sOOEy+/jEe6VfAX5DRF4No/rDH1Yf3tXZNZ6P6EOJ3VAjFQgpMKWv9ZcWzIkh0/3fSGZHJWOs1h9
yQPOg4FHTXzkC7rLMw2L88WULZA7L9zQyR59OcPuAQbyRsk7YLu1uPxVW73GtDJlJB3jRtH1yVCo
+DgoT4IDu2ZA1xLqgIWiWVIGBjwzPe+1BcikLpNnDw4v+ILi6UaXGYhCjjuqUXQAkgVkW5QRZeeq
Q3MfX9cncprrxSjupUwp1XXCC/Nf+cygxLhvFwYB28AgZ2lnBms71nFwaiOOnke0lwJvM+M7XHOQ
FG1kLKYz8FMBshgOvuYx+ZO9rXTF696jyObZ80jbCazHWO0HC40tZaEgFOxY/pKXjoyC1UDMrCZA
XZfCRO1rL8/iBfdd3REzVAyZX5dmcyBvlFDGhd1CZ/5X5CuoamBDkUU3dc8qL01kaRpDA+QnDIcA
RX0wHgYW3TOtlYijnRGR1i4FsqAJtYAtTPwqosQURPrZ/Od9cF1T0vgtGEf8o35cn5CbocSnE5fl
2kZy+g9qRz8EpNmQRZ1uCafvCz0tWVZET2RWq6I8ObDbQwqzYzwayRLdgk2PyQ9+AExPlNuN/cLS
ORvfmIrGuwhdpYZtO/SZs1DV7XmBsKyFR98f8GPkMM1w9SvDj4d7FsUiIIpMYOt/m50wg3POZGgJ
5THyi8gMaP/bLby9FBzRPrqY/xM+rN/sBQOqR2kPpbe+nXQGPCOCkWY4j8A7TZb/txvINc1U/1Kn
5AsaTYWLzbFAEBr83Y61sL54z/PuyUjlr5W33UG5Q5rpFE0fkLQRea6OKBUyiy9dO8yuF4boisN2
nICW8HZvTn+fAjIg6ZTh3WcWOsCsovLPdA0XaHG8vSGhzWTsMjugK7FTH7ATUXk/QJ/4nJr6HxAf
Hss0fBPLaWfqAdnPFNitw7bWYi3BMqk4PaZlfnndUxwqqqNq2r6QsCrAtE6b84DbMWajTtiYJts+
nXWiJR6vx4oy2gt0R2GvVqNni41Xez9UGmog0dMDVXsEqRa8sm28BgUJMKYh7V9iv6lrvHvOba9q
fbPI4BSxgsujrczVY/QRenLEnK1h3nXzowdx3IMfiEGMbnIU7Tdy3QQAx/uJnZok4UORiduNrUoV
OYgnuNkfUKX3GMoV+Q3aQ+MU664/bxNuFf8YYT2JQIRtbq9PnjPZ0OGVkWns1wsmlHluHuHt/UOD
6hOXrQr6Qg5M+VWJdmOzqRtzGHJlAHW9/uo94jVLi2Xkg9c2nhyf4yaRW08Beb8hiFRuBlK1dezW
iSIukMu9l3vs+ZqpI6XZpRYzWOfruC6943FeuhEY14BSS/Jw6MVxIdbq+fg870DUVyPY6HkDXsb3
Bj+0djruT0tk6jyoJQ/4+gO1ug9iOGbBXLLDlnVmT0lWcc+9w1wOgqlkfev+pgb4tjCf16EvBKR8
CKr+37QmCkJkg0FgSMlMSb46Jo2khub5NV3vYrWlFfiZO62qecF0peHma2QfJe+/XGbI/rEi+/PN
vPeE6cpR4VW8WQZHHIGUbcEHCtwiF/9zB9kE9o+mbzorLid+FQUbIYuDjxYWzHqQlkmONEEnMXLy
uXqh7Ctm/xk3wR9nAPTxMtrBKb2ULSdnj2hlgNv8oxCKgGoU4zV+s/Q/j5nmsGW7isYrPM/ZXekg
b/mNqbVBzbgRAywhrYauUYAJk13TdKy6U8hg3yY6MXxnJRpoS+GEouXq8i6kTklExdEDxCczuyX1
/CVu/NDhUbkV8aQ4dLS1XpCzrTnAxgL4bwxALfVKGqcbWDxlwavPN2PjRTywr8QDlJBj3J5niBxV
3eVF4OgTCHsDs5Y19bGXKrmLX1tCFTTJnOiSuOqiUiUv/xSlkhZYHGuTRe3cGJMzEEkIGf1MXQ3U
CC82uF/LMlZ9JLY0PfY+hHiqbSZRyExTOg6i4cCzUw1jCnoYjU4ZDANXcOm8N7Pq1KkeHt3fea18
TpPADgffH2N5Fdu+OhMg2rPUTIiiTiXdOjECTicC4PIdGP9AdCKQm+5syMCcMKtUhn8GHsD+GwhF
uyQPhacaNj6sMo3YFxM2jTF2lFIp6tylOjLRFP9W+yReGm4med5yK08pk1fMKdstFjR+ndzcM7KP
5jkVetVQx7LubrKxaeoOKIqR0m19096TwWkBKAlgTQ3Dw4EHUaPaQy4BRZIXbOMy9M0F7u+g6+Vz
rqYcSrUMA0PayS1sq9R4UhJKzQ4ZAl3aIbU7jzxjn0/JkzgcexbUeQjshF8vSk25+k+VS3AQ1iGd
1WIogQCbVaY8XXghRuRWPpSr3fzsWNPhDI6qjVgZtFbrIKl0NPZEiIm4FVzBtxHJLvQ45g9KVaC1
HwKldiKDpkjUBnWhpXYb/G5yDol/ZwupCvPCXo6NojH/Q9BVXs/GD5o2wgc4MbkNtfr0gbcBIES1
4tWhEGT4GZJ2JwX8sMM6v/bDVG7wBAUh9S4wu+ILkIaX7fzSKEIsI5iuoCc+ejbvNVISOArnLC0C
2YrJ/A9QRcupjTyhfsuKR9/WCc4OQQy6Nwv9lB2xOTAVFVyJAdxT6Xudv1jPHnZzAg7xz7YKrCdf
/o8joCw8enw3PJEjPcFIJL0H7t8uRv72E/PtRSZrsF6OvwP9AoLxBVdNUV/FTnhj4kic3GhDfQNN
/7KibehoyyTqKCxn1ZfQb3L1zM4rOv7VlfRag1kfn74+to04XJX5BzZ8JUBcIZpmYIpQ24HiZI/+
LmBa7w4J6CUEpJsgbm1M48h3QAO0Mrv40pdpPLpzhUGTe6yiGpa3/UEsmbsvl7/tCskulbpoeI89
i6RgGSuj8cNyKhThqmwS9JcnZK2eE/U7jKWDs+WVXKQAu/vL9678xK9BlpeLwXyhTh8j1j/II3v5
9iDjz62yAns0a6mWQHsRX4oXekgnNavOXckCegPZKkdpuEtZoe2+z/LcenDQNqlmBvEsyViGFftz
enWatWHiJ4zMpJdHF7VG3iI+oif4xtSQ5EwIoRG/PRBKpODaofs9Yip39ZtlzjiXdHK85Pny/ydV
h4SY9uf/xIsbOWXOV6d4G8zR7Fe+JUQfauW8ZeNpB4El60rpaDz47gWXu6sreG4hiqVg2PuFDKmT
3HBeYtGjrngx6CSkRNa36mjqATM+36aTLsHPQ32Q0/mwAEZngP06oEyWL5f79eXmokHoNCll0lJ+
jZ0kbMUHCnL1LCGaPgsZP2AG3OJoHFXRvGS5T5ySdsuurAw8ma0ddmpGw/sm7UAmK0nyzpVERZXL
VpMQefQUoNp5VjwE7hQdV63c8+szBu9EYYeYwVGPBQ2allDZxPZv+24p2j9LnsOgSIc2ZbzEUObB
IZcXCiCbHgMrHGriN/0u1MjQoSgdOw2VESZCpIyCOlhgM3E6BOU/Erd4I8swEdTksP6CncnzRTl0
SfZ/bxOD9jQaJDTrX0wisJQOPU8FmeH4Q7WhmVVjGm+indWm5EI8Xa+8Mbzu7ikHeseWhoS5wkwS
FTH0RyoTscJfJIcqMIHub5hok9cPIwosq7rQ/iZ2Ws/9m+LEUse5ruWDvnBt/zbSk1dTAZdgUS2m
fUXAqmsq8ZOF/iHAsas2jnXfaGBvC9oamlnw/mW8CPSG9VyYkIKwdeE68W4fDXjia3gxVMfx+gcG
Zmz8abdzNlCQDD8F4P67qG9r6YDm4rzGjpBlMkG3JmUtPVEUbly68Skb1PlNH7qX/DJ/D/WAuBVc
wTEnSEI+EslXk5djU0B2txXPlWW4clTpuwEnmsMDY35uS2XBnO4518HnTPGkAru1fBGMUpD4+Hka
hPKLsfhzltaes+OJHBs25KzqBJH0oJgOP+ID0l+QvAmGUbUQLkKjTXsSf/kH3fxjkxwA9GUMR/GZ
Cbz6H8iJadF8Iw5Kjco7zJS+p+LhPNJTd5aVAVBIYjk339TSbUwEnI/9n5P8NINIJkvdRhFz0WlQ
inKbTjnWIRZG7YCbekJ2PtuXob8TWG3LFfGgx+MRX3/Jp9xIRA+IDBbz4ZVYwF1HT2ASft20c4lu
CsrsYEFSpIZkkn3miJ93p9S5XdmlT9YNr43iIU1b9fEZFw419/RQL6g6M8HkarO7U5KuGfESHotA
0qsQxGfry0bnP+uUVZdJhMySeEi3LQeRomu8urW+QmFKdY4x4tzdgebOwhIVdM9KdR1STwtcvxwO
YIu9D3lYjctaBrpgZU8MDfzUnl3xjBHlmUwno2XICwTrKVR21FM9c9g521BXWjV4Jn9fq+WO4MYX
3WijuPIk8G0cemaoGk6sTFfh79lkn5Os4a+IWFz+aOyiOZupDYCtkdAwjgie1XYhqSG0MtedBi+n
0LwZsp0Frgtgf4S5ylx/CosrwHnpB52OtrWc+xY3MjYGKmk+53iPqMnyLE4EU3Pw8RERDqiUO6IP
1dukZuC430JiueFg0f84jhd/xTgA9GcmvEVoSFvMK/6WBJyzmpe3yh/Z6v6i6O8y3yjlqdiZPIcq
LG2AkEfatIpTUarP3hJDgKxwiP/kLuJnFGhf4YbnZ1aEZDe/47sqw7wfpwLqY32HeH1G38gg/w7k
NytFT28IPwxoHSyBoq9O4NJmybGlq6U/ezbMleh8JMrDrQwA6luDMRl3kSY4UcZea6PYbmkMPw2i
UNmsRCXvuNg35H8hYaKbaVRpSR8fWsNHNO0wBKKyqLhxOz53gu5bAYcPnXuMytAu/eaSdxNlA/tF
eFlf4re7a8auddHpeN8I218r4whwTmT/gBNp2/ITg9p5Xd+RM2VGxLR/JXzsT20d9uq1x31XF5+N
g9fKNmh5mgZYUnSgK4UO/e2IdkLo/KFqxnu63cADkO3ylUiaSseFb5sNe7RmAuOsW+o7HQUrxBoh
MlompKg8hYZwwAv5nYFB7SH2NfI04ol/AMFGt14ho04aNJMRyW3mIyn72gB1JOwgnV8EPdnGJoCv
AMW35lcW5/tgAfXYaSw2onztJi2LzdhhkBeHpcJ4dk6Ej2OFq7HeeNKhdM0WPWkjRsck0x6e6Zgf
8deXgPU3cbEXRk8c65kuhPgeqiblf9izO1WqbVp0b4X1ZKx0D87KGpC5qoDKH7dLFkvX6ZzUxgpo
hS9QEtUYTSU3IeFDDm1s9eqLQelhLooQovNCVGopgdn1swfm+mw1LfbaVvdR07VcMzk/3H/f3OSa
c3eJyNwffGR/IQMRTAFcIWflMywle2SiIXO9P7KRTBjDAYUqIQPWisQyMnWE3Nx/zQzIGs7etA1R
DakpicO9Wv7LpEBNKdyrsSPVGukOpm02/D9ML6Co3HH5O3oTITPPQOIUvK/MB4YjSFzn0+3LRWVm
0IYoSJBCkPIuIjKkHFsj2qkfzv6MJNBcPdxt+lh+SmWfKrnt5M6mi1k1KCjSsuKiByzZ81ATYIdO
uLumh6roMXSd8oypZ7pbomxers/KBC1fqB1S7Lqef3uRDkKT//ZbYgJKedewlvj3zrSxPOxPPUfZ
YjdZySdFkb3dWgiZA8wOgAhHPKWyCJJ03aMrE74Zk+MVbTUTxHIBfXHqJR8A9FTH8UKJaZWt8ZVQ
8BKLwq7LxisSjfcqYwpvg01V7ivyk0iHlI7aX7GOzTOZJ62SFzpH5cwkMVi5igqj0JeS3avLKY4H
AvPdFvt5JUefGMw9/tOFA9ITyNeJaiBuMLg1hmivk/uDNvnlrLcF9OoMcSwHMcYAc4LMzvz+++im
cZz00dPM+f5vb8xw/omyo8DSAff62129AyVc8eOe6U8U+o1FU97dWBXZg427DgQPnvrvQAdKDFOH
93nlhAdhb+XQQXblTVEFbgKEVmwYv8LlmVVUu0kGZbNCAjBw8b03RZgektF9ARZrWPaWsztY85Yy
RFO9wSdE1EmQVnSwU5gmp4ia+sjYgIQeA0m/AisLIVwn2uJjmV6lVFdaFZ1CnC95PFLrs2UNUOj4
1ll89W1JU3mFLfZVxY3YPtKOnhvEQPyxr4Jc4NM7/E1hbmZGPOSbYjbkZaIz0FJyYqBT68ziy61g
wyk/Wfyd9IkHPpQQsYaAcxhx/ccKAyLzjm/leg+HRwMey6F+1SKLdR59GCxK7kZXxM00lWKla4+p
xLe6xCgWNdBuErnYANirU25lnrUqdxXATRRE0X9wCLSlGk6EUYOQz1hphGO70KoU74hY0pf/RDbP
mBS1BjAEOwsIR82tuPb+Z+3Sx49piTAtsIPAt2vuMkX/Ku2PacIYdKbTWuTHGRHhivheTclDtDs+
n4yZuJu9BBsgOIfO02GElTqg3hmqVU1TsuaHevOPkC548GE8LrsOOwDTFPYwf6BJHxXjaQELxq34
pLdQhtiqN1gs+RQGijR/w4tD4UEoXYg6iIxIxc6Ax78tTPMsaQJp5tfJCaSGz/89RRrJqYgdW61G
Ly4JcC0ZtWEf+YSjhfb0Ku8s1jJ5qcGJhRFWTGkVkF4QgTno9ReNg+ec5UIoNPp7vfH78gA0lcOz
Ii8ubxqi2d84fSJYtIfNG1TTZVW0IUzoA2v90RpJajHncO/RUtrmjnlKR5lBvYz7nVrsvKfh+3mV
1zx9G3YSKGvwHBW3Iiejgws62qHyOt7RGBJxTaycF9oUTmR0A1jNWkeXotTzueLqqswIjjTl3GS6
1IaZY0FpNCDpEeKrzw7Mdk0rE9x/ve5StUxb4ktuniXqvqJhtZC2F3IfGwtLv8/mG8hvKtcpYSNv
gzuEq+sBY4Vdx3RZWOWDMbj7qPHNQ6NtUC1HM4rukma+nbeHtpXycCTUHHylcWyoBV4GjaDltdum
d3kEANnMuzxzAKTgy7PvgUlSD8gT8+GM3N5Iz+JCa7bF1IRfge7U2M5zeBQAYLAKWufEDVcqrFFY
UwQ1f6njqOqVfctgdsQYficfRAt5E97SoAN/dFV4eNBHCmYkKjf49L8NWaBdc5AHI0Tv/XUgsz7u
GZuv4AJSAjvmZIr4j7QivvikIUPQqjHTLKQL89J4Hod6afg6KDXsC/0jGjYaqThElfC2kZHYVygU
kSr3jE/70Fz2TWwYlDhBEm4KHuwiIvMUeFW2bjD3uM5tds4vASrO2seAP3Ny6H0TVtL6NNCWWD9+
f23KDKWCkoPFfXlOfEfteTvrU7+41sFVYCOyDKDuhrKXDzdxHZbyHjGs6CUep6+HwcU6ofkW23ID
pCf1IB5Bnjg4Atfra1s4K4r/8ZqL6vpXa4WwsIc1ZDhSO5+Jp2OGncd6r3X4GTrzppBwqa+zBpX2
8nTb+ZvzMqkpbe3DAXxqeSUa3A6pUR4yIg1kwUpN26JxtRGKMNUSK4jentqqjmTBeVIPyrsHkM5q
guO3QOQbo+tkTjeSLWH1Mfp4p1pljMJ/eJe/omCezvrt0WZvN4m980tcLJ3pGvGdk8BhC7I93xa2
WM8Pqob7Kdo7Q9pNO95NOWLy9xLFZdmO/mwuEHewYX8C1MDqDf/35LQikn8IdkNOVWzMJ0B03mfn
C0feXUsRq4lpdXTVcN43tyLZKBSeSE/6fjxgDU7QY9dnOgcmaaQSTxiDLYGMGzR/5+EdAnYbN5pq
ZXB5qCa6pioLIa7JrjAo4oiFihsWU1MFXD11AKdQG0oFz9q5EjXaRhapv1axx37s2zSlnWefZzOR
wV39fORiYVl4ko4ry2bwfodjXZ1Et9d9a6Aywvcqbvt4ja8bkYJQhmD280O5S1C0hxxbPFpLdtZ5
CXYjSQrP3DQHtMjba70VgHxts+98zpm7di+b1Wy/LJ94KS3MhN74ctMyFlYTCShOMJ6mk9Lexido
+z0Q98CFbXIdqVBBUBdYC8Z48Fc0Y+3pCs3Eiz3yOVXWttGNSVLsm3fEx9ADTI218274wTHE1UxD
LxM4BCzUuIllgfBh95ygiUH/6HBkt6uLGEJgsdO/m98F9atChG7mX0vbLKlVldGUDpJJdtARGAyd
K3vSWxNKx/Jfl8IY2sdlxWg8VuWuBW2f9UoKQUdEqvprDwBK4dVXyIzRU2PlGpxyHx+4FkPTaBhx
u1sN+gRpr4xAgogpp4XShTmEY8ZNBSIhaq18R2hR2pBjs2TksDNnXmFIGeJVxxA/mH9b4jURkgIu
6jQEJ0gUB/ipCbDXbJjsXqncyP4lL3P+zvHAA9jO5j16+hQ56zK6IwXwqXUOqJpXiiE6gXN0X/mx
o2A3NIPXqGy9/8/KdtGrbJJ7ix+8RVFHk3A541E+fA3mdu1HzO/77ajOt5arxwfcjhp8yruarl2g
DQoz1kMiRlrymCSsEAGGN3wYQuc51R5iZQLqSUKXuCwMc8Zo1osJj9K3lf9mVuNNI5n4rCx/0q8G
1tx0d8Mur24C9hsODkY8IR1XBj4EcfqY+a8WgI/uGCs4Nbagzhz57SHZI7nqTE/bvR5VSXcDLo/k
e4jJjACSEes3VkL6gkKEJJD7ckAHYQpVHmSA8TL3kfsF7xdi/UHWkBERy0tYEl0TVuZJ1UG6zfMI
2CJenaXzLp4B881EigHSzLEpbfXAReNnoJeZJZsZ6Qz/ZBxUohC0j9rf5U8TrQwHykulce9OsWeG
MXR4VBl1iqnjuY4ONOa3O6hif/agN0Zoia3DLPvh0nPZlkwZNiR2okXCSPxFRXjDna8B3OAMTXry
QUkXDkNyYVEeonARVPsYHYGiZthsLNvoo+MghcxrtSIrJ45mNDAdB7LmE6oKZLXgHWiQvvwSWyTS
truCsWNyasqE1fi87cJXyafuKApj77NPmEZUAQ8T4HFsFynR8v7dPLFTIKj5BtLUZnYbUIgS8l1H
yaNSknnygqBLdgdxGZYUkuHTBo1m3L567nPDr7zYpLZSHb9oRuN89IojUNnK7oJcZF8wFLlWmhDR
5UjSNTZ5Kx2kusuDIdHE1K/U7PlEx3SHeI5GUXCC87uUNoAtBmWBTHp7I//VKsayHfk3XCaVEYZu
JhyOVX0OWehQU9NCBSpS6JUX+Go45F+8w1lzFW15sLI2o4aMH7XEcHIVEErLIn/+Xur6s1oNOy39
oFD+6s7TKec9+nSsxrXgZRZKdkUi0BILx64ansM332iwT5A9nEDM78Pm0Zd4jScM56/DeDkfIq5o
WEw6KjNkwWc1cdJ7R7VuQ7A93An5CF8C3fzx0NSe2lPDYNPYdHsqgAs8MyK87kXsnsqIhGacDNaJ
Ik3ipaYa9g9RmDqs/5StLQyaqxhm5er5kDNLBBjH2uxianbUaSNfuhlNK+VzmHi3mWKkXGncvMEF
g6iFIgDTTGpxKGx3y16gZO5c/06NKMfC7VyGiQDb2mNhDvZLgJ6wjj0ohwXYHuOt++P8dZVABZKT
08al7i9zcyRXv7iYsOzj36zxMaUgPgj3hI7FTGJzcW7n7jxj824eQc8oJW1mhyJCsXHg6zu6lmMD
l3swIZu6/8rCNis4ucS1iAmlHqwKU0kQ+wd6pRdmN/qj7K80nbceLzyDmNNEAOQAd9uItQuAzY+m
sRXm5sA7isCjNITQTCBSOOYv3Uclg7e5mMXDZpEjwy42LIKNkfSWTLF7RyERVnx3wjjvdlqXg5f9
2yfHjM8hy8T2McHNf2ErwrBjd6kBpi1bE6xN/nq3jZjHsMRZEwRYWxMeCZG5CUZzEcULPXYktiLZ
5hK4x4/LP98iWM6//wM0BJP+rlpGa+GA7489A61JvT2+3Bh2gP8JSlGvdrDL86kBbEVnftgQ5gAD
47u/c+E4rbELDAc1Hf6LstXxdC+RNkgzOWANMF0GScHHUM6WqThXp6xT8fYBWjXY2sh5PavHZnBu
FpNW++ftH5PAp1wdR1YI19praDqwAXAT0DmjuMYtw1h69Q8N/QbsRh3otjHyFRQdYmsej2y6zkbq
SRumcEk+XV5Qj2oqUghqwuXnyKdrnsRFRlDHl6mcIe8mr96E8zU1ZYcXoIMetSztLt8h94WEhAa0
ts5zbT0KcsZGd8veHntPfUxxj9ixF5JRo/2rmQTwIOpJ1ap3OIfUQ+VOAIHkR0Pq4TsSq0+CJsGs
xNjCA+InKWRYClNmga+HbqmwAvbJcI7cIt9l7YNvzJ/TNZ/R7U2g2CJCaozvixT4DckqtmWzBpqF
dUh9XQktneZ3dHtlkL2xDxUhG0IlGFu7SyLBm6g6+WbX+l2jJf6bVQOtjHqyoGLA09ya3BIHAV3C
TMhFl1sbOxm9tHAtNVzp5OBHtp+MjKAthJIgJ3afXn6vvy232BRV2mBUXSP9okS6FVtGUZHYK7N3
kyUlN3xzEs3AVNHjKv9E6oMdn1VFPdmFLcXofTOSx9rKVtZhjKDAR5t2ROS7W7XPCTIz2o2+FTZB
ZhGPO1gN7m5iMvfxR79QEMEYFwFMBjHSiQj2kHb992OGglTjv+uFF0ukOBCT9NP6+1P1G0avhSIn
Y+A73hzk1WTXL6dQfDS/UFjXDulCfPvFkxbuoWyYBlZxXohd3idvHsTwUFrjjln3XVEZKPnewjE4
0eNaqD/9UUzztOwlCzUso2ylBprbRM3gu8p7sBEqEBeRmTXR7mgW6AkVroFvsT3qY252HmAYaA5M
4TU3dgQbTLqyrL8ByHedrXXdDzCE6woxvtAr9SGP10KUM1qGlzUQJ1QpyxTli5SY17r2d7Ls3mWB
N/I7EK+7beflg0Yx5IRaClJQzqEFrVjS02T5edFSgSJemi8dMnIIRxJg+mCa6W8x4NeRbksXZB/i
CEn/SIcY5416HT4hXMon4kHeKu597j5v6Hpu8P4CtfBo+Eq5xOdpmNQsqZvMbr4nMY/U2pymkHex
gEyLp7Lv5cMYeje3mzYfSt9S/kWl+YiM23ULKERZdYnIAsbN93+/N4Y4yfJkYTNKomMv4pBQ9czf
jAAbHEMvaRHyhV+SWyax60l7Y6ePlLBwtTNPBO/jpL99iT33RdxMHaLfR3vfEq3FnL9tgOatNIuv
EBgYXqxGuyVlFGKLuTEBhEnv9PQGuO6IZbBC/KioxojYFJOwmnw2qKrSBLXqXniDrnvAV9BgB12u
KtXbCYssZ6EoljBPazNxQg5lCp5lS4Q9FfUM1ZHQcjYwh255O05Ht4aUjnPaJjtOUUIwsibpbCMk
e9HM0wMwk9vo5gHeh+fmKesfx92ulxMc296jtFWneFtkl6IMrNzaNFa5u8EVDHNHJWxg5xqBqDe2
TdG1i6hffDuI4aYYxHCSBWTHAXBNV+9hwxZSSlIEhf77G5/vvJXqw8oTllxAffi1iditXXIkhn03
KKaWbKA9dfBziqjEfsLyLqRS/MfHHXqqJZ2DcmZz9m48nOVE/o8D3KIEidl4EhR7ChlbRzCxq32/
2wIx1fz4hU6kMR6S1GiLpU947TnhQuP0GU9dDMSQz3ZFGq4l1pbwvMUiXFb73QvRCmf61pVq75bi
ElfDrpoUlPiilij/+UQAPmK7zJ50AlM+DjmsyrnSsR2y7NkQUyPrq3oeu58icCgArI4Wg8tcQDV/
28awfb23T9i4eHxP/EAAKkU6aPythQiazIWrYMqNcbTXAK1zLQlbCNCnLyT7u78PNcXjrEvIAduk
cXMtG1MknbKvUgU2ZhtWElx5DQnPia6VZc13AOTXTUBkacCxljmpzhvxdLpRc+vK6ZDDrmb3g6JS
L/U28Nz175V8xjN6xGKi6w7vmWiY8W7lF+bAGDGKJfRJvMd32jE4Ir4BzIffHUtOb1f2YkXWtPai
VjddduGAvC+a6w+7GabdXzGeE2LoprrrAxNb5d1teLaPt5wWbySzcNpXGlAdVXPRQ+/x9aod7trl
LY14CYNx2IRqZGFcoqylJfQG1UB1/CE9vfyRZ9gpTRCzfk7Gx4d9KKRe7kpeJzZkNVZm5SmfFr8L
hopcyh8FuDbXySFrQIRMFzK+9Tf8nk9VucdJqUK+cswXsnCcTOf66szo2gbs8FiUYKYy8P/TnjI+
/XOGv6qk7/U2PslzjXrqlQDUWFEmgDF/pAFvhfvnMCB3IAQHqzbxUXLjDO7RrRE80vfoTVqXdDmF
Mtf3fzs9QD2cFJHJKzxRJAEkP6Oam0C4gG99YEtagbrhID6JVn89FLqzlABMkKnglc66pWDG66w1
4nqF1Vd1y05vIvSfltNprBksKmR3x4y0fhILw8wu/ChJ3HNnhbvSjG35jLsysoP8vXCqc+vAUCfX
8+ZnmEButrwgKKDNvI1TRvWDcmnnW5SGCFq3IfRtFLFy7dS8VMGTL+jaHB1ckWPqgNdqGSLgD21w
CNEts9nCGRDulxP4bnIWD2HmtOQ1f8Eobrh1tmDmJU1+1B23Qw3nsmyOtctKeE6OPk2sMgWtc30J
0tmKDcKKJ67PS0BnRpkDq2IjzXk+wHwQscY3zQLrkfg6VNVd2uUk4zY5NBqMnrNEybFrIq96OKF/
PN6LZwBcLgkrc12CWgdvU4qz6Et40w9NS8mZp0tFMfAjLgGV5Qtr+UBF0PSjbQgz+9/FJAEXvD8B
YpDwPRhwf7yPC0eQPDdJESaZpWf7FFQRshiRad+f1yRl/gNdEhHn4HETI//wb278/bX/Cj0cr/yE
M2Eys38E2TOXf9AtXsKdbWqBzeQ4uahl/q8xDO8KQ/FddqayWwOoPJhsD1h3GDMWT/znxYY6jMut
nK8niyFQGB4Jtzc5cAJK+hLiyLaXaNYseErJR0j3jQnpy11bK8I5yY52dDnbo+ZBFRECVJP3PD1e
kgBubxtWHnhTy7+/HNMsAnnt17wTW4s/GPa93Y5FJzFjG3Vy/MKdZgQhiinmvy7KA50QZbGjLXsg
i2VkDODiC6xRhOI0sNu4Af6l8fxwxj195LEHhZU1dJV14lvz254SsIRUpeXDYXDgSzyywIs9K9rt
fauW7eZW2MtmxfC0DOt6vZ5xlH0vR2XufmrFKEqx30mXdglTycL4v7ZjL2KviaZ4ge9fFSCFMx+p
X7nQbiXyiTLA3y/IHD6ssHUl9GwYR5+qgOEedYGrLdgzBnfQt0MnQ0Lhp/FEY/cIX0p0CjXZVYow
HsCObgtKSAg/KKYXuNuhD+D4ZQ28cjgnWEEFbZeMXqeOpKGq1nHjZMP92xbfDao3HMEuGvTSjnVA
EVvRwNuWePMy/gW2PbdGv3JojIe8eSnTJcfzMgZBVf+XuvQ5VtUpvmW0YbsLY26ZShMGI9Mcafp1
E2JyHD8BbUCdnfhbm4TeMlAA4Ui6wytsXXj1ONmWfyLhfYg2j77hel9nrR6T5vwzYD9SrYh5EGOg
N9rDZKR6HixhUVGDOr1a+8H+4Hso3ZQHiqGuuflP/yxm3Sv+tZ+1e/xLAks7TqVrTcpGeaT8IdUU
U+GjVyP0IOrrjXMEOv1LpOGNS7pTjKYH+JFJS5jBYmvl1Dctm+Ku9Ny0MYYbhrjUUhli/RWuVBwg
vxASLXhtRheBFQ0mqtQMe5S/IjmCIjM2m/W7dVcc1XGitWI1UD87CyDSnl0lU31hGMaCcyxnyxSM
OpTVpTAJzxxdvZZvpbz9OQ5OXCbarQvfYuWI3kRndyBUmAUo0dLshTbrZ6Kq3ddYOw0GosYV1lFl
bAQlxvEiGkRYhAUwrDjk9llJJgxuS2+PIEY326FBUTxfznqFxotRKok6jAs1uPVuuHsFAMvv9HMl
ODednQnAxi52xnL88wyVdva0VuvxY6kLF5pscTjcWA4MIOgo/sAOyFfCnWeCOi9ahjeVZQJqhtV0
4VcUMgACwUnB8n/+dD36BnOnnMFa4Q5Lx+e/TXhCWKwQ77m6aCujSFAEpZf3h5sAPqOGxoZa9UgN
mo+ZN8wRO9lm7VHoOcewvjehfwHmccy9TBY53yWDvRM5Wtb6mgmTceBy/ZRhue/ycPDKNpZZ5g8M
Dp2la7MDIHo1ncCNM/uTi2N1hst2k86m2vJzP21VoN+pz3C06GWozVFls+KkajHq86eCpXbSCtsN
/vIyh4n58XHjcEZwWOXCawNCIOOuKnk/shDf9abmKcS8TcHfexsIFP45gYzkz9yCTKO+4l/0eUL8
lfRJ7GTv1Hs6vXnznhq2CUPTdV+WoegICagpZpmjPDEUNsBXynLilThhT/R/vh4e44Gfkz4XwqXN
hgsI+WxfQFWOLk8SMu+aA7a4KXA10xeRwt/D8kyz73P6AwYQzoXOtZswrJWrXRkSzGTgb7NuOIS/
knLRLBiAbukzBBi4PlWA0Omvfl+cjel8QbTHOxCQXNPBK2fg01MR9L2mLXjlO9vNAg3CKAdjeh+b
r9cLibyaRqHohMFC2hX49rWYGdQ7XZ6CDQ7x+OOShNAdtBvKwaADKLLo+/hiBpvG5UXPaoZmq5J4
L33QViZbSNr5ievEYr/+PUAL/+mP0e9Z9XAp0QrsecAXvB4EB2tO6vnyM58GVRsg2gUjYFVccBaB
Syose8bb0Umm/j8yw57mK4FjK7rWbT3h4KQOIzb7Xa2JnCAQG9hIuhgFlBBD1KDV7T85fpvpT5oX
kmmIHNHMUBKG5Rp8Q+bC0zG2xzUvOBz6oeArnpJ1ZyJkD5szKyKmC8sXi79yGTMVev7xURFzZR9P
yxFP7Co+j83mAn+Dvg1ugVL/JPC/csX0/4aok3hrX+YQO5nSeF0byhwSXwMRb/lhc8mc6U4uNGyy
DwS1SMGZkXcVVy8oUKkvJMgxGRW2xdlsfZfTm9nrkR39z8oCg0qT5DVIKGLPT/o6V0k7IYlFeUHt
t49yek0AoraSCVPYOGl8YXdD949AHy8xZOyu3XSSslSdPuCgfoI5KNoqypfXNwXbGiJSHek4w8NL
3Rk86JwkkB0Ak+FxcxryIr5d8NXumOZ2Dqq/gOLPjOp7DCbuxwEQOCPNU3vYPkPLC6Ln6LqD7R7H
oKK3vd5Q7ZoEFapqPS9lq9orNrReWCFE2v7YzIskys5TTRpOULdSi8Tx7Wa0VZp8pczrXqs+7Q0Z
U+Bb8t6EYESpliOPxPRb54n7ONV+N2bTLq5RdTsdmMY6S7ZYKrN5lMfXahfu6zOQlHjNA3yKCGjF
i5ssurkWGRgVQQUxrWARUGi2DTzfr8DTiyFUkjYE/6U1SZIFRpu73Pmim4RUiTD5Pn+XuZFiYpP4
nTjP+o0o5tebCkXdcf3XcWbA8Ye4RQc7bJcXsTcFT7oRvhpO2F7xh9wtbpAdIrdposLhop7HR9bM
yuSCGaRDFyBUBC3pId5fwBn09xeRBR53V4eYu/b6/tDDz4Bot3j2yYjZmS94KIeirVqQWvmXXMYq
Ulq09skKoLleMTfKZTKmal9nV9vkN3w8AAJfnOe3hDSnOgdKH2k2Ye8GMtdYTfqVZ6LJzYDzYehp
j1oocsUaj81h/2VllERVZsbq4QmLfTe2+Kl9PShm1EbOeRN9ZHUWkm5qE+3S9REGOkAW5Eh7ddG+
RWaoK7X46pzPmFYSaTJd1UdDJTVq9BqlqxGSLOnuT3c1Zdfpr4SVyM4j15eRq+JwbeRhYBBDmH2N
vHqFQPJJIqPbhcPomG/hd9MlZF2IHROlbirQyf6g5b6V5Yd1ReJNQ8nsOWCO2Gi7bcpv70d+gW1p
zxezBgBF4kq26gbMvKZCUESYm3+WTRqigi4lJRPlCRhL4zab0qPGkwkbAZBHdyFc+kD6NRP1m/P6
QMQl2ci7pVFw7e7b2LcbjHAHi0yfk2wXyOh4gow6G34JLAe5g5P+3ZEiZKQ8s4DMfbjAtHORGEZX
y1ANVfbMMyecl2TLClca+VubfI/Ny4F+oop/sPvzGgjB2JJ4/SDlG7Dv6HsjnYlLqFr1tQVxRNS1
BAL6FOvQ8lf/l+Sh2rAxI6ZPT+xdXyR6sllFjvKH7L43ETbKvLc/lk8TFO9hO9t/QKHiGkY3cal7
ro3ZAniqlfvmD4MNmz/WTCET6TXMC7ZQjK1YCKUBpLpxB8zXO5nBxgR/N6caum6blQnYrTJPRBgA
VsfzJ86G4R5SZdUSiPTNT2mHmtAumL4DlJPd8Wok72oeKQoPcOuNtd/SL66V74otch49TKNMaZXL
FBRWURn+vZ2MEyZi4cVpIR3/s8z0GsDsiWE4bHk3fLaa69A2SZZmijJI53o6sfnneBflaj9Xyh4k
EsIRegE3qq17N/R6O0jV3QmzrvGbv6mhl/J9XucakVwWc3qwoijVXWRcrCBTC5Ycnpef7TCjdqvp
CDVBPY3MoRGxZBw+qi6v2KmFgH9GH1dXWdhZaEKhMXJiRia6gOfgfaDrV0cg/y0Ff1pMgWIEAVmS
evFWdISFinofI3Z9orkT3+zyJCVSuROvjXPpe4Umi8DdX1Y8/+TBaHzmMg162zEE06Bc1J3A6WAr
Y6hq/ym5GVMl2wuVKX033NJMIphwk0mR0YVMT+TvoCCKOi46WkzlWQr5u/hsIzA9HrKQFHj/Fs6T
Q73IKPW2zW+BuHWZRCqYPYrUpler3yx2PCTACXLFGisHcvuaCl7qE60Zc8WLLvfAbX6WSvt70hyG
4/ImaX41Es5SL/okiU7UOGGn3UBYRzRly7H0WxNOynE2smwyU19axYc6C6+hK/XxFteHFS4Te4PB
UocY0IlxdxOl/4cPSWb+o4Yh1iaj4ofFSHz+KCnM2+5VkCBV8AzwVH/XwZtJ9AduJg+RedKqqYwG
5WhFmdy+yf3JIJgoqBLPlyeG3U3RL/VbytgdNmG9rdWVDN0cYtsWrrD6TfccLT6MxYawTTl18KxT
IC+jBnUGyYGcaiP+rI6Zo/OZMe1L2+5L/lD58HzqgvIXJ8BvU5AN+fLroUAhM2bV/KV9IudBf9ec
YzWCF6Y7hZBwpROhQGZc5+uXMZpykyKa8QtjQuUO01rnPZZ7Ll1AtOJQLA4zVt3u9t4AaqduNLpR
sekh/bf+XPoRIOTbnpS19l7fHqJhq+L8E3OtpjBwcG+vpXtClRn3/HqB6moEuKlkueywj1U2y+o1
/rufgOgEoT/WuE2IRpOa9/Xtxf0otKWPqLTFQeA0Ofh3cik/uqoDv0/inrsXcRC/z23skTDYnxtA
IY5IMKqKgbNhOk1AuUWYyNMAZkKnte5b+JP9ha+zC3hL0wL6sJ4/GmCjQy9Imv0k9emUhpH03J3U
ZOps14RDRgacguQJk5C/bnu8eguMoDrpDVhmz79nfLMfAvxlY1ynVaJPnyjpLlL0b7VypLdZQft9
xyw/aicWsnQiVU8SUEkB35mdwqNTOVf5HiMhsfmHo67EtWuwGs1SmWrurLyUqMkgjS4+SA+GZPeJ
rR7NgEJmVtWjer6SywOdo7rxEcQt1tgi4yspTEM2Ha5H6Ej5mcXP4JjM/sH+mMgk+NGy3KlnbXqz
C/UsupAoANZdydRsQOuezP9WI08wJyenS2BgEIDvbD2/cZl/gBvkwvt0B3j1SRjcuuCgHkkXG1Uf
t6Clk5+IyxkM5/IY4lCxP8ZyipTjAgGJBVUc40j6Lifv1pi2jidsz5ym8VCgaOi78VxLSyzeqXgg
Py97clsrCsQGw9jPBfrUBnsgR4FdEBFd+ImDLH4kyHJu4ZMZ7pJeEVIp2uGCZbZF9ReZsRqztMUj
BeprMjaXdS55fw9j2bI9X1g3kEIEZziapJYhFH2Mp3r+sS/K6TRHDq5ePJmiPTKGREFsvsZLDLFR
g5TVjkuSIA+SKQtkA17GFek5aDH2N1qByeWDNu0NJhqjlLX18ezJRZ30YPxwEq0+A2jx2kDrdvD8
9QYrbeyUIVEMUx+r4cGEKEjw7vS79IfAneUW9xMaUGQEXgr3QLxOfNhr1nGZMHHIvHXA7YUdciL8
ZSStHyot0APpetrHb2iNAjIwFKXbXGuz240aqZbddYrt76HP1fSgAMU9xMRXEI8P5wUtu2E2oWdT
Th+MbmGG5LM3tSMCV/F2avyEeioz4aXns6WlZ9UDHM4t0VfFpgCcV6+1kR0l+kWNbpg8kj6CiTs9
Uvn/xSsyk3y3DXwXiX5nf2WVx20/7y27h2YPcIAWrcyH8Hd40JtnTJf4wpoABbejzTQjkjFkgtFI
2ql2+JO5f+cJmh1d/a94PeOwsgH0IYMLHlq+Kbdk6a257rJcMVrB5XmD4N8EuaJYRyPLAEGZ4Ycb
S7Lrm76juxcgPXeemHX1Bzu3MBH/T3QUNZsYE2xXJGEgmTrHHFSYBjySDeBs4trmbw5tkUSb45BW
z5HfBu0yokNQWsxe3Wl5TjqWt4oqXZxsUaGEmQ8QtRy9sot83mZYLjnM+aZdJn9DEBl105dEfgCg
m7B7jQ9Xn+8QOy/2kCg4Xr9xnNe9wSQ07XssBK4t2X3BnO/Ok2VjIyrPmvbr8cQ/+ETGlT2ic/ee
Wz5Dx8elQt//usXFYLeMwlu0LeF9/dBaz2l4/vmBqpJoELVcVuUYM+IOuimY6OPIiam/x4+KPCVO
ypXH5LijdkHiQVFaxsXI1bdPYXT5Q96z5E6a3XG0C/r2aiO1dB2eCqiruWBazBwJWJOvHsEq/WX1
O1IXZxdtT1hYHjQz8EfZwuqHBMq1hheLW60O6YWxsq7GHrKAv3qSs6rfSvTFVLJKP+qyIEPflHFh
yiJemv4aBDqI8KsCywJuasq9siTxHj0NSfcNwjle8T2gk27WoZymVNAH5MOk8CzhjzXHlFcLUILS
qYgNDPTQRGO3Eg11+GRKwaA9RTFUm2RV/Zu2jZX2epkHx968/iP90btttRhhli7FRhQw08ypnO2K
DOZadJC5Mimi6z4ITBLkePp+f+GslvLLUvOrciKVUKlj3hZWGS2wbn7FXxPnCV7WOcWhsFi7rSCo
Xd3zparnY9xzzrAsECZd/cfu4TmdKFJPXuEZu67s5SUcld9gczaTf2x2H/QOAt3UJjlPlmXPP57h
n0Wllyk27AE32W30hREOJ7qtrKAqElZNLqIbg0QUeWb/AJJaC85JgudbzUMWXp7G6hQ3FnbY0vJa
O9YMp2GDHM36iBMazubVZlXvEvbmAVjGywzfMAY1GQfJJxfxnOjklk/+agcUNXBary67JtjIGDgy
1smqBj8nbrwZCf0sk6RM/fy1fsEt/JMZr7zmvEPuJW3AY3SGxuoiRxhK7riM8gTA0STQDifUkixe
Do7nBIKBD1EzqqTCxlJDGHIHYzgerdtGA9o4kdXjVE1CP/Ii5m04Pq9kPif6zq1lhd/sosW/QJTk
wPV6KLJ/xR4plfdCqpp1pmVCMNSBSzfJLhHWi+9IPQqGYkHdDtHWCBf7DlkqAoJphiuHQV5aI8Xw
6D7R2jpwN2FhY0ElWGBYpEE+Lb6bWi2OVI4fFGu8HvNwWdvudH0CZXhGF7XCbDZPvIXdyM8pVJl3
nRt3tjxt1gN1CihLv865LauS2RMIZ4WkTiV58XN6loeowv0wL3ejZlUBMxqaVGkjvwBcIg0oB7tf
fTT2sDuz2MT9PiGIhMnvxzDZAuk1HlfDjcws16d2PrrVEla052Ou02brxpamRc1f1qLw4WBBJepj
cI1+KNuJppYD2hjihd4jSnPebpSN+98lNaHEq5TD1b8lzrtukoWo9TG734E9XF5G/8nD0m8sW/PR
8S3RIQyIlPbbeAQ0m+Cu068vm3F5xuGuonUGuP7flhXPiwKlyBQpahL0x69iHCCZKswYWVSVAdr2
RbN/4jq8SvRmoEiiUQbWMm+xOCpgSe/oQySzp/39LfhFeFtfBNPz7UXCTHS07IUlToJIrZfuaSho
UzTeGM0SKQVzOdqOIbFaGTapQg8zJVBHK8MYi5vBcz73XUKleHDe6qbwF759N4QtdZYgsmN23hWb
ZUpCKFgMnTHQhM7au+BMgCHGkHJtheDRWshFXtQlB2upErrZiCXtXdObS9Vzu/NBEjMnntHq8T2a
nVbHG2OWmZE80nt4zrLeDQmUhj/O1BO90rdo0t/78xhCePKQA/sUToyi9R2+LWI+/elQmv7PYavx
+vaLWa6w1+l1oa71xfWyyoYnsH6UqZyOxYAzAlJ35LXY/I1+trE8QuDH5QT7XSpTDhdeuGSKRqIb
39U1pGVbORMF3x+47mOvoG3UKB/jN4m1ARG/GbdSJtg0hQv621krvJDVOI9ApwCbj2Z9ByQk7205
+dJMLHP9MU8apVDjja8x8yJqbVeZnTCN4yAM4yYAvrF3ehgUd73uL0PDfHKlT+QjoYoXeN1oD8gq
IXmsMW9PmAZXkvgDquFfH7wdFSAvyD7jKX6e/z4yvdf/sSOBbo1jAJiCVT+zKl4QejQU7Z2mJ9cI
UFoIXPSLBdEOwQI0uHQ49tI1UWXq5bVKdD3hhz1edYKjl9jXHAbcI0QznWolqLeCMIFQ2aYcYVkH
sIsTH8OMAfSKPuSubvpGRAXOtBnhFHSMg7GZFfkG3idI7SEWAOqDHum8qdIr4wLzybJMgmss9how
PIKtphdN3dTUue2rpjkU4jEP9A3AI2TaFLyMaF/4nJQyfrszP2qFtZBaOgqYwC9/0BDzufnXFqbv
VFKbMNiNqYHpInz5sBBjUMGURcuG4Pu4QYsyUAPXN/sN/cA82lfAXmWVg5lJbAGG/W6FdkMpIOUe
5+IW9pgvJoG1lQ00EyGfSEGldad863L4AacLuBJ7UBI2Qbk1W3OkG+aJEVf5wobO9wTYe8Ocqs9K
k6vSup3JEhNnGJk6VOlF9FOxxQSe/kA3ZvY2zwHTi4iU6YLXAYSseIuphY+y57b59P/v8SD/zvL9
h/Si/Y7I6wThqagbLrNXNAJe2WG+Jz8/e6V5+BE+zZyyApWayXDsjdjN8gM0facZ9hsbrwMuZMjj
MYpRLNm/O4YBnNJquHkc/jJOibHl8BGQotUXWUlyCrt9gfDroFM5uW2tRjVfvkPvGMSeSGlkBbHI
MLpROofI5t2oGnYsPcRuBuBmnBdqzNrVbwnVfs9RN9bQpdTYw5yryW/bJhgbkn7CIHH4ly6mdlKW
ivpPziTkN5TsPHcSzdJBCj2fWeaUz147HAIHFJsTEjW/BU8h2+UaYb3fAXXRa0jbmnAU5eYSHNyD
6O5S3BgG0TyZi/PDj3Up0EC3RSjn8dA706M6/WoDVsdW+Bhj2Koa0/mnmqxRg2fDGwIn0yMWVQyr
ZdKTnq16GANCTXgX6AHiAhAEjJkVoy8KavByM+PtGISllxZjmfbDT13ht/4jmYKvft0KMVDYeM4H
NGND0i3Y1PCEhgYFqacNEVy6a71PzGyXUjnJf6eMkKfMYrsiYbLD8vSDcMgF2QpqGq9k/A84uHqr
R6/8JX4WEnZ2r8MUkT9ah31zNXIq2beSWzsOFWcnjBrA/twlNEyNAfgKQjC6nrr47y1uyLfzUWQN
x+WXL17VUEB8btovvsVXBr/GChpSe6uWAIMjQDO6mDvTSPXGodKv0rM0wKQjn+/EZjt3j0D2OfXs
9YK/Npoq04gjfzJyez8msgMxRSaUJkoKS5V8RO28siKPD65VkjU2kpC8CV3sCxVCEMw6Wbr65/RT
t2vPLsgB9DMHIVctLPI92x6AFDiC4UAIAU4vFRIi6H/lJXRqD6s2gB3+fgaw+XSxbXdaZ3Myu+DX
aVhwFc9cULBqbGUXJC5GpMBqgy6fIMI0WAALP6w0sTDBpfzLD0Qw15VuawTrcvdDY6n5/dZk0xYg
4fzfecCwjVb3r44xm1G+1sFni+nXPbnI7VkATS5Tw/shn0u7fjmWCZa91BUdxMcgrhQMW+FG5vfQ
fRZcI2ps60q+1HHXddoQB1OS3ksat608eEg++qBHBgk2ejcNwLb5mDcDNhI1foiblg+lV63vNMBa
0A1prpNPLAP8DFUkskOGCgVEfL7nNutaXkdNhslECnLA0cHhH1OANNJnVRW4/wY3sKUHTnHV2BsK
eBWugKBIZYRIxnfK06/svcwP3iDecDs9BoHbFDxjqFSNWF6cRO6U7u2nWU4IrJurjhmed5PWKrhA
IuOLo2Y6jO9IaIgrl+bAq3HqxmvhzuHIVsoDR9RFkqVC8bkvka7s6EXXJ6b82YKLVOSVQYFNcqLH
dBKlnchH/fMIdFH3r038j8wpyzmWHD3KchRnzLJHcr2a16KTlgqjHpyGsiAhVIysgaUwj+AM1xww
Bnf/kH4Lb+gNpO3MU/LSpmJ+b0UQnqW5eHmbg/RGMjlqo4D2NnRhYFvCp8Ydt9mUl8gXx/Kmohro
Q4P3pxNL5dLc1LVz1EzkGXN/9tzZVXx5uZNSQ0NTPGUgpzYUYQqENTkh2pjDfqTPtIGvedUJ6sto
q5aelQjkTlLpKJqT1wCOSn1acbIK6wbtSCIZ+yG32ZW0a8b+v4Vb95aLFt6MB/Q0SgsjvK/Km8bD
22Bsv6LhXthRvqnpZhdDqgasbmHcTtG2EJLrWKJwf1TNSPvpDrtLEm2hAOGABuJtbCK4cw7q80hp
GjBEETvE4Fv9od3eotL0i5iuP9aCXIf7q5vYJH4vCMFYhWsvPfUYP05tzWErr0GZwTNlTIkA52ZH
zY9Znf/31nTf7yHqgeRdPy7ddyQCi3d14p7IexAC7IP082PhTJ8uskcis7a2iDesrHKTWhOhZnh5
yxTrb9aG5pDDoz34054tlNk7wjEsH0Z5DQM9WSzPD2T0aQM0nAnS/b3Miuj63Jg2v+rU5V30AK/X
m1ohbQG5dpK4m81eyrdj3o3qLLt640PY/TnD8TxcxlHqyTYBau6wXPMNYFH1diJgwbfoTzt+g0os
epJ9FcgVtCAiLrf543t0oG/UG7Z+hNqdettWNB/aG3TfqVwxlafFOtgcqcFOEyUYsmznUo6+vw+z
y5P9mLSbP0U2LgS9hLFCIoAEZMhJ46UDQd+D9u56PIUTtgLn4YO4vbmgXRvLlW8ynYoRYpIGfH6Q
N4WblK9Q95E1pzhta1KP2PMN275ef6k5e/bSHej4ELbTQXZ93BWRpYpH3xvrD+oas0WXr7zJfnBV
EufUxM5LS3oeZTmvKBK1Anu/p+cKE41wKHed4j5rHqZMevR4qcRJifQahfJJh33qt5BsdtbfKUIN
HTsrfSkrsqiUQN/vx4R8WOxALzUAEQenAVgcSrgXE2WSVDBCSyv0SQ+Hu1PiTuTxUFZwrJnDA0Lc
i/RDQvUXb+VbkQqOoIA+zmhIHmtWWzCPLRqnbIIz8kCBIZfgMb64YIL7uDhW52wAwVFl5j1KldDl
PQge8a1PXwTeqmderB6wfnLBajPQWYei4T9CkCl0EUN6BH9bssPRUfQFybeZC0/Wl+OxxMA4+TsV
AbU6nIum6sE6Quf13Ymzy2dfGHjpaWsWuB3dU3HgpVypL6VpBgEL6g1tkcn4jdp9qJC7CjPA7xuo
+OPgZSd6fq1QgQpjyc/i8Sqy4Usb4I1Dydy1U5TNQbYN3f9PVMtn5er+0Cn273KA0/+0q/nVYiIh
+TpgR1Tvop9LyPtjCsxSlp26EFrPj4z6AYWz3d1Jexl6A050bWGf6aD9oASsGVqQUXM5lBDedzC9
VHIr1JmE9nVa6TOspL1M+A18Rxl8YSgq40w+JkzV3FGJZY6Whk+/OGghSawMFb5EFHa37VgYH6Bd
MqMyRrD/xjX6CS8oCFbzp8TRwzouro9pokuVyii6qqP+iWRGP1hVaCQ+QYIsmYIQ8lfF/Ivnrf7h
oRZV9Tqm89WrYunb0zHCfB+ENfY69rOVS/SS3+wyt3YFk3z+fFz8VCy+FtILDogc8eG786OuAWZR
Fc+Nt3Lyl5+EDNeaJZkuo+YEIQPe3QI8G/DAcYjMh+iJyaiCXVxqs1FFTyvESXgVixmHNZeZAoSB
Mjt7sUUrRaeACxXYEjd5CiPpVjtG1o7sqgm5rSoivTZr/LwaUKo7SP+QGfeacb7LFpp4Z6Njm+Vk
/9EEguSWL3w8LVVxG6TsjRVgaNrtekil/5EDfZ+HRXiUIsURmFCc6dGcmxMBNxME4uYDTih2Plgy
ZaY/Oqk/5xyEaESIhcNj2naZHOMnxqZutoYqnuHm7icusfPXHqOhQfiw90LxFXy6nAJLr51gVphK
YP4MJVgldPQaKygcS5qw6wPDfLVrgASEV6d/CvUD/DqVPFWbAdo/LBJcIuOoDi1KtbkN4U5Rc/4v
gC9Jn6bctxtBa5wl+DYPluTIaRJj41B3tSe2EM+jxmMsLiIQsNf6gv+IHY/2JGDT8EEtdGe+xgM9
46+n7saNXYeysk0Ad0oGA89wuXa6XTC1ojym52wY9KK9b3802rnG20HFkvBH6/I0U+d1RFRb3rHm
qnLnMTatOZDgn6sanUhsFT7W2mDECJlxemNmZvrSPIXCdxZjMa+Y07u/UvXtBPJmJhvkKdRRbGxh
EvRYqQDAQIT3LhiT3TKBfCj3Ee+le6Q/aWkcovyRN8tlrm1uEaYpeS3POnIUR8r2vwnApAEfMERQ
HWWwIkO0Zk3asyNWpKyfuE9DJptvE1v9NiUGWE/lZsuYl0CDdxua6SHeNRKKxXSIkFjOn7YX7sIR
jcBDBAczgYOPLI6hLch1y9/Fpm0oVI6rylJ04MPgMfyUiiZBuhqueDxK41MtBkE6XwLOhS+abfn/
MkxLuaKwL4aEjkAxWSVz3dMndKzZ6Stn9z+Xe15dhgfXLvpFjvxyjtomEQG9S1qC/eyTIv6/nI2D
UMM5ifhOfAiUHJXrt20hLoam/JuHY1OpLmoFQ8P4vI4yAIJRu7OuDYfDYjzH1nrylJ8gEn8H04mr
kqH8f6/UUBk2FvjZbWiYYXcrX8mTua0xP09Zr3MTmhlDGMiOF2h5x/1/U0qm/WlCZppUjT2ko0Dv
bZkknv3Dr7Uku8Pfmybbi4V0xGjLIxvEw8QCKOcIjKHEZMLenUXDY3CEJj9pKi+cB3pHWJ3s+/7V
A5dhM91nJZdQEkpgJ+VNaPf2XZ/5mcBODmMZ+JHaCOSWY6dvZkIh4J2L/YKYD8ud+EAS8pcSeeW3
Hq02TWLxpgewpQq3hKGJjBpxg4M4uIC2CV+gQP2yM7++NkhZ/PCJpP8+gDy3pDityvu2hqCUXQTs
RcVtsGZOTruCdEdp93/6q578NSHmO2wvNB9aO8zAVWn4gRvR0tpqtaVyqeTx3jmzVdmYM4mXLAv6
UQYGGOEMwrm59vmzNOjNpu427NZbxYvVD22aD0/IF0GaomMq4zY9QA+n2euMgXll0+HQwwlUmzgn
V6KpsYHgsxN54nriPQCDlal7IZqqjyLQbNiatPa3ea0a5dAcLJWFnmMki25tses1uXUOsnBrCO9X
hvWsa1GeKtbwa1XHVuTmuHi+M9ibK+Mf0ad9NCtIBMpB708buuJY+M1yND4dJY1T3FCiyUaygZPo
Usmh6PnNJervdChIjRqoARp4WQCcKMx7mzqar2VRVr/eNZ9PS7Cb9VpYKQ+0Sde3XaOFq9sK/5As
G4LuVHzL5VfbkKc5hqHWZKu1Gf/zK+4fjDVXoU9WPCrF/0eHFJZqbGqueFQK285wez92jECtNgLU
rJfba+59GzseGO2To1TrNHh3/zWvtvJbsVn4cwL7N3l7Tj6yagUfhYZ4sA3geSxoX6h887xYDsdw
2J8VWygknYkiNRP1dojCy7WdjpLMgmc7mhxuSZMXsNKb9YU42KDYJ3NHb/q42rHumDWeUMPX2Yk3
bgK9MHRYNcp/CygRiZpU8NSiZG/JPsh8NxW78I9Z5UHfW6W55iJ9dRq3MhrP9go8/zxq/54ue2WB
x0RtYaH502G4dollVIDX9KG2br7RjpS+wByaVqoQ7qmxbT6P2Ynr30CZps3MjxuWWKgjMSEnUCKt
LvSk5HlvmqVifz82qRf1gBMzZy6I1ilFER9mxAFkeU71JYaO72vyHAFWcde1Vo3xGaRdhQ9/lJC0
EUCVup3Rifr8oAk280UGY+ETaAwAwU78w/6qEhAdJeFhhUwoGEstqv3KueAHsRCWBueuwLO2TOhx
F8ENpEOO8JMLOPejOFBkkR4JasnX/ILRdNJAYHPm4CYsPhsFtltVEojH4+cuCMiS5SXpw3Ef+HcG
7Ut4EnZZkpXnXw4+mZjgYCYobREg1QJV9ImhSYgXJcx2i4SDsTcE8G2aKbb2/4qN5WY+LhoOaxNa
NGirM2TPHVRIrWvW2w4Vq1ZCjLsRZTtAMTOg0BMkP6MWfpNWD55kO4xFEz6tdod6MvHwoN3P/OFN
CU/pCQ6jd4EI9UbJDDCVLySII4rI87wULqr3lEbFzyCRv1fiPdOnSW+SkBeKQe2h7mwWO7EqCV4r
KFh2tB0XaOy1uHWmRZlj491unSWSa5HIV1izGl1+59JRwZkTQ9OoW1waU9Nfz71IYD2n5RUi+QvD
roV0wrgXHnMnJgv4r2bEAfwwyTzYZdalc89m4iBFro+FqCpu02eROL+/swaN0ckUxNcUOZQCs3ZH
pbVoYJf9wqy0rYI9RhIRrIC6KYouiuZofSVsnjJf2F7ZMBkz17vTXGR43Z+TXJx5C+dOtTnPEuY2
YbLCRm64AaYyiswtHworpbnDVKZPLYxnBx8A4uKFQS0Z9KTWVO23GncW+peJ9FKgn9MSBEgk2iYh
OyEt4x4DXdxRY6PjIzP5BBbww9GVe1F0JysTWI+J3o+yb5IRbNcNP8xsWq+6NFrHV+avcf8nbMSp
tsU1wYfBsKEyCqphoNT9vMPCx25jApQooIbDUmpumWyr7wS3HqW/9/RrkrMXLFr+3XyKHewL73h8
d3KUbr+qvLy+5taQfKQyyZYXzTKIHfvRIX3pX3ziAOSkupgZwTqopImZ++GfrpxUWb4rSw8B50hX
+dqn89slXbTw28lmPiJH2AnXpZ0deKciLY9WwCeCfWdrFdw+Dmyh7shRdq3/Qm6anM1Po81ceY9s
w1tiDy7pdnNCXFpYYg02t/760zTpJi5LfpV5a1fWECR+1gz6yU/88V3qyZINb5kqslXmsV52P0d3
bewKRMvzsCLaR00omslifwVlXdKAqiWA9Ryyqgwa2AmVVCZ+JrdMyv/CCURhH/6RKwBgZT2HZpiw
fDV6jEOiYsUFxQdlXu1KzeT0TlmxKOaGAduUHVA/0xihwAwwEFBNMuuHCbjZDd3U5HzRLI5S42EK
f7DjvNG/JIxWR5jr8DtYyToS9A6iROeHqRAs5LDjn1MhP2Sjvk4HIDxHDzeVk3nhPJG/y4I/EUfC
zetb4oIzOZCWMSzz+YyTv1LSUqeXVgoE+8MGJ5snuR+vrau0szra1bANJaY1HCLjvD16SRU8yyIU
Ijof9MVy6VzBoStMsey3wNWGEy9SQpwvL4hug6NNOuRL9hFwiZSqYXGhzc7n/Anq7QA6ngpSq9w9
0XmPIwkz9P+L+Y4trrj4Ss6Zj3F5KRECN2Z+1oktl8mXrNeKahN/MyQZVGfbAoKqYrBwi+Z7C8nm
jQRxU6OdCgiqmq07WkM9pBi7pMlLcC5dEB9x/nHe/pMRfGViDVj3xVAEY0F6NPG+8QxpbeLh3uh9
oCC9xYFkocmWzkJH7uYgQfk8hQqZnGB9H9KIgqWpbiXZbcO8+pDTeO1HG67BkDGIvb8f9A2KJzIn
Y74Bq8TrzPNVG18JkoPFdBC6H+87FyKsovSrxvsbdKsDPXwanzvrZKZLIoXoBsQVzkRZYQYoyr7R
LIqSwtUa9lqsJPRX7ypGE75uV9AKCTigkNOGbwtYzXvbP+nxramUFxAV1OKiHQHvpPIvDafbu5ki
JCTWW4RwRm4KqB9Pes0c6kisX6wDFEpJXxXzN8QMX8RnZfu1QmtEWdjycPjbt2/q+2j8gdTWmA+K
fLSlf6svI3c6RbU/BUAFnwDrLXCquIB3536FzKu2m9IEJp3KWn9yNzd/H9CjOtBaj5EhOi6UU3yh
4k4iYw2aU7HFEELXuxBCisinJM3N2DCMsoL5KdrY5GCsxHlFppU/KUEEOcKnlkKl15brhVCSPakp
0kMn0Lw1eXDjzPU9vaXbBAtPNRzdx111X62Wgfb1CGlSE8Zlmfgkxq/VqEGelwF/b2IrBMSIhcKy
pqKcgX6NOv2SBQLa46RqLqamqqn/Jok2VJYoGnmJsHY0sf7FQ9QEoUfs83Hnfg/yXCLJM2HWWSjj
HuqoRJtRzqRoJe3UC6WzbJpCHZl9qn6lo1JgqAtKGunCAJWXEmtRejIbhJusVqf4b17Q5+EFSnyX
f9YXYuPmCVsFHHXOEqN5zcUC0T0gfVQfm6ou6CU7Yl8JayvebmMg3NXF9YcPlMCzc/ys9GiRqTVP
BU5uKuageBsgMBl/B4W/HrFIGyyr+NQLRh83qNiu5twsDJisInSPCjV4FMDX0FnPnVrUVQa7P2PF
rAiiYoRMX0u/wms08zXA0gZIBLVnD0YWuLUWW4386hknORC1toxHlZlrN8wen6GfIWKZuhBb8IMx
Qgk2fQzbs79z41jMg37IIbOKuRzj6pXwwo+Ho8NnNF+LONpWfYQLz34mwTTBhCbtXeIPbQ+4WWLe
HaEgPU5Ww+/uMwYN/WroNcdZh0/t9P+3CbuzbFyQf02cfYW05yS9PB8grkC0Fa/rlrRCjchcOTKN
VIz5Ng92rUAWucDcCssxUKcm7Bpo4oNs9pC0Zrr1AiXy9kHIjb+0TMtVo6aNQHIoAhwIx26gG2/d
WFcx1w2y9LnSIUoolZU5MeDGWnVbndxPZL5yPaOSTFHb8u9AhHiXNn6/cxgT8J4P5AyRUV6PnXAH
qi6xsDVcjv/v9+9CUf7TfNDDaAhUuVREpD+/g1R6gVm8EtFkvV7QnpjVeshWrDvbtNXb2tqBLxIk
UbA2KNCpkjXQ71fGOaSzcd+jFLXFxXjCywwPZSH4kOVIgOgzlRUzTpioJ91p4luZInBGdShDqkaO
AzyqLbeQGogbBYeMF+Hz3Bn0CbceVumKlwPuOTZ6vrQCZ5vyOySZpzbkiy8EpCCQ/ERkzd//cHxH
fr9uoebSuueBRLje1rVTyMBOu4me8YKUCP8H/3qRWA2MljEr5B2NFwzagJwGS/LzPVH+f96lyL5V
aeDtRk99Mzouml2CtaAGPXpY65s4/u5VMC9Io16XRR0UQe4bOM8K4zTd5oR0l7+kpV00QEASHgtx
mtX+eHBmzfur9ZPynEe3t8Iz6NRK5bHtUXuHwWqRgEBVRlE9UGM0FoIbElR3BPaVecdf1D9G9vmx
0ljRVOqoKrREm0aDobXngNi0fNwWCmFTRMT3IC2CvBAzTxJZfjWFHzjphadz7UmlZWkwpM9dj+qV
GF/zkEwLDbHTsfhxFMOjbrXNXC2ND+p1t1/PSI702xvDr4xpdDU9U86niIhuJx0UYJC7sYQgGWAz
VeHWETNMM6EZLzY8PrC0c8N0b1l97S08t0oCCypc/9iiwhhAkk45y7i3aOqATuuDjIcR1vJpTYDb
Xr9ZEID65lNwLQ2TQWnLdBzA3XDYlxBwsqjl/AYXhOce4QcC9A7UH2/sjlNodOcRAzG9HUWQ1se2
6XApUnNwQKSasgbS+bQSFMGnayuAGtqXdC+cXMo7lTjO8PTuDIwlKfEMRTzWFr+CkIHu3GBWYwvE
52LtamGIMN8NGrg3cQt+7M2U+RFZmCcqadKi/LO9SfxJRc644rdk8m175vuZK9dpZ1jUloRq712x
XQUqQDqNaWEFbURLcB9YWmW/84LN9Btr2qQTrs++Kog4EcDXIZC7vp/r/H/7NX7iV5sfs+TIBizq
AqdGXzUO9AO5Ea/TjgsbYL6BzUZi4VJ7qWymXRUUY/7sZ7XOEGH0l4Q4bZC3MSA36PxBPdEG1ddA
JACf1aYzDBGjf0R7QA6NmrKTL3dG76ySHTIPwjSwT79guNZi0bzkoRNp763U0MonsJU0TWAiWJvI
FMKBxjq9dOKqw3OWArxzOsQYX7YzCvdQbNJVHLlkQzBW92FOI+XFv3SiHvURO0UdvZzDu+WQmVI5
wLQ5r+Zr1CcwiVBlvIv6h8AGYF0htK2zg5cBZe09IPCDKGri7l8sF3OAMotHHZso/gx1v1CqgZGR
Ln0iI+Xu2DuMfcenPyPFI45WPMz7rrwcXkUS5YxusM/PUpyNN5HbHEpYx5Oqijm+rAMm5TErz0WJ
wMPoEX+0W4MCQy1ZEbcwyCGSIrO6Qu67eOnYX/FOUeawQ3W1C0fZiN43FqV1QIAdlQMp6UjK7Rgk
KlmMoim/ovCeQsH03z1m52bQCF9wVJji6K2JwBQr/8iaZC5huKhUPdlYaWoqvO/u57MZOXOFFfqq
dAPKAc6dbSFXMhArCb3VYqqYuCUdFxGy/+zm5fIoFRDWQmtMdlDs9MKo30DwL4pp4KLF2TD0tzX8
z6kdW2nxLDL4sCv1O9astxBVBdLaFMSIIrVHalGG5iwwnkm7Kgx/l0miM00Xz7+zm38Jr+t+Z5kH
c+6sBPOrcXy6LEwwRew7S5SSo9qYez+w0SfY+fGAV99eTNacgeapjhp7UdetZcMG6J2vh71wtYvB
dnFEDuyRnuRuCqxHmzT9CVrbNRibxi2hrCOpRZiIb9qyNju50J3oFiS8AuVwcVrwgbhXIRtGKrTA
XNzV7AJNT/bmL2xGoHUfTuFD5ZA4eOkrpAd7Ti1NN+mwbnn3c0mHq4FeDU6jyz+FrCCAylhbjT0j
60LrftY7DYrL5aqLdGGwiEvxog/64Pfd48owMtfJL/HLEviHp8Pmyron+oq5bR1Y8qKmQSCVJKPc
4jK6Ws7ZJPjwN78WyMTPI8Snzm6Jx/3SiHQ4sU7InmuMjZuk67SbjamwTNmilXF/xAzMsjHX+eQ7
+a/5aSlERpD4IB/GUXIQTgxg5b9XSLf7jNJbDGYjmheGGazxle4SCW633vn/u3sDcF7WJTCW3nYv
mxpMzAgmpCe/SkAnmurn8mh8Kjm/Q+F+QJBoQm+4/YxjnkODAVkDhWuDD8RDNpQZAfvATFWHZPaD
N4CTWHIyBVnUjybBBD3QI78XhY++vSKuRqAWnRKJz4fqtTIBne4DDpuNCEj596Udn/IZ/2zB7zdf
8gcKd0vDHyfiGJx55SAu1EC0Lnn0MNUUKiUaDhHu7jtVa54pEoj9mplajs1VJoE/OZDgWehCAHSM
jZxIA2z3dg4Cha7hn0Zpjk8CkB5uXI2vkrvpEU6Ct7MP2nPwrVDkIsdhJI3EjXEcgcxfoh44ajBu
XhWZ6ENw0RVoU8tyUU0EL8KU6F6WWC+mSi9XQBfj6iJoHoh3letOEUPLqX0NQVzaTMrnPoCPwBzy
e63OH37lZOkddmLR/ta9HKC9zKx4fBfjt/V5W+k7ado+ixjykK80LOIM2SkNmSzm+MWME/NpdDfO
LJRZwGtA8fCEY5r9foOGodVN3qpAlKUHxMB+J6Pj/q4Tw6pvFtvjQta5Bybzcq+a9vKOYwXw66Tg
qY9VtrQX67xw9geeMqcPVYwI4AGQ5ybiauj+A6clEOe0iseatVtG8tQSCms1gY/8RvXbVt9UxFkv
ziNwNWTo2XwJjS4KbBhP8ALKu0cXG0ysy/8dvgIqjTKqEnamdixxcvV11y3oXtWbzKU/44WVjSyU
bCeZ0dZMR+ILkE6TvJSMte5ciZ9M/F/eat7jXbP5MjAZOWHt9fP2cW38INTbAeJjTvCub4i21zRq
rf3Uf2lnHJz5+em5idZAjw1igJhYQL6cxYzluKkR4E0+JRu+Td9aUek7RGtISuMYsVBhfN7OyrZb
JwchjcGrvxuHnsy7ehN2mxY8Qx90aLfHGyRFxP5pbD4mD7v4pB/0C+gMAc/kZi5B4efpVJ5X1lSN
JKaWHS21AiaVv+vHIlzoM+igPaOv1Pt3yuJ07RHisuIpdz1NO+KxTpDttp5kNNCmJDpE5P3Ak8e3
cvUucyvoZXWnhJcJidwC5Yhs3Cs7S1PyIzy5JwTf+68R3lS72SLtcC7k60EDNl+YmPsgsgZ/YsBD
vIG2LrVQoF4lNaz++NQZr+RMh9XbO5sTDwTkVhwK9rg9DRnbUgzYkAdMaGU8rqSopPkhjOIqlBJl
vN0Fn+EzaHxYdUf9tkbpbwzpf7ES5KKC9qjoaE0kW96nsR2Cb7ijv1Cg9eAyZp6KoqxsadSKEjq/
t9aPDfWUf8tWDdHAxQM2i1JTkrW/Co03AO95MwSbHV2GCpOYzfViD3h7fbPHP0kjhMoqNO73ugJH
2ebN3CvEQoRiXgtNNRkzHwBdXRt8zoZ2bphSoU33vxTwexi9RuCaLO4kP8zjCOkpyyNFW7uvIqaH
MEv4oLcZLR6jbQHud4v5pSOmGrH3u/sGKfprYKL6QSr2VPwqs/HwCSBllAc+tDTT6NIqnJ1FklJp
+ghb1K8WFk98wXoK6mf3JzELC6UtzSFJm3kJstR00Dhg9jSr/5xUxIXqipgmUzeYL6zu1jdvMbT4
XWJG7UB2rNkFV4Vxks0v7aM1DGTn5rNzBaFNGdNFSxj7Jw340QBCTrWwQCbItG7v8el/Xc9K9Y+G
lAdNdrxqEuX5Xx6o3Oe6wjGBWdJwKicMgiHUBKfeiv+0ydz5TH72gSkQlqW7foOjmWB3w5mUMztS
5PcrZi9Tpa0M4kxFekWapL+u/e30nWolvz/B5gvJhqL1ZjwihEYPZFQ4VCjqc+Z93ALEzJ/Sugtv
KqzhOjc9m/0CKA5RuZhL2922LOeXL4o03D37qp7H2wbaWDKx9Jc6n86FvHMG8cRj6y6FwSlmQ2Mo
NRJPJR5Afb4bj+/GEm4cUOO2n4sSUUopzO6fUYgDTKk109WggnxMs1+7BycjEH0dxzJh4EPuUTuH
byCR5EKIOH6RANwMdK8FEVffhTW88JrYNsowaK4k1JSIlMqeelfcMK3QKHk1++CfR6n5/oorsuI5
EoJonKW+cPCaeiXpJnSb9nq/gflRGZCF7QA7cUj7Y7AO7VAtyzr5Rp56KXkTG+bY196EtR9lVTGk
zgXxULJ6j+waMjN+VDS2ShW1gBUesXXeGvOAmDk7lcMQvBKMaLcYXJdHz4TxgWd1F01uoqZjZvGK
QQu40KUKRCw2DbcFQnNDj69VqcATGWEhyQ7a+w7gfr/z5huzoAst23nZl/FNRwNYmHOPviSpNH6S
N0zYL0MvEz9/qSj5LbCnnRUOe5xO13odyj3uxseKX/+NiuiXZtXs9/HtoxAuHeDyAnOdl6ru88Gc
FXv1uYHakw1YdXvgGe5KwA8mplIz09rHluSMEvGfAu9Nu5+yo7ZVk7dZG+QErY5W1FC+Ky8pslQI
bGUI+kuZY5tsjz0X6XSY4c5283RrYGThEekRYh+0Y7bJA+DUwxzBFKCLoLnUhJHzyJZQScRFACrS
QSDP2Ax6JWXPa+i1LHE7+cZCL53/Vo4yru5qkxn3jLMjEy2kd3J43MiDbeG8CYK8XlgxRGKUwi6X
dGyqXFckYcg7QUy2/CMNxEuyBcwICW1cwu89Nd6iHzXKEX1T28zzhonFdjeLioxm9UMB3nbL0rvn
owQ0mVr4D7Ts01W+c0fdgeXuA9b++gc5gc0jL15YSpui3udGPsUmrXRE/SwmqQkQH/3Og5PSv5u3
AHnvexoOz6Ek3KCXy7T8xyLHsc8056BQby5vtpYcp64WW1mCu2+M5tRmyrIYD3+wIEa7npwioL0Q
VqMIztRkhsrGJ06P8SNM4UxhF/vLuVyzJ8v7ruYB609Bgwsz7RG9MwkRArH+7rwHROWeHRb9yODS
yo8QgjpgZP0PSgWDqrD6QeADxuLSlMtx+A9M6ohL0huJJmgxU2flHv2KUBbRy9DSrTH3/2e+0VsG
GRfpxdKnO3jnuUl40VA7Au12ob+sJLOaleA7eFSAvJX0q4SBHq5phQMSSQVDS/rNdINgUVn8k20x
nyA/jlhn0RvR/TE3DYpoovGjNwHoKE38wbkiED9EPm+li6vISN8nymD4pXEYa6klcVy4bWS03/zr
b8fKmr+pQ2quzJ1Zh9P2KgZVqfZhPL2AgQHebrlLxlNjvrxGcW90pZ92m2C7WKw9jONdlhuNyvRd
RLBW4uG1qO4xM8IQgLXKBvQgoOpHPpO+5z5Icr13/Z9PyI6YDtqv0cnhCjPYiOPrlhH/PBM6hMwQ
eNhp/jOLxO9gbGXN7ki1f9Wzm+/8xZQeU4nvZpOkozfZmswwDvBUCOcBqtTDrmGcns530U+Gj/9a
mUE060SufK/eDMjeRSIXJDAOoukLLINnvFz266/3edAtf0ysiesyO7wxoIh1NW8RrHGRN0LNgWhq
g3meKsGGsckylRyPy/4ObgezNFoYnNYt8oHlYOeR3MNr6ryVtOXebHZ2q8Vj+gLVmvBkNeIXkua1
O0xOJncgcUeUszaKKfa0Kr/mv9moxM9hdFzB7bzNaZclQydxdk5xYzgUkar81FA1Svq3vqnSthlG
2tGgmNjuFGqItOQc8Gt+iC//OwyK8SEFpTmALQxIKQ652UmaUGvEryJUIeavQPHt71MHT0K2mGPi
kHXN15LRkTAoXMHuY+YtExAindXnktN2z0O78AQniHHu2Cx7W0YhuIDfp8igUJa8JPQZZKXcPEAU
EyYs4ZXFn9R5kJaFOcsFgRQtt4NZ73bnZGpD5Rv7c56WbjwNDGZN/i/d8lh2nlw7RkvTD6OLKJEq
rMM72bJHlo2P/vMXj/K12OwD+0/LGm+Yq9cMlcAiG1DAAaTRasN6ogmD5s9Qt+Fxn9k3SE1Ad8mn
TTVPWDxG9826lVPk9IBmekIPjBISRP4omcTSeDP/0cHU5aWK0svtGVTykYTeaQ8bb0iCgpMdspO5
jUuvsuxuw+4oDOOC3j72NnFaIUyhU9OrOZsT3tm2FonK7Siy1/nKLn1HhuZcZDNoppSaCJ8FVzuL
tbummO3JGSTZUYp0rrkDPEdLjRgDxTJY6m88JRu+gEvSM/VSEpmT3JKNgaa+V5xMeGs7RhCWg+YW
ZxDUH+g7Pm0mnrpp8IMW8ZQO+qF4PE/M2TMoFg0NXzP7SbXRtIPMARdetjw7CVWAXOY/4rnMU+NI
Eg2nE+PAFNhn6WCKCStrH5IQiuj6ercIpHwGeO/nGiP3tk/IwQs8u7hX/pf1vcxQegCG5/2hwV7X
Ai3ADN9CzirszWxaGQneCo1JRTuARb2gwhxXsY4sxVPEmlW5jTdf9c1RLxieEkMA6q2SyJZ2bzt3
HX6zMTxo1Y0tQ1WzddPZenuc25rkMQwd9cL6UrOKd+CMNKcVugjWV1r4695WbwVij6nQWzv8pXYJ
sAfnj+/mn9OmFYlOWT0Y6wAWvSnK+xg4IYSF/ZOt9LMYaACCpOqjmUubMvzSwz6bFtTEcBXmrW0H
CUyCHDlkv8XVxN9UhfhmQzWNMf1I6X8Z1mZHddodqP8D10MoD6MwL6qt/9gklH4bG3diftwUWLBP
HMubXNb96RGE4POdU1x+tTTzq/fPpZqmO5DKR0dVU+gl3DNJLbzmpA3LT/28hHSdMm6yaAuE/gm7
ufct7luXk8vsrPuDAjeeynqoXcT3rVpVYVZPEoMMyiHhoAuWQEbMqh59Sfk42eZR9Yic+ROwhYyB
FWXIzwfVWPWWOvJdz8qKhh7bAW4/3nZbLrGiYBH1zPO7aIMeQrKQxEynPh0cEB8MMCFB0dcCpzMO
M26W3wqUeQ/qWaz0xa3lSPXr5sPq3eIUX3q26lMYPIFFnM8cDu6a5UduBErc+CPq2qWYCCSs+kOH
mz8vuW2T+lp+CpPnh82s3yOPfzO32bYYAOMnc0cyrRAH3gEPGdhnk/xSLeNY/XWXaJ6OsYlHeezc
24Ki4G0cLqa8SDgYXrrwLJuFffTJFI153yF5q+mueuJcpB1Hd0XQBC51o1I0ycoR6cb+NOIky+nS
vEe3xEzYgX1YuD2qJVrxeQJrsyR+q9bIMZcslP1g8zoYEnpKS5vXm1heOrUP11ZbKG2lGH13LPts
NVqcovWISjJbwTNEm7FlS7Bi/iBRBhP/K4hjYSDcoLwFkxYA/dyQ4lx5tF/h/nGu1Fsaag8O0ae+
uyg3+pY1C7y+4tgpcnw/wJVt05kfog8eCewIfBFHVrroueaaytc1A0gWCz16pzyN4KTaerHBcAf8
y1klbmGqrAhGqsUAK66wp/QnVhlvB/PSpiTWvtS1u1kt5S3+m0e3QNp8Y8SLdC5nc5UtAM11+FGa
r1KpWriNcqpAMZnJDJNqPkrM5oPhy1x6jgg3Kcc6E7FWS+VBLSG48OpWftGLwxCvuaCGFvWMWXSE
esZxGHqahnYGATCftcCfnWtHaw4Tzh9qvcMFfKxAxwbSGeE4MbQyaXrFFdAquYScWa4kewa/UQ3O
yyws7ImHU94ChVN8O1XWIWI3nWIaW66z4VficfTn0tAmnyU4dK8zxxC09JFRzUF9T/klMIPXttAX
BalS5IngGmU8XSRy4b+89P7p3iOIWY680ELr3x0VViXYTUZWRxF/57rqDYQdDoTeLGAEukCcl00x
SbKiL79FeL+xoO1TFdDKf553OHxAmtQ+5KFg4kOG/xVnIUxp3Pq62O4bsZ+eEPcghYg5pxsh7uUb
w9ZX0pI8wPKlRPvOnNPcSjsrTriIBzAtmjvpXE8tz7kMFDReOpvZoxXnq/r0lUeL8PKC70hLz8hD
hzEvuWyLHQcp5dDJ6rscq+1xtA8hfo6o2QyZcQ5mQLWyPuUiptp49xh9uqYI3/mILLph7b77xxKT
06H25UVnEqkOKvCVAeEFElT+MD68YgYuMOYTkDrWASB0R/bwReIizZHPTVgpmusIfjrQh1lSzOBL
vVuz6OpG0IPfBkpkhnT7sK/nmCjDKMgpeORITYo3SkyFAwxeEX/Dm4NUo9d+IrGlAOAQFN+TG83J
R3RsmHId0BAh62o9DILL50AzUdCYm1nigbTs2jv8E8PvW+zgWoRFJZTpALY/haslI6068Fz753pA
ZBSM7/OMTL5Wv7z2wyv5JabAN1O9RftIU/udIKkIxsyAQ8hM/KHyafKhu0ouwhJr0TZ7BPiCR1ss
l4d0cITNN6cDAxCF7V0MGFj2axLDbUYK7/yrt1nr3kysMlDZ4bL+pLhlveKFiz6rcIP8ldVBWJ/e
uKAnEzbReI1SMxQN6pW2v9Xkjn4eajFv/rMn6OuUf18bbzXX/qiH39gRMDMvhX64nngZzik2bh87
q90/spiR6784kosjKpZ+h3/n6SJA1vswnrxizANNYjVbWfdlqsJAVXrL4OkPJMx8Ln6F9O9fe1Lr
zYJyrIrjcwKLYsR4UN4oWqKHP1POwE3KepDjeyh0X8ErZSFCEzIEGBW3YnUfJJ0Nxlg9FBCPfkAe
mrQ75Vh5SZ7zg9dpMBk2gYwcUapKr6mjotlolnCIngHv0LTLhi6DSZbmghehno4W8Lmhf42hmgnU
QRv4L7QlD5g22Zxyi1+OVLIoz1DfU9pKm8SyA1OMAgtdA7AK6pxGIiLqRnn9d9npaKhSBmysVws4
gDkfDagIEV4Wycfa7lZLd4W8+isYshmccASBQ/ophd2VwGKR7p7ZA3J8uHoBgIhTOGjBmZWY74XV
EsHtEIQUW4FDjct5DAZU7tP5gurk54cBbWqQVrC7llJ+3rBB444rxzeEnt1d04imA7DCk/s4Da8u
n0wXOcwYuBYUMFu5xtEeMAMnNua5Sb7HZ84YN0Ax3SPhaswCusLpZen7PtbGzvekYxIHHH1wEPYC
iOgR4lD/fnAwJ9FQuN2TXxReWfYCXTPYo/TIAIXjR71fpJMkTqala5UgdKlAZw/rS04IYqliTUEn
zqIz3XtVl1U8jnhHWYlbzrFupNF3XW8Gb13Cy2UttRsDrXMp5XQsbVgsOFaBjHGE3ezHs1QMsfWt
e9YJBQBNUMTLsxxx3roD3/XNiVed4A8QiQBMLEdMbaVrrFQCw7ZT3qWLby9wvU+l8CHMDu2TlZsM
FmrTxOpORX717taaPllU3siGQD0dp62YuwG9GAPhSAYSTCizdNcGOK5tO9LnUJVuRUJ8mZnnlbUH
sJ50StHeL59AqL5PJZzjY+Rml4fFUWGh1GnpDQ4j8A/JTugRqC2mm9yw1BNXhq5WVmH/S+pNSwbA
mz6l9aWgP+Yh4aRzA39Jwm86LFBkPOrXtDomOAhwguPe1K3l6otfp5dpQvU7I5vrBV3dh7LcvnGj
8ksU/CKM9J3zXr3AHMF8kWNOA/x8VNkxiSrFcheg+yHPgK1IJhoFvTGqPLb1TcB2XQhMZcHniZy1
IACALJRyFeOj2edAlD4wZUVlwl70i3Wf8F0OW0FqV86iy/MdwkgkevDNZrbDUuiCfgq5Fu2jhScy
LQCHIFwPis9gMS72N/zLEZkmNKvlav39OL1IJ+PvGSv/gDgZec3RXmspiGQX2F38EZwzzgjuGJVa
zlInrvcGcGa8vRjNXY6w5Hq1CS5GmNiufVcjgj4vmoB1JpC+tVQLyx6DXv/EzmTuHkZHBuXm0oHn
mQ46rv0ndeqCNJkdMdTK/mVhxtDd6gnq8jlv6zzZ2LDLcJMdq7jrHQ0HMTS/pvVz5QoQ5LOTOrr7
G9VTUw2/+6cix/WPr2kTf4aLUnGTJ/r35c9hdvZKFDn0ySIzfHb6qMfVG1DB1yqGEH4XSmzoiuh+
+pdujK6QBmSIh7qrT6aztaGboW3XHtkPAV4HPyhr3Vd8q5av7NELVdRDqaPhmKDgtMgoi1JoTNEi
di0/kZ58mG0Sc8Fyj4o5HHWaP7xrGZcd7EpjkXNTCbi5wbzFGPCqEhGtwIHt9hL7ofbP9M/1uRZg
muCt0+Kua1jlCkyfN/YfeyVcPM39gU3OLlttrT9RKIMcr5pNdg8FvqzWkiAeKc73ZaLWlsvIOOo8
dZjof/AwcEpmyn499UEskXpxfn+PIqMkTOXG8JmlKhZ8aOdy0gM4s+WzspatAYVBiRDnSPpbp4Nc
H6CMX1ZUvipYZgobNIg59pyBNik1MGJHmz9K3UjiDfFC3HKlEQsXrtP5ud3s8klKTmY0Q6L3jADc
2TSijXBvRp3x+rrzLh/VrdZ0hb2dP6cZ+1472y6DTU6NORdb98afZh9xjIBwmi2bxsrIjTX/xlWE
XWxLjfy6UUorwPshXjnasxt0hS5i6UvL4F0tE28qHMeGnUv/SZ4muIxndXAlxqHX6SyKoBL9WCQn
V5K5LbOSKS+dIjsS1IvfOrY23ufBDdDCfrnXKj666HTpQ474OvQizXN0JJkd6cvuhSAnnclL6qIF
DLleYJGxnLocexpf+Ut0Z7DefHi2Aj58OuwhWpTultRc5hKBkYBrPw4NmLyD7wplkvdT9ekQLSUA
lYuTmX/fQp/dOyng/enMW68YT+9Q35/+d1WBam2+7aZsRbfr1J+yFbMx/EeATDnmTVTVQAi4aewj
0oTVKynz70JF7jxtdxckxHe029FNgRw1kH8HGKFEC2ZosOT5FPhX09y4RbbGarDGpIDE2/ZJCpch
ppS0jtxhMUiB5wkZfbWP31j5x5X+1m+g/R+KaMrzuQcVZYcnNkhG0C3QHjdI6KK+GrGcx+1Plp95
b7GXg1oJoLAmKbMYM7TKrdZSX4fZrKIx2R0ZTV3a612oQOXNwoP4inzN8ushq0u0ASQjjW/lSlIk
HYzI28/O+5WPtB/0MsclHcvQOlGt4um+t3K2GI+ISeD1PePy2pzKpWf0WsDJaoEPGskNPjDLjY11
zqabNXKD6sKOpzZ9mNwvGWYjZ1wwezpNHfM+UmC41FWQF0XRP1NpLLez15m9RS3iiqxhPVCJOia9
AB8LmrQHjKhOVBTydhpx/H/T/8QDdOrsz9ozmVc0Dxp+xJ+Hap8h0JNh6HRLhXGU+Uf3td5ARCHT
abiM4PyTueyyzrVMrW6biIyHmjM94BIZN0EGrQqKqx8MaKfUPDoSfvDvtdmo3SCOHNA1waoDN2Pu
TI12OQBOS8DQA6sB/h9V+wX+K+QwXhHqEtyq28iaLNZkephFi8GTYT0hiWJViD390WXAdCubeZeD
HIUCFy1n+6zuSKIZO/ZDN98ipywldfUHJSA4/JbR5je5j301o9eSLXobFm1bPx4bv564hOzCOWWq
1ufakd0AcqspF4AVUAuIDXMXUv2nwCrtvdUfHxbHTsw96miN84RNbXvHwXOF9dC5YIT+SLMNmAFH
kuEoZU2cldxnT6j3VV5MhpyAcrju4A/6LL9WkGrXki1n9uFadOk/SsetUNzzYatv/eaXtthPXKUd
eQzVa6sZAaifj/6bsrI4F43NLcPgeuiwYfB6nZ/WoHD87oXbc68mFOrMCpqLWqsevST6/4Tj598s
hchMvdtUZ/RMz9SllkDBI+zfHGGopEx5eu2aNgFsJc4xKukDS3bDSDfdfdVVgXtzjEbQct3AjtZd
IHi9Lj5vHWF+s+pxFwZMYV+R1UHiLBsjx2IUs/QaEQfJFjGmYRTkmieNIkpk3WeKre2a8Vem4juV
Rjedeuu/pbPZca3VtpWEsx5Hw+KReGb8fbExcP8veDMKMEe+gAd3pMtepEJMKbngN4IiMbPydVpI
Lvi7Ns8zAvsgTkQgXJlj+i/l8hECqL6Cu+LK9N4DF9JNCU4sm/CWyGiYUROniMGXsenaZzZfms1E
vxznvF5zuoGUbpPpUZeZ7biQy/4n6Ya38+X9yxBU+Nk0YcqIP+5f4OfKcwHDneNfaBYFqQ52GUWE
Rz/mcc0mIO4404DupyuIAn1JbrvCgSUNPNj5yKr1s1abAdjv7V5po2vxDaVOrQ2G0ROzxASaEJtM
oNw1FkuKajWfUN+JwuLWZLseF1MEkV0QQnvR87XYSZhrvjjNJBZa7Tk5ZPLqUJ6oS6WnzRM1a4bO
VPTCR6oKQ9Gp9XXMV7F6g1aCKWNsUIXayA7UOdiJJgn8uTlh7fJnB+91my7QMko4NpF1/RnPdseW
r0ZDn8sT49EmPNWR3EjC52aPRMX+08n1YksUP0zvSudbARi53y9ZSEAR0Bk6etxWogBKu97ESFd8
ZBORWc0mpPMymoH04lyz7TfaAvmeVK8GDBLeQRwCXKQ19dywTEELwMizJgwTzEm6BPCnpS/4dslH
xvkG2SauqmMvMsDVuqKMYLeVJiXwNyLiieJgLpWsQC3HXv/O/+uU9IoPOmBl7hgB0paUqdPT2pnw
ioSwTlYwXWSHX41FtWissvoUvGCzFtr8tMuhH2Lue0jwLGgd3quIGQnWwBc4702N265sjhakYobt
Lzuyzkp/3WmxFuIZioUAan0in3074t93gRf/CT40pcpztMzEQJOI8LrlVLGbAaaHduQ06dd2T5UT
rwsrCMJ6bRDAv0GU6jgZRjg8CCvApoQxar/zQpD4/080Kp65Dt+cVo6/hVrCOE6b0iA1e+VfUefm
IzJDtBeW/YO7e44zh9s23GlLhnEcYir3kOFCwjMpj0KOtXlJqL9KxE1dFCTkFeUlnMN61AhlMAOL
Ah/0a0RNu4ug+Sevwx8bww3QOXyWs4pXfNXZgxbXed6aY4gne28KcXEBvnopN87uTfHWdFvVVpNT
wIFVW34s7COw6Abdb6GCp0rJ5547jNoZdfFg9EaHueovdJNwbdH/YkOjsFtyiUiTIkvzlFByhgNt
oUfYu53lB9JN2e21JVyQn3CfviFH6ulXf6G6ZI7vQUSWB9ZlgFEQfhcq5qrOw7bHMfZZAPp9RmMg
O8H/om0dVP8v83HEv1RJCFelXd8vb3DeoLDh0eIXDrwr9Ae8hdPOVlrv3wt5FPQNsWKaiURQPf39
gk5AYqUxJDfSiOMeeoaUk0GgGYOFOarj6n0tmk6n/GoE50UZjUbaWmcd2v+zsAvT1wwMkw+FS9SO
jqN2j0/6u+YJCM9gOHOLqmsDC3dHgtO8VSEPgcZs03cQ+1qC0Ncaw+zsBWx9IrVGV6Il7NirhJvA
4NorxoOkYfNC9n/HIODzC94FO+OzvSwWqaIztr2IS404m8uXTvJivTTUNSifhwmpgDI6XxXDIKlY
8tFeA/Xke2M4ptzI05oVJf+YN7Zm8jajY7ml+4P59eSBXiiJhsdUS3c9/J5fC1U5jb11i7wuuMYe
7uT5Reo6Y3PMryUVPAII/+y+pd+BnNiAcBBdK/9tnzkKES5fEVs62TnuGvzNoRpcLkG6XskPcYIt
9AJUITcDDZlmySjRXJWGcRfTIZvxnP1r/oFXU/WdyqB5TxW5yx5McMtpTIO7eMoKmhmPX9DjHyVJ
YWS2BLq+bvMXb772TKWFbDjX+UGT6NoNX4dZ8Q46FRpY1a172824+8b8YTodLXbXKtsCgiGHyAK5
FKSoHl+QkTb5TZMFJU/YbIzk3beF44MrxDdKSP4/Z28wWQlc8hr+6l9bOVOB8FZM1S8QX4xF2iMr
p3Isl4i9zxP2uJg0OYdWXTqTuCEw0OAyJTr+fwsQ5wjeMqdMJ5DI11cfSOKKC9zFK99apiXP7FCN
30bew84RtobmckAO9k4sqVPOrYWbm1Rr5W2e8sRvPv5MGUOXUiis9Oz3m7HC8POqApfs2NJ7zrr1
fsSIB83wIMzcZ4LHCDO2tIuUvXXcWyzTnsRSoyaHBS9GFvxRgf3Qf1BRmxjBMF/G5liTmei+uVFc
FzaiRTbLHR0oe10nTnEjHGPQC6CRNwOTUJhxhuo29k+Dlw3CxKLfTaZAGtp/vW/Jgb0MJmPMKA26
v0zmdoHl+VhUdl4+PghUHo6oyZo0m6AicpWIYl7o5sWE06t1eVcOdosIa5mcK3sRU7Jr6oXEpmt/
75YFXZ6Arl5eojeMtjOs3wvNWFATL5xf4Kvro2gFl2ahGThmvD6rZAjtflAL6Qw1a0QxEl8tCadD
vGjqBxJfr8r3np2S2uSn3aqf/dvdzitPG+j9a5EwTa4xZS7+atWX6ab8Lr4qAQmP4npECMoufLIn
TF0z9BJuMKfQT9IiHxxTlIBMvTBPdCGndx4pNtjXtoYiiCAorppl5EkOLR4sEAL/BjfW9R1KSplW
1bz3JpzTthbBMpFPAVxRzS3dBrziTJ4KfmQv9xS7ITJkJv4e1/hxqmxGzNIraoAxavqnKmtLllUH
umfFrVSz4l3N+t0/3MfH/gswcSX3rUeyLIWoVzW66IyXKirPNLrjCToVp7Bmdywudyp7k0rzSh/P
tuCLFgLmN611YVq3CSQXZuNgCKvnfgJDujv3i2cLisRP8X+woav3mZRBQeCgvJcZD4aErNVcwlsb
phT2Wr8nV3Jp57DH95FlivCRixpBy8vA7Kg6HTYFj21mvM9nBW5gdDB25aSHrka4Cg6fn54u/eON
hCQLoQpWa2RfchI9PLDxz4+6i7FTSg8D6lfRiTYwOire2Gaz4f4x5QclQnURDCLa1KRTEDxmbqsA
MitjWTvTMBNt2wknfgucBCz4zjinR6+Khxrq2szGloEjN6fgcCBNqchyIpZDTwnmT5NVXfEPgPl7
3M7gd3DtYyIORjghdIiHm4WBodwB6lM1xQZxQn8vjC8C6wOG5nzlfTdXaUd9iz3gZ5UWs69hISqq
ZO2tu+gVEUB/lpjib2x7tJCs8CW22XUs6UP+lHIyxThxb//DCt1ho49/WgW1/ERh0Rooctil2Us3
fYHf1patV/QJosDTIP7tISCjU8XMk6FQMV94G+CcPWuEcr8vQhxVueO/hiTKutbj1DlCZ81UAbCJ
9GmqA53Lc8HTXM+3z9UtscsPRBcBSq71Qj/0YEVfWRdAV8pRLqAk5KupfDKJuZzgzdcb5iWO5eiP
BJnoLC5DpqLzwjOgj/8wL8vCFMO//YC9V/VTpqGXFJDtb4qwUb+XBYqkCdJDO7LnP5IF9iPm1RhD
xyt+N9F5qH5oyfiO6QHnc94jZEiIMM5kZaz9vvz5zU/pxmBvXpYtHMMcR6gSjKrlL1Fy9VDRx7RG
PvJT/6phC7dJtkV03+cL1efvtnxkuFYXGxhor1nZD9dChCdtENe2BO+qQeRnElQduCRhWbngLEl8
W6Qp+DY/iGUOcDUtMoFQXbc1e+HtJVKxVkTQzVe6bdYgIwnXCBoyFaJAFgTWZz0yaOyptaS8Y0Or
dmfYaVHFGii2F7NXcTW+hIKMuAMBYgGNvo5Rts3D5jW4CQVGdcjqdUlSdN673vzugZoa0GqYNhKY
XMrUe1BZuR8YnYIjj+/DFD7jL/hSlDANimuY5tKN73ZnOBXR2OSgHTyRq/JlIU/STr5Xp8rS9eAk
pt4yqS1Qd5zCz2mtw2drWiE12P+aJe43uSBln95qHwXHG+wKZY0gINBv1xYCq29kIYYuqWVq5o+z
deMLsiZXgU1D48QHbH5ghcS7Ip9rRMbvnmX8+/v6UePMPgdqcqstDAd1zU5/gioSCjyxHD52FYvf
SdZvjniFeCTP20ph1LrCmZB3JJb/jxyKhqp0/mLVtJorPuWUS3ogVF/LT8Kl8ilnDW6cvCxqhPzo
zwj0MR8NtBZtqN7dA3TYGcgrA0L7R7fRk3HdB+ff1ETlPub/LWXuQ+tm9LK1SAc6Z6Ppf4vBGaMy
lZBS8lb1HnIAnbvgkOysoi6ynrcUGuvMG9buX/OjzY6FfbfE5A+lXRsD8xDzhPSlhNk+mAwJefUr
Hh96L1G73dBlrC3+XSXHvrbre77TFHbigwc9QwTm31ToFFY3b+qwVjOB3k8Fb7dpshScc+CyOvHe
QGsSaySCkze4WUyTvmypsSBJWIknckna7ZtQE6YbXg5J+BzgPv+5olw/w09SeYAIwvPKIAYAvnfT
2zKOFLfL73WHiKSpSMda0xx6GglMEAlAk0iwtK5SCRBnzJtz/ZSn6VE6R517COEwil4gC5PfPqqf
6jC+ViTQoWvHX4AKYT2J0IFyTvaeGchYoeKWzLqMrmRGrncpIFvY3b89VNGXSs0x7nljBKKsej2w
SImXphkT84Ru7+ODhHZ47jfia+YhRNGdo7r29qg9g4DQo50oSaS3Pb771wPZkX2qHiqUcRvFMCFH
O/qPLPe6C+qBxZjEaFKhEyXiRXSOGW+UTRyadXCzXSRUdpQrtFWR6jF3nDKIgWrASDrW7G6NPhip
qzw3vK9H/hOyJTBXOkpPArf5Gg2aWVmG5qJf0mS9lJd0vbv9pc30mqF5sXLsiY/7gylNr4ou2o0b
2WcsN16FGiRPalIK4OdCLScVcjiNU2Q2CRf2a0gTRboJ+w2a9fkZBSEOxdCwGPMZpvig0uH7sJbp
oh1rQeHgjhzI2ghheZNhsSvPbVYhcqBEpWK2X+P23FAhuVtFUP29qM/0bBOEb8fFvRtfDyYu6cMf
2LsCou25Xvnshe1WCL8w7aTjgUyTzJi0lfQ58MgGJ7/1FFL7Zs1SIGMdWJZkZEtDTCZWGQmctR0m
ZFfz6RTc+JGYPliCkmh8CK15Zboi6wF6uU2MWi59/H0dP/bKnYHfztCF7riTxeGZcnrMeLG58fpo
PBJLyimeUs4zlWuF3zes94wQguN36CBqHqEJ8SHBdtJ14aVS3Twt0WX/tPGZ0M503qfAT948xb4p
Jd0kia4btv7TFtWE5kWwj9kt0C0jFLkXnNuMAln9zdG5vwo3IejJ9hL6sRr/JG9YepJl9Y6cH6y3
jV4fnVMYFmfDluLgk5RPu7twhiA5TTwBy3jOI+vzqqxY5603wVbJxJIdXPupKBv195CHaf/Rd5sS
ByZVrKzrV0aVtYcEAo5uIFIpA9uEMk+IgVvMd62WWsgc8oLpxYhoSm4C6cLN4EXN1AeAJPa3rEIK
sPSA9o1BUd8Hiu96hiEh7yPWsyW9bMT7wFuQkeiBVuBefefSjWleYa4g4cHYWEFbG9Skh9cZUwLA
uTA/4aofK9jpYqvL1hYUjGMHtzZCeBaURjUh3C+5rIPWlrkmUGN46vmaq9oqLwp45+r6ddjwLSIh
/tsQzPnWQsSXlA5mUSuTrUNdOK+b/hbSEiR63uaeLBMXdNbvjPbwbjq5EV0KwZ4hUG8wXEYFax4p
pIGdbbfUKI6m2mhlbHGPA23HupkJfzbcI3lANOMmoITXDEPS8kfcOcer7f2u03mgW2OpE4Rad0gz
Wuwuhv+FX7jCP4NT0/SC7ipuEgo4UMu2jJ3YXV6foR4AXYC60CLH6Vw0IyOQqQfwK1K7q9S672/Y
5AUMUCjw51i+o/VHOH4HXve4+wCAW3T7dEGMSjDPKKj4DV0QXowz55gKHilXTpHt4RAPJZOAH8Tr
9JbZdSidFOqXgedO+dEhnFc2xugPLHz60gLw6v300XfcskhgesJk2AmS8oTs5gC/j6IWKnek2VtR
QIlnLlOsEEFAGX2wDHMz4NN9glm0asAiej71nh/lZMXue7IH4DZZtXjxZU+rV0z6OTK2Ua2wqNFQ
JSOdMKFuMHOtO86WaOcqeO3S5Rd4R7iPUr5tsU/JKbuoDZj8crhjeSqz5UE7Pl/gfMZ4PP2PFRmJ
GEsGNm9LSfpM0W+yUeko0CP0lIIIK5XS5+/AEpTrc8FJrI7ZpZQB2othcM+iQ1z8JFRlBvZhNGzT
JgVe/ad8Gzdh9/eeFYKrn57wr4YCF+++rEUoAOyKKFjk4vxIHkPMWVcAnvmHrN3cfKzEgUS1XFXI
+5I8hlfjwAZkUhgItUZ9ueJCnGjUORHETm2VclrEAbI7N2fGDksqhNi3GWGeMvjubJnliShQYxN6
2aQmn7whL9aD0h3a7Hc/Hzt0gzoEiYeyhYMJPDndrZCF/1UDDqq3GYcUIJeZhZOCB3GaoBkC2UWw
65KntEBjK8JqV/gegIyu2tuQIGvTwj+NMikAE3A71TeVufWlDbcNm2iNYKFz++iepivue4MZ80rV
a6vWgQpyMyTSLFu3DC/TZzXTJCTBY6SgYNqafhLm3bl6Slx/oJQA9YX8cXZMRUUjSNnFgEQ/xPxc
7tM351cw4f+CNxfic6/DQYhm93cklMo+LFvgdh+xAFNRS8Ttpz6PSyZ6hJEPtvOYMiOR+x1G9dRF
c4ODgjNfHR8ipZE8ZeARCXDLbe+0jecnE4jUiLiQOSJO07+VWlzxsKUE7DwOOsNTJvt65Hy36Nrh
Tk7m6HLjy/tfuEvfODsBPyezNb/hpafbFvlwifIx7OxjZDTQHcQwEIA/9Ln6v43DjkiSpFSHs7OD
Db/zrela2OjwnCb512X1z/ikLFOqkLEndUTfTbnWyLTKkT8u2Alk0oM8IhkdT3bY03KGCNAaMLgE
wHCevis4PZ+4avz1q4CwWnlfGnWf59iIaBXkImSbw3TcPFE59UcOlWCYv8v/9l+LDLwHQSsK+Vj6
VKRk86evDjsq7nIeQSB61tlO0bMC7wudhKCz/SwoXGDCs6/6xzOy17xlj2mydO7/gUlgdA/GmUpf
gOICFfyJzCJE2bR2KYWQGUqSfBh3xxGN1MmK04j0Diz5k/m83CHLpTfHsZa2uhE/5L3YsKFsjI3l
2SXhaqnrgYgtkKkZQTCMmxLylDtxYTkOz5CCOzC8z0pt+degk2AGlsPCq4EvDe4xdEvNKf6SwHhl
jw7vcekug98bNrF2ZDSAma4HQA88zCCX4G13YzLN4pfyfd4gbcPglluUeEM2HZ03WvlT66s8uTYQ
gg5lOoDOrWzexc/6KuUHwRAupb03Vusmo3oSebYnAgdtMv8okDcBMtDCS9wReBdV2M4Zh2xZnjXq
JgGDCeHcoUN+4kHTcwocxSTZTrVSp0BMHisoZyuE7YFvXaPKTau4qcLMmLPTii0wx6/70hBlfiVg
JczD+sSMgFuUkqZH0jjDuJ5PnrX04qicDkS0E4JsDdPkRjAOfLYQRMs0GDY/CL8Ei8IQCzETfIen
kL2jCfF1Du8wcnqpILOy8z6EyWsSwr7nIs1chr19pIAwVFnmS3gTqSToyQNy4EBlKwNtPUWD9S9y
GcjWZcVdD3efsJ0Jd+gTU6wptDdaprFL8vukAZmT8myEQVWyFUS7WHRNsQtl4RFcd6xXC+4wp1FW
m4jxRTAKooeAySkDSH5liYykQfHX4I2fDGZJWYQtVCyAfN2ifAiiAfEYYlaGX/FgrV/1Isjrz2C1
qpsb8rEgop1+uZN54TbUssIi5/gnibjIUYXRV7XSTs97RFx4HyAbCYvUDS1nuwiiN+Dpif+VpVZc
HvHpoO8pp29jkYykdj1Tw/JWWY1RPHYLqz9Em+sZLRLdlLXBESOjYN+ky+KIiO71LksTN2xC7SVF
8diItA839MW654noPQNWD4uTOdKEu7TKNcbyXGhY16Lw44WbyGVeTNGlJF/WgQIZkY/nNrPnS+9R
f8TFFWWTyAFdY+C42EhA0sLsDJ2w0xH+YoIu/G3cZJSqapThA9IGBl+tkpzUgG+o+1NklfM7TcpS
lPc+t3sQx97nFWZNqLD+WB1/coBAbIHfWXT0TB9t0WXOZgRjIUaLyUMVRk6ktg/I84x0mWQwv0xM
1QCLEsRxYgMdKfdKu49NnNcApPzjlwMp5FHaoCeCyOLsN/RjNek+moDQEUKhHPBAFNhkw6Jdlioj
dMdOLi9dwjHpEBAe71ZhnoF3PwEINpgOqmqEKyGsMj3tvw/pLmBum1aywZa6qG9Y6hLPooyW7Byw
pCaucC9nfolGO6FsAbObyX+A4zsJJ6OcDvak34S15fr5+9/HkN6sUUZUhpXxOudjpNHdUUL06ZPn
OXbHqzL0rEbM/Cxkn2HtLP2zM03Rs69rxQfB82YOmkSYHIa4hN7wgvMHZNtfsAJSFcTVW5JwatMY
z6oG6d5CU16Ff9xoGcZ369qVo4GWVnOUGygAr8sNQao6UlTCCP0+DBGajutFPLKqPFT/4FPQEQ6/
2B1IXjoO2tEw938B0ZItSIXkSbSpDhirxOOVdoHoj9B92KNAMvo9IWHfMF++QV4wN56hYwG06g41
3hgh1xp73yA5GadGQy5WrfJO9Hp2b1+z0WFK65TE9RoS8Gd1zDVkziFWipdL56vmrNOMgVvKuDJG
jo+eAJ/LEk5RtbN58CSzpegfrsRdcSupzAhUR9yazAoud+jBLKK5Cj/y1OcjTqdgWIw2xxLs8AeY
I0SlD+/O9qVTUT98XIVR5F7bsHJDIqFChoHzPk8Xvp5YRdYnBoDPnuUxA86HKUtrdZSNlyKLlAdr
08IX5YnLpWTb5hPv/pIgrsurs5Sl8RknEKTcQO8fUjyzupbMFOj1Bm1j3/4j28un49kjFdecEvFk
mIufKifk1ruQ4M6HJTYzy/o3CCvKnKIIa/EDPU+UJe05jlAPWuNTpOvIRgdcrZbGquCvdk7AEfuw
mqp8MKGvq0zgkorlVQdnSJPOS5N27d0iDW3lsb33Rtw9LYcENTQABRyqwVWEjxp2lcIp3+coA7e6
Kt8u0g4JCIzYk2xPubiKDgcWCEgbzc256VR8PkbSIQpO4e6jfVbaDqCgiT82dzuJowwPnHNNpM7s
0LkC86tkJ+Xwz4NnF+OdvzTyyGqCcEDZGT7sihw8hZAqyy7y4VbHqQoqIS5uuqGHCh6NwX5htPDf
qjVg/E7+OeGZ4SaWhZEpPXqsE2Phknc37GXlIwETvHchB2n0BTvnuKQKey8UjVpAI3JhCL5eN26W
1PdH1rpxMcGd0JbpgRYBUDbP5Iy1HvmX5eosWwUSDgxDOKxZUOxgw/z9ockLVdo4GK2Iyv2/51pz
4ii1If972t+zcv29Cnr7gVHb98/2I8fEjip7H5Q7CsPVALfKZw5O2tJK1xsn1ZDg/PjpLOGliZyu
Krs9ayE8/KZ6V5TcGXOg3InQjbGGHsVHCW0GlzH/lngKRhzMSKp9BYMxykuLMEfOP/ntZasIy2d6
Yte60TTxnWTvVbsJQli3Uy+mVFKy87nheHP7XyXwt8kv6yVkX6Gw8U7/ozOufMyDHDQr7NEY2THe
m1RKI6zoHlkR06B0pOEGQdcMAmsZvaTCDmNrnLMRlqwVvEv1f9aJkTXIHpz/rjauBfwOkkC+MDhy
2B948pfjvp5Bvf4CI+syIefM4XEuB9MyG8eKedUiyjtaOw5tZnO4QuK1KwGRuluyLt5A2iSckElp
0oWSZIaYxmXUYBBBcrRD90g7x897jvIPf5KCUllQlaY64XsMWOlujTd4UdOIbKVrthCYF7yYelF8
NvZs4wR7GKUvZJKn5687tft83IPAcGLDLUKvKPbWgwFPztERuVI5qxC5D1Ypsa6ygAPYTUJimcgT
dwbnyajq5Y9ppptM6w+veo3SDFbBH1RFl/MRF0LArwAWzzWf6U+O1GSkAuO1ZMDS8nN+coHyQh4O
FBGzVnEhJ/x94yN+UMK8Ud3tJYxqQS5fdoyqZUtGXueMiO6tj65+kXJWqBugAe8m3qqBh1tqluIe
n47ZjWQbfldo66u9IWsWzrxzPM+IU9SZMPjf5s7R4OGs5f5VNA5YfkwIlVtQYu9+THrxNnnBR+Ks
AR1dl5TAQ2+NqAhBcv+hHq6aMp1zrFG+jukb1R5nSgjANuuXfRVCUqClkXZDbMomkH1vpaMrt1Ds
NoIXStpaAUT09cdq0AyFn482AJ91iABB8q7uf2pgYAvI7VlioWP9lz9xwGIWQiDc1sQsraN1duTm
rR+HLUJZGYuVHDVVxWNArLSn3tHommcb1dbqrwzhN/KG9hqnxRQjvPF1q2oYzMdTvivzapY1f2xF
4MZKNcjObQC2lH4ssYwYQZiYiwOZMVR+/FfX6lkw0jZRhuNI4hXHW798MrDfpRMv+x2WeoJfvoDd
P8AFWZCicN7YSXuxMHZ1q9pKX5p0FgNOdtdVPKr1DcSsiutgLDpM4tt+DCVoBOIJX276OImHEwrN
0i3U7JklDaWgfMqB11pLCAUtlgWlbPzadpEvlhliCpILZ2QlwASLsE+VAXh0YZVKzF8n0Cej+MQI
V/VJpQtYZZrdmIjV5PTQ/yM+xVrX5XVNClDeXIf/lhMsJQ3w7bqddrUItlv4dqiencW3IOdUuqiB
5jV9W3MTwop3rv9ku3XSjfJYZn+RZwArR2QMpxE6LYvoribJJmtnwtXKL+jQY4OWxfcFCrfW/de1
MWaBUHLvskjJ9k6C6hQzUYqtzGt9z7FsZt5ln6sNun9sKT2Aj0IFJjiRXlJtRR8BlaJpylCm0bOh
KMlXZEipgxcB7Ve8PfHSW/kxlD0PcCzKJFSa4Fomb0BB0Ovy1Q1OwpdBUqmaCSjMFs1tu4HRpaYO
QwW9Gq12aC0QpNMCyEPbIwHS3hLPdtK7XciYbCyxM8HtqVqk79zaV3nEgHrbec5kECJFeSS1OFUT
EROlHTIcAwKulFTpQqIWIJ+pNhuns1fMhExQcQhdE6V5Js2MQSTsuee0oWYx9El4J9xNM3MEsEZ1
eUzD5OA5Kd4q558fq1W5gSA4rEKtJ4Oi+D7Qa0RQMn4ARTIO5As0+ovkMeLlOTJQTTWZviqQR0kh
1ChWRN8g18q29aBY8RBv4QCS9XC2SMTZyEKQo/Poo1xtEODubwTFBaGRT/o3oiXk1rapAmKLESWl
KSAvkM+z6EH0Pv+pxKYqd7p9JTwB2ji/NTSeL4QMJ8MPDo55HF9YOvLCh/a4dM8lh4I88vHCZUK3
5qoicOrdiNxm51sthtl/nKI92xmNtEGaUPmyxZXuxiSVPuVVX3L7eSOABlM8V03BLP8umlId7I8b
hAzAL0t4Qg+ZQgJ8aUQmckMDwGJw/N1S9RNsMhi2ME2DeaZxRwMWDNOBfr+kRAqw1fjOByrLg4k+
1D6SNHKQ9Fw5Ux4tHQAS66FZ2yzrzFAulTr07WWorgOIA2Onyci13fXF1mycfgFRm86t0jRWgCwM
9V6wkY/y8PZUENHzOqwFCYlCG16Q+50nuIB6HFOOCFuELEDSiuClNdfu4YnH7iAWVJLiMeFVF6RA
QRweE3gnXwN86dz2/NvMKRjgq+MjQr3C1tHZH1nsXcwsKZGXYt9plxAexmsZs0jeKvTwcaub3Sxs
LWs8kv6pM5e3SOf8mqBtgrITMcwmRGeYvn5hxesKhLqdc8nDBgevMAubgBte1CEJqlMDeywWKFYH
HU6fxppLcMnCNn5TONUw2GhbL1SUVLVdqZ6QQ9xNVCeEQzVYDovr0IrbNZG/YG9WLUlL3BEJSVa5
Uh1YDOFSnLIBXT+A6lCteLCfzjaRSBmgBYcGtasrfNNbgVq5ihb2SS5c38mRARodjOnP91RzVdo/
qBjsIoosE+NmAOGRLVpOlEVL5xeaC1C2IqZ45+Tqk5+pZmd8Mt3YlQtmZumy2ylgoV8DBLOojHiW
DkD5EhwQyTae5qBYDE7JQDz6qcBF32yyug4Td+W/v+YGbFw8qkTCKW+6juV7SXKEn9C9Z2VjndJk
75b6f0c+TaQWfAoyaZKzDNMf+ZYTHKZaHSzlGB92R3qNRXytWU0fQ3sSqEHPzCVkkbY7y32By1KA
dyZyNYtdmX/iug0q6r+717gdVPNuWZVWBU6BcIG52+HzjS27U637e4M0kwcj+r/3mYGbMVM5RrBp
mEDo/HoERCVpDkncfy7J8IaZ4lr5Cv6PlCH2n9zijE//DlquhYuzFwb9TComSYexxAElqyjGOx+Q
LHrYJsXOgFDXMoT3PSxJaCW+N4cYhvw3cKZQJfdU7aE4o5KUVHS1By/i8CZ3ZqR/fvB8iKwmWTc5
SezMVlWJNnwF7vVdUCoKL+ORvuDfdNzebZUo5NjGadIa/lnvJPncvc4ZfjQrShlElTTIS49GO4ro
38vN/tEJXpxJ4UQ/vYgR68dVQocwsvUP7aFEwppyw7e+BXHkdKKOM3Q5JJMLx++P3IAalm0bfls3
Z1ZLvHRjacEzcQfwZEMzZQpjUnhYpY4jc36E+e127QaZVuIJJbu1/logFT+WZVpabCvVOTCsTo/3
f1fwOsa4ohvNprOJmxa4pY3LevGvpYUb/8oocT3z4vkZW/69josqSnJd7Go9GdMeXOP1wzy0hggC
o4dOanKXyijbggiMhYOXzJo4+4leHsocWuKM56HNTB9iW6x9WeF62sCeUsdMZYnoZVhegQwNcxNq
fRb6QRpcfX70KDQKDZWVMXuzK07ysMi3Qy9WKh1TG95xaOnojRVIl9aL5F5ki2GV94xVYl8uG6U6
/BPkz0liDwuhsRc6+yyL2el5SM/+DgAVVvTo1reuoHYCKgB0QN0X9g5ocqyjuNOalnz8HzCDMZ43
Pq/5Jc5vSpxtbOKahgwSlRqTgMqJeV2vu1SL+piaPzWiaUljzzqYJOuGq5QuicMWEgxPaCj5EnQ3
+oqGF4N8Qb7QzDgCeeRlRniQLloowHfDM25sP7Net+azLCbMBbtLH38tYdzSH7L+6B6tPHnYTsUH
8E2OxduQnmlyQqeOf6EsdvJd18ikFAagjisM+RD2OU4vPHnGXuWFdAGonK6mKNGFl9hjr/dI8Xrx
b6ECxVA8QyTwThGGGyc/GnWB3YEv8+XouN1mYp3P1NXqkC6wAsviXc7MkBBEmiETlUHvlMUG4+vn
Y5h9+0k9BEb6mzsmfsC/2bkohkV6eP7RNYn77ndIGBpAAAN8CFHO9kdlagWPLe5c2MGjdgXwxUk1
Gzb6QZCWPTxog08vKthRv2SdGshJVscQGZAjpCMI85tcjoTdRYiPt57s1u3bPnAm83X4P8PwyxVN
8t3yDm/1tBX7N39QYhRPihMypqO0/45xp7mjB51w0HjYFAOLdt61yOEiEGQT6F5L9SCHv/P4KVLL
BqRhno/0er6fi4oK3lBIPgqvxlDc2iO6Z4Vdb8fy4KEOYC0cDGQ+GQzD9yRuUUljRfcDXyUB31bT
cEYVUt6GO9T89/QjX3JmcP91GPb8FjQk0p3sL/6unQkkzyEu4Bsjo/67q+VEmSZrGy7Ah7TrwDhL
9hTrmgK4c/JGq76+S4GBwmvjfQJ6AA4p0WYU0CDDGntM990Cr4opJO3uUBtDjZshJIs3oMIS4pPw
af1JxGeTXf94kYkKr9vl9OKs3FLSBkr3w20jUQDlJC3tsnM5AJU2dQPGKBp6idgjkIx21v3iljXe
RbRBs/DeNCRZ9aE31304l0US4Ii72GxiNwGcK2Qrt3XP3bqzRW2e0UOoDwTaR7ZgWJblsHMtDhNT
QJH/xwH/mUr4k0RdjOidS/zjHTD/qIdOyPFs+p3SE2m6jl9y0LhW3zd6SqHjoKrK/bAAe+tnzI0Q
dPl1NiF7ek+P1C8eaz4ZAvUDuBLqMlQdUGxwbiY8gXnC2opcmYcXAYtRrkTquPKClmThQDAdv79A
a8V5yi4Jb01aEPOFJA4og+zDr0QSQPDUvn4dISb1vwXMNkVJVx+lgUVmQeVMUkjqNZAmAnYCdWIz
GtgkARktVhf4oc3jxd3OiT4d8OvY0bV4h5GKbWT0pfPpq+I4TUpzDNFNtEK3iqMUctxpRCm/oXw3
LRblA2Eb5jo5cngJ5NdBpv+7mxYIji9Vl3fogjabWWcNCy4vd7Qg+NNmKcjO27MhrScct4HJwa8K
cnwKjUDdvzS25pGOoKpPE2xO+cHdjdxw6yQzbndbZ7f1OOJO43mdtaNhqgeBPTcmr3sqXYS+PIuQ
fa70SCfaQNXoiqcyzLfY9l5Csxifd3wJZSQLRd9y/vKK/ZvZ1t5PnIePKUtgTW89o5U/89B5KijO
7yINEKir/wv5GBFaYnsmBfoM7BBLspJN2Trs7ZNNpEuicoJntsS+fOJD+U3u8EqA3A7nqS9EPmqO
/0h0ZaFpvxMZXq51zaQTsBZXqObSAHlwdcYtGG1rtmIxyu9fNaVgO41yMPpMrs+JOriB0qNvp54U
urKlK3PZoT5kwG/k3OkSwfv8zLVfS7GbV6Ts97MrMARuvgK2kRrVTZ1s2DaP48Ep9gkwTKmRK5rg
Z4BwjeKuNIEOVydXJOlVxPOOM57OA8FP9EYMl4vr/OSDxSXO20bDcI2I23ObwiTWDYp4iZ/hTUEj
n18BkzVMWCv3HWVfGHHogxFlN26endqtTKbxHp8Blvx2Nfr1TXwVXAL0egvASr6Y6ZXU6zjai8O1
lN3/Z4ocDt9fiZ7e6hiYzSO0WvIsP8rxiEeTlP48hEwtxNYYiG1EQ/bhjPAGzgxFDbucK2E9bcW/
KgPw8ZLOii20V4tXSg7RNIjysdtw9EuxgCUwVtWG/iYH8SeH42A3hMqUGsx9Gh2ZIw27gkkOrFPO
9Bnf/JT+qmao5YnLMNhmVs/LDU0XcVgPzrfUcSjQoD3IKMlu7leJQfnDY6XLclgmgtwX5tyZ2H0L
ZrPh2obUlNYfBuivQKOsup0WBmWoh4VVSL8LXZ+UnygT86eY7NkJguUaiST0uqXL3Sx5ECnsFfES
ZUh9YzxgBnf02gFLRHik0WLyWNx4tKouygXKDhEi/CI4o1rhQnMyoWtJA76QORmcMLd2bejqi1uV
LMo7xPxlj6aCCaUIJSCq+xxlDVMMii2GAbXaxJtKGVBeUZ25eiorPxmtZfYf19FgxAPoB3czDm6E
Vy463rMJOtRjnwNOGrCI41sBuGTl/Q5xo8IJr3pNBMnisAeCciDL1eZdJT2sxcsYk7kQboAdZ/q8
sOp6W3ziX/VUlTKpp4M9wHJjUuH6EavHrx9g6a7omwr3PXQCPF6pabdgnV98VcJbZ6VJ0EINnsJN
F7KTTElaG+HHZj0joOgxv4AGSyr8mnNlYsUVBsrWRSsQTa6v3ak190pKgUJxvglSHfYmeuuTRhpG
WgzuLZOBEqUjfwmjZBSGPHbVT0BFZqSWEHkAV57F442r56kghP28tgnfjJS1Up2tpc8Ff/734LOs
Gya0DQ+30jGTaLfy1JysFTsU96bL88X9SqzeZJGag+FquaagJe3RlgbThqAgrDt5vJV37AeG8qI4
NDTAj0pDU7QP/y3FzWfbITUCMX3VQ5PMmQoZEuTqaCoI+7KmrsWztjmhAWu7/WnKkKYMD4MBCYIA
6aIgT+u49iFFGcoQwjsvmKAZtbCIQIBs3yEAGYx37z26kbAlDCVU4ie7acHYYQVH0VEOfvyLxr22
emMaBD8tx/dY+VQewHVXQYKd6T7HjAqFkkUsiTht44HgwITVgKgVi7CLXPu3Rb1wc/G6uy0wNEbI
p6aq4XlXFZ9y9GOoX89KvPkPDyutrhnQ0k3sHagaXLIrH0Hq+0AUcbUmuNrdiARVka7Rh6jpFJrt
hqXaisg93QdYLcvaPiUdvEGIuQdR6D6vYDCPwizZtxRGsGnkhdCRnY9PVwNxFApmL0wG9j8yTUMM
vYO+lwOTKqhp/uAzobRiI9cNPdYn9T/gkJ2UqYQSEStDyd6x30C2H4fC/XL6CEM6eDwYoIRdAy82
N6KX3yP3lLYddi4gMYqPnvP/s7waj7wjWccCUI5nyCM/YdbUHPOkrSQstzzTlgGhRLP7Sqh6AsLk
rU1K+MgQAuiSrw7EbUm/KhscYhV9dq5M1iSyysOX89zu+ZjhREWLdILLJs1yGutsE1MczrxIvUmf
ow/+TPuy15mvG+KqUP2PQQeQIUYTnuaoBxVuDiMn8L+9xYeqZtgxgbmHFL4Hi9VmCs9usXj5BmHY
ooq6gsFI8yvk5kpF3oQ0+DuilKmpV3iLBf7w89/e7lp2DJgdyPbNutw9VGrmKgnNyhw/jyVY+2cY
8VxAu6VmDfBQfb7uk0lYgNRmlTOeVbBCoyloX7/zecNJGjBQXe2PgsHjfWMTBkZ7iEQFMefQkKhC
9r//SOyQdF70qG+AN6FBw2PalmlSKsDR8vqx0Xqf5/20fCVvYjd00kWH1DuWFj5VreQ77CCc/kj3
kghCF0f2T2XJ64wb0nKojzD3m0Ye3vda57e/6wPDEyDjF+Vopc+vC7QQJ6ICuHijvUKYGMsYQ+nu
kMQd+x8Lv6h0j4EP6gj2tcFZfKdeikViAuT+77C2Nv5QHlbPz0xvEtDiTtKfo4coLQj8+F0NDPNo
+HfBIfEOqFADD17oPfN6gldyjNQJo1vqrPBmA8S0ybUIWAps2xGQ9ecAizCDZsgTKNl80Y973P+d
4g3kNbB7EjkAlwR3Km5T+eCh9hVFy517+19MYlwTZ6pT8r6ocZK19KmGh50dl/ri+qqpK708Hotw
X6NPJw3cKoGBVyqJAk422WnoJctP41ZHh7EJIAmYAkBSMtG1rWdVACsLRqXXWAww1U6SRfXz4uz+
wDcmmF/z/c29EX16b6Qp6VTkMEGJsECgutiGi9iNlB7IjrwSC2wSLXainxL0betaZBQKyXz4ausl
7rYdWlxa0t7zeJ9Az2ON6D8oiysykerJO/GpOXRRAb7TPf8HysMrNCBsSDY66wMkPEURu4vZtsXq
hbGRYJkpEf4KF3iP4CIzS6fi5YygGQajhfKvvQ0oZlX03TbFBGRQrE+Pp4j33uyjs8nmhXmK1qdo
mUv3vIvzwAouc95ImcgCO5a+sKFEfWETqB+gomMB90//GMXOojyGPQ4YI/t0mW6t5lqVUXLKO2Hb
TOcv2k1rZEvzuBVugHJzVKqqSLXRrxBkoyVi/MltFEShPuo/re9iOdw0Kr+h53hysGrP5fylN2Eh
CBTEXmHNF3FAnDMteTnRVL4/hKFJLCY9G7wxN9JRO0pGw1vrSBkKuY4myx1LCuVm8Je0n3Ftsuw0
tW/b25vEyjqR5eReBS+5g50UeUz4dooWMokoa2OuCUSS+svzehXLhk664CsQNBzKMdljrqHPeEdM
kMnEFibvIIfUCxMOY+yYYTAPHqoaqpHw6IPB5QEkxOqocs3OE2qb5fCsa85nh7ojl0V10M7wyurD
5IaarXR9M9RnZIKWjoF0bBqB1IdsSQtF6sg2T3DSdTn1sb/W00lffGnULHe2cZyKeU6D01JfeJbK
He8xkOn1X/v+VuT80+IB8bDPwvq4WCYvasMQBATEiHtKPKeUzlEoeOf/AmpEKpbYFK7Cw09l62Jl
FicPfVlNRsVkB+2xefuiRt5VXLWTbXO4W92SNGRIWeeDJ7BiNIxkk4LenlfJpfr5eB0Y74ZRnXt5
EgmFBPwSgiD95mCAGGGGFw6J9bWw8v+pZTIwbG0rKb5mpBS28C2yTmS6i3ppOBMr2xqLfijNrybr
8Z7FPvt49zTvdTzYd8Md67OMJOfUwbi0Xf7QW+saB93YxQjJcS8TcO3sJmhVHEyCyw80TwU9SahO
rqVd3hkZd8p2HwxOJfocq9qC6msdJUCvnaFLGdTQWrX/pEutao2TBNg3D1CB/jq+J84tD1rBZx2G
iLT7lqSMV8Qt7cHDWUXeYawv2FP7UzFXT39MTAP4eca36K06NaS+jC5ZH2DFRVRy+i1I4EbBy65g
4BylUssiAZb/vqOR+ID8uz10MGf600BEbNca4UpltScyQ60dNN8+bK4XZcauMGiJHkz4SoBdMwuL
/kaHVdMXEyvhfE3ljwK6K4V2DDDG22tltwiZxpIwKIeTNtyQC1oCcRvXu3hLUGGeF/M1D9Ofkbxe
DTYUUvhn0+e3UP33ZxfQM4yzOrPwO01qk8HH5Ko3sZ7iO0GGDuwWhtrOP8beWwtN4Bsnnq3ytUk6
rZ8xPf/UsqCF3raekzhfkEcxkkI/dkt68ZTNqcA1nhe9i+gP8jn1+UTfyxiLirAAlF7G9vFY3GUE
+2/iiNbelhL8ZdnSDed+Wb0ylVN1kQWrurLJQlSmxFRhI0eVjJKXz6/4yItvguTOSLcYJ0Ho+afl
XKgwuWGAlsSOubZgdk5f+9YgXG2VE2g7eGmZxsZaFvrbOvY4/KiSgES4UiJ653h62cXwpb3eEEhS
ixdS4muCLQrVmMxWGXU9DMsePd7Q1DbrzwrwjLihL6bMW21F5f7rGDFYuTvfRMC3txA9WU2gdniN
gY3ZC4b9CFyt5BN9HT4lqTCkdDx8VRXgNs3JlQz+kLtlHF1L/wKqf6tsRYZy9dIRyKRf7AviSAfS
xSEvfDZdpp9ctNOdd2teryumyTDFTRqNK92yhgnBmXII4EUHyaglsQrz2E/aN3ZRxZ228qLN3O69
pb4rNig+b3lb4ulHVORFrhS+Koqc+/49DpAoxAdIS+GIDovNTcTrFGIynLNgQWx3s2ZDQ4/Uci0n
oz9P4tGN3a4azwZ8jBj7Oib+D2iXf3lwLUlV7E+cA1xQWcUNLBLo3d2V+MGGl3bvcmhxmo5zJm1f
MCvtgpix3cYK3CHd3TGwbcGgxuWlcJBjKrK9B6AQlvtGHYE5S70t1q3COWMS9Tfsgw0TkmE6XXYt
dQ8qDo/myfk7Yr3NGM0UL3txGZTKuVmfOCGEk8UQRaGn5pkzWfb7Ass1gg5Wn6ODqFB2IKzSdRDy
m9J752JX6NOp+t8dBaVG2f9CYPihIVAzgA5lrLrKw93xL+e8OVn+KZ8co/p6sAN71AKZcbG8WXbm
sFbRoBw2zERm8U9qPhQg4OZ30YFfIar1ZqUwuSfq4cCDuZtuy0x1svTnOMsSVbnH9YHn9QKfZi3N
evwSNnYyYXMEw02m8B+1w5B68eCYKmG5PmlIgFWkClpGOZ+YXqybSNUnnc9Du5am1Gp2sJPbmjyN
TBtOCSw0bUKQHuKPS7vTgcoRmLVs3F51i9e7lcI7h9uTiFhEYCutbXmQ8npxIs/04sTsh2u73NwP
xogHfEY8Lf6jMtCEzpVeegsXz/sggRFshBUO3FfkvthpRBOf1gVFwhIAyQ8RYKo8wlZ3zp+f/aqZ
rSZWZto6yHm8UkcD2snSUX8EaOl89q6kPOi5dQuD4b9hmK6PW5QqKeTk0USO0LAgRBqp6uoB5GeR
NDPFOYzVqsJ7lm33ogPFKeezi/eOK5IedkXxvLB5nuhto/CrJB2ECMHTcxDmS5DfDUIMIFAzyGXp
vv2Xj84ai458oACCR+CMg+JqZIv+FvU8HB48sTLH9KB0rfL5ZZvUb8fGegPaFAlWaxfPvhYdcamz
U3pqnr5Ya3Cgium97+4Px3f5oIbTHaqDSMj5YL5CM2F0HUsDPz6C2J8WRMuT/ZRry71caXJjl/29
ezF8ZVGVkX9OxLnWHM0DhiHRJSuNiMDsN345p0nJT3/gqssF6aAXEJVLP5nf9jw3rjrg6bgw3TJQ
O5Ec3h7aDvfHxZZocVCbrFU6Gbo3qlOCJBtnXfEOrQGTHcIxdG+t1urEPiz5lNLOiFocgghHPVbH
+FQhUam0LdkxWXuEcpWOjfLC9TnBYEWpHPCw8zT6Br77lfCJU5ZBtyrw5zyAtT9hXJY33ncZrwk6
JQBrfmrcXqsmemd97dZPji5vsQtAA8ySLDwrv997E8AHyCsJ0ORuqbDHuJXoHg43Sy02+KN0djrt
Rwpu2gDPIsRdPQOcHb43IzIBBFlLG0SJSl5prUHJmsJ/bp8XjrA8FI5M+MZa0oUDZy6X4f74VtDy
c29le6zfReijpNFTnsUOp7OsLb8mQRXaIgxIsKxhDDpNdx75E3LusapRuRsm/oXgcICgSHBTuwZw
m7N13Dwq36VneXjp5szl/S9k6vfPvurpfEs9lp0iuk5ErTwPSMCK27iPpSzD4rSD4rzFNsPcCw2v
yqEbSGiWSuQdkoMkn1ufYWZNl+eBNuXBwsOl3FKS9DTuNjwfDpBpFG/rW0/bzceXI1CjAE/LkSBV
yVvGwcyKr7bmCG689S9vJTU64no1+jemg8VC/8btFr3kZbaqN9OE62zw01kBs9C48V7N4NTcmaAq
NfBUBGOUwpIew/C/EdNbDUcBEpI4FT7jwy6OKWv7zSLXCQJMZcUchg3T1n9hLz8smHKBP6oH8oD6
J8uy0BSsjlt4t6W4FqrhNo+AH/3adnjOIpOI949kHBuzXQ0Oo+3iiK3vH+HN1dSAdtTVkjgyawB7
Rz8Q8L5sWdNJkR1ik7daEOMAaYFnwpqeVCMb4q256erNU1iLfbZIKahyJUXr5FTKC94zV3qMfTk8
e/w+V/UoVNyISp9OOW5goGX//+b6UcDW5cFcuW74OUoQXyF2ZzrqHZoRhdy519JZ7G7SBmLi9+JC
uwcd1WBWfB1YHEHUeqfJCQp+8isbAHEDhl75LElJE7MUrc4vMkTzjP5dejmJf5pn/A+lqakTljPb
IvAd+miJQ/X4PZ4JJ8KeknuOxsb8LJJrLojnqLs48n7cQTAe0MEPihVxltuOtUdCfB1FRsoXt/d/
AKPWKSbvLEACHeGOaV8V0WN0vc5WoT/zk3If4IElfnpTcoQ9nYwPO1H1ltw19spdAEVCKN+b+PJ6
yijAPmiszviLeOcENVNLlxAeI4Fo/U+IIZdwYJJZQNNlAuRGA/zdr8RuSY+oml/7y2aIUFvtgYsh
IeqZipx7IerLaF7xbjcL3NAKJWXQNvTuAVDOKwGKX/dZzLPUg27vWYsul+YkF0j7pW1mVe5yIspc
2xrBJptZJoW1NJgmKwgtU3JV6ffzXeLeP6lSLvvuFw3Dn04Du4DNT92xMENFGZvN3yaK+4Wo2bIg
c1MN45JSV+2jfgRHbrkVNZ8uXFWwUyElKZ6ZZa+qKF9hNcvn3PYY7llYyYqQt9Ws7/a8GkFx9LZ9
7bi/f5iWjeV4+nuR2hua//GOsRj4StN3nCIna5ksVUsBKGae/26HcJTZoMaHHypC3fbN89DWL5xg
0lJiz2h5KRlGdMkNOpqnZdGTxZKYEGdoP7Wo2sjtwEdaLPNgXgtHI6rEtF6XxppRrtspHz6HV09z
9b681eHzBeswQpdhXEhad8ZhPEpowbzwSgfC7+QBx4X53nwbPg71NDrjHF5wsde6HuSExHKcAyA3
oxGQcDHMs6bOpUCBf54n+5UdQeuOt5ZixsT0e9+5WxRFZh1+oUZjxkaxnNfftrUdl67T0bv7cPqp
qplepXcr2QHuEJcxPrT/hfnVi1/sO2zkpvp6OZ0DJGX2j9foQQhqq6y0oDadLh86SM1LAJHK9S+l
LPx5xQY1yAbUBpuBgVGvO7CCrebpHUefW08KnbYxKLqiMFoi5OGu+ecbBF2HCKNq69zrdbHj41+z
GEfn4yCWs5BXTI3Rj235YLWQswuUzyPwOG6y5Q70TqqgTBM+pSvVYg4K9kqlOmZdsxqAfgtSkJmF
PZl3ADy9O1JiAvCxYm4fl1h9TRJM0WCxBzeqnesfzmniE91UzoilM3QAHgP/I8H0drgVxGU3jJ4g
toz0lMtUOhNMTwX4LhZI3QpnWhmdp+lpU2PlZmcrmcF84SlS4hx+nila/sshRvcC/QMH28s/noD0
0Dg2a2oyUk7jXlwNXfaCsBicoT0hIn+NDvnsloPu79BY14ibqYrS76/zDBguOlTtrbt6rX+v20an
ucyQruhp1Dg/Y8UeGLDvtYB5FjSYR0LilDQQgHnPcFYGRoFhpJ6kh1KrVJS9itYr6fEn6+dGqotr
6CZ3BtzVgKLsoF94pmn+zBjGurCvR5SLz4zNtOdYGJj102NekNY1ic6ykKG0ZUGzkR//tbUKCF6z
PsLpsxJIwK0hcvRiLxilSocSmRqADmgSc6JIj9F11d7VPOgEc9BWMaKoE63/b4hzGt3wcu6+T1Cc
3wEzjuxlH1ilt1fzFcluW7yQxAiLoK5eKGBIs20iL3vU4NRQuAcFSLvfp0YqpVQCuw5LkDQaRUYB
fxDJJttuuAs19M2QuEmB1IxfVMTItFCj2u8Mr7KY+VC5hPbRrV2gtbj0qUdQL4vNnMl2FghGfWlR
AUUPteY21T8UcZie0vHXDFO5CBT2l7OrjEKhzLt9qhG5evxWty/6Z7ox+SIR0CWeoAbSiKOx+Z3N
diSs6ZrEnuBhxX65ygVzqbIRZGHF8QMbWoH1KRk4K1ddWuD6+TfHquVjsXAhF6oXiMTD2trbmrmy
KU26NdPujy455fGX8T2QSPKzolSjXJETQ2C+kw5kyJzDFcWM+vXSAwyZNkUfwL6ya/VDvhcxAq4f
XLaBZN9hpS6cmTtRywMtgfoK3W6awnRT4coz2Y16oepHldII4w5SGGACXS7pX7GRl26IS3q4kxO5
Hkm5f+01R7QEGiSUCo3PmQFjg8bAv7bGqqszkKAlzroDpQtzI0MqCr3IRFjFJmDcLRezFX0WTX7I
08/oKEVC0kQXiPEORVCGt30a8Bz8ODI/7l97wBwiYQWpVgvXyOgljwXoMPWkYSK56T1mvzKuS7SN
8wcD9gO3YN8gXBXhm678sZc4owNFvwOpSrBbb0vhW8qtrx+fjVtDMkeviN9qpeb3JUsbkpqqVsgb
SyQGaANY41rh3I3kUy0jqApuvnQqZkNp3WnjphV6RODy0PthU4d0vJX1CFd8EI4VQEMPgVEfIerm
sjZtMJwnrZcSRPaB6swXT9InbW2lbT4ienTXyaBM4hTm7vLEepNCJxQmW2LYTuJnpuaiokkelezV
xAaH+7bHln0tSI/lljnPdhjzV93LedQIeXOOpMQUgWH1WjXfxXHHL0ozygkX0T6vjVF05BJAZTdZ
iAY02Set1Cu5rOmBJNvNCBcygAZb0G6+2+YI/bgqG8seUqZHz/1kMqJ1T3yIEKUQ1TrXi4AFxBtU
vdIEsFJBqVJw+gp9xLT4vZDmwYdV38e2SEKavpoVguxGyhpiG1oh2hSN0t9Y3v2eBsJYP9PYdG/4
EFA3tG+AsMrC/tUd3toDmbUwPmQ6UdBrpc14hwg4NiK7nEp7zvA2vPjHA4Slh14LU/hLiFHP6MZr
OQtoEq0W7oIjxI62P+h3rff9o+RhyZ/r4pJIU2oRVWaMrUFga2gh4gLwuCVQpLdvutEgerpwu7ng
Wq9OTaVwZo1P3dSgLKnDFBp5r5h1aoVtt1e240sC4iR/r6I29DvolRiLVE5Hn0i4ykfwyIfp0Qia
xTRdsz55uz96+Xo04MiJZeicCCvMnlZxII3SWZXVU+ResAItt21jPLyo5r5Orvu20l25UrE3HNbN
hub3WMEohVjkAWVN9/jkpqRU3Yt8MPNpxWmstXJQcxJqlNl7NWxe/ZRGS/N1NmchfjsWn3CHaKgK
hDC1ownJAG4JLEoDaZ5Ujt5SgH3MucCjzfIPeP2XvNEe5FoBlJ5T9ltpO/nWCLozY/Qob+CXYXVW
Dv2Z7JKtDUA51y7SGRkGLCt3TeOshw9xI7JpkFH7SXAT6AuFjJCJSzWTX/GDve4V6xUrO4fRv929
Vm71TL0r38jXw35NfXRuhrvUmts15yqFZQ7kM9fUFkXY4Gra1AvetdMZhVmh74NkTXotiH4vf51M
cki/GBkJjYL+33w0/Ex+5F3kMRPKEnl+dqb9DdlCdQs7GU/iYONO1cyx5dYyIP1LLqHP0+HBa5f5
g5GL6K0JkPo8qBWGIJ6TY9EZcq+XgFbPtztRfv7NACieC8MljCfO7o70t6hx3hui+paC303zq++c
2pf2C2VJg4OpYrTfFQhAoZFysliYQdPBaLaSmiqeVjsxvajl1NHBJuD9yopHtFY7nej8FSbC4Yp2
gmhd4hBjhmZR32s3taD0MJu403AveIvCpNwwTjzaA3zmMfUVuyzhMyPuBAcNT8ayeBvvJ2MYVDdK
3+mL70dtx821s38YYQfBv2C2CpRJLsJ5JTJnpRuqxSxHo42uE46pgQUrnwFoWHVZa/LujG8oplUx
cN11DeXSo4JZNeFnZOL7USFZCMEosD1DLCf4AsI/nUdh4f/uLTxXx2JS/STim92mr+1ADlDpVL7s
gBCMuV2hxVq6cngl7cJqnUgWV/wqjTMngfuOkdyCRvOoiyTbm5D9c3uO2sHM7u80UGqxubm89dxl
TCo3Woe7LmEdnWSaBpQDRhDBqKdvNvYTyuiqcc1nj0BJ6rYvsNEtG9H6GJxzmGrBL+k2EuMRziTG
HKFM/N0QS3BRPo3CqAHgvsAu4JcISc6DW06A3adL7gjlV0wZAG/PluqnzJup61bU9PlsgyXc9WsT
vW/8zhTBURVukrLrNm+neZ7/ROPYeFlSoj2vuQ+nQBK3ABgjl0aABnFRcZ9zK6ZaKJMIfXvsmNRF
tNYvjKJ2m8TNQOlJ6zvsCc14uSotkf6EeEo0U2kYQVWhswPeYIuvIbXcTc6WJii/n+zZFJmJcCpg
Urum5UC0mzNQQrX/8tr5hYYVisEKMo4uJHdPYwUkCNg8rvFsjBidmARo6GMhArz1FZwF6pyxoWyW
wfqzcj8TLD5YLoF6VBMPH4VsV2fBV29nFb4IM5X4zKKefl3D8dt1k6+FQN9nqA1edKz2eOb/U8Ox
UxISwqUZq0h7fdlFS5sK+lI9y/b6WHhGGGsk1yst7lIOtTgXEqDAZZd5NUL00wqqlYuXgKQA+zwf
EkBT/nrNtsrLgOwfJKmZY4K9uTVKwF9H+V0MuQfoZ40MthBpLMZwYm43cPEtJXHzhz3oGDJYuzrv
XAakZRdXVXggOT5zYzWAtF6EP/3zRbSb7Aq0/QAbUXWrcthPX0n7duuSXmC0jHmKpTk4AVpvy9Pt
9f3CB84Cs3+ogMgXFv7YPi/zcD8UXVn6Zz4fuAq5Zhyemg9waf7d5Q/fkgDhjVKokSF2wNvjbSEO
vgcBZ4vj/EIJqCjvvDBn5v2OKjuct3WkCApAooJB50imlczUEi2lgqrkXEqW7i6JVdGqRy0VcBXt
XzYXHj2YI/W3iId2yIkR3nu8SRXUX0yGC4IFwPDIy31/JzlRT4y1m9VPrVGwtn4cx59KHsnICrtC
YXOinoAtQRPOmy8/Wjp1I/3J8DLslW0a7gZOfjrCQ3DdNNTS5XsdfeysnGSRc3W4REGMRiFERKuh
76BPNwdTV033mdU70bBreRKsNkM/VyzP5JiuXjHfFgCPCSuk50lJmbBBIdXLuD4LXh32VLwoy03g
KKd7kdJ/ckCoDblE4TwNxmTlj25XXddfw0tcWbUih0nnILAfsgJ5ROcZm8GmtvBS480FpFtQqTkQ
uFEOkN/IEzH5tuJCGJHWrScp4MpCiJ052vAJY+A6xiNBvanyvoxVbiALRD3yZtTcExPvuXm1fz31
nhtjSKbx5yZCl3wILagMJN3QD5WRjiscUIzNyYgkDqOBucYfORiX1LlRWt/WK3ebz5oZ8A/K73oI
vvAMZyJeP/mcfEmzjQySIaT79PLm08c7S8hlR901Vjhv5CNsGhQkwZ98IPrGP1usqDvRmD0IHyxJ
c2F9ktim8wXrdOets4rkbPYGk4YzYAUHiI1sKEDCtxOUZYG2wpDovoZW7+oAE5bxlRM6ExZaEmBJ
MQi5qKqGQJwS6CJUbJMInAmbenPWecdVgw1rXUXyKrp04pkD0EQ9U5UsQk/46pbaNppfEwMAFh01
J0olP+bBZr22ygT4UAp6xpRBnO102a4ctFpcRKanNdipy47YcZV+DXvflb33KEDcjjNF4nUJJMuK
sLMWcqIRgHDlWcMJfCGpTiPanpye/p/HI7BPXWZOwun6cqQkBv7nbuYKLqdDfxl7h8rrwuIbXvID
XBRy+gteF1vbIMLFoaD6vREK1HH7BBj7P7KOQ5s/vw3DK1wOzjKmy1jSM0gnPi2TFPwcImXrIdB9
oR5XAkMaF5ZXbj4ScmcjkPvij0l4JUa6E37Owy8Sfvc6mnJKtHssR0G86GuLJKpUhZL1hlV5MIOG
kNbcprkGUmi+6JNNlcyze0AZ7v7HvVqjDR7BgNt3PR2Ujnx7c0nm+fkbY2dZ2dbZjQk2GrIcmlLF
mwIqitRaJJ/TcnNde0532RxDfbynSMhxGcddeP8IQ3BneSX1uGSqOFSSexXNiy1SCCJ9vXx3TfyA
AcYUbjNEQImVFv5j6fy51scrWhDIal1/hFgsXsFcd/GdMsQbVcCj2PuGRaHnVUrigZoBji4J2iUq
3JVAm1GSR2z6/Hzed2DGzLa9pSKXmu9jH2acmGEKqveJJgvRxgmhU4Qg08JfjP6mnjYpAxqNrZwo
aZNJ1n3lfIbIAqlQ5hRRDYtdYWw5/jU3+rgAcey7T7T5S/XTlemowrbnfvPz590HUCTet7+h0gMY
UJkURctJfdhyldY4rM79y5HtcK2VqS8avs9Yi/1rXKwTeigpw0jHj0GtjqZpF+kqEb/yHVG+dw8r
/DgxY8EhiXHlgxjrYBe9sxK7TQMx+r64kxv6vu3F9VIh5C4R+tXNkD+DiOrRrxl9S/lj+nQdHhA0
js1pALVg7Sipu+gLh+qBO49tHFvzBGgpo9maFJIAMZC0pfsVU1OhwUnnDtFytCA2KVZA7LaeI6hI
7URuCG89w9E9jjUnObnQJeAvWA2MsXoQEfYkSlJPeGSCa9VOJoHIZ2/Re/ENYlFdcdoLhiYUpNaE
kUOKFQTqWhR+FrjhVlnnt1Ba6jfR7ofwf2SasauO6/gjCn7Q1BhgzvdjJ+jhjEaJYUqUPVUxu/lh
6i2J1TdBD/9eyW5zLy1tLzp9PxXtfyzuuhTgqfCIKMKb8TeTkkNqUqHv47acYVTCXZq1MDv9Kt2A
YbRbYfaAbfxgdOp+hO1CzT7U70tsxwfTI0fjphtx+n3pDPcu8hoYrOxrUWWbYi4YhRRFJ/fl6LGS
u0xKaPNjZAxTPyKfo9WUl4lS9qWrf/jzEE85JVLF8M+Yl2sBw8r6X6gi6yOLIlFL1BAd9JegNIGw
01YaukOVVvVEX0Vu9hnjJx9Um5uwnGpgvdtbW52rgiUq6TgMI3GMSLkMpDGarlPBMAuZ/Ns6czr/
k8DM0Cd1ZHf0uu7UVh/taRiqIfyj9Vn5VMkW+IaEOHfNQwym8Kx5ZNoD7w959AEzbpKLgKvMOLhY
RvE92axSyzZvjdC17BmfG+1G5VmuscC7NwxAaDQQ4LBcAErQGDuWktjwnhZZrmYNlnswgio8ZD5N
ksBAN9gL41CVk/NGB725VQPt5mugd1B86Ueoq2WWfRc/96jMt2TdSC+cZw36nF6qFMNjp6CNqpmU
QUJxcGESMOOvBqSa6AkpuC9OrE/nG5npxXOFzK/k/l4vbF6ENT2qGK5FPm4otymzIVVtqCoYlVx4
hOQkNfWsl3SUbgVflXpUkw/llHn7APdRSDZoYi1W3w/cTgjeWjAwR7hJ6+T6qfSelNzvsr+s/mfO
tPAcX/JtWtEXC/2Wade9lr9YIpyjXemOrusj3PfGtsmcB8XEP4wlD7MzftL0WKg8DVrVh7DQbhse
SfrUuChr60nMlfl//kLD12nKfyE3Wx9lMpmXLVtBisqhk5sGnNVeCVGHc9D46iLs93KqIKOZhIC+
S++qTHlXeALWrSoPL9NtEBL8Os6Gq1A6itOay+SwfUqG7GpKEHb4lPktWK2/mP91Bi0c6449urA6
3d9amW62y8m2F3VHFJ3XNEKX+AuocOXoyPFah3jpK8hW1sy1O/AHL8+DFWFs8/Kbs7vN918tyB7l
7TwAnJYqZAsu9H74SPMLFwzcKNmkL1MrFeB8A1fq0wY8ZDKdtJB81kr1PpiGzeoELnBZMzKpIaun
YqlfGRPxi6yLvA1gVrl+unTLSWqXZTkRc/pscfhvPiIA8Me+eWXykARyiRuTMNaMDzqPCK7rXwhq
OzsfFPKPoJHoOkcCIRjCTCb2BfbxmrDdTOv4mFeXnRj/tDjBOYnmqau7AQHZIvml2naT24sm7rz2
42f6hoIpntoAmFb4AxbGtY/y3HyF/tdRjGNtUDhn1VPXxieIsl8kME/ggpTez9bzP1td4JP8K/5C
F3b4rOB5wo6kWSYIhYMb2ObuqqqP49d08B03leJTXuOvAflM12mU7NVkOOYTj8SpIVdvAfUL9vG3
lo1ZOnzV3bOXYj8VC6qT5HtTPVVOSmnepghTv/lv8R8NmDfztKnOhEokOJB69yuWNTgJCRIkGhGr
YiiNKud5hsWpubOY+vGLUxh5k5N9nBfVRZBCKlA2ux+TY1nWninKjuiChc1vslkpIXPovGZBy41j
L/qW++BtgbngUkC8YyzWnuIHfCsXBRju6yBd/xUUVH06CLSM/MjScHBIw5Dy+IR+B06SgDdb8sQZ
2tdzkfbdwmJ18SKb6yidM9ciKbf+2p6HgIKHmMmvAzoblooME7wD6gn8xaQKb+JxJQa9ungUxBsV
7Fe0YT/MB6GrDbeQSIC9k4oGH089ZNSvvVoA0vw+IBzOhumAYEPJkArZRcVEusqr+lW9fkOjWYNr
j5ioENTJk1xuWnGzSoNVTOdNLjlON8WJLNuCg8gLRYp48Y8PatxGVPD6cJGrstzE7sd4uvHN9XyB
aanDkiNLn/xWYP7mKBvvatAL0GnbncaepQsricwh+QzAMdonHsm5yg/VjtBuMcbLGJOhKplNxjmw
VjPt0csK4myRYCjf2ARZGFuk/o4C2SkPsCWhLpZQSO7xk7NK6SU/g7R8LoN/p1LadB1yrC5EV8bw
2fJCORusv3Al5h9QpdzeYMdN7/vpYgGs8Of27rfLGd50OIiZJo3Jg9dNzR9DwzxAF2NWL4GKADhO
rM5q78/rPACW9vU1lq1wDIfr6Ats1dmM0+qbAUNvh/OJJtmNbLe8YFXNG7JCH1jViitbCiPtrmio
mvs7VX0kxac8v9NfRUIpelnHwbBiTVIpFG8hVOpivlahj8FX9GtOCfu1gKO5DUkKhDRXFh1+RTC6
40dAshY+AVIv4Vgg749641fvJWx0W4XZ0bwj49AauwJ00HG2k2Jd/fLSqyAk3Wh4LbVzYK0YaQS3
tbh/cgvflnZwZwx7CVCdn+JQ3BtH3bVV2yetvUd//lqoXzk3UGEa7KGVrf+c1hODjQA6bEkLAbRo
kRqMHUIWa/P05IIWUBfRWZMWlqRxLCcC+68vUrFJQZqoOLcyGiqD2g5929Ifo88ofp3H/oquPwRp
iR8ujQnZ2MOttsT6gg9lSOzOGub8sgAyUgFiGOmet3Ryd1rnyvVc7yFxMyFio0Uw+ANQUemRK/H1
wgLPAuiiSgmYNIAFUFC+WmQwoTCsShKy25OxOZ7LRb/BFaXUNgGOVU7yLhJksdN/MJzIOno5oT0f
kkjDHV40rdA1HL9MR2J0K6RoOropoeyXh3236//TpKV4WFKa5lV7/r3qZYehG5yU76PMDJEsY/Ti
FUCzNvZpaxD8H7mnXTyFMgOo5giFksQ9kZy1FtHO3DZlEPWfIERFsy/qe7juHA5/7/ejQPFcr4oE
XmE0n/Q3oEDt5oWLPuylZs7VTvAUXmY4RiKM1T/+zEgzu74eSHoIfFZLRgRI8jDKWUdkbEQLxXm/
He/7fM49euKQgZisLvhK12P5bdFE9//jn33U6QSbn88dv2ZzqYJiO4PGf5O07/OrrBxHT/eC7xMB
dmWXGN4Tn4JitZJ/liUtb9QaUNJYJYTMuBV9uuLFAVILDc27VyiRdqFtvg9EaOe2mkZbabGtnzlW
O8ZorpW0qwBJTeFvoW6zNR8cqP5fD1/oY4BRvhrNtWU4qGUscyBxZGozhhs18cGU0D6jqsLdsDQ2
KBIAGewhmW6N+qdvDt43LQH186CEKPWkCOriv2zgGnbt1v58nxFpJlDV/0J1/zPM7bB964D4ItFv
XeC/YSn5uvVUi86Ww22jvqN0bUXac4rKcIBG71A249w1X1WnE2NTbb9P8lAKSXACCZeBoPOT1Etk
3ryRtjrbL0LphxxxmslKTyEhmZCrsBVP8GeWCp6lHuhG6oP4q/F7did5RIWvy6z5BxH6lqQsj4Y5
0f2FJAP2zB/3+bE0SVB4sCfEG0GgXl61RDfMWGLYOK3YU3c9WlatDIDBJMXFCRrFkSVBoUFfyXkQ
xM8cmGlpvRreMS4C9VZQV2oQW4VXAliyxWf2ooQB2fIXbdbDFhL6BAZ3BbVm0LhSL8pH32966rLY
Mm0CVms8ASTmaA8Sz2Z3IJ4oY6Oa3m9UzRiNi1MPzzSAgcaUFZTPCIjc9+RZD9sF3R2Kt8swN3E1
9ZsRwkoDmG4uSKXaqHeYV6XMjkzLBvMOiZ7WjDx6DAQelr3YQ1MP4o0OJ/cZpoyjwuPVomITUKnT
569UOjx+9TA4+CnMGzisfpUgBbHQXsWgNav2tq+qDVAs2jP2ddj6TM8EjwUyE11HUhcb3Teclkky
Q01mFZoBvu51DhkJw/yt58t0nWcoXkb025KLNUf42B2JHcLV5HvwOv34mqsD5Cbjjs/DQ+1+rz7W
dDiJMaqpatXI+A0t8kYZGu4efX243h/FYE4NVs24TekABoUyK0yoEzft6dwEmYeDZqEHGa9fA6I/
ENsr/VEAv4ZJssqIxg0zP8nIS4G9AVwohnvH99isbEp6ndPbAV9Mce81KHdrM7ixfC71ZpEM9jp+
kCrpCEKJg1Z/y+CZA57Z8j+sd18ZNdGGJI4NmF4qHtYsgDAK04AKkyFKQ2gag2MlBmel+M5f8uJg
rp0XVmveHfwtG7O+Aiy0KVBsTJHAMOZRknpahGhdeNkUOtkAK42YX1jwY+Mx13Gr59IcxJK2Bxco
D6ginqc3Vbk/8aE/U+oJdyQgVaWdKszbloOMb3grE3yQCJ3zeF6/ppEJos/5ZiNYV8jQaw8iIBsp
J5nUbeCQgkTUbdDo806THLAu08jMSLP9sJJ6mrFzmY4S965sPnOSbIwPYXppGCOsoMJGDXO6kykK
HQ4MFrSyr+epSqMcjDtVURmsRwqFLUKdEbOLiShp0ZUALdyJVLWNNIt1GwlHeoYP30YczVBqFmuK
WSy3Jtmyh8DMCFMv54Aw6dkP4xpSdf6Jw/J3FvJ6tjDIIQHSd35S/N93G8n6GoK8DpL+0N9S7EKt
UgGfpgPxHwMvHfD0WyNA9CA3nFiw/6MBhwCwd6TcZa8sZDbY6uMEAJ9Y1CMqfAgCGMVqGl0tg0rz
/awwBhsHXc1xyxMii0NWtdwAK/d9qZw5G9kql11LuS44Q9ZmkLRnFkm2+gO1PvLmqMQBWJ6gg1xH
pqYxUZu1M8gkPLK+w6wol48hztZ2RgQ7TkBmupKzC2JotSWubALTLkhP/rJIdT7Ra09enZMCZZvr
vnpH7zcxb7fFsTguvzGg0qudB+u3TT9WjKeMutC82gmIxxbJAB4Xm1o856fS0E2p8hGdTXxMV+vO
/Bx+aYXAUqp5vOJOUbDd2YQzyAYSWJqMW2Cfk7wV7f26Uz4wMVMoLPW3HPlyMoy9Bl5oNz6zvl3I
+JTn4oyaZBWxn64hT5qdPA7roi0OJHv+BsvvriPZMXZ7sWqw2sJjYjl+tJv7ACGaeTerwNGvsofS
mtczeeXhYxPfW3hdKTRFQr+mGPaMFLX+eqVkNiABw2rQU0BlqG/FFaRxlqOwBP92E7oSVh5jGUh7
Pl/uWYNbuijNU7nU/FmGi4vUmf6PTIfsDEFO4b8rcLrXjn/ZRpwRJliiD6P/S4maJqwMmn+bzksS
8fDW3M0o/seWLayHYIAMhR/cjtWLLyv2J5F3m6fPaUVn74h30VZp9doJ+EQcNgOCGpn+WTs6tOWW
v5roL3nE4YhOnLXGL044srJOQMVZeMDn4uRcplyJClOA7Ot7N3nHh6wwpnt+3VdQpnyjhOoItT+I
2d2yjr1LTpHKXsO7qv2wD9VKNita58AhwkX2Sp6DnJsDyJ/PWgvKJGOY/XNjSnvPL+fDb7oLv50w
wtJ9Qer0UHTa+DJaRbQYGMoDJibGue34cLBBU71XaHTvlCCTwuY/WKNXlSS/Lsb1QmfRWWRAkSsG
w2faq7U8zVJuefibadQG/b5pKXTxQxDYAvs8KoaWi8Ikd0Qv6nMjlsO71pvskc+r05v8tKKPiRYA
W1rXuYHLh6zWscH0o1X060Uy7fwt+e+Mb6D0QNKZdHXoKDnu0XlJpGBusIaV7oLQmzn7I8ttxnGf
mR7uGNsiLaWYn/I3AFkjWgBAxMd30f44ERllMc4TKet+4ijOVxHxum4AvFdaR29uYAPFD+utunl2
0RBq1WMjK1esz/3KBpgYGyYlrkfNK5JBwb0kOpW/Jdy2eFIOVTdJXFFyanNaj/5ce4wzIxzy+Ger
vpgJMlTEJP5yY/xcn1ROz93VphN27xKBjZ1/ce+c8ey3jClwHh+9phBXwYVgZcx+SJz3n4CRhiIe
aIDoDhLl0oELYnVk7uz93mUqThsKxXx89e+TzAfefwndHUfLxqszcHX2cLB0UgDlh7G33q6Nu9Mm
mlnVVmpWw+91mr2sAwUvNgNDaGFzOTBtLpWTXYt0XlcGlTWCaXdd76PwUmzeQLFVjRcmmHhpYR7v
yucyIEgDj0Hny9m2InYdVjjFSZTy5OxZsH4OoomOsihAG3/892Bem0GTMy9e03aEcwD/fcQqIMBT
plMKUykuI8AhdbVXEmNE2bDblBxN6BPEclmfHjHjqGOiDWUWwq55rbGnkXcGQA+f741jpP8jqNiv
09nb6ckH0EUu/wszptT49LhyMGjyRA1t5bm6+ikgjMS0h5VGEQuZpttwx4Op1Syv9WBDF+9myWRq
zHVZ8RCpB1RLc265eok58V1PA1ab7KhDl8esQEQDr5FAH9pb6oBlrnTAZRBgjoeokyKbAufrBzj5
as8QbXfSHMndwmz3HwabOWC7r0EUMMTrIyvlE4WMfisA7DPFwLXPshEyWeL1GM1emcQ2PcKucu/T
mwnj9LdHUj93EL5d0flN54cyqmR3A/yco0Z3PKytod1zmTMOVPhjJ83sicWYEqbLFKGkbvxKTNmY
N9/TcnJXx48nM1hpqAx6fhRgj5ImHgjSssCkMhKusUmbzwS7U7frX+JLnapTZmRBnavPff2q/TeR
ttBjaQFyxDn+1tmoya9bCMmEVj/pWP3wQV85cK097ES0oXsg2rqM5rSiK7R131+wek0CY2owAfgb
vx4IHZTvmD1akSefaa79FNCxwBUBGmxnURC8vT+B/uRn/8oHzf+Uv/5QSCknxJ6GtUELMJkYYLjT
l5l4AAk3JRKUzTXPtnHf9nv8pWNBB3cUCoDOExrFBQtidXSW7bUHotf3jULYtHmT9RiBRoJGVgCt
8VF9NSQzjwXV86vLqJ6VjGC+8TcP0zcoX+e5KSG6rbJxCIlCP+fTIRyBciXhOg5WT2jqZpaLbxRX
DHeNZc2rkYmJKGjjZd8h15rnrqnxNo7dHar/TPQCLeLpNPIc1POWDraJmJ6wLN+qEKJIOJUoYUoW
AmhoQcD5J94CSAtufGbRN15oz1xW/62URNf5+eQYTvgyqtluK1zWt0QIWrsotNMRUp2Q9RRmitXH
g/Xgkdzr3LxShO6C+7lgkrV8GkpcsSkufT+6wpKZvt1grA+OISMEmHelkEOidU6gLT66QVsXk+jS
LM/tYqHHvsUbo+yJ7tlsCvMKv0fr56lw+PPC4xIikOuDOThHW79EMbRKI4faV1lxPnPWa5lLoSDo
qqjSjPdR2Nrn2ZGk3BsYhi9mfXx1VpijCYAI/3HLlYnIbIY7QFhcFDTZxzbGpdhN1/q0Yjz0q3yZ
GuxpPafhXIdsxxE0kakawC5Ywcqot/4q1VkUvbUY+IsyKFZMGi6/6257nv7sYfRIDZxgJIX9BNOG
OLvhYIkMtjcqSZFdQ6xPHUptT6rA2lxFuYlg33LXWjAJpPixqxeQIXsRid/q3jCoOcYHBEZ8njVj
4eXwgxKBl97Wxadd6cwuUlBnpNMOHuEJ1IibgDsahqBE8QmDjKVMXV06BpzX5UNj5dhOYLdhAV4z
68Wp3EmdTzlSe8QauEPepJXZs3dtRWtwIE6qoSAnPiAOCRGpRebP8MHV5v0Hu58WtgUFVayy9qx4
kMQ6EThLbwpTqUC0cua0W5T042h3+bcTSkb3Zvu3HrPnM6uCf/5mqXNxxOt1FKck1Lt10Y3k3jOy
fqDCHzsWQradNy4b5f+VDMOJDsM0RDyJ/fbrI2KbaYd8oMlHyCeTZ2G/2J9o1iQfQWvOBMI0qdez
df5BIHfUluTrbvEtiSdFo2pvb1hxkEBLnfZWPJKNpXnxvFyrJc2zlYKb8ZTohdxFZtOuNt5+lPKH
VrlGj/vknQ8WQSndDdQ+SLn+6zQ0XdjGLX69lRFxRdNlhWPc4RLwgnLvxTJFe6Nf6ANuKE8SfI/q
cWlvkVj9CzQApA5xaB5wYLhYupZqsEQKu3mwFCM8jW910wNWhFppILsCV3WLs7CSocjgi1uTo7bF
tSq1m5IWmqxuxlA51UGR94AbNIygOnN+GJ1X3oIDPP3HuZj5rSHIgeoqhan1pINOjwMwzMMvE8VF
QMj+0LW/98j74fKUa3WAw2Kob4vOHUtow2TRMvjzoB9vyDD0/y1aNDrMLw42VbzmO7QCZKw1Y/uA
JYmazqw3EKjFG3hCH3d+X18nxfKOWese2Wi7GH73sWGcKmsciznXd3OibnBMfJRblVGL930JNODl
vOTLwOlLcC7e+l0nORf4Tqe7FAZLjcWoeot78wiaQLaOvCwCesmlQR344FAH2nv2vvTujijt6VAi
EbCU1CC9liruTra7oTaSCf++HVwK0siOj3yBHQIQPOTHqH1aPWSrOMmIyJdZgsIY0C3MWwSnp2vN
oxgIsxui0JIwjRe22aTmogl4WsHcwm5A4tMgksouRVk1e0Rb2GybhXqQDOnj3a3px2UxuNBhP8cj
txzQYF5GEKeeim2TfV/2rVoPr57PILOVsdWK/RFcyR3lC5MwVsajeqV5JYSaBDCje+skDP7JHroU
ZnNHxqbH/OUM3OJY9KlZGhMdpD8G2lqBjNNC2q0WhMaBVUVk9vwq2stH4cbz4rTgBDmI8VEwEIDf
ACqH+JqkQp4CWPuTqVwtnBfP98TSUjUsawYxKKGnevO0vMRdHT81c6rEgN1RDg7hJTaYBUz9y2pt
4Ti+M+6JVb3w0OsHgY6TClii/qUE37/VAq/sI/KwYJyMykEpecZSJHFRWc2SiLZSZbjgoI5+ln9R
qbYzhQxF91LKx4ztTvQTVQe8SZqMjk/CJELaHFTIhKnJBUveffV5hesmYaOZ7HtRsTYVdth7qPNz
rg1fHMM8x34YapxF+ZuhB7nJvvCW/NkABthOB7+LRXu6DQbRKAeH9gErdBgy/x5xbVqXSVn793BI
Ezt919PU9niqkPEncgU0lYAqRI8dIPtZCFFqoV/E0heZfQTv8ifGb8y5ffsDp04uqXKE6iHb83ug
TM4FXBYe2ILb9xo/etaTvor3/6W3KuETdbKi81d8mrKLzGnnA6B78Nu6mKHHS8vtBjUomnfIk2vw
DbMa0PZ1LKTD/WtEbQaZxmWHM1evf/KzQseD29ECfzXfaAGY4Tl/Adwgx9en+2KZ3V4T0oPgSVdv
t3QwUh9OYYjnkZDvx94hxUrc6aVmeO4fK2axvBcGguzQ3M+di7gqe1qmLcb4yiZQyw+UsU+4axky
VGB32jN9Xi6Tf/UF1H9KctNkkbovQo09DC27cLgzOjUAoQylnFrUgPdm8BTHn03kFinUEzGumYK1
3MUgX3LHo92iyInD39EObNgIXJnsOXNH3mCgbS2DSaz8N2TBGNp2mssw4gBBDSDLZ6hA3YW47kdk
DoekXhmlKsJnxnACi4LJ5+EVS0FGjUhkjLIvaRqvznmw7Jx/gYczIx4EBW5kRXwlPW8myFYIafSv
MqGADM/09vonBWqPM3QT8sMDNXngv00kdGUC0gLVD1XAVPs2toS5ZBe+Bt4jG/hR1fB8sjCzBKEQ
E5w5eBh3hmeh9919WqRYOr6MZDq3/ammr7SlROI2VCNbeQtTCpRRm/fP6La/YP/yttnmmjP5P685
h61ss0qoPYcFpVn/lv2hGlmsPKHgMp+rtqglj+/kSR0RkMre6BcQJvyfaLcdZnYJ9Kia7Xa08u9J
VdxYamWprfq17yIQaZI5gx6mygRLnRM3xeXcxCVxywlXc3OGnb28OjcP6B1q+vK6VOfQpDvG9khP
cms5iNKCQY2vPDyTNsBPGR5c6+5rU0/TRzh1VY7VP42cY16wCilEmTEmpoWcirJ0RbiEPXJzIhNE
YY9gc7iyrjIW2wSnDDvqjSZhgrEBQQTlBXBvvdQLPf2r3Ii05cJ8y+00gRa7+LYIOkk80CJDpWpw
SdfuEDXfZYfsZNZuP3oW/QJu5x6qJvzY8isfoTM//l2KG2bNk9Ql2bEWzbFmNd4o+uobqHCnDHq7
NEIkne/32GBqZ4epHMWNFePMckDXWBbch43cKkdAWbpwAPZb+CW08wo2BrsFkQGoiaEdpMu6LxrZ
bVAsx9v2EPfbcyvhNlMhqFUkYpo0PXwHjC1dpVtcpzUz4r6vaeTWYxlsOTP962zfqYuybD4PEMBG
ii5+BBOgVoaFNFoHTZS/egHdMaC8ycVucBW3jfo06heZ4B58e2G2gb5/tx3rolFtn/nzWsCqW/MW
Jbgpo5GV9HH9uH/94BhJ5IM/7NeWk+CcuLNcrWMQRdnpRDs/Ox1xkSMrkwCFvXf23O551EZH8+d4
+RhdPYlpvmq4+e6mU51Tg4qs71GY7xKFW9zZV7qZfYACpNbe7oeTtTr0AgteljQYJaIogVaigohI
C6wOLf7Cq6v3xABnS+qQsug/5jwaa6tn20AkQmUkSDbNznjq0wpD6JhdzYLT/d8OoH3d5T6cYgwQ
4XlBQythXOcuSib2n7w95V6TfH9tWIBZJhe+rrneywVjQlM50ZWrFPUk91mixJaoUagnrhd465/G
9rN0pQ1bxDH/E0onitMLJLmPzuHAxSDjDXN5G8QQL4gclUWu8TZGSq6Psxy3otJMx7poxefQI+O+
qkkl5V1zpjkJlSGTaHHvR0JPS3m+/k7/A+oiSPmdMCY5fxXMoYBWt1WZjHxZZEykwLJ9X7bdDMXT
c9QJmSeyP++NfVppGDD5Ni480w8JJFuQJk2fYw0M6XJEi4q0HEdJWPZ84b0O1wtPFNKP/szDNDbu
IdoU6jn5zbfMYPUIe78c/eDg7s0yz1dbuOH3bg3dt+4mDW8iXl4n2T50BO6FC8N9yfdLgfG1gqb/
KXE8oOb8qV33Wu1z3XZUziC2p1PP3k8xxsGO3Kh6DK3YaagFMQsbbOK+tPIDHpx76ABfucs5zt3p
MYHdseOXWf+xvKr2IuSJUz0ZvUOqVaAjzJIsCjMAr2780eLlXGMMSBsQl2W0UludqBGA5IilOAfk
wurlvgS39MlZQNf3L0cCTAdFapCTl1B3iBgu/oaBeMFsiSFdyWc+bhlDAezQ4tG/tzNXbSjcb2zg
FNJE8G7ZYLcpUzIrMQIBQV9XKGaW5v1TnrA6WirWIzHS3R84F3An9h838Ta/3MUAMvR5l/l7N90P
0IDLANLtC2MilUI6saId2eL7RUK8obSp6DICF60jNZLnAITvNl65Ve9yPd769LAR0C/wGwNnu30/
dRVxtA9s8jFVRnR7LLU9QImw5BnhRfYOfm6MTeqKIn3kkPLREhDkTEdN9gIIU3jD3ngv5Sy2CrDg
K6Y2PdbnDSepGvazKeCTntIGhH92GKLoapXhDb/IavjmBjqXasijePiuW61ZovRUp2EPowo/NRKg
nJAyE41gYc3bEFFIgfQ0iftVtft5BXRXEGSNv2gfNFtsIlleHCCZ27B0EjFV6wnSqxdWO+dMCljB
SYruprLKMoCZmkBiuxqrz3oaaV8hl1Txx+QN3vLJbjShXjMWE+PAfPKPDNd3mGU0KhRLNJoRIJ7e
v8/v1hSYXlfwQSuBGq3qDzAyjtNmp6B8w5W1JQbcK0/Y4B9m8tj1QguuP4iHzVWWDrZaC8Y7yH8/
lKl93wGw1S2uWATqmWeHYIjY8RGISNiNJIbP3071N/ekEhCtG+Z3XLdYkoMfHuJmWniBq1tYo5XF
cXeGSNJY4fCYJfJdkuopGGe5cEQqYO9cKORxnWD/z26hmCRBGB9f0rcVNIBSj3fepGj+cZxQ3GEw
W3OjTlduO6/mfNt5+SmSWL7sAv6Ajq9I8VQbjtLAn/JkRg8qnPOiXlwugH+stiJpppEkL4ieStNY
9bIoKsv8CDwmRZxLon+ItePeXG1L3akay7wnTpsxXLpv73HrIxkF7zFNfJdNUlpaPh5UP5W5o0oF
KbDTZPWQBD1iQx+YWLGV6vkYLNcBiRqzzIATAuauc3ah4HOa6AMBaYYghFmdPssIbDCrm7NgnUiL
2T811s2+PpPUwVi+qVl6gK/KFIDOMOi0JzjULUuYsFlNLZgk3zp7EApb9SOM6EcjGkMAOfP5SK2V
0oIa9R/tu7D8ZIpPlMWNjyZsRoSgg26F63TkqP+qnuH18Op8/PrD1fgp9Jsjp9FvMj3t3pRp31KL
uefR36tIOvRtoYxIQAJ2r6fM+SWMPER2HFHQ6H6VoQ1KwSxHPug9App+3uQ7wsGmU5ShoiasXCqZ
ghDGby+skD0X2l6UTAvANy5dVaclbwI58aYQQC69p3sCqWob6kFKoHLotMmFRCiv+A5X2GwjLaHZ
nR3iHCYKmlZOOMXTSXeZ7aLa5rAMAlJzIeOIsqEvo3W1ynecLDo9E43OUcWvVmZoQIs5valdIfF8
ZoIAJBUSprrvNtZbK2/Kpzypf5JCJU6xA24WClQu8OZj+W1WWn+aHNSwQjrrnlkKlSs4AEVI4m7I
0TpV08Fp99YowgudUSX5TBhDKomBi2Rd9bfREBC9G47nMF7w6SuKKace2Um8OKHwHvWqVAJrFUn5
My+EXFawSxiFyNCy6KRrMjRiHQVCrA/9/vpPi5ZqZamKbdorAxkzpbxH4ZVgN8abXfm/nl0/7n1Z
g3oY3+wbZuXMuWWSqtDfYXyaQbuTVVlsKB8ggDCyxoxdXOxvr4gqhIyRu+1QWKVgUjm2sBP6+TBu
gH+v93q4cqeNQot8E0TlsaqOIZyswNo31RXTmWLbaCiF1NF9VKKw9HWxixO2cl8tHSefaDNlnOcJ
hHAKEw6UbDH0zbuzhY7JnX6xl0Pq+9Dqy+2EymqU5hts8SPN2+XmpmHyMD8XSUtVbFd5Hg2XbH/+
lbAtTQrOr82tWgLa+vkwoH3bKMJrgGp0J2o2cnBm5omMb8z93qg2c0xfmH0fYAgR1EXXzKP+K6lQ
Osyp4xdx42iQ/PdbZ4n8Ei8NBNFHNeNgjmY9bvpjDaeOdMXnpPoCsolKJs0acwioVEOlXcHHuT0s
iyWRtkYEkiTmhTNAceTt+DRg+dW5dzEXz01EemKeJ7uXE66PDs6tzd9PSioiUq1m9de0opKbIsGd
yRRd/gwKngkO6LEwVjEQcvf4JjjyedIRlqND3pVaBkzuwm8Yrde67Hx+aJsXPBpqJOUTCDSG+knl
qDD1kB03XbxR/DvetOsXjY1Gf0LxR9z/85UVb1bPgmNRs3PFql9WmQgSHDJHKRJCTdWirHTKaqk/
YkfCkSxjXqIkmQsD+gMnWqdgsOULekX0RXJHEY6MLKpvhmuYbWHm+bZXJrxcWwMLyWSrcgyaviy2
pu/8ixJuQYou8r47KJJglSPlImyLAa/jcOM7+jA0S5ehf42ihv1eGad+zmg16ktGaFnEZIb+ZTgX
C4KNlmqr1LqQE8WwRJNEIUNBEjAcWDBygTmoTtODU8WESC444N3h9IUkNCJgJ2XZUI5UhTxAfwOS
fn1Z/p0io9XTeWhoqslmbXn5tmo29wOf2W3LRr5WXrKg1h2VVC/8+1rYG6joGy/FSJbE4VBBvpqk
8GMITFF5fHdeRPYOPx7Zj9tgqLj6K8XVUWMdY9hSr+BHDnoWMqwGc4NxC62xIIASqiHFtEzuKZTv
LqCyZNdqA6IZBYdTrJ5sbtSd31qFbRpUq56FXcZxwcs4949bPo9HcisMcXaJ92lUGaqgxhcq8A7j
DpGJ0AxKZ94D5HDKXMhaZ+K0lo91hKr/7zbCseOWRfsoKzlESKUDD8blMsqqQdu+1sGIfCcsJfr1
aHwkWIXlLzpyW8kLVTGfOQ/hdftnJQuCYaRebHJOAAcktdkQ/5iff+L/Ahxx6MqJOW13AFfTOvl7
loT7+NsxUqQarLZpFlE1WB7MTQBdlh9Xggh5qLifj2kzxbPFaiWCC6gpm8zG7Yx/tEWCv68C/Gmh
89ztI5qjbKEv3IqphFnJGUwnIndn1B4aQP7+su4s6lX9oc1Ic7/KA4yVskC2Y+shkNxaHyhX/Jcm
TqCW3HZSxWXozXEU4vtHhbQHSbADMi50Gxqe8PND+Kkp2vX+4S670Vk030XPpmO0b0OoJGK6T5U+
zPxs8zF13A4CekdHRYhVEbKck1sB1nqN0J9JRHsFYwSnC271mK8U2MJ57gVKgq/dxFBbLbDHIocC
3PuaoqhvXqmbsPtgkMwRuR7S5aMIOOWb+GhptewVygDnL1PgvrAWGdxiwSa517Yj7LxfwfupmqAM
we0b0E8OQ4KegPJG2tpGUSylpgYna8I3+kN/tasOSApvMPK7QWQFPyDqY6pNmpRqzggQnnqecbdI
601Pxumh2WdAYoVcsVpbK7FQQJSBBT5/hyYMn9tEhZg2WLDAOU4Ef1Ouo/oaShyfb8RGc43FaTAe
j6cGC+E+NMuZXlTcSbh4qv7nqI6WcNqUVCGnx0vZ7gOseEIGof0v8QUjbkMfRNJQT61vx8WsHvCv
KHGUVxuUMzHLsaJ3wKM03hn/A/2cXNdjKv/mpt7pOTeR3kglVz5Zuo3crIxdZwBiS41ECiUrsqgK
kW9uMW3cwrs4mh07m1GmLkuNj8npUksy2Z4VH2PsZFe1NzdpsWroof+MNl4qwvQW0QQUdvBMBgK4
gPz/uxmFBgdffAVERJriCFKVj6QOMT+viKPxbRKT9/TBOs9r1LEkSVVszUel2yjzjwERGZm+1kxG
Zpl/56Hjp7WIGS0q6Yl+n3vdPJuazLtS/U/XEEZ9mP2mOWI+YWJy2DadQ9Yq6VgKW/SCIGmu0/Vp
aECjlzdGaLwaq8S270aww0HeHm1zH8y8mZPRr6a0qzeo26H63RETcKWGu7X8rA19IyCii6YhKS1l
2XyNXcWf6cqz7ovlkeT9KqBlvg98bxIaB4XeGq9yJe7VZ6rvLN1pX0dljnYvfyg8H/WWuNUint4y
/4V++uByu1ofRQ5jF4N6GJIkoW5Re6NxfMjqSwtZYBHWPq72K648Af2fBOh1ZoAdXEQsgJnH5ixz
1dkHjfTg22PrIV1o4YoIF6yxXEMR5649PlphzWilJD61S1Ftrb9nlAPdPoUNWxqZildDXBntMbUz
SaJN4VvNT9w/pb0ccVKqSYNDjvJKgIKfSpjIC54L/1F4I21gkwZo0og83Xn7TLcIIrYa8i6Xw1Na
+mly3wNTfV2eemfg7ZoW15SZgCfLITjnEl6vvHXQV1hOqI0O/IAcGujUwwbmFbW03HJqsLgMypM5
IXKqFWTNxXerDPILU1MTjG4Mb6TyD6UjGwbzQFctzWrBl83qqcG5zbYbrnnq5JywSX+Hcbm4H1eM
vE1HvjDAZBMfwFb7cM/JSoCIrwNO/+ADNbVjewPZsPywjcACwJrLvwjqPt7Wv0at8g4h5sKoTNPT
fjlRsBHMBaUmfNrb236YkfefXzkKvJ1cwvoSTClxOCibWI2xLxIhErmyQn1i5P8gLdJkktkUbMLQ
QIcJu2F2LPbihpX0dlnyHr2URzPfcTDKh5eZONoFdMNgaWXwc/iCnE+4lilC1VF7Ygl8PX5amf2l
GF3c1QdBUVskGd1fJaUESA49kL9/Z+O4axnbB76IacuouVJQ2OHhFq80vmn+fIFDSejWBfWDabKH
xPKIaI+6o4q+anYNyo3X/LY/XaVunn7Hd1NFH1TyzELOBGoNJOOTD757mrcPUOYr2OropZs5yj/Q
tmquhlG/A2+Ugwy3zQl7JTMmDLsNtIGbrQQgC3A6kt7T24KfoTmdbc4zf4gMvN215MODqZknC6/j
4M98d0YojX5PGZfYwd7Y5Dy4HtJ9FyPXGlmJtAcbi5YYyhgI3mb/vQHKHEE3slipp8twvWM3Elk8
3NCC5y2ftoNvF4PqSKjJ38+0vo5izebYdokRmw7d4h9cE+yh9NUd/pUsFiisswaxKCYk/EvWFDhx
GEMXH4BKaIudMySSrZ3LLuEZdq4AODQHoSBZN9WFgR4kzTG2sUG2I8nWcNQ4IFf5EGPifMIoBQPp
lgeVxaX9wl5Bf1x/ZmLsMDYFBjdysKQlUB/1Hgf8Ig9GdTHADPXQABFEzwKMDUiHqFqJ9s0jVxww
Oy5jhYzKYn7WXheyN0yC5oE9XxjtYdCNU35DlA+ftAOXLkiw9EV2RpRD6jQNCMQfdzdgNUZbghZZ
cAz3EI5Ww7I/1K69r7EEfCTW/50wNv02LGqFXZSeB3tX40Nt6Yazz8+iFiNUgvJA3t3eD/L2r1gp
BW+Dmo762UZ3locfKS7ayfYg1lCA5jG4skTFUvqh8vqQOuGRiQs8DzLGw2USqeqX6r2j91SggPox
9gchtgIpnuw/48V/KL9eQ7vYI7xP0/TiQyYPYSPmKq8+sipFpuojMjIzby5bOVSSXkA6PzNczJF4
mtnV7pkUV1OTCkQX7rWBoSMeXtrWYv4zO/Yxphjgi60ZRjlgCa00MVqNI8fhTslGJqmCjmv+yrrR
9vCKSUMt79D7wQROGMA3c8DyhvcWDEEi/rTYOZilfUR8oxBdaJjZ9rqFW2yXQe2fE9JRtLjMPaS1
fVSHVatoOMVQZ1CdhdArSwMIXISRqXsfxCknITDsrHLPCrDbp6fY//Ozqk3AjHC98LWiuKU7ZRDm
FmzLiO6RC0vsTb/7hJWex6SItcGcuAloalpqmgVrBKCfVMpDgr4wX9kWgrRf+TXU8w9Obo3YbBsj
6vileFTjWLQixwQoyOgkHnKtYto5z/ZJJJsfG0EmGaBucf6jQ8Mbwgzs0M6j19ciaIcbljyUW7Mq
gOy02LEk+Qzdz6HSWC+0MeBP0Pd3YcnZHvnnmqK6RwfN5uhIrWtT/RHFUnP4xPdhhAffqSrminAt
tX5h6MuV5c2eGF8YCrMoUxL7gyja8jbIEpcKLaVcW9CW1CZXKKrZ7vL5Y7zrw+eRhl/nWVFjms+t
ojVJgX+T0T7rfCpHblXU9TpLsy5ouuAXiAvNjtKHfFwW2QWFdgO8zylfa4ITNm75OQK8/qJWcwAO
xeixnXCRUtHs5SE2LfXmPcwHrYVav+mE08pMn3fQ2UCSToiiGwUH3p3vNh+dvwsVSxiCOCMRBUHT
FEuxYTDyYy4Jy9j7gz74dvb9zxFkebBZbWWQ6crAWY5s0UyQafEKxfPMKB/nhY1msoK/ZhSNyNQ0
5yXiDXRgb7QWnWf3GgRDPgI8EMcKbBkSXy5VZe+J2XmAfXvOjpyBNrdU3zb19mza5ZI0IcWWJ51I
EN6M0tnYqRO+jB9x7CyeD9p+pRHQvwS1oCR9mGO+pusuasQdVOWAbpWSOC3mD8tnxztPtr5j/otN
MBMfv4LUnicApc9I6D2UQHz2QyIcrN9+jEe8/ty6mdT4TtMBQv9pXBC/d5Qix0kAB1ftyGOgSkHj
yKSeXz7UyplJ+Cor4eaLdqDqA2XDYlrJsMIdkvi1UcM8B6l1ISCNKrIqrhmgp26KbB22vHqSqt5s
urg2VlRrAp+jNS45v9q0Cafc/778BjnfxUeLvC7vfx4UePX1xp0YCrhYUuimvtjlJFyhIpn31GVT
1Qcn/j154UBKFtRDZo/TB5Yq6ecjlOUEbnvc7OWRl5RHqGw8xsRBdr8LRh0CkiC94FRdF8uN84bN
kBWZhFuz6eF3yT+6Kr9T03O4CihLU/RUdTmJYexFZjur4+C8ygiB0gYr/GjlJAF441yfgNrsrRhT
dcQa6W5cXI0cwYjCWTa1mMZXyzcl3SAsL7NmsyW38Goexu7110oco5Lox/kkqY9rNQ+OBqhCnelb
KpSj6eqlmrY7KjoE9jVhS6qbxzwXqq5GMimG/H/U2bBFWs8ie2EdBJQ/1FuRVE2Z59D4bK8c5pgK
Sp2EkQ+ehwXLZW3aItbMmi0w23t9DRxGR5kDj3ghmoLAe0hclzfJoqgYat+J9VvYFyksGenZvxHq
z7TbWACTUYPDu3ZFv68tQSqXQo4x/39+4XqA0YAUHnbxxbiFK4QyCNu71NVQ+tTg05eJlwytIN88
yRbQrlTTgWJ3ubs6I+JXP64vnnuQayAEJSxNMYaLRCt2lp2S0d0RWrSAl40HFl3B1Y9p7Z9DlqQn
B49AMEp/b/nrQ5fBh6/SlUjYWpAL7xztG3GR8lrTu3y6ilESHSouGfoHKOTOt5+rRS0a7K0M/2bw
Pt688YaY8EhR41rLfwYsljqE7oslrGerMEUpXgkK4d4uUcZVeXjS1vI4opyKndXxp56PcHJPzLoJ
4DL/LlHt35Ab4uQcgu+vq+KigniZpDKCTKmS0AqUPjALlLmjILHLJO7c00cstFwhsMLzr8rxSpfY
zv57gVCBVRONaUmUygOwBfAcKmwFaumh9p8XLn/cUR8QPdRnxRfPpoFCEJsat2BfnF0Sn7tUoyNO
DWYw1npWHPvFKfg3bD9ctKxuYkOlpt3EY8eiCtvQYBKQECW4xcyQCC9jwq7/PMm4q1dNQouanY+d
oZRwnMX+463YSwKR6GAIIBvvYRYSj5fuU8M+5s17HBn5uDhqeX8POChPA2s2KH7wqD78RBIqL5ww
sBSM36wSRIERdksYk/L/2KEhFyMQqFR5KoW14CRHOUtxawSGyJrR5vYm5hHAiQSrOrsKPiSxPU+0
fl21HLI0WtViHuhFZnNnV4T5IxEbXWKEOIQ1paEai5BScZeqa4egTXzvujS8pqmhw3DS89aMgxK9
Jnc6eeoSjzyvM+BtZVcIGcP7kH1/Dk4N4KjEGUe+GUTEXzr9o/MeKX5ZdxFqx90efju9GihQqS2j
fqKyKsU9zSZpp0iW8SI/ou0uXSyE8GBPh1yOVKkYxFY0s4B0ezRYl5A6s5t+/lEN5oInnWoX3fLK
AIqd3o9mxLja0ZK1kVSxkzLNwxi5+gS8zCtpL7Ztvq+1iC37JEgcpw9xFiQUNqhZY5159XGDa2Vs
rzi/qa1Z2ZyF4JXXGzfUgCG3ju2yraw2HWv5YomtqUBoIyXaelJtSQh7yFMTEO/yUgqPTJcxzKtw
Yzf0LArtxkIfp0neW+ppUYYyg54a7t2TV5Ri3LotTnbv3qE3bmiJM6HqZOC9Zb4sy0kNt+C1hTiY
IxZ4hS6xLe+HGl40wJHtJGul8azyaHWBTpB95It5lV4TKYsxL/CrNLGM1PUEpWZ9KB/IR8VJwKWj
BljVZehfd/goXA/e+bcPlCs4E8MSa0ztgkMCm+TaARHqWqOq4He1Uv5FKxeruYMW5pghNiMNDSc2
BSslCFfIAvH4CyeD+xg20l+sX1I85dUoINxc1Hp8obgEVrgSSN1n69fCjnzUC0UYrwh+RJ3Q8fNy
OY1Sx8IpZcbLkuklqasdoKtXkvdVS2cz9jUOY9yN+BOo3BrFH1B0Cwa+u6w7R3jK24PVorTHnHCL
Cd6CA/BoCHlZSgZDOKLODElJKOOatspzQElMy6TuKDAJYTNwF1R215x0+IR73+aFyTVLrb/PXvnl
BOfRXqrjY6m/N+4mABSEhdAzqdv17Q4xUuA0+G4zMEj8q/1SjsKy0nME9MjX7pXAV0F3ozKnO/1W
QOGufYxqYbRHyV6SGhP2LdiLgW/4Sw4V1lthugQLDnW56mni2M4Zo65JMt78XkaL0b1sjGSsMj+2
sescarjtsSrkuHK+cxRQWMENY0e5ZzGfNVjFP1qTVVcx83B+BAiJfa8iHPnEml3yITJGD7EEs2wq
jG29aRKdDj6f6ZysvPRqF6vuGQjr8+UY8Lm6HaOMoOIgP4DJczok5GtzsZvMXxaL+tHLt1CKVHLP
mUTdhCdbra/goAWGegRT5nUyS3WBMbjRzO2mGwgpY+Wvlhkvqin+69VZYv0C3fedIIhI40BUWPE6
UQuYDvXGtmCRzCIz5ONUrC4EQjO/rp80EIEf57Mubtkot5F9q6GdW8KX4pvLRetUZ1kLjsqJ/ydq
1lXaeybam1lWlIniISOl06M1JcrAzcYj+uEo9mBUPi0ejeXmHWKbj5wSfQv5eeIvVlGwnXK+SGMs
KUiPXJ/UfR2AfUvCNixoGwlkl2A6ay1p1omtZnmrrVarT1A4fdpzFGfCB4zfDi7XM0Q4DwwCpSzZ
gk/STLA9isLXw6YQfydZPu2+HX5viZGDDD3mMHJqZ4nUf7DgkcDi4m4WKMz7SLVKT3kEvl0cKFJ2
0lzAg5bMe83XllybyZilBC7W4Jym+PAn3NjCEKTAC9AOh3mTpEwXPPVo3EF5KtO623PU+CeIbySW
36JdsVeUge5vKXSK/KGRJnYJVOlkAg0aYqG9hp/dEQaNFEd4qhSASOls19+5pk3i0fLB7H3tOFdg
/9Q5fPH/+WxiTzI2NvOtsgvv+iT/h5qNiz1eqacLC7hbS9e+7zeE1vi3zGHAQ13766dXt1uPeSQP
aBPiqms0+UFEVSvkmOAVI3V9DEHHrECGG5POsD/VH3SGXBTxLxLWZd9giy81/qSOSomHAMBNvUVT
skrMSdoeiXGbql1u6Q9kkQkJaWa9tQgtzlKzLPoV3u50pw8yqmDcdxb3PllsI0IQQTVky14Cv4Iw
I2u3iubYhrcgroI7gLQj1saDibXIwX7M2ihL8Zrz7NvBEo80ZsMum3laHw9Dpce78MpLRsi1xwHk
w2WS1cKYGKq3eZFr0hLuU+pjSElJCjZNWj3zAbw5ZRx2wUPDGDBjfwMA1yxFRJ5w46oWLCICgx2U
0h4Xj22omLDSJ5PjdBanHTaA1KeDR1wNbh6hIszGvqLeF15aXqsw8JXqp1EXYhp7wsaipSA97N0S
zmZFxHeNUKInXkRFp1EnY/KSAOlnKMZSv6vpYXqAY6dyxUXUa3QFOP4kH5ixMHyrGNAtzvowDHOI
X9NKwYz5734N98LjgjwC/wRJ2YUMuVqIIkDWhuwnyhCjuCBGL//ch1JWDZvFeCvtMDsRzwmyQ1Er
Ur46cy+dvHyJ8tyuVedlEkM4AQkNthwWSVBoJhCI3UtpMDlyZID3lMexIODiZ3Cq6se8A8gjvgOa
TWEvvgmLl66rbVJdZLJnML+OOQhspO/k8N5J5g5OGV6bZ1PQfyozri2pojObjy9RdmWnb+OJi1ma
2DuKuEWXLib1GrWD60l1wFQbOQrE5DMA0rF8OlTMNDPg79SfVuCeEAc5yk3BW42S1FTYn/Y+hDCc
Ojp4N79/ZCmHNoFJiYFSHHkO69huoKzlcergsZ/ZWqWxQbDvI6Aj2o8/2jyM29Lu6DjXgWTJKMNh
/KAzU0T+aQ1cQBQxVHiIyfq98GRzNEZPUf8wT++DTIHXTrF3TJ+cTFa5QBKWkewExlhdz5wAoZIc
0ceq5BsGvtyF73NM8OoR24XY5NudmQNk4CgscVFVyYfDHGFkttgGCgIthqfxkduC6Dl//I+dzqpG
UsVGiGLxO9koFpO8AVL19sbMjtKxLbn6tI1CgjDZX86zxXkp1dX9cU76Xm/DhDLpchz6BUkbaGYd
85ijQZB+z4ETOq3tzAhzN7ZwtnAAwSu/PxEoH+5z0/SdLuQG3aNOt1NnqQrDDHK/Qy4rDQf6jsQ4
OOgFoWRaxyMGbhOoUo68kYSw0cH0FAiOXy6SCfMBddt0i6eUgId4Q9025yhh5G4yPb3qlIODLEPb
TAFaT9LUDd8T3FlrnSjBBLHndH6CzzN5HPUoRzXUjPQxqg4FhNDcYFDxmffAuKW2kihTH8vBeByn
bl4oLs8IWQLElisw60WYUKoNNwkBL3agfZ1LBFWBkkrH78IWN0JoERFncvQupHVdoNq2nRFyWSGM
x2eARY1XPpFaDPtVxlLuc/jw1WRzLgWII8ViAfMgb+jUglFcZ/Kxjg8qZj9cat0upHogFTV8viuc
DC0iqmcvPKbjAYSyqAD7/iLwr9N4zM199o2iLiMgEzc+xRkSjHJ0RcQbcJEbIeZDGslOx3TD5Skz
6DZvzRV914HEQszHyKp2rQr74cYl1iRqOYuSEFyA/jF8HcaWdhsYyDHlVKaLF8BlI2Iw/KJU8J80
zBrYM74xq+icPD/nf+HeJVVARTlyKj4OSTqTM81Qc1iG1yXk4hwb5X307dlNPxsCh3n5r2qt/8PA
Z/Q84JL6X5XrzARY7uhHJOU3t+lTrqrddyK9SEWdhvCGc6oPEBVDAdLS86lIrILt2o7sRBJ0WPGI
n3HpNXtu90lnlaABWPY0dnpJv3OkB2dl0tFHnurpg3oqI60HWw/d1V1W45Zs4z2/GFcd7/fp3GW7
PKL//Q7NQifC7NfvEd5v8nWM1ZgVn0SFHPfNE2pCR3NvXUTwtiKoAqEF1ZezBqXHOxu2OXi/ECUF
IyN6lA1AI4JLyI8Zyx+CxKyG2JWKdWRgJr7sH8Og0M6mszuHGjjfFw9UjvFvd3MUG7k1aN9bDy6H
tZOR1DA82ulD5QMW5lKGH5y01nokmUzxxuUXL1HRTguQKwVuCtBcpmcxJGaYkg8wHrCFEAj2WQkv
4JitEjd/CzGIUVQ/3EybpoZw0su+XHIUbZ35DTCGHB01HMCgcQBLTGIrVDO1IytCUje1TY88tGnt
S5LMnPMrKDtala4q+lartNAyS7Ghr2IAu8oC73wJ6YoW8SwiKCJ2shfwZRxnOUZpcfqzG8rF2MHH
eJUZO9RS6H2Ops8acmMgJ/N3ZohGQhOyHeOl/AL012G7y+bL1StpDubQFPLOU6u72sDPwPDZ4pNs
WPkt/xBjDT2Gv/QKHOm+a3tjL7WAtlR7lmpbI6t9N0UoE2n4YY6kC5lLSUL5I7C2T9a4rT8f352f
uRxNgBSb+A2NxSRZDPCvl9AH7i6najlvHgE84ZHg7B5AJJ9rSx1iQ9USmmrXpP1qW97l8JyfKXpx
R+rjozqPFg1C/iTkSkEBNrA/rhLzSG2+uRGa4IgEQWqe/Ezg6rk2U8u9O+sim+yq62ImlJUYGSgT
F3g9cLCCDLD6zS0cKXuLNTYG3ThxWALOJHoRT693f0A2LqOA0f/R72trTPuEEBVYZAZn3NYS4YVb
jFZt3qwXJlvA6Fa4YiJugMIHC+uyp+dArPpCuCcjomHZTlXRnF6hqmzzuT2Omy43Ya1nsPjuXAw1
COfhTckI+hBRPGaADnV1g6MMwHyQ63dAg8nmEOnVKtgybxwl0R3nLO5iQfGSk3lm4hBbMWmX082S
+LN8+d/tCgRZs6X2jIYekZ4J6XeOT4a6Krh/M3LhUzeZO/BvXserBj3xqGswSbRNIi1Nw9yoGBGr
/S/FV5KJXj8SxPAAZWxtULdbB3HXbacC7RFDRQuulMauxDVoXKQY4H7vF15/IRuU+JFOtXuNQhQR
7hQRPttnCLg4n/prLCsORblWULPEqf+aKUa/1iSXkUEMDs/JNQYAmX35DrjxvPT/B9A+CdCSLVzb
jocJ6zYa1fN/EsyletCzNYc9OMo72zKJ6afNXGgoxoj/ZvI9LZd+f20TKrImypueUL6XBFiyQvX5
vgkO9QO6ki3Ew+pBXjcmvjA7xDhUtqXZ5Bbf3b4h3OFDhfV3Fuy72WRm25Hli2nWEnD0/dFiz7my
QaIiU0g9nGJP+sGEPNJSmm2asZTNfFdAHpp31Ec9wQTZ0UQbWd+G79lYExEzBJlLqUC9xBDoI1tG
I6d3Rq3obDsjYVorxEE1YDTjncBdesF4hVMmDoBDAJKvtu7F9yxQ7vVn25hL+E0jkNqwZhx/Ufe7
Qp/nBOvcbuE4KK388G1Pmsvg2EdRnCIJJ/jdHQgotWrbpG1L2z4A8uAqfxQzmCNMVGLrKzZYWRRv
BQ8Lj1TYMrTRT2PMQnF251uDZtUzoLrjfbP4vSTG4sjrIq9STFhD4Q/FTrlJXd0AURZZa4VN9riN
uRWq2hbZKVkOJVJdkJFDApTjxiQkPZ0xWsSk5FZzifF4Z9x7+6lzFTkKBSNwwmDtoEXVGaEZNx9h
gWx2sOecE/+iMyUUvISdtJAYEHCfPXPV/qsRXH27WCsnCiJYu4hFTj1XSZHGr/M1OZIuM4Df0ssN
niomtEg2QVA0m+QiK1ev4JH3a/att9tLDINcj6yeFhd7fTupnsAy5LrumQVdsZwLkykUMeVxQfbK
RYD6MxleO9kuPrihhsSAJC1PXcxxVywhk+ZNcaNLksBXXhxdNOjzs10188bh3iDieA0WccYbSu7w
cQtb1Z6q0lbKRTM4ezJw1kRGLw4kCwJR+Ikc76iVMMVUDYKtp06SikcwyYO2z1z3b0sFJYbKQXMy
pKCfEvfH9jZCqr3jcKDMQfvIkctDlAVdssAH1YC0Or/i5NulHqXffh/8kSZpNquotalIs5VZgwJJ
10D2SAXRx8HU8aYdWcqsEUAZJp6ojwq1PY7wECivl0D1InMt4/5iFEWWEYG16OafiWSvS+F7InO8
inLlJNlCDZ91stzf4M5Oe19a+LimEfSEH/ThUGgUuzAgzdZ2WwyuhEdGBZQKR5zVk6odsUOHByRN
UDQ91pKWwjmCeG3YciX+V08PhDb5DhAgxwYE8CosPGi3nhmP6WZEMqU0fuLES6hNb24J8BJ2D8Tm
/O7LOJOpP8Sfqbb0n3aWnQ+IsIZAdQB2V/EzECFWmkmqFfGVUJAf8381+McZsMoVpfxrjrroOxgA
IhPaLhBi2Qys4jrCK7WjVmD4PFYgO+um4JxRgwL0RX6YGBSeRAeOVUl3LV7uSgtz4XprOPs8L2E+
vQCdPCU26P0FpR8UqFEgs6j/C5Ums6u3tOUwLqkjfwVjv9p2c07rfD0VQFcttZ0VT8qMe5+HGH8s
L9qC6ulE9YlxMloBwPdZpt13LMMRj0cmpS1XgZZPM734F+LWPTmlwBk6907NgfdGZe4TSnz5Nx7U
Sz8x9+Z8QFqcsD8QGjvzCjwxjDVuwX783ZvspcXcUA3+QcgMGO2gtwaTo9lbBrT0QleM+znfu3US
nxKpNb3HF/xEdBgHYsemfxc1BFx+15uOjAag+JfOhBFErc8wwsCcYDCDK3qDSGlKyYpXa8uacV4A
dYxOLePxzvfP+HBYeEcuouZVQB40xu52xMrq0H25u6kTKGnM+wFJkZz4szYPTAnypQQcJDSqUq72
9I9v2z1lsruLNfNyFUMMe+J5zbCtdyZGc8AzNd6im30Gqx5EzSbIlmLBqdFabccM7pXcrbTan41j
3i1sQS4KEia4lbJEv59glt3iMabOdiqNsep/ApGELLoTbO5OmEIoB8RG41bzjZor+lKZsUrrwiJI
j7PranDeANCX9NCN3vdpRdYrNfZ37F9gUceed9piAqsGre/3ESm5dZugQ5YhDJ2pqrzt1oHiarKH
TTG7dzJxLz7ZUhPRA3l2z9MqNJiGWkyx5hmTeVyevSyq8R+At/7Jz94vk8rZ0w24BNtSQ5oAhtsM
WhbRu1TaaFI6HRsShpZSA+t3Ot9Lqs6vSkmf8uPbm5IFrrUxlxCenOyQuww+3ca3WofIa33Pu+Bs
4BULYaSdjlX3mU6HzOrBGTitSasRanCn7ht+XVjQTvHrnco9TpmWGbZya2D5F8Qio30Xel1lBIh2
PvOAnjQSTWYu8qTcm4lGj0bGDjdbnNMNfkyQQ42zZdUj0JVHR9Ax4jcRA1RzNb3LFyMawbgMhPF5
J7vF9DiJfRyHKCd3z0vIuZNMud0vNdjYGdtLcU3plk6CxqoFJryFuNWjKg2u8ErNP2GBSJIWf5xk
OlqOa/DOkWUZNZTivirao9d2YqNWrsYikThe/fslIpaFghChP1PeYH1Kfca639rBf/REpQetWlGc
CKAZVa81BF+9ilRV6JilyMoucyUXBwtvxp4w92sEyjKMVeyvtONRiirQp6l0gaEAkJh15qlUrpJt
K52joEev6GZQhRiQB4Zs0hyg3FfRzUEtxYCqhJHvoJouO+UrZUZyqrlrv7SfrVxw8xfsHz3qyNes
djBkSdl1Ut2ioHHqib63t7hN6c0nNsCOD8fhYvu3MlsIE7uizQIfcbJcY7JWwQbEecB35UgXRH/k
LqdXh+9x4J35QfhGswEhbIv/k7fd984Ucs3elhaY+nS2q27vMbOz+l3mk85IFLI6EdtyDMfYnH1k
0aE4a13iEY7rXIKWef2EGTQN9JyjGRb8Qj/wye11HZ9d3kt/i7PxEFq8iQi0XwLLakZOXtW6WWo6
UJSEOOwJRnyVcCttgELaTTknWnEmGj1a9azFWfNe6bICZ3P5AO0OlxEhmz6CIV7wHH1M0cMIrFA3
J1OBRV4G8/2TF+ZN+3XHL1lqhnIMT1Zk+va/AlEH03ZqN/BfOqa255wb+OthNC317rnBKFxsrQuG
XshEOv626fvwsgGzioSszJAQIr3nET8+qBfSysCprXKoTOI0bvhwRM0A5VjTJYzwAR72duhIBjIx
I6Xj8Wo7iwEsJ1q1f3jziZsIFCopm61P7vurD3mwgl0HnULK/+znqz73a5gwPfnAflXAzPAby7vo
ArvvbaIKs27JphMbSP63ENw7zJRvWEX1/EnNj8WprHdor9YS+JjP0BgU3FK7jskWxqD/lppfTR+Y
FyUOie2SIg0+Q3PXS4I1DiDYZNJxvA5ST/JFV5WKaEMEJ1VKTFwEXWeDE9NXjr1kgiJANruJWiXZ
ezt/E8QhpCdwQ6xVNV3vexr69GB99Cjpc0S7aYUnzcT5tIoJmF652dgSlxfAq2LXwpo4KOrLiKxp
rCaTdFcybXtG1Hjprf/ik/vZnTv3OWSa1b/54IWp+kdmF6RW1Ec0+KEHL/Iqv7rSajHbVE7u26Yw
emJv7hYVsSJfEm/qnGvVgrF23Sx1+NqwE9LePrDOEEIZgX16INd78BhZJ8XAt/0cgZ4E2Vu46Xuy
PPkLiZ07Zo3O9eS0R/CbQL996h/8IqpEM9gO5KqxR6JawvgMtyy5/pMQPThowU6UuvuJbA56wWDU
PD13n15Cf8tJMhBZy/cTD1FRZqYP7DfSjvfk3WzATRKkMbB9GehCDGtjobPGz7yN6Pzol3J7MMPm
/nvcfBaemiMS/Sj3d2CNsJmCY9vCPqP89HXfda+HzmpLHoNg+lE0cQ38NVfit+sHTonZS0lzqmX4
FJwvCyNySJAscF2Lg24h/jha38YpW3tpjiZncdHR0u+HuEufGtWnc9gyd7b1834CfaPLrOAl0WyI
pj451iE0zssgzzTvWRuiKt3YDLzeYFfHrp+LPxSZxrgHS3eZ1sAGLpAF57JHSu4Zu3rcB6WsLhvR
8M3CCVN42zjEeFAnAT/p9ibMmlC8LIelA4bT2kK5tQeVIkLahZA+nVkniX2SYdxO7sgzAvBtS7UN
Jaf8TQ8SyMIM+N9yFj0p8LPHr1gNWL0/1R0Yly6aGxEuH7lxZ2v9TZtdzG8Kuvf/dncxkl044nzD
dRy6yUluGsLQxbXiuRd24zIG1Q9KCUG+7r68Ec9KZADfH4a8hAfGpV2GZj3XgHlm+CvAkB6sG+3/
kKHv+CQ2L/MHWPnI3DLKhezz/VqHj7dyGYRqmSiojWadJqveZ9c4xp0iX7bLeAnzRFBJA01/sT9G
itOvDZPSq9IooamHHR9neraglgCFPW56rHwaFMlnek+hP0gR54ol4v48t6789uqKfTw1KlVwUri6
RirIz3f7Tv03e4rviTCchDq/GokK+ny2nsyjSr2WvM89vkXPa+n8MrnYoNsyNOClER5DrSzAT5PI
/dEHZw08dO1e4JiUUyRK4mJW9ObetdBFR57lqVOxudAM387EACA3BxanphItV+K5wdz+dJM+rYGG
YGxx9j90VCQsFAa0y5DNzrPR5nrD/daHFyyDIPQ9S5+xATmCQrpR2S8bflUiwp1K+x5YElNSEtOI
DJ8tf+26aRcbnnFdBH2C1VhpZj+S9ax/6M677kPIrwj3sBNkg2ibByPEMCqEtk8IWo0LuMKnWcnB
by+fmi1Rth4Q9B3tEnM79es6CaI/Wd5JS4lcLb0Pu1il6RN+4q6Cutr5eHXP5oOCJFeuPutJHkDN
zFSSq+tBWgpfC0IG6fZe+07ywYRrhoId/7JKnGCpkgCNf9Ee1ATQehxeLhlOWJTQh7Mcu3nSBDEa
+4rzZa/4LpWTheMlDdtcK3tUqdz2d2HQct46May9w8/hr4jfMazP2vH9hqYtxG5ELb5kQcTVIhCu
WuaYTeAA3SyBPl8aR3R49B5UDOvdqKUcRJrFHflORxm6Ta4IjTy/T9uIX7GvVvA1gbVeQKwa5Z0t
7Excujfb8IHRo5MbvTDZKtwUN9K+vfZT3RwAqeB5GPaBJ7ppJmKCgOgecQ8H87ECl+psVQT3rQ6N
UrQLcbz0CPDnqE8QD7m1yjZ1aDFiuD3YCHjGyoPMhDouI7v45t5ez4Xi6QQhaH2XziDKB8BHsjMo
4apaD7rQD7rjwX7Y7eLZJClBVRx113a+hlY6tcR7Ad1TWKrLGe8lctvfdx0neiPgkFnWAGgdZG42
Nh9mKLRkH5pI8OIFRPZqdxrqp8ySAxGizZgH633ey/zNNe0wGPOGEIAqo+0U0eUViyD70AVM5wnl
S3fEMhlKC5dErcv6Fjahx7XJ2HsADXhTeq5u6ibPCzZg+aKUQbvq7jlPpHZcPDcRURlr1CwhiG+A
8Rsvb8Wwv6+h5PmHMXx02IfBgyyqZaT27RvgUDYfWsUaEXetr/uc/yDFI0JLUmLclcql5DWRBbZ8
R859wxDhzJcR2RTwSIlhKQd0QQ1pZNwYHWH1mDqZatLSsyCOf6OW6xPHvarxUjhiyAOo7vALiT9c
BQTaylys67WN0z02B4OZJZwLSL728nMSZ8UrcjOpooRwJ6NHZkigShtJNCemsocY6zm0p3cEbo37
bryc3iXoSYOLuLuPFdRs12BtArM5180flx/vvx6z/T4hIB3tR+HQW4gmQ9G470mvf1gVItQpFIMx
fMw1XGX164pFmNrNxid5nTwIVkpikcgmNB8mEUZJB8DhzqS/4Z/4QYtFW4fi6sdplu/Sh3shesvG
LlTGQAgu8HrmAX6WaMVDOPnL0PJoHfZ0faijgVfwBuV9wAPLWZn/kZZBouVJLw6CUgXoqXfMnDqx
vJlEyyWwaZzUPEeVj1dzsyRGsfn0Taf75o4g9SFiAS5VNq12jZVXuWGPVwktcuHfq+mmUGwlzN9G
GnZmdA/ZdIipj8w4Y9MUzsQwvPxEbVfXbvRXRKMfwYDHBQhNBdduTu+NXI8kn2DCgTKoCeg8UNxp
KpyiMsqchvINLg6GTLZ7WoSMfaOkCg4/1volAirGEElW2AM6p20SFNdLQkwWdkqpM0x8cbGHylcB
e8i36TZy+mKVWjOzO/soHSF1AyY9b3zB3QlCmxH/wiIa2e6mMDlXV5og0OZ34pilXNyZnZ9yeyBh
3iwwMvY43xKtlWxWAastlRRazGM3TIOLyApf88K3K9qKndyMTH+YEkwNIYG0qL4Rxh9HegSalCVu
ZeRn6CNz7aHCUPc8TGXmR8W+9QkcKGEDHnzAVG4OZ0kNQBClwvrLLjTzj0FANuPuOI3A+T4OiQrC
tiYvm1Pa6EnoEYvrwJ0uZpefiFOnj1oaUgW8KQhKDJCbh360wT61D+zd355GsmdsgRCZNWHOUNYu
40QCo8Vt9Gqs8ZuLFVNatoo85n6B9LNRuMYg7lJIsqPwPnkkstLde2FdIG8d3gTnhJRmJMCKukjw
4T4+/NLgOmaAPdadXFWSO5tzbj8+EqgzoOKuoLa72ZBo7Wb8JxdoIYm1DV3Dtj+kKHaAiUk3viQm
9hsJqpZxVCturaXBM/CnKsFlYJAGu8ihA5FKpSmhaxABcxs8B2BHRMmmY0KqCNSbXK4hdbHHbhNS
oEmdXw0pv/1QVv7eAKCnFa48d/gQBEOCxS5vrs5scFAwhJaeVZMfQN+MfnIibYAPAiNIu4rNaQTX
Ww/gkgDdxx+2ZwyhodYEiXxx6Odbd1hxW5XZIQpp35bSuETVMcGeVwiloBst3Z4rXlkVw+tboKhk
mMK3O3wegzR0aLDmhs/0mYLKzxDYZnptdcclZMIbf95q8DFUFnQjDIWlTNt6Q3tvP+SBkR16EOcd
63zFPAt8ycnnrrumaTv9+7cXjLXFXcuWtogiF4HdIVXeo74bYUBbj+WshlFWRhh0fzEoMOL8BKCA
FcmUm3YPFOtSR07O90mzK+V3sj9OO+0nmy+4fnAOo8PQGOOvdAhWMUV3f4TkPokwFIh23M6ENvrG
QRFbWjPIcv56Jx/HwaygbdHSoIVF5cUIUALSoV+ZM4Tsqrzsg2OFKgAe/dtDiu0Ca0VSHlICRgGA
OUj6BLOXtz7+apEuWXn2O396cxu9Q3qfuayUPCAJYm7JNZwMccNIBrwEOgu2ryVr/BRaOlaiN0DO
lszD0Q/pP2GgxMZmgWvhdqdMcq5B56FD6gs2CPO/j6oCb83TZAPW3s3W+x1jDMa1esqEW5VszS3W
luiuGhAhyI0PxtPS86VwZAMHlsrSTJleKajjMdRR0gzyY9wWsuMPxiJzrCAGh20/kMLzMpPdtUJq
I6K+iEem7YjLvli2FYxSzKCCruzlrAESPoUQD4XV8BGnEgdv4tLZ3S1qhZzz2ds+EViMe5XRwHpl
DcWHBFOU17YNRqVNu+tMpwfX49jMwko8MlFg5PmtgWI4vVMoV1YDinfcxO8NOi4Vbx7WiiXcDXcI
Yh26oOXh3msSjAMse73LfimQjZM0vOWUCSK2AFDsGAcwls6RcBjzP9tLIE9b5MhBmP3+iL1mVw4T
iLLVEuHEdVE1L+7IyI0lpCDUL+frVUdBnMv0pcLFb/GW4VIVo7UFJ2Y7nxfDRfTpKNKiJEyYqB7t
JAsFwLT6wpsP5xuBt1JJ1etvdapezcECUbGnL5ormQfpnjrrxdY1NXy8Lgl4ANWSeJ6PMrmBo7hN
hfW/j0oQSpoyJpXExddNqpWdudKNEGP8PigQGG1OzyM5ImJVngYngQXy3OWRtMf5i0WDb8czEpPF
u+7UTvUi7pyZQZzdIRbIMbOWcq2D0goF9EOOdUgq2q4ktIzx30GPKyPdpVhBKiaMHYfAKQBdErq1
oX5ZlkkF/YdKZjloQ+kJUjsfxGhx3l1pDdK766Zb7X76V9Md0rmFi0tkfb4BbB3u5J8BDTnwtYBp
+ZPMX4zjvFOLYgxRwUKtFrXZgS01TDCCW9sdmCXRDXCtwCYIokY2TMzWyiKDtySayrPy1eOrxRxB
ruXLXElITwemL1P8xACeMNL4vZZQJZQHfaUNycybnMwKImFMlPEOk+SbzmLqRon+nIv8xkQh4n8s
GyUNbjbJ5ZOOpcuwzBB6BUCLk9IvCVMQhRF2/hbQMm5GtGh3Vv9ZMGCPzROkxlRthDY9bWYHOrvx
37Va1IHOk6ge8T9x6PJkcSoRPiT4bRQvDyikGEa6znc0KTs6pj+7AiEmcjWtSshp8Vtrc8IsI9bL
ncDVvT/VGycnyYo1MTJI+NX1QU0/EhBRAaO/RlxZWh0WMr1H+4zBcV/wWOFvkt+gIR2VF9FuaTK5
uOhhr0piowlJ82FKWq7aW3Gn+Ehbu3eYbP9eogj4xdHp6ioqSmALKBtjrY3p12TkM/8TFkrwCikQ
MMGbCCe9tVgKOQe3XrSs6H44PnKiIOt8+23x/TPr5hyY4hf7Yd7ft/+Yco9HEqh6oADeQbkjoRA5
skreO89wZNwUy5gY2sXX//DZ2cpr3VjBus3l0Qqd5GSdwbslQ77AhkwtNrA5Cj4Grk6fNUI7RukQ
atBOBNRv+Eq7tBExNL52CH2dooIhTgcZ70K5DbnXi2l7a+U+hEXFl+TboR0JtoGhm/PxAoWxYtZH
DKRrX2KVt+zfwZB26tTX4rX+kXTx/Em6rKVC5clAdFqGLM67xNTnRBqtWZxYjqrZ8ORWBwF1ZKBb
p5KzgChJnIf447n7Eh0wC41WU39adB3aeywIx/O6zonx0jgqAfxlH3D1GBezo6OJYv1/N5tZdYSa
vVV0UwYr93sBeBcFeqY6XQ3K8q+BFaB8MtgJjxRS5bFeoXAOjL0n4C0pVuQ8jTFBvI+/RmNrOPSV
uVJp1TQriLpMC56o0XqDUNLjH5adydGpqOnhafwhYm4bOxBR4fQaIjhWjiIsUXd+fC8jaHpFjGGP
/2cl+NpED5/zLp2FMq0s91n+mGtHQIp/uAG3AzFjUuNhoH9Tlm7QdOkid5neauvN5ndE8baHENvM
f35Eg+LEdq93qBF1ufXXUGO1fO03bdNTVvDJKFrXBi8Ey/2dmj31r14kwQDgEtRD56OQiNzL4izf
Hj5uy3bXVpd7bNStvYvMKbY7x5uwZqFs1DgPGmYLatczjnnzKS4+wKzdF51OBPiXaLWL5m+kL/ab
NXhrEZf6HnDcPEQGqk50JlW9FyUFtWmduQeGXTmB1SFxlH7+XhIY+J6QIQQI3u8LASdzLRbUbafl
vYVhtP8VT3OF0ic41KruJ9GQbol7ygMi0y19szI5Y5C95c0U+hSJrOzA4wdEADGoaluwPRInJtSu
+vmvmGJPx3rvSk8lt81UZJjDvbya6tIELb0TaJVOt+G4knvy71HD1vF7KTZMHd819lWmLMiwoGEV
IsCI5tdoO7GvYHYBruY5A3rHqPQ0LYHL0R5xRcjB0gfXg5WiNAeyI5EtgZWlxq9xdcNapZjAbc5q
6Ap61OcssWZUefesJQxU5TYGTuKVbXpwRNiVgbhmBdtq0eYh1k2o8P6p43f8LxO01VZd9fdSHLrx
vVlMIMyc6xch7AKZovR6HPIKrUxYEh2YY43yFlhbYCcyI96Lcbb/H1Cxm+ldsrs7Vi20m4n32cbL
b/kpmeoiceaxs36QDmA9Djby3gguOFgcKZ/a8cyA+nv4Vqb8WxoxS8QUEDSzQnuA8YeAaqSe0Czu
Q/4SGcFpLfTZS6c4fp+M8wYucu1bJhze0VP4Hsn248bq7c7oAesae/bPivCgFPJ+bkOXcuWVLw5z
tGJ3iuP7bS30FqEalaloFCjkCQZTc8EHk6FNikGq4rLuISqTCTiFSIhPdWa8/Ehkdop6MhMFgNH7
uJZ9xjA3pw2pTwWkdcw/QyONAl2EjpnLtv6q1NwQpEcke7R57HmMJEPZkhqkAjHGB9KSyuQTNzyY
5Pr92ojR6yHKFYSoDXhw86x4YsCukNH7txcgOCr/QYD7Hd+s1GiHHQqNOYM10/PHYwoUKr6yGz+h
VesPV54TiLj8V0ejRgn8MalII5N38YF1x+wWDrk+fnfdUVIzI01lbdrafkNjwrSanC67/GbI2EPO
XCyG4PoRqquEJ2RNth5AItEit1SnhSAwZRpqKSZTAShobKAvnY/jmAaiZTp7GxRwBko2LnZPfrAH
6yjn0VCYItbLH8XToru3m/3zTB91bnWjXlEn2Dhq3RdZUVgFq22MlFPiXEZBlWTQPQ8W7g85f7ze
CIYaOsoWCxSEe1joq/0z6HLmxZ5jsg5UPL7tlQcke+ditoVI14KCkncjLlz5Jw3EXXUp0POwMcxJ
KIjx3aRQYHQTVBBoDQ0sjgdHlR6yXf0YBgkzaLiMW1GI1mPcXV69d3g0FmcGPqXPIt0VraXoiZbh
RHhJKraZUtX1tiEgWMqHl//yCRn5F2ZTop1ccN6TYS6Lb+XVI+OhAY1jOamaelHpodta8mz/AVap
gtprLRYS65H14UHXknX6Hb+oVItfnxOkAqu3COe8dqNC8iBMB441jRH8O1779BroV6sBaDJS7jv9
7w89HkGBiq69s137AGR6ODhMhUQGhTEic22y+MMaMT8hk8NygbB6d9zMa656LE+aWZJWsh7ZkJy8
jiiXjOtqgyVJxW5nbi+0JgQzyHn+/4ngE4LzHXUDMveK1jtSNU2Wmj/fh3kMm1ZfkhG33BGL0SQZ
347rDZ1S6601giklev8eE3Wc6KDLs94m1ZYTZxnkUJR2aPr9bJRUhfNuIzgdonPS3O1iqe32Cahg
QEiyQmgUrzoID+W2OOOuAsNJggzfDxQST9unw46QzttZMQDak9JnbZHFWsJ7lo9wUjL+DEWIHGAw
M4x7HiB+xhzzn+siPVBwJRrwQjQU6ygKT1f6zTecf0sUYJmu+cXx9ojSHfs1ZV4TzARKz5/ttZUw
9cZOw4stYV4sE6bDJ4l0coCACMlqDRNe+oajrXdZ1mQCwjjcRMOPhLnTunb8CNkXxtVdi649cLHh
pIB07UsUKb5eoqXFWXf4cLvajJhQsZtlwkXpX7qDAu8mneDDGdZveNpi9ycI6vx7o5DAAHm//den
uSDzwL56A2HbIieOUOfQQa98BcNHvay4RGCwIvKjaR8m8BROhob6WrDdnW5s/AbF/afvhU86o9FY
v1LdvuE2C6VYv4ZZu763LGWGh8DUg2y7OtXFSRnofSfysPT/EPmpuMVCdO+xh7HaSKNBO2zV+tzL
karC6rkRiDXwUibC/ipFN0XIB5VXrMe5kFF9G77VXZ9AJtS6AHBv/kUEMZ29SYhenZWdiDyuZKds
3UqnO2kMHKuHofd69g8xzGEbpAfdMQ8ZYe/SGfMMKOq0psN4E1skOllb0rAFj2CvEAApnm/56LrX
gRWif+wvn74MQQIHjQY3xs3/bQJj8h6cVdHxqKc+ELDMQbfXk/Kbs3fx6LLZRFE5orpGKYBNyNXT
01Ir/sFMOAfPxPyI8sisdVmvPzt9joad6Kik59IpHg+XTND840lHxx/KEZWCfgwLdXjm4c3EMKWR
a9j5mYwxJHsczS9s5GNzgcMSJf64HZeClXsxAaxOQIbby1FXmLgUUcLBJK3yQya/CJDcONJM7BGR
VVf2BBJ1w/cacXCUuMeipWPNr6mjx+omQqTduWOiHjyEi62FhVMfm7FUm8UUnscOSjJBy4rElcmg
2m5rIkq7owHsGzTURjLGJR10fc0oFUkrOFxMXj2p7wQYt/EO3UJ0bkvvOtPAz3Izl4lIA32+5Ova
s6etqWGpUuWbhK6ti2+DC6tKKdyKVJA/IVcRQ6WJQoSylZCD9jY7zOCv0lPcFzPODMQVeKtc5UJR
B8w9ROTaVdTDmEtD8VbkCQvLXfTSqWpsl2EwRw6GLzoeEi7kgipI1HtPZSgTRyOZdQf7MUYcsPCg
Y+0nhLFg3qMhM5G7nB5DwCOwsGPmMMXQCybBlF0qP5tF29k/5SxeD4ki6EVZyqh4OVBQ9Kc75Nx9
zuFcb3wXQNRr9glx15U75nTPCzHO9V+6l1DVP4bbkzkhHlKen81s7fkAW7N1chAkOFbN5HHvkpjg
Q7sCTG2U85UK9d/fy+yQUwV+EGuuNrBdy3w+sAqchwCK2fiZ+x7KUQ+bsa/7L8CTAHwLqamBB640
EZscNyJKJKi3Nx2EQpyF5tJejSH+TCMwckHkKNn3JPSR0pI3JB2W45Fx59QqRqmt/mCaZe6TQHOb
cRRv9c5PMDTxTjvsx4mpy+dPXvwSARxJIZZqmjIldqEDSr085ZGOyxsch1yRJkKb92VJcbOmw08/
PN+HmRj2hRY0w8JtdgI8Q4a6LCzfKqvyzh/X/g3qK84TVlGxcnDXgEuiILJ2IpyF1QVp5fDaAtNV
1SygL+Afq7cTAynOfHN+WQJrR/z9gFBG9zHsrY4Kbr2L6vfwDnsqpfHSnppWucSuRjLC0UVGnPXE
bvndhL+ycdUcsb7Kx3YA/yDSZBO+YiQwqbM1zDuk9T0+d1ZEFQvlqlKtQiXpUlGSKodoMoCOSzV9
XLJRN/q3btGSG7WUpvB6UJGiIQ1e79ITTKZvRJsGc4mZDpSoDCxNbGQ/X9vsK7YbqLdE8ZHJimzD
hYuVWdYerZxnyHc+znr8MURYjomLkiGIypFRVpsKvhxxFSLwa8PkmcPU3RCtBmjhw54VWHOzIhG7
uGVsaBa9ltQtlYsremyiqLYARRlKTHTe0DZT+8POiQ2c/EM0bLKoAnYwT4AoFeNNfjs4x0ng8UyC
+CkVo6B7ekO8+lDdQj0d5w2k7fRJFdwmWrJsdvgVs2X6curqhoottHG9WhL/QWVmnLiwpnI4ikJs
bAWSdPbJQYVRdGVvrzP0oHAUmkUtbvtTqOjaBJQTOWgeV99SJ0a1w63PA+zwdW4qtze9QNl7oTyf
kbNHAlAMC1VQFipMAK5UVffP0tbgqkcBJy5gmfug7J2DnAvzcgVdkJSB2h2ob0VuCWJB184Lf8Iw
lezOwigAni4Sh5bNULES+hLt2kdtJ5yvtsqSJlHAqlliNoaHR1WUOYRmms0Z4hCjH3YJPF0b0tCH
ZuxX6LMKPTy77U+4mAZNb/T1SPvLyH+vQpSAdiIZXV/fMsUzu8qQN6maCblssvrKPUAWzjx17Mjw
TAQ6d1HCXvMj6dcO8ebTgWYIdwUR3oj+oTQD7ItQ0rwc+mTBS9BgsCergTlsvZ5QKBevSJVtoIgO
+m6Ti0SqVeoDGUz7PSFwjHQhD5EHyZMb1mEg/pBzLeyRGtY6H787sXFj+dzjYLYFwFjOTVR23Npd
QIDIgjjAb/dMCeXIMQR6isCCJTP/dp7lzeGitDNuiBhq9CZR4/27K4ahk6jjvw957EkPPIdBpyud
WLBTR7ZCuWpRtt+VVnlqXIoo2kezkzppXdsBXaZ1kvgKFEHdB8ThRhnFOwlzS+YOwKKpMdfWl8CY
RDRnoxS/FrTtDHGX0LSrXkn+pIUyGvEsCjby/PLbX9OaErbKcpZcrThLnCDousL/GzLOuFCMNMMH
ZqmgrJ6bfsudImnmo+Rb7NzNdEeARFf5SG/r7/JkRciO0RFOkVysPxLeeohqh5sFMTcVEEm8dEav
ybmiIMX11pJHCQDwiHHLyHCXf8jc2eJrr+E5vn4OyNCq8ko51VFGZygND4ctU6IyMqT/WvsVHhI7
4Bmgim1klOJdLC4584Zkm/taB0oqFJg157DUvsuZjokQt89GXeItvoRvTYhf4zVVaOa1N4kmVR6V
HMyborkitWYsPE8qMwpKjj//2KgbKgFwDmyzGgNLp+ww7tC4zTmSZ41carTqQ57IAeZd0T9elNkL
3rorD9nCFo8+DfaQG6i8defghUxPVGQAAudlQXNnB6jQF5Srz9LawPldaNHaNz3g/nK0fgoLycuY
DAvzj/eaRQnGiF9/F08+qzJdvBaWjo0/ei3OIcukUZIeU5mW1zETCZchsNVOKZDW6yxgKryQ8R95
V1O4xY+NUx6PLG4vljMKGeuLqIS1zJh5mvYiqhqAp82CsDKGQrI0YP9vS9ixJOXe+IJBNIA/W95q
7YoxGcg6eIAM+c4YIpMuqTdvwjWzYQxopQ/ilkp7ZDgeplk5YsJMEi+1x0ixzJcW45h5WMR0Wsjm
9SuKgfavuA+bZ7FQ1dzul1mKAzBLohKSwN4B93d6hNLySeEg7cXx3ogv3z+I3AccA16PoywCMtlg
sgljcG6d5ts8wbEsk/L9VZIA7LpgwsTqosEdLrCh3buFECQ8id1OPXEZ0DJIf4S2zDWN2Ptrfj3o
fXr+MuLvpfM19VkJVnvuPuGg+QC+g+LsvbHikGFtM82VTTv9HmhAPMa5NgraCAnhIfJd9RfU7wNL
6C7V08DsSNrVolHAyXzdsQ2ppscI+HXi08aegMGvLBEXLu5yX36riYTrzc49Ey5XmhunKVSGO3Nd
q2WtaDZJw+w/76uuXzHr4s1sA5rEO+7awCGwhfkBMDK9u9C60iYsmZ4qLOCm+xQjG2jD3cWlRwmg
EQYzSqVE4wo4f1bxg9tvaZa2MSUsW/cFnOB9DWCXrqgVp4vYI4R0m/JTca7CEjfHUjZ3tQ9GIxJX
lJqputry+bCrmI4zxy3jjkP0wO8FNao+k+kYroMzeQgQb32ctKBnhsxMRyM/Y2JcPbQJadS4NVtd
gt7Gul8FLlsyChp/yHwOYmUKVbQyhdfgMt8PchKaZtdlYCAfbKGAAYuFHB4HqbDM0ncyaU9cBvdQ
GWhZyIEaATIDHjp6kjDBhtd8u7CEHHktEjA8V8hcNCEvO4mS0tAZTIajuCHrm1T8haYvn0CyvLeh
2AeK9E6bn1RLBZysUG0mUfmU/pfaJyo5q/hXA7y5S0zuym9Z1PQ1LlE2fsw33BW4oLeP4fg6PK6q
sJRC/4qsD9xALO1Irp82W/8UFV+sm236c1g3mSjPZaAGghqJgqb7rjqHGu8UEjd8YhsPVyc3mJ1g
lOpGDXcgHTb3aYag8DnArhUI8/lzPnhEdwbUWVnQOHEz48qYCxUtDHp5i1iaOkRV/noC1/kAoOUz
atHTwMdymphSGhIV+5r50kuLqqM4sTH663ZUP+appGQFlg9J/+qsVIKAr6ER/qU89nKx1mFLU5VZ
/ObOmKTNDB+ejjmkVfVdfHFQ/+wL+IVi0VtmLdkNiBibI8mpnoQ70yVvlsMBt6dMyhhJoEYBGfQL
+xZZusg/M8xu6xfH6eofY1RxbDilvQHHdU6v182O/T2h58fv8RPkbKHIP0YoBOjFHsO2S3UTOUeH
9lH1Os/WV3aNrB17aznV3ofybKp3REWib9HR1DD+5hNt5jKyiLUxyBJohqhlXFO6EOevMUeS0QEc
1d2XVHVpqxRhHes9BCrml7ahcc8DtsNqrOIqfCpHkXAB8eB1EbcIfFXCwnrU6efaewUzH9FW/iIc
yFkWk9c1G60oNRt2xhssAx3SZm4l8SZIWphMJVGs6owtwC0+UoiA8NB8/y8XpIm1UQT2Z6nYFgbr
5zanHmI/sW7WKhy7JD2Yojr8OBz+9cVktsuRaPnL6wcQW97zL/u3E++/oDESoqUvzk+49Tr64scU
4JJR10pIJ2eVEj0y+4rjoHaRZyzrxENBYuXBInYUNC9yHPTN8d9O/Ngm+ux4AiC7vMJsN8wR+4DF
CyStjfCzDTnP09I1injkytQyCsRWIJzT4StdvZATJCKKrwz+XrIGcApJ4zfs3APubmIhWg0d9qNu
NljBGmDFkV1yJRIr9k7WW5O1mnCsbqB+VKU0tOQtaHG7YR5kiB6KPH/dYPs5mrOYVT2VvYBdk3Hq
U+XaVADoC0F11J08aH6ZN6VnHlkx8WJjqeLpHIVrTwckdHRvcO2xTqqMB22smUfoXQPS+aV/l9WM
KzAM3nlLnrLjJwRA7d0cOVaR3e6wz0wybDdfsTyrEZpL6lBpdEJkn05ELgGd2LYFEi/FhG9lSY2g
OyD0Cf3upL18NtOD+LmdPnU1Cby5V/YFKBmjj353kxq9GhFQi/TftZhU9zfpbM5Yrw+W4MGEBkbP
yFQYxbT1VlP9qE0OYvWCDKBlM4MlWp+/OpGIVn8528bNykGDKriUnRKu97XlwGSO2RxflPsncUNa
BWUZ959yUlHGplsqkggChtgM8eK4I7QLZWB2vpOGvKBOvZSjzccBAAjZnqdfvX3919qT3Jz2DMmI
owgWwFFEuYebhI5ZnYa8ai/SSh9MoDeN1y8weD3L3Xtb9nyZzYqLYr7/Ujaw+cusItW6quoH/8ex
TajCm8W4LWZmfY7vINJJI2Gs2OYItle6dZZ31X57XHZty+p/366A5CCCThMR2A0lXLY8TbgAPW2s
FUBkF4E/HbT8oSXp/kuqw3ojUUe/8o0E/2Le9B/ChvamWlNJ1aUDl9BGK0PSm32O87j/T8FkRcC7
hwW+UxIOFfXPO/7lBO+nlqwz7yko6g2YgpHyIhq4UnCWrTlj685HjovUJaRYJycN/D+F1w/KJ290
URtVaoPtta9AYB4+BLWGQtDXNxJgVe6QskAyagm0g8dJobNBEbS2BCykCGUmS4mt+T0U5yvDJZkR
NEYo6t3cadr2+su+423svizU4bul7uidshP8+dZ/dQtkAXHQhpgFXjba+U801+/Ej+A8tNpnlovd
e4O3zYueqE4P5GvKJjMnt3u73t0PJbk2OyhKQL9/TsWxuc29t8+VH8CoY+ZHID06uQJF03cU/lF8
WzFMs7pYP/giDl50CckEzPkCGF6oNt3s4bKzPYJHLvobIalpfUmx/q2Aldhmabj8Erw8Zj8e/30W
zzfzsTmir0itAecwdamVI9cIr++HehwpOthaurExIz+2rz1pfFdDPZdIco7S10baPM77YGrope32
e78ebDp8jF5ZPbiOSDMLWgkMPzrco8qjytXu1mYsDzdCjGaKox92R2uuxi5heHk+Uyu6chUI0gAG
3V6OLSCO9SqzWSiyMcvCB5AezAA4kQtSZPinQ+6gn0YzyQ1FdAPmTIcxHTvA+3shqUDGYeLmoO/h
8ye7/My9TrFUdSFQWD5kRat0QW3X8qlLPHhWYqT9hl/QDjEJyuHLV3UwZXie7BfRqFuZJmpwlzRE
AtoVOXIyAFeKBHpjLJyuIGvLdF8f9KOiPc27PD2hlUvWua0jHoP6eHup7yKy2sb18M9B8dvJMbfk
EP+54krzanCvh1onVQ6IqEOtooCLjjyF6oyNECHjlONjL4f0XwoqTfvbXvpGeiboLWnWhgLyUDAe
a/B39/kVgn0GpfANIxtdZhqH+HsRyh5MwF2eQYKEkwIvxDrnPVXknRA3Mby8CMjYXULgY/gY2kQ4
p+5qfy5yqfYcXDqHEvBrfDlDPjGoyrR8VJgNZGeIlp1zxBLwzBr0mm1SvlBopB1m8JBG6h5RRO9u
bthRMbweQnFJ32Wc8sEUfAD06E0nRRqBK5aOrFlm6PDK2YpGSfSFhaQEUr/LBWo4XcVWWtonn8dD
+/sShU3ivXFCIjriqZPqA7Z1no8ZvWh0ZMpoAMu3EZaIfd/ezS1fPfrdtlEgnZKQA8gZ0xp/cUow
uBRAWYO3BfIAJaJ/6hMAL/KIe++UYlIYr9TzZbKBlSw6UC4o0w7hMUGvkUa9Xymsgc6UECg040eA
kh1H7yFsXvj6u+N+vDsqmkUJAy1A5ziChpp/kQw3JP8XHHp2eqtBW9rGwNnfMk/QZXfkeZVHBBfa
V4RlqunVx5P+AXCh8OPzBxrtB3UJ6Z382B9eVOwgdpUU4hC3Gn0K40vPOfot47yxhjBzR967HIgf
eiwLe99uv0aOcWHPXhnF8GPP7fSfsVHZJsaTkrysW8fUwU7RVcP6M7M+dF8r3rFTY4OsE8QP/jlC
iywB1L2wSTIEN1pxyuWF3uQo3ob8JcgArkasqbhSFxtZ5k5OMKwQTm4ncE3UqYqS906U9oentK2t
QiOgOmxpA3I02r63uqAF/ipjLGDKWB5f9sG/k1z3KzXFB0F9mnSzbYzrmQETEWZ6H+6s+VsbbTc6
rylpos3SE9KWy8xv9gTKVzRlQn+QoQD2Xuek3r0hCl+KZ37AHrrhVGm0iWyJl8o/JYZ2mRKnSuPs
GTPoo9uwHptFSq0hQSHcIvGAQM8k096+twZW4U1jywoKJJ9ZhJtGdVVoLJfFm+h6YbB4FZjel7Nx
L+EjxbiJZzV9ysPR8Jd5c4GzI8Jwh3sQV418ym/4dRFT8JjcGB5DuakxWcb+UXULil5y3q9Ew0tz
tz3x/zulYxDsYV2hAKluU9olWd4HmFnPVeWhy0DIfTPoUWdlhqPo+Mi1WHpSSUC4+aghPKXk6HZx
ujPwr5Sv5DxZwS/tsPRHAb4+5jWPuUXUr7btz54y06DiHGpk1An+qb4Z60ZtmqjV3y8gznZ+wtbc
2F28XzZoxtJ8TXKEAKtwupxeIEw5LfYP0yNywHid2mAbCB8NgdzYlyzPTOKig7jS0kxkX4fN1Ksr
dWHG5rLGeBUSny0pA5BxGd7nCYaqhc1cyHzK94n7RibE+g1T/6tzOu03gavuvayRuM65kB/oTsJf
PUttKOL/HZam+PwRsIc9CcRAUW/a9W2wZ1ac1dMOsDvMr1iBLcRe9uuzwC3hC6x34tKejMXfFM11
DBrFq0rI+/q1HAhUa6+iwmBW0AVw7rrPqi+GLaH3hv0KjBrY/UzRhBO+vuSD+OqsGNYJFNRyT/o4
npE3kHcKifabBoDR35lzJldjqS3oRZr8wBo82kj8afeZ7rw+MJg9e6JF/8noIRS1YybZTwt53HqF
pf/tWfa+RiJ9kxmOsZV5I2CNqtsmAeAuy6VyrvWjMfyAmvs3Lswzy04LA/x4pbtwpEWM16geqziI
9CZo00h0rapIQ3UUOM6kQcJNGrSQ3JTXp2xZRGl+LwcBq9yY+IKbn9VUKr9q7nGoXGHncQRs7NwA
w+Axx66VN90790WG6tDlepmyz15J0KrDgvwsgTMrWYKEOUkYicwkMS+H/yOn6kT86vrDObqJ2Vuk
1IwZre6fucAk/Aqd5ZdKZwvemWzr6/NrO0BwhwETtTRj0jwdOhaDsoQlC8V/MPUPFYz4AqTNTEVD
NCz85ZKcv1Vit1sQBtkDydeC9zG50X0pPwKgsXyhEo2IqELsxuXO8fe1vmxNQ99VGZL1cF4IKIkC
zkTFe3doUAHDF83Z0thH99v/4O2m9j+WPlHarJtyBEzUYCOlnpJM1LvF4dU6KiAG+bWkHZltuIWD
ev+AtlKGiCuCaGiCvLXbnXBgY7WgFVIToCLCD3Nx3OEF8g0sLPZQ6E1Bi8eIPL6zRHI8MTYGlidv
dGDzFal48RWsV/qdpPdR/vLfyNPbqaSHcLsviXpamUcyB2kxZn5ZrERtSTvX06W+RS3cuTdwYXd4
mstKQgI+wk6Hr70AMsBB8pujPQT+ceu7p6p191S9rrrJZgCWfyLdABvmI15PAr7EzpVxxmr4P3KY
hZ80YOgZ7H8l+j8RskIBHpU0ejvMOf6y6gjWveSBDdajhvYwJdzB+Lr/wkL1jUgi17xA8an5B2eK
ptJVPzzl6IhFAYBiEwX2nmipToolKpFP8Z8/8cW2B38JJ3Ag9DGJpnrdvCBIpBARr9srrjvkHq7o
83CKMrw8ZRAuVGFUbEL8ZBMCcj22PLqQhndo6R6rr8tbN8hzgiLneb+AWGPT7T7KU69zSPGLHYXk
s/H7egkN2wnxMM/xXZlahzryp/oB9XHgUGBHafG54P8Hv7INGZlcWhotrMqIM+ywbn+nOVJY01tT
fH6qYfjDTZvD171cPK+i3ElRVIETsn7uPWBlr8Ci6GBSLyGw7NmmOtSEhstPwaDGuZ2DVSxdc1wo
YUj0zxqtqNIXUsEVzlxpDx/gVQg5IoSpkyGShWyope20bPl5QuceYjgVhTyOJJg709ZLgaIRIZRj
2x/1iMGmBIdrQEMhW7cO0ltTuQh9hnLsOjNFld1/6xqf2sVFCMnh1ntvVvqGDuDctgyIJK+wBoVI
YxZ3NIDwU/tQo/JcvbVzsLGensK+6EUHBwPFceTpoUrcEXMDKzBEGYZkxS0dcjf8bYKiktrQnwHx
WXjbQQ4zab4PDqnMhK7KRw/64vDI+2R/llzR3O6QV3S7DwFgOwotQJ2gLTm0WLtpRigaF8XZu8xt
nJ4y8dkCldBVonevegBbd1BS3kSR/XuRknPy1W3rR6XamL7cxkfbUkVdgaRTE7yfSE23OJ9OBowQ
xG3VqDfwOsbM9Dg4SX7VlphQvfbTzG19fMSKeQ9kHcKHXHJ1HwJH6v4L6JzvpIMNCwiwbqw3O5Lp
tV7DvtQWoDQm+2AKqRAydS19w7H4QW2AKL1ht/AsHf5u3/MdXz1SuiBXkBH3J1xq5Tyn+hl2u4EZ
3hCkGWlt5v211t1XRxIQG7wKwTyJzuKj8m8Ybfksu3+JgEIE04KiXU8q5y7aeL3LQNUARFMrDZZC
yesYtGCQ5VcdmAvhlzNUmbldLnzDYZemHyLAHQlmwYuQLSwzlPbyhVEpHIWTfHhbkb8yjVurletI
3q7ve/l7Ufx5XSbUsTQYddCyGc/2mduWVBKrHVRDaAhA39GV5TkGcEctW7xqp7SORLduCD/9BP+B
VI9z0gVvPcjuesGusGEK/EHwP47/duHBTbHhO6Wf6CW+BIdzYbLS5XTpGogk+SoQLvBifsgFvOk0
blyg+/9hpAQxuIehZMW4X4eL0XaKZM7qZLVRerxbaIIxZ8/aWObUVIDfUAwdgluGHZSOoqjCDWZh
u/r+2CK2YdtoD3Tn+9FGDx6m2ZTh7Ajasehaqf5d6Om0Z77p7m/7aZQ0Okp51VtgYIyR+UzkddcK
uHa30brjK47V/fGkTLMYyuRNlXjgXzCI9abr9N4qWIQ1aexQS3sjJ3/kUaHclFd7I2JgKpVGKUPb
BT8DQPb7oW2TyKCbCAxZ5EQPKN4GdqtDinFAub8apOVHeHTXGMN/HUXKGLRU+PNll83xhNKuabHD
qoMFfeRbNravsEYnDBSQl+PSUkvjKIARODrhSdS6rzMKWG5W2KE0yAW594uXPupjwWts2MFq8Ow5
SvLES+PFn5+PSFIR7ptkebilv2L8PTyt3Y1CbOF985MyyvH/N3rD2SAa+hpGPTtEdEQW2j3kJG7a
+LOjaByTcSgxEBITYeXTCdbox4VXMbfThkk3Fzs9blYq/wwXmlfCV7BRr6u8BC0F8At0+pfChfu0
wgxv4Cj7wEkiQxgvAJgDzJYDdushJMz7/AgNGTDZEIhbWFQiaYd9SsayAZhuXxRZEVlBbSYsKany
rVsnQmYUEd4xsfdfUqu5bYROidVH1RhEqeAvfqQEv20F0sDerWu8FESBIkrD300CxdDQyP85cr2r
VuVbWu5JmJKKsozJ0USt0vLpaBvEvdPRvpQIiQ1zgJRRQD4BtfXQSJTCjnR+GcYuVDBuEkeDGXfz
GQ0jXcC/2GQ6F+Kc30gcWCePfwhByXovKOqIUd8nf7Kw63wATaeoOrG7zHrl7vPy3580NBTbAsGz
3Bo7gZXQNAcw2470irF6B+kfYxbqLc5h0RKOIbgn3ic9/upezHnuEbrV3ou8lv3YbJOyRHNvcP71
6TWRpePoObPHiXbRhbc8pCF7/zNxgj8gUHmgsQVOh55UCDE//SeN/ACyqMAHbSYSvOeh55BSdzmD
nFrXz2HIruKVhWqiu/YpSHtaXVaVEOBcvH9193VoUb0WvyB/YANLm1YCqC8yz22kBoV0wlQ+eYAw
ck7rz4DX12aNg6L5rLkxkqN/vB3Sx4v/IfavT38sAbmsFMItR5mLNbZV0bpSVst3duwZf/kSIbX+
SdTAZvS8BzbeFkY85JwyLwVoG5W8leNeJr3T6AvWZAOajgGPQJyE6BJEBjmpKZPuKJ3uGR0G66Ns
RK4YTm6F3yOgeyQHNuKB+kTGlkO4xPZZVus3pTGOvi6qN+dBPtR8Aag4iKL5LVjNzAnKPv6hsIiX
3ZMKKADDpLrDPCajrYXuBMRS7WDi5YmBTifD7iuMpFvfltP07VxGK7SvvrF+9HCEIvh8NRRNmKj+
W6mSjtlXxMxUpKLXmaWEEJxqHd/c+YwfyIqwb+z0fZnbpypkLOar+nTvewRQc1aPZh4X5E3FQrFu
R7SQ6TUp6x9BjNPR6KKyssX83+ADNMAEzuAPmOfwECL7qBF8lzzyFrp4S33OJSM4FNauT7jycW5j
KKVlgSNrYi74elOB2n1KGw2d3naKQQPEpvC7ZELrta1pTOAFtITO6Z6ryv/U00cHik4eBOk8a7wv
uNGiu/bnL4euK/LtRIISdkNx2kFt9XTULeDWU51nb58BY+pnXq9U1+dg0QoQN9E6n0r+E8I+T700
pFCSfXbeiYWLMBoM76h5OiaV5Knj3Ltuq+VrQXzezWbarvkaUGhf+aNKc2VLyiKqhvmtkcTJApMy
NHPRQ4NRMrnhLHXCg658S1Mt5Ve3BmpwuZs4e4AcxwNXk8xE8CwVAmmEY09p8HJyOEUjkL/eIbmG
SxIlUm1Qx5arKJBPIZm5Ge9rWH7XXEZnBpvSi6PojNcSGVV8HGLjbeFyOaoU1xQXJdTx2ywx5GqP
rd7RCYD88Ys1D6lgRo++grjU9MKd7auLVuDUvYbQRlm1n3P5KJpOXFN2t8mvQyo3rUPdoDb5I6v1
mj9SLMaYASHS8cBT69Syzsyp8mT0WOOyDDuKw88RcaZ+SrDKpeijZmJl47g75Pu8/z2MB66ed0kh
ZzbyLWlwuLSXB8wbucPHEstDjLAUvcN4Yil76MUpwvHoJ3SD8PiJYesxQH9fA0c3T4UBuQWxb+Pp
hNRZkoPQBlbOnnV8RTRUBPWSd2vQ9B+au35V6kVGxQXGHJtVhOsSYuWuXj8iNf55f/d9Q6oSq0nf
DP73AYlmy9a8s4AFh+WbX0pBhjO2yekTUdPw3TXS7bbipMywWKT1ldbKIFvRQ3mm3L8gJpu5qz2K
QCfushXKlrBHkaM0iIn6VjM2n2lGSBMvsFNRiPJc6n6lzB6tmxV4PA2Lcb6Uw2HekU+itf+6OgF/
FOmvLlxQhwulLs+sMqCH1JjNkh13k+torQIsnUp46HDaZ/+s4LuIDJy9vhGBiU54aw13ljHPun8O
tHtv36cPtJDXogGyFPqm/fcXGdnkxfWL6zHt9VL91mzMYXokenWItHY22Ll4BVip7Njyq1Nlai02
gDZNuNqxf6U8zcr6M4R1iDi61PNd2Nyt4iOeVE/OMsn1gQkL+ixkjnhzfmq1sLIAEVxl7bYQV9Qd
26o81hiGpAydeqnxiVLtezobuTa13u2BOKZGF+QPzGJdWn11bYpBe5JYaKYeE0XB4JDVB9NaID2X
yn2cWfBZPOwrn1gNu9NfBccbFSanZqozi6yinX73SE3+1d3aAAD1xxWiBpfOVDFeLLGp6o4BUd7+
x9tLHbViWQNLX6dtekVKh2n/SQLquIozEAdnpVyJRbWkFkFXc6pdgG3Qz4st0RDatzTI4SfUctsb
gHchW+fq4ST9Id+s5b0HdIJjPUtYxOyiZmfC0lcyqKlEXAimK6ycNvgGQqZBNaVaERBbhj9wkT+j
hz8U6aNpk7VU4bI8gQ+TB6vvP9NQ0qH+jE/6m5OIGUNDxXrFth4EDbh3PpGSE2mWSy4JyUnU5C6x
VJ0xzKDv4vulo66zN/XAYxjj+97tNGW7zX8sz1u2kzUEHnzb0TugVxuqsl9b90FQCOwtlof8gR+A
CSsm+Pr9FbpsXAQ9J3SjUVC56vD9JB7W/m5CNoNVpBmjGQCkVmadg0unrcIpF6YwaqworfNpTvsP
3nRlLCK4P8nx+vtg8ysxkrY76/Y2SDAM9OqSA20+ffBnIJuDN0xKfNvAsVugO2/NiOjjpwhEAFHG
qwpJ0nVyfdgeIoArXPacE25pQ2dNVBt2V85cjPNAya3W+PMVnPNShPuhlRc8miw/7ekTLd+e6Niq
ZpNElRSvmXM0aPyvgvc/qLVlg5qLddw0lhN8EwxplOxIReHUIKd7TJjA8SxXdXRbWKOyu4K7UgZR
x4kJuZ0WcjWNWRh5P1OQxjExXGW3SJSeZvbAsIRFL2c20828dFjsg/NKuUV9/y07As/CyfzHnzC1
ChQd5ivOVt1u41h9yV21rBf2LfFooDQQ7+ltGh2oyQF6vxHBB9UyHK/hbT0iMaa2gMqeEeami3mR
SRDb3MpB3Nt/cBygprlAAMazUbNDl0V06u97NtouFQiZliU8dxITxJfEKSvttEL3HMBYMSQHNhTP
ijmY/J6L6VcGoMoW2FMjORDYVnWkRXIv2QkIFd4jh6MkOPdAPWlLs2h6sHFauJ9QXJ67EladiFcy
vsGZ4P+bufEZpRQMmf7H0Fo0+MzInXgq8YWB19T2Iv/0+Z8A5lyKUblJ91nAbBmvyC1h3RXqOqxe
LCqnYH5OXUMORz2jcSo6Tq/3xTGfOegEK7p7M0YTCbWJpUKnzsi15Xk154ZKDCDJbSpWHjuGZ0BN
uxW+rXTpnc91Tqh/6tua4CgQivDPy/z24cSSTbwfJvKS17xDRWjegHJZoZ7dryn0Dk0ECWqCiizJ
xY7escT2cxgWIPsGXf7c50CXayR1fhVa4yodzIOQO+5xpoeEBXrY7vRbXLK5w7eHbyWcJMme2MNl
W0PL4leac9bRzFwwHjzLr1RnA1wVGAL2VjKnSP4fo1KF9SuDl3eDc9o3iRyYumkmmwmABIfRo4uw
cRKFXg6RasuYmM5xTT0coRAqgjbI8XZGd1O98ld7RFcXzcA2IxvrPwev5H3q4c9mXIaGBzd3o7A0
jMCO8N5hSKd92gAj4tR6mLVuxD09a1MTzg+iSb1g83YEj6lU2TaeAl2NvD1NmnbYs6Ah5o4klQJn
mHH8eRApkiEDUe4h+aZbKKCS76OFvbKB+Pp4k0xEEZnQmR2Pugzm2l8DDtUXI3tSxGLJe+H6mJoK
Ov5P8y1YUePUqKgPo682uoMJcQkEQTOeORbmCYNc9y3Alw6TguElQUY6JWzvdZAXljpA+L+PCQrK
GPq3x93/OvRQ8IgqeuAA0yap926l405Liq0oluOxhdjdBpwpe8jDU1o12ITTkqFXzGhA6mrh2Qbt
aeXoP9l/kgMPF3xcHyk47waxoGnH4KhYDAyk+dF2Gj5XDBlchgSUVq8stpm+gHosdCce6xrTjkil
jGfXn+oi9Tl3zck+RPmtiLT4A0C2K0aa80/0nQVOZx80YEELrcYe5QKbjmwO1MC94PydMNIwaVik
qR56a1VljIAUfnS7OUAu/fKeplzxSl9A8oVZB30Qi970Bs/6bNv+sFw+nCstc6sgRMKG6cjjTreX
Mm61OSzTARO9IfqqmHQtoNhkBLFsa81bTj1WUrAJTRx7Wcglj2T389V/urNjhoPDSdpyxneWgtJE
AFm8oUsfKJaqGlrI6OmUaofrdPCXv4mgZ1swzxXWnqcCS1GzS4FHOK8YEMoP2KLjB7gSNiQR2PBo
FYrutPoe7/be5RuXBoN+26uxvLhDB3KWIZghabFt9XKgk2LtP0LRXJqYA/EfloMw27MWN9rSvOAl
umAeHC9JVhaETC2h6ZTXkK219yPnKd75V9DS0HyVtK9S7tWXSffmICi6CGfmvfaPBiu1W0WTKh2N
hqoIgVOk2C1MB3uuTmHa3i540LsHgB5fSfyFCBpjJ0h1m1GT0/SYvw7FDF16q0NfLmF0AsrdLEzo
ByCs+pztWu37cRwkVPQuYAtNFqGm662srhn95uDHoxSMsyeJxjYKAsxBRe3wlXuOckNpdEnV2xgM
WFoF/8XAVMxgYKElfVZRA9EpUIVe19sevOf3G5qKfOfMlrC+ZMZ5dR4IUL4oocgn0dQipWgPbE+8
VCQiGRrha4ow+mItIv1UNU2g0bGDuZXvp0GblEix7ZiUKFZ3mJAQvMB0ws39WxTQfOry+sNnZ902
MiVhQozSMfXZU4lVEudD4GPjDTHtpl2Ev70uZ0SFI16zjZToSDkdwtObkhjgaY7+nYVipFKnCJXI
2zw3ZhKb890M1Pr99Umbang0/CQyuVdOnQdxlWN5vA+Q9hhvJy3g+rAVjcxu2YpHkyZNkNpsUSNJ
/hYHtn/7Xi+g8OyU8s3xd8+PbqlwiqgSWWDoQ8ijF1ZIznWwR+tNe3/h6fhesdysx8xF628BdE2W
d5ZWL1+sax/80upS5EMMwmRXTijwOdZ/UzTbtiuBTup4lJcdWwnco0pdhJ0XnanEIEHU3Dx8PD1K
AO2xrRcZP41BuJG0H609Xh0VphkPkkADLkbxhTNYKpuyvhieezPEh9jQa8HT19BYvENnVkVV+X8E
nD9GbY2kmkHmpurlkbTaMWyy3hJX04yIpg6SIQArpbX4r41ky0QmtG8pAv6nGP8x3DVeC/CXbxOp
hFuGxoVmeKlpcuO6GVhwoa3MKBE+YKu1TLpDHznKkEH0Wxz99GrD9erXGBuSf1ZqK2Du5/78ln+7
lYkF/xcqCdftM9hdehQd7H4Cm/gPz0ZEtNRLxuZkUDFbyy5iQ2XtQEaK/Y2nA0SobDZO80gTLf/J
ehYXn+NMvwom5hbiodRBjUqge7F93HQ5qbd9LP6+cf15eE6JqwODfFJ2+6HYNDgYmXil0uJxHTV0
JCzpN3rba7GYlsGnWIvJEeE3EU6qZIkvqFkaigt6kyxxCBezQsOppBAcN22i48lX3XGx+11zj5Eh
iDQ+PDaBLnfL+ThFJnMUtuaPVOxwHLwIPK+po+/UufRHFN50ANd3FcqcZnB+uxFjbaVSCox14PVP
BbpQQcZBUmObBCilJcei2oLKJX159iEh+Th3TwfAJwUbg+zwHr8uUwMDDJ0l/qyz7q9pCbiFa7m4
6MqOtwWZHUiLyT6x0R164p1M8McJ0EZ4cZTKisXkzYOkDxknEm2Iv+6EZLKrNghc9hTJX7zVeCi9
WLAPSwntZZ2zlmnmgKKgIkGqETdnALY/d+W7Yu20uj+McoVgHpB5YjHYjgJlDdosXu69swySTug8
GEjctdNuVdm1g//3YfRIkMj+KMFWDCZMewivM0ml6CLYu/LfIKrKAz1boyFAdpT4XingqKwdXvNm
wHan942dyh0I34t4g2pNwQOaE0AyQE6RRQofby54Zc8znfPIoaPawedw+WM4szPOaRn7cmPLrXqU
PU1MvU89Cl06Or8Klrz0sXcqZrO3wtN27TnM+Tb8L1deamK96f6nkrk6LC6VCsbeXmMXHpu+T2iu
XWK9FwqzSyn7EAUpUAie1Ec8ZW68yZ/bvHp0lAJvIq+Ginjgvs5fX2oHvl7yokXPCsOJ3ZuJFiYJ
73ksMvyTJFcrF/XW/XWaNToUq6fucDxeAsnUgbZQssEpoddc0Ql4n7jf6n2S6Xyp9nQkL9NdVE+J
/AbUFtOh1dTrsXQetJavXTfGTFzMS+bT83UbK1d0nHj4iZfnZMFEZiI/YQBNTsiXEnxaA+TzAUJx
jOdHDuyWgN0XOLaTYi13NroY3snmMdgki74XSHTu4LypVtNZeT5B9hggUztQr8VC6tWID3zqZMMg
+TkscOFS65EMfYlVrMeWw/hMWAvzC2Vl/uPKukiIe5rGfWG0q6OTz+NtLim8dCiqhJ3PqPxzwr5K
a1xQUUB79lPsgkM4ZhejEpQcj5dM4e6BooII3qfvb27xH6FoLNQbOGPwVwjeyftdZIT7GsAdKjXd
zw7ckFR7wN3MHZVuFjpBJEdWgc0JijUdC7+NWjVnXZGy6rUmfNWpu6p2xaGZvCPFLXMoVNGLe4KM
wZ78E7EHei/iFTdQR23ZZwreQj5usoWiYFJQ5s7b2qVvhCqmpUiSkBOyl56wOaQfy0rjI9Kv1V8K
a0/l/QFXOucaD4uyUPys6ktXIcVakZ1qxTVDGoRLFG/wKaucgx6hCtKT8zrHJqLzXfNxcaUf3TpO
WvC6zv5+1N8ZlF6Tv3lSUA6hSwdtik4WpjScnc7L2QF6h5sNQv3XFOGyTr9kmw4wyOdZkfCUpHIJ
5RkP4BxsteQZbbn9vqFxvXUJ+DJYyNL4jjt9LL4UK5LjoGGicYObNOdWXsd6eBaDFTL8EWb+10Z9
QJzmWKgvJitBrjhjIYBLwycWEspm1qYdcYaSOCp2lsaaIuDklN/zJwJfXrb/KG1RUKB/0NisSIlf
xn5KceFXudEig3Zq+vDVkLoi2diBWk2njsaFDTtmPP++0wXugQ6fOr+cr53haw7/GIQ5odnHbWVs
qQkFnEObW4UxlY0dNVghUyAFzzcMxfD2krIdxJbw/IcfRDXoS4BAC8FFG6ZY9WaTWsHFs/Izn7f9
eU6VBbet/6uisE5ULu9wIXYHfps0ybRZKSLnkU2ncYhuYlES+CI1qWV3fER0mwhhDtGkIpL4ke4C
Er0ov8o77jeTQbzQ5KfxswUMesje69duXmvVCOCLJAiE9NSuL9UqPpJ7HFfDuUUQU8jV85GKsEHL
BRoDJF7HzvqOH1xzaO79VyXhQJXRW6RrQLIdGdDcReU4N8GxK9l13z0aJTKgvoX+e6r8E2BWuv+h
Xy/PpFQNPbsY0s48l+YC0EL33ym+rcrW7yQTVpdeGj5lNAoenUYOaZ2DndpvwsGgrIZ5OznVxnNm
57HlizG/A0QShAZgL8BqVKI+1GGZIl21dKnIyFWDu0aZTsARsbc4FAy4ZyfbQIGKNbozEH/PsHPo
dMT09ucc5t+XjVfoRBtH4tbQ+CIzOBV/Ui/imVPcSUxLvmIHHvooWREi5yzrqibQgQ7c5lEIayPy
KZuS9gXZ6xRfGrWy+EFyiVHKIutQ2eA14+MuWBNQCoHYNbbnNazwqrJdsIT7f/Xb4woXOe4Xma2f
HezWxZ7ay9jIffOhQ93QewDQxpSl3MPmhH8grwbDKeV7WBlNEWnts2i12yr8futVbMv390k4XvN1
pHYAJgdbi0ctT2VlvJjNkODQqya2alkbN84nOucNHfjeWPCWG8nq8vF7Z8urfMEjHSzaB0VuWGyh
1/mKa9lyo8wdX5FzqKEeS9nMh+qpBzr641yVb3/YV9Kl4FYbfUSbz1QwTSrRSFIuuWKz19a7bt46
5Xwy2DgmI2MVrMA5xi1OGFdlfxo2xibCBsVODlVi4UX69w5RTkYcB6Opa/7pCjGF6z7VtuHxDLIQ
tHpDRMB12Y07o7lGTKYP1sECzDM6gaptNlnj32aSJzJBD6b1HzZAyqjEQSiuTzea72wB3tmc6QVT
JxfpAxL5OJfQHbx1uXHoQqeVJp/JyIgajg6XHjIhaqj4ytra2c6W9b0wqC5yeDC5mpbdy4idxPx7
1CxkmMYETrnRlg/mm9hwGpntP8v1d0DayJGHV0xabyQ6I0sqLTCx9t3OcfzriZ3gbNYH9QMEMXyy
D6UKJfOZ8TT6kqsaA/YXZ6xmw+qxUTi8mDetI8nlEMDndeRKWYgGI0MB78Mj4yH5cW7UDLFJozbG
LbTBaxHYBHAloZgFIUW28pmGafV3Vgm1PMzNqQEEY8QhdEm+fMb3rvnECC/tHtH0A2crtDwYqO0m
CHISlCALqc018iNcW5U9yIQyj6aQ6DrH6Z4usI/zRFWRsQVBlMcuBl8yZw3nyyKVujUFLXf+JX7b
m9KPITEOXqahpbCoGhUEfCU4E27GEfC7Bi95vaDbwffITTGvOGg0eQG7v1gb/9dItwHu6690WOJa
XcWQKvGhxJsAOwYLWB4BKyrI3xe+nA+kzlvU0HFEsprl6knMkRvIh70KM4qs95OW/zyOg/F5qDro
WjMH59G5ntlRD5eH65XzvkRZf5rwhiEtroZUQULdgnN9N12WKAP0wEeZaJdYXVJXUTJ7MxoWYNVN
JSsKIkCkswG6sUd+QDWzqJSs21wzUTEwnJLwUHjjimunf5pidUIMbuFZwt4bKrbsz6ZGaEVHCIVt
ZfLCO+1BZdAVl1QJH75cUuRJOt/nGTt/6J4wsnZGCve7S/z8yZdz1oOOGi56dzmt4u6/H6mWKU44
k6vRvaJR1jKWvK32qczvhvTdYIn9WwxjZF7r+EBIrf/3LqsHhju+ILcFUYmkEhyGjR4DOsSKOQ3d
wBdCcvHb0wdM/i/srXaEZhbJy+mkZrjsLhLliQ1utcA3atZghoWofjfKuR9xIFEhr1ZihuXZMvQx
lbjYDqyEz+Wo6lLdFX36nkOm9amVbsjaQjGljclmTXLPVHTbrYy2BVStLxWpJ1X58CMZkmD6yWnq
wgSf/ufr3/mJVNHwN4XQZP5ITWnXIHKYgyp7aJVO4F8tMtz4XHplrC3w9exuha+r0SMWLi7xPd6C
vNlleCF9mm509NFDFo6qR+edACdWRo6gXQOt8Jw/K7bteWs9gkGhbahRpcoddef7rgrpOfH3ZsT8
RrFvsZElfP4cqKsTvf6qmHECEjYLABHA7+0tAUlpmEizqUeH45keelvdSiEkmlbmyqkVYGlbXdK+
LTmhdxaRmOjf40zyykyPFV9+vx9MdIEMTtDNT41ZDIkrDPlln5rpWgQdZFt9kIEAyy85P4yDbDaq
QFpZV+FjBgzSRgW2c/I1fPMuBvauBfo/7F5kIKmHximnBNCL7cri8FUP4k4qKHal43R+o8FNsurp
JmRUGNp0IRoKhil+5xozh4lA0kW5I7pPc4zNtuL8N1erw2LAJdRFhZ2bnhVBtmRTLhSkpvDb3qDN
OplcAQgkvI4TptnBUM8F4aTMn2zkXPxDuAblngDIsI9xlu2DZnnA2RmtgCfmbFN2qKNIe2PWETKu
l14KktBiHoDYwzJd0KXBW72GRLhPSa0S+V/FdZx4L+HIsKc1x/MX8bJ1IEK6pS9eMbAVBRFIZmHW
nkp8Oz+ngvShECtsUqxzyAsknsBXY9CdT61MyPtXSLHSCxDGqLUuZlaMyOcmH0P7dB7jMba8nqhv
q9PRbChojGg+F0U6bChEYeWddW6PUXYIKt+bM8gtQetz4iswry0QWhh3cviW9J1MwmL+RDdFpf+C
dyvTEooZ7+5NIH3ujwrwGpCCRV8j9sFkCTZqbenvUXIT/cWnAEv7ERf2zDerZYyw81WHr/7GvQlZ
qdGDj7pGMb+47rvc6ELgeo+zj7aBVd66z3xRmJzC1ckc52maGkZHIzD7Sw7Dtm+WUih15sDXNI1K
qSHtw8oYvTl2qGlI0pWHZ5R+byyBupLuNtCFmeOcvN44bGazJ01D4Dx/2GC6shYig2h7q4qSTb8g
9W04ltp+jH09zb7GKQJ8je6X8mz5PjKobQ6a3dUUqFEKiVNIAcpJVZlXy9DaaRp2K9r84+Xrf0LT
araBfMrEz/XptpRl8m1C1elbpPUaQGSmyYr7Ja7KlDkIOyvJdVaA3epnqIG+LL7y6exG8UH4llR4
RUhyIdxAuAeKz9pD7+jTgdQwHzkzRusuOhzBc/GHEeCm9SrOfPaybY8jHHB10swKNNlWTQAKbPZ3
6bA6P7Wqk/tqcueboYl+Gr2ZUAFJowBHTwzrFu2L3QG8kinx53sm3ig5BbwH4ueSlbqXqL7DNaNE
Ys5DvBWRNK+G5yWnPQsiN50MKAArjAWUnvB6rO+3U4RuG0ly2+jF9lxi/R5EO+1tGT8FUQ2+1vfl
j2eqHigO22BsDD0JmG77VRTsWvTJbAgpgBmYmaf+6TdPTzxFvRVGQyOtTnJvlZ9uu4XjZmEYwPNY
Bc4MLUtVPU5IU4adMtg6XIEuoJxNhoBno+8wsaIrXy9HdUqzsb9DM9HGXqabeVleQQY39vgaR77C
9vOm1b3gSRwIQwhD1NQ0JJyKhoreLPsjg42Og8JIZUjTVqQJXaR3fORyW63sgtkjo9PjoXyw1nUr
hUAI9u9+hr6z8+awgmwiJrpgsqZED+OMio0cKvjw6tRR3drz9NmTKuHUV2S7329AHkFylFUPuunu
/YD+wwfs98Kxs49/yEtyZprmCH7v9F/04ZiQhMuKg0TkX6oV4VNSg8jS3Tq96i1bgfESDIlEir07
svPl4//4UhCCD86psaS1wEltIyRPnJaMVta+aY6P7l/ecmJPZtyIGaJ8Ks8zpCbi0Avd7BU0dWCH
Bff//68KAcQv7PG3wK0nX3/3WSVasG4SW2OcHFhMjyNr4JEuoUrKH3HMYpX3AB0BWoT8un2qrCsq
8rFFgowqOH6kenJX0q/3lZEPisykICObfTxxsPSCtTB+lQ+kDm8VegfWHNpDdzf2TMeu3o0QU/gz
obQZKOscwKR69tOYvKq68Bfa2TrlxFUzdyWBMu4juKNciTx5N9TlfHTZdv09O0JMeoXNsqmSgYv+
M/wA7qeFthsgMWgPjpZsaQFcMSzkw9q+bF7iVh+8DX1rFgZNZ0l0Bnf0qgIY2PdbmOIbLUehF/co
6szmwfB+HznBCWUEPv2qpH4OStJwewlTVf9lZeuy3e8xYg4gii57J5MOUYUz0aHtULW1CXAtOxtj
MFSaQbTNXTkMyD23hom4xjs2hT/jTL3Q2jF3Ib26KnsTdlQFE2M3RRF9S14rHA+aiDXmyeupI3K0
yATi9krZUQg7ImKByoWAOu6tkywvudH6Q1k5+3VWxu80e6QVZYhutXmXJRaBsDObxDvLvnvltr2/
1uKXTNX1Kup2pnxpSR3pNQb5wurxxckGEJwJl8XiDCRiopPNMNqKN0rVezFdKq+bz79Kk5QmRCWY
v/Sj3yy7tXWCja4YagwJjAu5ALQfCUG3DQxxoIRCpcJXCNw+TtbEkuF3WLcf7yXFJGCyqofgrFuj
pRc/R3j8R+nJfBSHRBtKl954vJFSVMuY2+0cs+4CGcAUu72Gq2SQs5PRfTcAiEKf2JaijsQH2W+5
Oh2++lDpaa6UnT8zRM1fXLB67iW1I7+0hh06UfU929OSVcvj/1bOVP04fnY7//+NP+D9sEO3XcGM
FbE+wky12MbtK1/bJf/hbVVvx6eHh/Dzw4RXd/dyq+SCg97GINVXxBHMSV3DH83IAHqUwh4bTocP
w6XoF1h9QJFabJRzxGrxaHttvFreyYQAFPJDvmenG8CAKSuume+PrLrTONV9eZF3c5JwraJUWpkh
H9N9d08YwGf64cF0xU/laJrdDCgciMA7/PVF/6EKGYxR/Q64PEsupfv7Jw29ybEhzHLaLKzm6Yg6
S9VPMUveOYCbcrfRgAjwB5uCu07JKnQ0Z5VdClD152bbOiAoWcnZbuIn2L0b8SK/Dtwbl8L041d/
kwVLmjqOPp9WLHg77LUwebNyUIPMBwW0Bgnuwo0Cbq+NNYhIhYFDG2O8ortsGMZoiE4Yc+6QKVyh
LR5/IqEpko4nwf4vLts3b/vLojj7Me2RnL29nabPVsaLQE2IuWqDqQLZPM/RzHE7Rq82QQwiKynJ
/QxBEo7qWMVo/EuI1raK5yeozMhjLkYx83qoGd4InJ9VFobjgfvwstuyd+YVWeQ77ax+JSLIiuUd
Wz8cYofyTRFLyaVlEXczlcOT1jlBhVuyX7kjUnFlhmVmgKthFaFHu5LOzeCTAdhgeX+EQO3fpzuK
VaO0iJ2AJKEFb81YmUXc9JOAX5Xdpq+e2z+Zc4kQUuowvBEY1JiTIyd+tlIMU1tL5Gio7MebbYqG
hvXx5v7VxODcqsEZ0Vo96KFZcPukGGa2uVRlMi3zTvFUj6HFEvFwMxRVKhTryXIKVYKHDlZ4SZqU
LDpxLROESlEGtX2H0yJ5U0sYnJZMAlLLJW3AXhGn3KIt6ZWZskQU/IAv6pIKhXc0En9GiGo0zjPb
J5k6udkW86LMDKiGKlkm2hd1xO2vyXzPv/DKDb9dgsv8QUlNx4SUB5avSqF9ym8KCRz/2D9DMe1J
snklQ7jMGxZxY43JgA7CTlydlWfX+gqVfwC6gfpWDWbHy6XkzqiKuxH8+//ojtujS9TXHhgUyE5s
kq4feVxJj65SLY2G18JSCWEnFCtZmZ+P8zq+pVs7MaUV2eZO3tpN+feeI4z3/0mkIJIKOmi8KQVF
dfFhHIziUu0lIlthQzOE3pwoCMQxjxahG/vRJf90H+PMrzB5Y1E1heZX3DTdmxJydYOiYUbBV3b2
sprGSkHVwLr2rSN8mmFMszV13umdLZptMZ+RUtXh54G1tEZQxyG2Otqku9Gz2JgQNfdraCOKJiri
QRPIIYcfXoCio6TrmljOCa+4dCrwA5RYw+0XMzZnTVQ6RfTj9fBIQTQJM6rdFbuOJfGxwGZvaMgR
Y2TGgrsqnXuBX3roi1i9ZlL1aMXNEXg8sI0crCbuqxUDNx/Qwil2Ce7zSpU7bisfEotL9+RPD2Fi
eBkIK0fz4RMD9t9y47Y6Tpkqjy8bkwGj1miJjjyMPrfHd22F42gBvffjuqLDEnY+QCOQAgaVVPmh
aXkGetFcEQswIzEel74tjaQl/SSsdE6Lx3BWqkMOoVV5uRMG5xo/4IJulnCVS5gQ4NbcmUVGdl00
ZW61kwNnzQHX/a45n/VdLhycYeXlTgH9oflrgvTfbQke/g52joeqi/DTXyVqxe4bc1EW9DPMg93A
AywDpa85z++30B2E8YrdLuwu5UEtAkWIi9I2bmiLGKfVMReJP1JZ7+wN3eHopeD8Cr0uyC0753R7
a+xW3z2rvwsLl4SoxLU2NrRbS03krzbMcdcX6BLxeNSO/2tVxx6v3YLC23b5mTTVr0YcXmeEC2WK
7zvViXuKcNj60At+bUdaNrxHuHYA8WSOGBdGXszNX7zQzF9fVScncM63TTiDb7nqMh9A95UQfBxb
MwnO6YIPbqftFbdJCv5IE76YnEzvX0xB8IxRF0RB+tLLD/tE3z0rUx/iYNsSOZFFpqNhHjgBRcOd
nDWvqh60yV1hjMuahtjB9zr0zF5lceo3KpOjr4iDbSDGpmrdCjaay/cViFaMAFS7HaQCDmpVbXRo
v/CT77L9yR3dllSk+FNJPAEsWlWceljl8cnM7Bku9OFt4FoMmGbUEsSpA42RxyI/vyTFegLZzf6j
u+ZqcHCKRz89KTQNj4V17tFm6YjQHignYatf2TqsezqZOWIeMRjNbINo7lafQ+1UdswDK/8qXg5e
MDMpbvY5lyF56N5t75by3HSOReSla0rh/R9+t+rzsgGvYZ9ynS1hnmmce8Z8eOMj7R+VnEepcmCS
/LijchBX/Fzh3YhJ7W8XQv0wZv0R9M4UGEhdaVyY13h1fTf10bCkMFH89Hz5FfkWSrIMqsH2bsoi
pWGOoXA1QSmxcBM2cM8/0I69ALSjDdzYuYK3TgLKdEZdOQSKlVGiqpsiX4IcP1PDJAAPHsTtbIuq
HOo8gO3r+1c0ceRAfzVll5nRmmQL7jev4R9k2/dT1UmfV6j6/7IA/k3hJn5lf2t/159nnTTpH7Yn
A7GUgP+UwfMlR+tXcV1MmJTBSR3d2lJdnPVaTJge8hvGCJPGb9Cr+nEoZjd+X3Cj63J2glkX3o7j
ErYG6thtFYpoE+Y1TTZC7LaFIqo1VOKMjqH2H3Db46QKhjiH4/ilVN5UGPO0uxmebUo/UPpK7wIA
l0f2ZdBW+5UJz2UuqsoLgSiudXfWmooiiVOcwb5TI4Q76hfqDD9iREaWPsN9E7Ls06RpAGaitDWZ
A0151N1yBhByG4B+b8mTZPHSGEqaOHtKkTdNy2nF1gWoJ6Jv9jXrto53a5W9Jdj2SuJsZEEmFo08
6KzFYIPtT1kX6jOw20s2Sxgwduwm3eTc0ngRB9qKycQcUlHWfuQeVXn+VVy7/AZwWGio7FlcOg4L
rcMcd0hnZKHLq26DIZ5dFDpEeX+N6vboq8A2i1l9GTk1WNDm1SDnRk5oyuG3fxfsiEZUPwS07qda
2Y9S8WuOQkPtrRjvLnJ1rzNwVdWFMXUXVwLKy3sbkXgDzMMHjm3BfepziMySeGvfUv1hAUV9I+g4
oZg+72zkGQPZcgdPpTqrzMHuBASIwqwFFClXH4Ovao4OlhTOl1niz0jxkXGPifURlz3Qxu0yTWvm
2TKKkFP3zorEZpqINydJXwUplnx11VYi6xyAGGqNHEQR4mCHomfwOPIzYXoTv3OCymJXexJtVQR7
GeGu8H8FOa88GMiv6b7g0Uf9TwDVpvP9M11r960VVE4noN31RtZYlKW9K2Mt0MvWnRxVLng/B7Xe
mWo/GcFVWvjLZpFW631FIzZ2kljC3XWdhwAp0ef3obEaGFzniANlUtV+QdoqS/nMBroe06SW7bx9
8hQ7+9hDCYe2JTATtngaqpE1rsvDf+T/G9yxd5t+0/x+hDICLf2C65jsPU8BdLTTAIaq7xvXzC1K
ChIO0mdBcQn9yWEn4CrbUXHBhtpWRiBUMiUpDaSYCUY+Zt6uIHwnnE/tv3Q50G/uu/rdAKQLUsZ7
JxmzQhhwQJJaPPJG2erUrnDl+zdZOajnxCj3Yz8+jFkAYsmHqbG9H5i7smeua8ZHdoIyatCE829Y
ACUwQXT7wlADF5eJyWAEHxWHqHdrYp9EeRLdxn6COAdTolVMZoEsznFGFk6GlYAToRt3VUbsjGtb
IN1xYND7CgbGfMzkynEg1FcZ3p8qd+eEFOMN4T1qS/1ibG4QXtGDXfuA+uzBuR60vopV1oiMktLC
C0pjZOUv62NfZCV6bWeJjCLqnbMyGVUA8WnszpGFxV9VLl6Rr3lFLzpCbWf9QIH8/vbNZ/F0KKoN
TIbkdoarBe0A/v1q4Qzxkb+z6TUpCDF17tJGAA0qnW1xTFLvFC9qjoTw2HZV/AJHaHd+SewRdhwM
cl4lLf2fSlImVYqFZFhJZsa/uT2VWjTS0sRq+9UsoQjyOok/8ISzx5g1OXo78MrXXhFf0uGTTNf0
WHkCJqYD5yQ4aKTgr1yoQD74TmH7yr/SzFzcLCkryNDlpA+/2WoKzsv31d/BiL45wOGy4EBEXyjt
WyHwk2RgMfLsgpuDM9gcL6Fh45dhwCND++Uvmt7aCAsehy4oXwxOZ9dQPFFt1LKeVjD4ZICYOYpT
KaEChqF3jwFoYX6pdfCm4/7KXodDq2D1d4LA+zFYjjfRRZLjUpx5VcQP+tKrG6Ws+zmLDwEQ57nM
5zJcFLw/1dhk9J4Y3vvOMovI7sSDTCUVjYIYsn4JjhpDUSb23fb20mJkavbSHl2k4NBFWws+C24u
6qV1wMsSjyMdItKMGjiDEPKrfW5rLdTqMgai49pLoBTrZCw4ATWBNeb/+3xJe/sCE9Cgjn5ii7na
Fp2w5Lb3MqM+EX0p9a3yQfN6tPQOjUjODsbdjaokR1XmRbP3Ha1UJ0GzWiXzDHWRqmN9vOq1BLDR
Jc2rQ5vFB0irGDCehWZf8uD2jfQ20X1uI8VcsvNmpRScy3yZgmETHdD5eyH88Nd0j6BZSDJG9VOR
gL6D4pcSV4hlorwkL6epkOTbnIv/M+vdy876DvIllpLkty58N30H/Du9Ry2kWz7IWgNZpQxscUAs
D2/+m5I9x65GVvMwdscyFdNXORV8p6/gm2DVToSx4O2J137I2LcMNxsXtgiLrOlny5NGjF5cJXi0
AwdQGE4Cf6Z8X17JokyjPOFGKqMxLC/1Ui8+hWba7BTZZhKdDQYaAh7mhpn4+quNMpj5+K7wYMcX
waLlunufQ+2FGN400/8dDSFFaKW1qIrwzhR/7e0RR33VFQZJxmBjn24hY6yjwmmJvFD5ipoYol1q
R1tvMGh/XQQCNVV05bD6ubb3zE5SYXbxtU47SEbrfOR5TBlBG5P1tYLf+vF4XdEOJpRwSgLBuOg/
AnXAJQ2EJoM3nHU3s9e5gle7glto9+CCcPUVzFcVn2zeoaLJyOy7sEiRkXdjTSbInOgmw7jx1EUj
e7TtPLzD6arv8zmub3OXFWd//Tt/m40zGwizg3yKkSkvjN/UgfeZLQRJY05U9nAzSNaNnpJ9gdAN
eUKwU3LFbTV4wWBNPclU2qAiR3JOdqQUgSfeQ30wJbkjkbKMfNg4X5oeaeJ5zH54WimCOV7L7mzm
FPMUYQzsx6tBG1ccUGYy7VBN+sTuLVz4CyFTrf4OkzqBWPE2vfFJmTi+Fn66hB1aol/X5lflsPb6
yk0Bmigo1gt8gdQWBVyldpXat1wIxZtwwwyg4RlCvtK+rCPdCwevt3c0q18+7gDyucEibUMujxi7
/SCF7VlfbHBRjkSaHzi0s5sZeQ8TICbbei+qosKTkKrNSfcpL+tPGOG8BpjjhrX1lV9GBamTOgG8
rFJlb53vD27A4Pdlen8mL1KXhamM68zP2tIxJq9Cg0vZB+WnKOQl8wY8jHYIAHtmdVyDr0fIWYg6
qhfkj9I3Ai93LEnGXvSxSVmT6n6eqgHp2GzBcv40L6tyRPfeaZb7GWYoRqsx92sPmoJ1eudLbgX3
TIp+hqJllfcyDxjKb8ptVP4nVoxXRmcXoZBbNBv/lE0ugSCs6CzYh4FQwvNsGiGHkb75LFZOAx9H
9vvEpNH2vp6g1QQOhNcd07WUbpPOV4U6VF5iYtHjnN66ewNKgNGbiI0AN4oqb2VfwsPO1Y/9kLmv
5VDiG046nhHiC2I2WwpADkM4m+PNgdcBW2HO34M1XV7Z4hHmstIxTAISSYKYKftKaVYUZCvnwOrL
R1+k4DCiI+TbVbTPM2r3ml+ecL/zlBkzSzYQuSxQ3SdAgk0xzrzWZX/dWZUlW2QhCdJP8MKcPke9
d20kr6pnfzwQTNN54t2bZnDmTMsNBlYidNlv21fw9TaOr1lTm8/YBvGA7ScAN6NxIDFZsf0jUSnt
8o4DuVyCrww2yQE/nhx6Ba/hgUHzu4AqIPq8fKV3/QmQoR7lpuFu6s3bt2DWf+9pDtcek7+Q5yJP
mjBQyXzLsmbx6M0GGQCXdqZuKfaGtaSzoqhblzEmlNO8SQ1rHD3kN0vPgqvFXqgBlfSFE5wr4k45
VXF6PFdEohBhuqxpDXkvpt0RrhCPZ9lDg19lw5Li/hC44+JLWo1XcnuW4QPHpNFIWJ0oeTeTldj7
LCeWcIoB5x6CaS4PWBtdUlKc4saLio+ADXSezwmcouVv0vF2r45l2ZGmGbc8VIKfBhOO1THc7KdP
ev4xxU/YWMFFFVzQv4jYvhQE+2SUFYcwd7N6i3/WBNDskRMqyuCV4hJNLehuBmzUHnhasrTl+HOV
fU+dzc4YkAKr1F3yskFAmx0CYSDtvzS4/3eQj+ZgDeAQiJRlAHgrW+jvkeDg0ikqSRlDHYfcuAc+
yYGRgINA/Fw5zCbkHJ1TwMsHu9Pn9/2nbm4jsSjbZZfF3MuIeKylyKEJr94MvbW/LQQlweFdG0Ch
t/QKkkN6DbUBCQ/pCz+ezLpG19J45xxKHusDxiZ3znCP3WbTpATh5tchPCOJ9jHirZmaRcEJVJTx
XH90SvumIofRC2ihzMeTQIfrMwTF/K0CXRN7/ob9WDT7Y2h19ioXHRou4MNa32dCgDlKVNq7gXQO
3zzvSEe7DU78BExykMZNvO/i9L+MushYNSvl62qmzMcGDzRzsg8SoKJZ9TpdRCg6FdOk2cptyRja
HtUHGJUvkdh+s1+CsRA1gnoLXZ+wJLbiXOeWeov8aWd5hQZmXyoODa+sUchqEmSEpnerzKRX0SVG
m7/JpzCDAOXC3POzOrZMbH7WfiUd742i3FJqq/nuTQkvUROvQZmL54pvSanjCqXWtmoy9XrjnUvd
RVh3acepYeGAowWx1oi/PyfduC1Fl3PL0D6bnHXWVV+PXVeLSi/tzd6d0DN4BqzT9W3tzq4KXmyV
kFmYMS3u5ndl0yY4kOyl9nsRmBPWbAoTvnltCsVZ/9XIwKiQ96Zge017U6G1DROHIcY3xwBQ2rGX
CR9q2gA39AlrfYKzxk+DUbpamC7rCBhIPfueoCnxd1uL1UHky98aP6+dKL3iceGJex1GQAGzjRiJ
ll79IetJmZfvscfdA71HMi0YpaQrLOARN7K4yZNwyIPsNSbC/mg4in8JI3uJwJr2Ia7BOiWKCeJu
o+AhwsFozwBVeo3IKOwOJr14Jkg93xVWbJDdhlCTyEgD/bIr5kWOVLCgDFGsZAkaseUM3Kba9NEF
Zlevjv3hAdD+7da3lS1FNQSpL2NtKEt3ltjrp3MHWsoNBAgR0zseoK/Sf2JdUOs/JTV6uzQ105yG
x+NPDXzlqU2Ag9ogbtw896VdqpQZVvt9aBuXM/GFTFCL0xt4h2jEsHQBiIZJ94nwrYdTXFAfHRE8
I7VseTDpW2CZWsHKSkcQa46ekXDElUgtSbvIqBLGfDbz8qQGptpILMEl5TexI8X+Y5WbDajwdGEh
qW9fSWX+eKPnKrw7I8rvKa6aRsrsT6Tr8eMbmdNOqwo9fRTIKYXGHkqI/nGr1TwO4T7IOpaEGQ9F
VulVJKlDWfXsxp2SPtX8HWc7DJI/WsBwvnMOzO3G0hjkoJS78/sucSNkVqWg2t+Pw6AlZ0BMDbMK
DUpqFECgpnlsTjzn1QqEQc5lmEG4J2iB+qhmJ4Ti1wfcHEALYyVhH/rwuuaJ/+Vlg+ST5KIEI+iy
BbbMlQ8wLIi4vMIOXKe3h2swSd3L29r8tNhF0EojGjmkJ8Y9zNw/zac0xZRZCigLE1ahY0pDZW+O
yix5K5LuvmSSuUik/NqKmC5uprvK4i06RpQnkIqMKf9r02oB3pCcxbp/MdYiIjCDA6laXHV0Krpv
wiyet3fM3ewvfN0F3J7D8+dRAv3k7q3wlD3HGwD4Hp+MCv1pKeCfJkUYkPNZuADJWQgWuVIv+fdx
XqcJruvTBzoE9vzOXVSV9ebNqw01ZmRt4u9m6B+m3k9mVs0zRvOehGZOJngNGPBBKVNAVqki1vGt
hlpSeOSHEulcKvzITNl+xErJgQeljpSKLWY8gXJyHxnForunj1KJkE1JdGoKGA2YunUS7Ldky9eK
EhmHcLk6UD6V5qudQ1xjf/+AKqhK+3e4svPCSigt2uQYexnVJ1zr1bHwp38310MPxKLSnkW80uUB
VCfW/FXeNstAJIenj2DzQlnd4eDM2vR2Onrw+fRFrRdVl7LfSXDyrmOloC4s/wmPKNnZMud8xOqY
yb45TIUbSbeIDYUJDLM+HeVGdHXzDa+SSZVgSwLzKUU8txUs95pQgPO4Eqh6Li+9jwCgfBJ91Ytn
wROwI8vdI769zYP2JM81QUCwF8IKdZDNgIs8HlyKdBnwBdrEoA7PMaI2bfXwZFtxuT9VY6hCN34S
I2QnPKV0q+M4lRHVJux1tAxsqpCndN6STs9Z7zB3o/lV7/koh9vM/NTQqhX5cYL/jtmnnovuspQQ
CMuIKexjtr001kjQGMhgeWE6aWi8lTIQxKrSDjtmTRJaWbyGT5ZcNAtmUfuEr9HUYzUXjFUT5myM
pEy2UZBjH4VQM6JgZx7UA0LQDKIG9VWyaDpCCjf7Zi6AOJoQ40JdsuvujEC90Yvj0cTMsaWJFFuN
pTagYM9DvQwwvo5L47KMdw2fKnoVyviKSERCJSdqf5gCxyQX/OtYhNGNF3SG6HCzDL6CnUaA49yQ
lTdFQapI7VaQ9WOJiIkCKiF55IPYEJvzYlLqgxBl8OOfqNTMmWSuwky+Xoz/hc0UsIP/D3nxSQK9
2na45ucVR9qV7AOAnHIiRUZ7OMS0m/3sFSaSD5Oy+QyixVYMAvJjFa5zVarNIiBaZEmtvAcQEiIO
4jrg3Ifw5qB5+WfP6oGvTaSmw7sg+BIvOivAA/gE7dvGLDYfZ9kE0KNDftZbgi+dPQIa9Y8yDPG/
0hC1bJDD8liO9FPnQfVo9pJd3zMdjWauLRd6vkiN91Mbl/nK/vO2mIvPY/2sapHbAOLRq4Xthgmb
U+ZKC7EMsUOYPi4J+5i05cEZkOUcNznVnLXKQnn+1rwFTupdcPKedRb9hBhfWssopzkto333OiFt
HSYY11v95+SFz0WHKwuBya1QvO3T1NCfdseyXAECMa8x/nK25Tbegxd6qfh3HnX804s+uao+NvUe
2ukaZd97XmD2jTMahbM7E9ug1goEKp63rGo3CDDVeSAczmV0WBPQn+KAy7usAfk1NKNG6cDco1OS
7xK6IEuWNzIymVAYLC8nKt7qaF/ABuDDzjziJUJpbGHh9SNQTYtISX7ge/bkw694A5hU3KIKCyN6
JbiazGzldeUpUyL19Iy4GI5mlsjm63lHelT6ff0pxUgE+5Lx+S4+jcXCowy+y6zNfH4G+4wRm/6r
+E9QkEabP3lrXIbtYU270et6XVomAdZ1fF2T3H+nkz8Vvl/VSh/9CwjVKaBm0oqZJdSB6VdbGDWl
8+Xi9Cjogdv6xq3Pln2LfP6KFdUfEqaST/Vip3ZtQFaG3xx21eSBY0BGc0SCwgDUp7SsRgyfbGjL
Eg6JiTsSTrcUY6sAHjlPTYDuP1jCc/NSck64hDgmIfIx0cRXRxrxJ737jKPh58K/vhhzAcBLaTuM
Y8k0Mfym7kMAe/jRSVTWzoNyo1/LOLsezEAVH0YaCfVxBoa/M+esMXvYqX4QeHA1pFVzdXQaTi11
faMcVOhDh29A114DmJ2Dn1ADwd5RLknppth0g4lp/2OJUWuZ/Nqh2Kfh/BTCYTT/CEmZYSgxWaQX
ra3jQytTPFBHNJIWcVTvnr2G0RzYU+hVQFYlQ3t5a0Bj5d9EiF0eU/j5p+J5FF1hZs78XQOT+7PU
5nHORjbrP5Me8F6XF0FpN3u0WqgtNskLbKlHtYQgvEGJtpt77gELs3fSmIl7CNhcQKGXCumKf9WS
YCThq5zPRS2KMYbce4Mdjj1DdlV+sXH0HLPfmbcS5fSAF3aYOOFcXfwlRztQTxyu4h9UXtt++0WN
n6iS1gyGqE0iFoHJF8hASsnM9iaR2IC+n8QdKwfgaBYPPcrmVdRYmyeJUsyf5zJ0K30UNig8Gqf7
gsJFVJJ9CeWPPGkvj5bhm0qicv0C+MEPpu5PST3f3+iMNPoF4ASmGGGSN1pqNVRFDzI20LzHQTTi
BFRs6m6IoR3fL1ASC2fe1ZBJMxBlxO3uePieqZbypS5whnFfxfbo3chQUU47dsChqSyjV9fdimST
zbsV4yZaIxqtpOSGG9gBdxlm4WxKRPSAMRXfF8osj+lMLl1hDRs3dNw0OIrVHqEnez9YPnkARJd3
YNp7+xZCJ/sw0ZoiTov/iO64IEsWO+agBTSrVkbZSaJxKE+GCzascb+CWGk0fBMLEGTF6ddbnvaK
tpNVtlWp9NhFY18uCpkBlLY4Ip9ocsPQwmgT21MZl2q9uYf6wmJI008xUYXp8+ak3Lyg2KYln4Js
qwzB0QPGpFfS8FfioxGpdBaRb1Jy1kcRnOB0/yRrB4FJwhrlODC5ZNxZ2DJ/nsIfiepazpNopGEn
AIyEzDd/RB83LId3MZ6VwuZJw+PHOkfo1RXaJDp2mEhJecCHkCPdruldNNDGVM/xd9EVRmgsa+I1
yMrcB/+8EVywBlq1dSTe/CBxK5bUFIJs3KsJVxnUgGF9u7l5QklYFfVZqd8WGfH9a0cHSA3A1MsD
NEjfzE1iHtHzAbMaAw+nJwkKXDgVjaF2Dp9cEjRmcz3iRgYwxdzct4spdnIv7ztamSnlKIgQmDYu
f31BOvfrove39ykgf0eqSYESRYY17+JVgPb2paRGjYYMMcm85xBV9UnPM/zE2JoCvxw6pwvddS19
Mv9PTUMMRbKVuGxJ9vjhhSb8283W0h62KMs2L1P3IdtbaS+tt9G4XTUj+GXlxd/4f/mO9VoPRV2b
OpItBnK4+4bVuUMb3bFFt+D2Q0wHZ+V1CkFaJ41mb09eIo4uuSSzC774pUrVldKOuCF4Xz8ik3td
mM7YRvGl6IwoE5jXSsBpC1m195rC9VMZRmOcDJKu6uAgSfr7YwphoPXcGl5SOZDFZGQ6KPYZTpCW
TKliVFGDZVhOuTWfvDisrgA5dem2egJ+lL7kPIuhVQlyyyVU2Lpku0+vtRgfgGD1qDXEchyJlLKu
LskOBpZRrW+mkLUiSED0urHXPwQJAB3tbjl+bf/hVOFYb0zOhYI+39oZJQo8IyqqFXL7yWQQYLR5
3mnGwCDQX/LV5rpCGULktCTh3TWatujA9iKztXrA9R7myWZR3B5FV1flvLXChjo5L+OrYabexcBV
pWyAXbCQ1Nk4FAK0sBeDA+Kx6nLuj66XFhGkW3saZg8PJU72t5SII9NDA18sZQiwNW6HNHHURhxM
NplbMd5vygQzHw1lBYrzy4JGdrxV3MW5pNhQljobwK0VypxT1aLlcYnTGYrkUMvHDdZXwc9KKsHw
9VMDZFxEE+C6OkOqZp1DwHnWk8NSYCLWg2pC0rRLKtBDgo4j3TadnKutka6cR/x+khvK54aEKnuS
zqwCKOBHP5gFIz8l7E4ouer7gjmXfqmgOmDOrZWt0ESTWOs/LLPVA+AdIcbyJBgpJQY459hsYrn7
cNKsVkDOqL3w3KxhIN0+knWHlhPYtFYHVoPBCQhFKZ+Xh8twJyQQwjR2MPs9Y5qBzQd+NErfoWKr
Piq9GRI2sqokGnf/r1adPtyzF6gEW0o7b7KlJXdxUdLGI/KJivSW5/IQz+ZB3lVvRDBK2IriLcs+
F0fZHIBri7g2EQ/lnXyV0flOeBuRCc2WdW+C4w0SfbZxCuMto3qcYSN4UaDbl4qRgzpmzf5EAiij
RQ3APUZwS4ajNBp4jWvaRkxp+lpPRm1uhkhQ6XabZW9Y5ZhpwXP6Amm1mBz40QslTef2SVSMRoSD
hj9/w/ffNZ05Ip27o2go59WY7R8vfeDJb3vIHRq+bDoFZNmxw7VvNKE7aFI3dKgOHVSPLd5m/wk/
m9iwIxLNA63bKH0P/sWsl1CNojmUiQF+GojtlyWmC+8WliKv21GIfH68qU9LT8Ay7sKufxEp1bxu
S2GweiFTH2d+T635pLuENY1An7zBKAVx9TgWjeuLiVRBrPV9AQQTGCS/PIBPcgND90movO+6nx7u
K4TvjJdrCP1zLozj6OPCD3cNsgnZEPmA5WCneOk6yIOyDdaul8qGg316QJRXh+HOEFoIBeF+A22Y
vrc/6rfsOxceGSfZz1duaCnEV5CZlKf5HPP9WMEFEnowrrZeDMZ/krl50nXY01yr2M5sUnTV+RaV
4KoIfcln2rBs5xAe+rLCdtiT1wgayT376WW6WYhpCrVTU9dr/Ed2bxHZyy2rypY2fWtDzZzwE/dB
Y3YifK5fAr/JG5edapLOewr8mlIXWCcMGja/k6iiNOBHqMqZZr7ys4zGIXYVDUmiVLojnMqm83mG
CPTrXYPA1W+YZ8tIC6MRHo2L2P4iuEnm0wP+62l59pfBAWt9t1RFiA3oUXsf7R0AlrTPo5y2jK78
SHLCvs4mXDrs2C20E6U3CjfIY5oFCebi57Wqg2xQJMcqAOo94H8KvAtASp5p7TL+X+F0LbyIxffI
oVfX1UKHFkoUpna7fboFkpz7kE+5yWdyCx4pxOqERw+aBB5K1jKxDaDOi3hcWVhqSVkaz7xkSAhE
nfrymspYABmeu1ojIvC0R5d65G8GW3B0y30Cfrb8HZB8FUax2o7GUVEvGCJEGQuGcYT4VmjPFTB8
rd0P7x6YC+M4o9iF/a+zrcvVg8sERrGPkKiKEsgWslnrqpFE4Q6fA+4I2g4AZ62atPEO9GpSsXeu
NCYrlgxRnwoGGrG3ESRjB22DXQbr1pISPDFZIfZh9sp/YZcv6P/V0gikhbdJEzVLiuQRj2T8PwIS
0TsvIBI5KZoz7Ru1/b6G57hxxIU4xjOd4MaqdVWnRlXkRsV4EjAoSfwQR9mKgxJJDGipWN7kIrJB
J5c1/vR9CJxoSN/TCeYz/6a1ITYO2Sl4mT0Srr+qR4DzLyH3aTEtwPA5KxiMw15OgpmGQDx+YpE2
jqBQuwYR0do4CBd8UrFZGpZSDhu/fPR7P+x6kuiBhUgiZVseAOL/+eCa5KYg3xG4uZzkvvQpNOEB
wykmRYo1zCAtpDxTf9axA0TjP8QuHDFYdAguPy4Fch5GyIPgrB6uk2dogxGNY6x0iYVS6DoHdSCF
FDKSVtPXRPxLAtuDWF0g5h1z17shbVKBxabUn2krySxAuNdk0IuCu+zsw4JcEufYclwKIDtcB3BO
5ExZzZ74+vP5SIaXQVIeKFYFvQN+jdY++nQuL9+zrb0hUTyldMAASIGNOFP3vsi8uc7kYtpFDX6N
gC8tFRDreeA8YoO4Y0DGA54r94vGLYmeCop1GQfdSNSxoqS4As01ML2GUtYzwCQFJpl9DeWgLrfZ
VaXP1OEPB+gocReN8mCgWKse2y2cYRax8nF1s0nhB6c9M2cgddvg+PUaOB1uZYmEhaQv0jBYErXC
I83uAZzBOTWhRms5raIlN8qTVVzdjgDiYRwVlxJENFqnrbH8FhF75Sk+spiF9Mxfr87NH9frEFYv
92+1EH33puUDxS599DCqrosm6DIIIg1ONnlsol77FnrdD4NbIG4TEZFvhSrSsrl7+xTLDN832825
eLJUG+OjECSRhJ484hgWaWolrL3haPvkjvcpZRl3UJIvirKeUkIJq/veHtqkRaObWP0gylZkUhe/
c54IoOK91QNsjGv2msgrRUPwG2UOX1p3niOOAywvAOJeHil8HCh2ZgxmexmrDL1HcFC8rCrnNE4A
sWrp6f5dX27RzFgjKAGp6ltemQWVMZrAUzFMEDMYJxUhIzvmyZHkbr9mtPCbdS1S5XcMsz3UBWUL
z6HSYgNq0nK9HIAFwFriERgp9LpbnVEx0Q1uG7ldGqW/0GS5tAi1xRnPyROUtmSinaWCXaG/Z4sy
2wfxF1V4UQZZB/RZocYXbHsI9sY8oWs6Kuc4jZ7VYHN37xDIcB3MNett3oBHHs3kiaRNkiDMofRR
uTjlQIDRsJcJK5gbeIhntKN2aQ7PLa/p95S7jZJ6j9Gy8T25zALTy3/dM9VA9R4X92ASboIGUUGW
43jwr6LDoa5IR3agOI9lfCm3CRasiHqxwjieJqSPKhwPYphJ3pnINdWdScKlsHOkbwuC3HUretai
Sd9pHc6jZGWtD/uW1VvMEIrkYs4BO3JI3aOdvtV2o1i65J/t2wLZ4yZ/pSZyfXiV/Iv5PZjsxZ//
LfZsYsJsOfWLs9+DA864aYOONNiupE3QiDEM6AvWWBg1RBAskdFy3wciXzU+Q0FS8+OcLRC16YKi
2FEYy6o8gw9iJegXzdg5YnmJPKxUrqUhn18bQu1TRijYKhn0Gi+F2KYbqekxlEVRFv356Yd2heGH
68lOF+6q950hLmorr55a6wdOfe/mC6sGCJ6pAE9zjodQXZGbhxupZuLkrluR4okZP30nAZ9J2sPQ
w9E79nuVDkYpnER7/OOxl/q1zk0vBzS0HMU5ArAtph3vQTQ7b7OFWicdyvjktsuDHaBKIKWbQKu/
Fv5am4iElH3LNYfhurzA2zVF3Wgl/qLSeaxPjlTee8iURQVxz9fOCBGmUgRrFczn9u2+YYs8UpvN
BScDJdn6uaXSBOllG+bSGKUDxBWxDzJWu9egr1Lu5NxYE3zJ+m+sw5/8lixtUfZurs6RBM8RP6q4
CG8iWBcc4s2Tg1DdST1tOs1t5YVFUJDF6NZApKnzMGKwDo9i0upDXGqzwDPeTdH7tmWntsjXlHgB
hd7ijZlDon2iT/eJIGY9knPO6uTQ5xHr6+urI8URT04GJlQKfCwQea2CJFF17c4qejieSkAiRMXH
1PQ8BvuSCEhC3Btxn5jQ50HvhWTnT8by8WLyKlubdCJeiH2AZzNzlPdqrCLtoBrJOoXB3574PNCH
2Olhspf0RR5mqL5q5CCCA69c6qrTkqKkgDxoOAO+D9PfS9eFpEzbyE9oErTbz69ZTPgQTxTwFCGR
t2ye6VbX0lKTMP62it+Ry8+1tszgizf5qNDozubDAmdDoR/c0XKwwIE9y2yisnHH5iiZ4vl0j2cB
IglBg9Wotn1SEJoYpy5CUx3vhIWPW9YMHK9LJnViGp+RiIWWRH/l1/MDoc4WIIFVcombQY0wDWBo
igNh08ol2+h+Gxy5emxBVzaiSwxuIgR09XLqxFiyCOmFlZpCqdOw7gAsWJYl22BtwnbHzgvyFwNq
mf3zLl3ymHLP/7AK5WKiKNpFWhFTyxhQb+Lhft6ByzGqQWsKrtUUWfouLlsV+qa3rAsR+BIUAyVB
DucpqQhsPNvHjKQa630Pzf0VJE9nbzVuQJqTzNPD8vR6ECpd6YXRiLTwEQ++/OYm2Di1MNljiu97
A4J9K2ibDyKlWFulVkdOr4uvwR7wMvI6g/1CSxp+BsQDaaiShu8hmN0Dc4fH2DZtqetdfBZZiHH2
vBPLxtAAu6zQl+h1T7TX91JxNiDf+YjMWPOCvRzBsYuzip32R2OLhFn2aWBllxI75X/M4jzUVpmk
CU1Wkt9n2srxXzSJuhpIbj3lBZM088+YOMzzbQ+TpLC6FNAze15dqgXFE3W5coGZJ1ANiQKSiqVq
Jj6kKDG2Fot8z5S/M6sOTGH+w8GmIQwjCjC7gb6l6M/4VPcqjK8OR5zcMtml6L1LqrNmyoOQixK8
ibUJTdvRZmXb5aFQQ3fXwjelAJGot7ojlWbIfehAZhAzbrVPRk3NM4klLztgEe9olQytcZcVt2fl
GNMg+GWV9yvY07784tk+/j8LMuomO08rbpts47gsFULDDpu/wzMzTCs+PKuihHA1lzWs/ejVT3rs
GDHCmyVFTDmjHrFc68GtsGekMFZZc+8rziHHNqy0iAdePCzr0d1eUSII+Cw4o5VdR2YouIb7m14A
Ruade/hoge9sMTCbVGzC/SIpm+dszqAM8t8t6MQk+iXu4fJJYnmYs3hstaOlTrcqtHZkjN1Z955C
EbIPNXlrOLWZh0YT1cLnMDM3h+cuELI6rKHCjk6P981LlVKI11UAeB9yqZTnoRv97D0uaI9tRz78
omJQNKlziYwmGwjTDNJveF071g89eFrATV/09tqac2VpC0/8SFpGxO++xgyoo+JJRwNIXgWZxIQd
8+9uBTTzjxBcvQPRTpB72VNUAIDbO2kw0Aa+JTfqCTf7+KlGB0ZP/fwus6MqGc0QBNJ9CUzqFKru
eCaQ6QZUOpw9a3QG4mkjhqUuy1xm9bhylAL87bDWyTH+IUV8WK5n9Z0ECjgVSqxXgWKzCU9R0WBV
CILqGZf7pOK23LJ8HNclafbFj1v/WUPYWgor5MjJHoFJo0udDHTvmrSwqcd+sngmQPUg6Bxw6qQa
rCjlWQyEgP5HuqayWcps5cOCfiGD/b9Q1Y+ng97mNPDSWpZnNyEqoG+1eoyJinkTQzJsP5Ylahp8
V2X5TtMbhGXzymSrtNvloDehBsJOg2FJNpDIxI9Kt5b828nPcwEAOv49xHWmKBQPY5/k/DWHyZYV
kUJO2bZloHL13CrtjD5QnDHlbMJ49GaxKXdq/12o+4Wc7ub0kmlV2sAkRKFXbZkr1DWo30j33V0w
4h889//F7kanivLlZFWJPG9fYTsHGOP0+wXMqhMzQFaMP2x4e6LEF0eVH8YyelY4C+X0f8noQWVF
FSbCQnEJU8+jUHk9gfNx7f0D5S/AVXfoJFEp18rY4jxlgNgjY+VtmEwFIOxpHg80iKSPBUxB2OmV
c+KArAoYsDGGPbKhPdduM37YTWwjIZaLrDN2meLDWC2Ry/Y4DOsPXekR2wkbZ4/Dw6mXV9K90owT
v7hPBy5OnUVxIlQ3Ravmqb7tzzfekHsb1zvL6eWhY8Vpw++q/S8q060OOyBf0ngANQp2wm2dLVxl
NpkWy3MaR+6PKsttnOq+Z1FSV7FWZVWShN4xfc0SXmUTEdBzZDOg59FfNA3NDhAdxnL6FJFIa66R
RXNE8nqvd4Ljft3JTLzI8Jje4BX2vmV8XhVHRVDzBjpOcjsNean6iz3uaa03ZIIaIMsaIoY4IBmY
huOXyf0JETPqRNwyFSJ5YaaW6y0UVis9/8p3qJ8dyCH7wK73D54uS683GF2bo6Rs5djzEYRSyTsn
6sqH8ZpLU79iaA4+xiuhnddVqMzL9FjTRa1mBmoRxSitsQ2bVx/ASdnM9fXFy6YtJj927RfxkrEd
INizTew9dI3PVaqqcNbacwB8sjV2Y4QlmquLJDCMuMH2vENGcpoQ/putuSSkn3+DdiwumwPIaseo
9Z0mPu/ekzje/0fEzSpfKB3hOwByy74j0aj/hPmxy42r4d+cT6Fov7ExIO/rH+hh+PHaN9XfmGGI
LcljTHiJlLFVYchIuOCzOYGu0Gm8v9voXulNAN286VO56AZ22BVhAYEVqXR6mM0ITVZM1Mvv8UCe
+oY8SFe3mprUa7Gut91YSFYNYbD/7KLra8wxWM2aXJxfldkMuzI0GS/CvawUzzRijtSeFUz7BChr
f55/qEzScKuTRLbSmwDb42+Na7Y0L/LcShBSm90a1fyVnWE9kOiYNwj1HOC5Oi/6Lns2HRX5nSTm
+fKaDZv2FvC5z6jyZutRVYzF7PtMMniBC0aI8Vs7zXhpt4jwRIfAgCZAHEAo8GhY5n7rnnArB9SQ
YTSrvkPobYYk42oqPxI/+tobiuDoSIKv6jK7Bd42R1ZSiEZUOuSi9TxZpzqboNHx4IILqon6mEWn
bb86kdlqTwatyxE7SoXHewgCGirdN+AmW92GKlWGO4prt0Dj0HaPxgKi8e0+rbsfpMcAzFgTFLOa
x8OKn16mMHLGMTzQI1PracH4HwFd+FwcTqH3nTo5PWicYVotw5bjcSrZh/dMbh6Q66GnPvmdPYsH
hXKYRsZhIxcU/xTkP6dABHlRHeXToVehJ0LR1lg8Chczbei4aQt2QfO9kjt7PIpuK2ktxcCZEY+v
8avrqYNzOXG4os3HDHo4mKJhc9rUZaJ1KGNp15+Lmrl0be7r/WooONq011EHflaJP2Tv5hropMTP
ZVfAjVcZs3Kh1Gs1j9oRlBz3eW2MHvOzsA+biNxXSn2kUXbgDkEavZNl2IgPhnxA+82wJJCxbu6s
9/8LFc7pLd0ptUjPd1pZ/tje2v8Mkz0/iU14I9PIrAjkUBPFrkff005hUxsRfuKB6rBItR/bHoXm
sKWA8Jn/JfHfwXhq1i/6W4LUbqKLh9lY/GQj4g5l2o/cSt4MiNyCN43tWgJvYB1hQ2nQ+OZtJiJL
FmC8XuDnb+mckcvj825CQC9pNxTNleFYJC3v0iEfmPU0k2VN/edsgJ/nYNqfy+FeXqEBuuC7ozFj
FgHnilXaSMLgFvizhFjxdULLL8hTFZR5Imy81n4Va1b0yvB2hUZfpCuo4Fta4W1wcc4Jdyosy8/4
wNPx/AZJi0551U+0v4smvmUeyCWHK84GjLTx67pCmRId4py86Z74W71UGBYMPgqOMjs3U6j2sTNy
5chl6qtz+k26v7Y2azc8TmbVRO/905QOFgY03IAwwwJnreqzcNkxfzKMC20VcccJ4VnYgjs73Kd5
IYBdkPZrocWN9FDYXnu3p9XBFuSrOPyPHAuOhWECjlNE4bLHI8xV7ENfiWQ0BVUTCs86DSQ+DbnX
+OfMwMn/OLQqZUCnKRpuTcfUbGw/TgIKyUZisFDPa6u269Ve/gpBaZv2wdm74OVOcwTlkpgwHlQD
XDiBxb6+6NDWczy+91F4uUYz998wI53CqgsywNTnvZzVgfGqarKqfpAsftxylc+SO10baNduXzRl
yBQFnv0R+ExtuUACDhC0kJ/k6G0/njjxJ04JVgaz1YbRo3/iGu6P3bLfQzEcn1UL4P8QGnAYwpzv
zph+nLPA/uQqfo5P4yfpVq8MJZfajh4J4D72mj8HWOecyMKxd5IQeM95Y4qN2H4KOeFuvER5UhDN
p/5nbIbJEvh4zyGF12w0ca8LM3aX2YF41XOIXOG5gxFWmIS1a9OYiRgF9/lhnCwa4rgA/ktnEwgm
RrhLCwFV2wThCIMbNtt+/b6at8I/uQYNl51uRY2ri1QpVwH/2NqNya1897njRO2ZoUBIFeDUzlk+
SoFJgazFMDZfTSf3IvbCpSqt/2IHZ6tGTK4rts69TdaHZdOAmD5Z69hPqakEtqhm3HfzMthCoesf
2WxwNC4vaf403nTsUHKCrUqZJ7QB8zgcaSq6/nu3DCsuLJVqSXLboQeMTWJqTjN42/ySuOz5+peW
FSr5rHOe2whYbUtvZmEhPOinMNMVGI2oyrdhE2IIRPjd4hYfdD4FL+MCcWR03y+temgs928KP/xi
16kw4b+aGHqZQhRg3W8E+EVMCJpUz+9/hdyp5rqQX/x1B41WUid6swDO716xPMpkYWAjyCOGrcqd
OUVFdZU7sbB1K7PNjTiXOEChhfg3OGwLjJODsM0yQu/FWPuTAPs+tSl1gladaYEQ9rNR/bo3VDz2
iMNQInSmFJKezGXulO/AqHr/MC78zKAAlxFTvNYNpbqjBFCVc/28f3plYgp+HpeETgEpGHog1LlK
L2qEBhJpYrhW+v7/KtnPOlXzxHwXWo81UYaMz2B0nvTqh3CX7L+78lCbJ4/3OFl+qwLchGcxBVmC
vKbT7ASEn+eRrz5osyoXsy/d2SF8wDS+MUv6yGshPmd6Y5GagDTEJ+9dapebL497ur3M1N22P7W2
zMqxx9rDKLKmQy1NgiSQZaMc1FbL8SHCu959h86VJ9El8kCi8bHuHS24Px7KoXgOIBlLMxtRV7ov
LPlHRYaSIeigkiw8gsuqDfiTNrnX2Krfg+NqxgDNwOeq+nqVI6vuFgcM8BjILG4toeRFwTl7c48T
5RcTJaU75MM6Xq0WiAWWAEV/TGxO9QfxihiDdRDTk7ZeCHaisfLYFpTzo5wEhOmqwBVtVvt0wT7X
P6lm29QZ6+EgSEzrLfbPNJTJIQ+/gfyN2fNFpm2W9acov52nEJgCkPrdXT1aE4IIglBjFUZkr+xT
4Ph3br/afy910IX8Wwi7zLEFmMn17CYqud0pfGDm00AU2CYr8eXsBT+TpkNry6nuuiREABp6vO2v
kc/3U33eUz5LMOD59nKSAufrdnVb1yRqHPzjniPZCFbl3L4KK0HTMiXhfBxfWAPcbive73o/z6Sf
mYTZzlld28N3bQnGxV6paRTL1KJW/Xs6Gj2k6MAzeKFybrMpALuVypExmIn80MudS9x81OQF4gru
CedTnSBMgCfrmZ5y4ZDFMGmPdXOm5yFYBdaW0P4yvhL/1xny2QZG1r2x2IYwpfgAryZiOdMqTlG0
Oz1BczEpoq0LvXTRdgnxXx1v+PI3v6iOfyrJnpBrOo/EbZLO2A58XYy6KYBmsM5SGZyEY/182dx6
zKeuSRo382uR+nzVQMkckxbQz/gAYKPuiEjI7Mb1VM/RbsvRxu9IEKH3UTmHlu05++cNlZj1JCzZ
NLzcAdJ/x5TgSO8KHdu8LBtfLNUnKVWtmXlv7Upe67GrG2iCExpWX6TgTsVPF8tSZg7iaPNoZ92B
MiI7wWlYBWIV1KG9flcCZChDUojdzynJFgNKLfjwz1hy6acxq60nrXjs2bCzke9u8aLcLV0TZL+g
thxGID9WsDnYxr5HTay/kA3S37ZIIWxvTdweDwTonUS2euFlQqNdaquEJlGv1FfLtRwUOe8QRBZR
xiMetcNQnn0I8DFR4ysHVXAbqLez+X2M6mSC2FUTIgWFUGNQSQZJ/DWgbW0mI8eGBHwm3vley1qC
z8udmNZeBcVfl3kstmsUWQp0lGjCVKxI1MoEJKXIH0kho2OSjzJ9UqUcudossbEPNj9iaFIVtPs7
pxxL9+u6Anu1FaVFX9qEPIeDmj0+jxTCjEDQCpvpS1A2H2dHHO5bsXpZC4LeyXT58PmsG+HegXZs
8nUAYnPmPehFIbrHJs3he67bJG4znhH21XZuXXs1gGDl5rEPPYxcDkj2HV6z7mvpcVlQRPx4MJid
m7IoZ4JKezLY8/jY+CaVMoeKOgPpjP9yDzAA5cw3DmQk0rrF/7XmxJksnidyhHlj8CJ/nC3cU6JT
I6/MAS3dSaYNPyyClA8GeCdE0MpK8rfZvVXc8Ep53nTwqYvt7HndsExxabye0D8Exm3AfvU+R53N
sdTZj/zf41cv4z7kCUSPTHqBc1BR80xPBm/dXtbnRv8OJ9+TFKaP+8jzpdgMq3ywbRXUM1QHiQln
LiXaApEHUFoQo/q4hGmgI8UKUY4JNEAnq7obsLykyue8IUG2u9fFFpTsbsM69uECPK9UzXAM1Kit
kLoDs43kPwpg9uWf+Tkky9+qjeDkYzMaEtNYK78U2CCpFaF0qj5ShUq1UUYmT75Ntor3qT/KRxpS
kze0YpurjRBvg1Iw6oIz+KNjoPUmcbh1k/Xn0GtIwfgcq2V3UV/9BqLTsdC6vpY2xVybmO1BaDMy
sWREWPLwFhPGi/JFjT0DMMz2Tguk1OmajfHmMKlj1HOVd35jSiPJHBk4mSB+cb9oPu4rDI0aDNnG
gz4fwIfhWsKCH1PCLISuzal/qXf/OaI4vn8O+FqmRQL8VuAvbRarPMVotQG6EJLumpMCAUK2EeCT
ajjPhVIe4XQspQdeIetelvzEOSsSbyqOC6khsRYH+gaFDuhW/s4EFH+VQ/CTkKWwNv0Xlt19vqIQ
V1qf9vNQGksJRHjUpaxzROPsvqmBky9jK9TJoE79SJ1hkVtZZKo3vC0r/7fwey1ILM0Yj5FeBbWu
1vgUOB8IH9/CosBfSUNicILWVp+6ZW9TSN2Oe8Fj6wqZbkQe57Deqd/Au0+uLoPgHpr1ki8d3kA3
Gosykpb+NxyOszF6w36t81tEMoc6bUcFw7cGgt21BBybIuk0U29tRSq2jfE26c5HLbCBpYviTX5H
3XdsN25coZtBiCQGoZdUcrhg8RyFwjUaAsSsT4sSpo0y9LGjc8pRsCOgUwPH8bw8MVxBVmfzUzc8
rzR6EMq3qBWomTN+EFYke2gBRoQEyzQb6/mGhG41H1YeOtIc0mSYI1JUdTLXMOvOV1p4c/IlTq6Z
BTN7QzoZEKzmmErF/lpwKAXCh2Mf17njS41/JcMpE/6RZQDqOOrnBT5O6Xd9vadFGAVnYle3QZel
HniHABJe8o0pTH0kJSw8LbzekPgVEux8Sm+zvNkj9+Yb14Bu8DtRMIp72s1b52EWwHt/mVAXLiF/
lhXP//2358u/41Iw3MEfAet2Kxp6RSit+bO7ibAUS/Z2ebyF3ciGl66yUUg5NLRA+0C/DnJIbPZc
ruThcbaWHJh6meAIEGXE0rC8fKH454ge8jb6cWKo5jCrzCft/8f3XG+DLYCe24P6iZDvhwg4SUrG
ZxCpBliuUuplACxmEiKp2ZpQMHh5OmqesiwLkMa3Wf8LmGEVZUCE5QkjXBreM7IabZUKrcEuwoEU
npdt6ZsHx9Prbh69ZyG1p4fZikI2nyAK/olBmVkc3gnbDz5EniLnRRpPVRvO4mU0sm20xZ3Xr4I3
VUMK+xraQeJ4mYh4dLj7JfSuxVU68lKMy2IYJFiu+MOPrEaToVbrGxr0ZuhRcfqW1ZtcHVEogbdS
xbdD99R9qRNbPrMlhah83h9BnxGfUos1V3Xdd1AYujU3787PrZCQCF0sLbQLJZv9E2rhrsv3oOl/
L0tR7C2oVPKYorYCJlxaB5++B5KBdZN/HzxhcXGfQtV7U98dV+bnMqFI/bkHuuI9xBOiMUqpj66b
EpQb4rHtAwAJBUHPFK7nKsxxYG5nYLyZdihI+rq7pD39n8hqktYSlpfKR702dgfCJ0gmajqarIJK
tlbfl52Xf80UWMumeAtrB3pzBczWCyaWzz944WTYYFiWIyG+x5hVW6fWtUShcuZcj12XDwYQvRp/
qvchOm1DdLm4tCcRSXMnNjYT4NDfYo7fcOV4l+X43G2EGggMJJO+0GABTyvfGIHOA9FJknBXeMng
FLmhyAv44JSTnlaYrEKxlESHUQey8+LBfN7tja7k1pleB0ofrTAaN2zArAaVTkGXIPgjgzufLFyC
aO89BLo2v+EbyurTayVyBz6ngcN1tE9vk1i9kRkd9APsQZln/TJV3LK/6xQjGtAcYj9Xp+yst2Tw
PZj2pQ8j1slL3IcdcorIY7K47QHrZ9RjF+Sb0EZjAizL7ZxqFWsFwC+VpqNK/srch3ubCpAG+aDY
UhZK1ZDdsCATU7gOleVJ80rFWyrI/NYkfKu2OmYXPWPYWCOlKudvqWgyCeHBvMhKMN4jJtNry3qR
r87RQ/Nl83IzSgYqKpEAsf1prEtAAnjnxHgRCrE6pNPp7WQkJX/7xnG56rKR7m3q84S3fENYLl9L
iXy2DPXj1pa2FtL+NSQTy5Hep4PfhqAHKV2vwH+un7KandUZfKmYFL8wzT3rUcnabF2RArwoeTa6
g9tEavHEtv9B8IJQ61w7URkABGphpLfUQ4PGCBz/4RqckzjQXMZbc2PBu2AWddwE8krzK7QS6pRp
Lzsi07ZkRDOHNPAi0P2pp3LEw3aCuB+5Z+jE/p+OQGm5OCf7DZ5VWmdgG8aziR9HUl+bqrccDmqi
F2J+rj+fih+/U1K/jkHZByCDqriiDwsjGzc3EpWKRmJL0HvOGbD2yBchvWP0Kbv3552Rg7f0/0Et
47F/ZIKJ5eoaF0SrExFcALoSi6w5LfuP/pndkSTK11z0bJbOmqp2yc/4DumvNyTlzApl763hHKRS
TI3OWUi8LVuYDIgqi+PVOD8tsi+mpfAS+d9OmrsAw6DOZU442o7ScrsVOSgOw3Iokij2OoI/RxI8
E0WU3Cg5blN30s0CGAdB6/Yr9DRmZgWkhA9TMfxiR+RVQ7/LQlMCfBvKw1k3fd80rTu4TQksfRw0
tva1eKqHk3DtwOGexXTVJxxFjNHJ1/xvWoRr7vXdjEokQZNxZQ8CaHnsHy1LLegTA5lBtSco3bEn
ONbsj67GBNd+QzbFUCm3dmjuzlprjAwuyvgxbCGMkb9ThTw83Ps0ldh7evebCgZTapNYniHwarWG
5QFRI6SiTRm6wTkn/oFg7A25vwYQDf/4TpS8ZtQp95b54wfCMlA7sDEo5/UV0BrjqDH7sNKT/o4r
5oePgBDRJD02Zt1nHCb6seclL2nk/73CO2qWHw1JJG7f2uVUdjFLvhQfQkv1RDPQepY2FzsZPk/7
eN/P7qgi55HwNxAaMPJSTsqBy0kZJHyycQE3ruLTNkoltVNpacdDHkURIE9//IoLIh3F+0TwK752
8EiKq0XHB1GieTG1KKGkLefw6Ee6A8FfErH9OCNHpVu35Rm+8SbowWesoekjQj6DC/ZijH5Cm6Bz
WHXBEJRaDwbspAkz6IbPW0zam5AwArWC9VeRjblrz2Mdca9W8/hzv5re1ZNrvIQInCk9DgLmxIDd
8aK64rRYPvlWEXjqosBhFqCrT+HNgL3NTauTBmI+ZQeZdZejMRlRv5TQmVudm/J3pnN82IsHvmzj
DvENCwV/GpuTfjhxGFEZsSraKQSxGLfqRHXY8xDeoW7lD2YYSanerVd7HqX6FUHow+4oiNM8t/Dq
j6LuQ3Ffxr7b+2nCa6fh1AOV3l4y+FhJIorSLuBeoPvk3zduQjygGyRXuNRFFEAWsTvC43NFebTS
yvcUQsT09twzJKfXPJRtqynDBujqJxMyXHlPO/V6a5RDqyoNHO7tMB63aCplb5NntadxXqu91Pxb
X7mNUgiyi0vMDUcKUlkMAufd3g7uyoo9XDJbvWAQyuxZmVIUGskcqn9UvgENOIfi1OOkF6Mt+deb
a7bgJqdWnj9X6aQFP3ZHtEbrzTBj1DKu18dyZ8tfd3aV5VOD+CwLbvnCx2HwckwA4jCcwk/GvpMO
u7tLnNTo1t1qkBjEqY5I8+a4WnKcGwXgHl/j00AhAVc0UkB8Gbu6qpCJc3+zbh2H8vA90sFHLTVv
q6CXJDq2Lb/8dRkbphEj+cD8EgdUpeLAvBTuuWGIG4S1EjUqkAQ3ylp2F+FZZRLNrz5fZQA9HIyD
BQVF8u023Aiw9ZXiawOvisqjsfKxOjNyZWaigKF0T2sDI/OvJvhph9P+2mRMh9oLZWOhZ8NqOmRt
zmrUYOmQ0kw+TyARo/KWO9e+Q39wkkc2tzaWtuZ6GX207ViswaPMWjkskr+uhbJ5cNkaK41uBLtb
rqWyO8vxqICCAp5Jl+2L9QBC0daGz75m3sdwJN4XhW7BYC6FoayU3ch0Fdf3UdRk59WwBk37InL/
snaXjt0oPhyyAkIqFNwpXKM/DiIeGkpOV1SrLBFhHRJiZ5Gomwm83SBpRT2SoKXZQgE2AaLARE4q
RnK/CINj63kBbS6EYjqokk724IH5uncFo3ZYIjAXMQsF28DfAu3VeXpDQZCa6eNpblifwbpmQRQB
UIWcylPit+xkQNO90N4lZJOZHJEMPWpX7zyWFNLNWgC2cHlLLd/imqzmP1imkbMvo2U0i4DZazip
QtwJfQZnq0KwyWjN2L83B30LtV7kPES8VoSweLQBUGE8EaWtObSRmgdDLhM0PgUMAKppPtEKwMBM
r8AuCbdCe+lILfqkfW6eZI52pgsx79v9stOgAb0h5wKuGkyDAIigofx6dRJXAUh0PU7dGb1FX87y
mvkcJ0oXltnstzYYDUPWVQ8TkXoA38BlFVWpthi5Cl/88nt0+Jl7rYcnOGBV6aZlOvuKL6djY4Cj
FEkQajvS77d5CM1ptL59eSJ0iKMOhTTNq8jIR77lHSpK9igO0VZEuR0wXJjR0tpUViHiIW/S4d07
dQ9C8A7M1NmZwfovwGxP0ZasLB1qhQNy/hE3Z7i+QRtJC1wChuHhDs/2ux0aukZkfVOHSQiyM5rI
XslbvkNrsiwvyQiKr6xfzQAkMJM9OEGYNg2mPOiSR1b3Qaznm4ZhuBqgEenEgQ2ZCcLoB8rJUeDO
tttNg557d4SLalkV1LCbPUUVJsP67h5+kxp3SSOY3T417f747AsQaeyBf2CAbwmbTElfZrVjJkx/
rAyu4aiqGDHa7+s1tyhqpA5Q9qmoEb6jwPhxxxUv3LVk+FPx6K3EquFGQRpzcbfBIKdGZ68Vv6Ui
GyNoYGcprVSQoVfCxrgqkAkHb3MWa1V+1xB7QlBSYX191C5xTpVpRh7/qYRh0t+6XLr8PkadIr72
avFZ+v68xbE9M6xuGsqzyJrDacAE2lztIWWSsznBKym1Lt3odNyWp0KeJjjm5tr0xhz1yVdafyff
l+gywohQ8+fJ/hBCoDrxEtZYd7Ve9MFcYRwIHw6RZU3rj4jqSJAtHW3eb0Bluk5VQ6Q8s8aqBmQc
OouKz8FDgeXTC8MzsesZXfuG0HdJ4yw7XjjDtxZ6+2V8x8i30AoEvT2gjzcHaTdHLStraa1B21ok
hVCGi/A8SWauiYM71WPGxk1oJXCuvZ/rZtUfu8jQwn2Jo4wLOpiqMwncgUZYkyfkQBBBGdqKaUSD
AJvG5Hvxv0pAEAYEBBYyufl4WHlzBGTYLJQCIpRto4JhoFyuE8Ew6rXvenaqrsSc8Kn7CBo2e+ZO
tqoV2/8f5AmyaePoM4IliyuY5Dr9XGIyPmnfYZnCSmCWzKnbUmdfYtwAtLeLg7/eX1HYDcCXTSE4
Ww1SZC4kEjG8OhmwzaTEu3pzcOD2XrcI0NIFz0BvMAP9R/xfEj/zhYElZdVgqEQ7z855q9hZGujE
tx+0o5lzNnoecfhh6JJkzSxqvpjJCTuJSNSbtXq63Lr/4QgqJeJ3hkxWG9TXYmAgwgQNnitFYxkn
+0cyvuIWVM1pF5fyjOa8wv0TDZyrh4X+OiE4wymiRZ4QbSV4dj1hNwWlNWijgNaKrhIddyROmJad
zbS81unbxWaxRvN6i/NHzLsWACju7mhDU0EMajSCpdW3Z1cT8TuKUmJPsjh6XxBKiYK2K63mLB7t
8s+tcqAgCzL/y2i1scEyi9KtwQ1Nl+w5EyuS5I9I0GQX3ToEzlh+O78VbYXyRt6GiMsoACRCQI6l
+4mIKlwPuu5S+ajWkIqQHR7/rKDjEsJZpQqJFTJyKyqnoBuGmMfJTh/SlmXzZLZeLwPnyRpRQmP5
b2rR2rqQ91c+QbBix9vMCaohwLuNrWUNqnf/45EmX8i5VHEnT2Ah8rryprxKJY2RwhVgWVMbYG19
WvEjYxEkG7KWPxxbDg9ImNJ4RCJ35lFP0AJxmMtu+26RDBmIB5JypCw2XeuQ2maa7qLPeVGp/MMY
Quh1AWsfIqIp6CovWxFBuMsBCQ56XlPTIq86TGyACxu3O1PsiPadIp86vSo4746q8S1Q7pDLYUpj
xyTcmIDLZgRUR3RW6V67eYcNux7TsTl08l4BVT99+6RaMc0J/0XZYUu/2E7gh3SGYHACecFjtS4u
AltVjPE52rQatLiYwkBzyhduX4L7DlKzMMEg59r6rTbsxpq92qJ1cmVyETk1uPt5MRoNsPI/BPrk
ydfsFnqPxEaWdheC7fEq8TGR6q2S0ouFpmQVQzVnbxwr1fb+a2bTwlX71QayX+MUzYDIPIE+C+9q
WFAhIZqbVcwaPj1uJd5AcRR7BTAQ6pKU1U1KTo9hqmJHJTAVXEzfI81GTmQx/33CvUb+NR5zQjHw
Ijke/5c+mNCfgAu9a5gOBb5pXKIk9GT1VO7nOnupvg84m8tTaf1WS8nArNDSX3lFFbZAof4JR2YC
a/Ox71Z4g6XkByJrCqOuKwDAdrm3MygwPZa/Lj0XMzIvyULNMkUXG7cjzP6vcHsfB2dqx8C2kAEj
j6Mi5+5vN5NzoSSeYiwupyyOA7yH9RKsj9HErC4RukWmz7Wt9N+8r8/F5uuMt2YrSBc3PiR3gy6K
PHoUR1qqQ4Kz7lCkCuqRVsrklraSL8My+gjveem85x8TiTALuqbNvvwFWyNhnso/GzslobxhG0TL
fJhdakpPMtaNUsXI2SGC+ffrhVsFbf8QLpZ31E9jEQZPZ1TAZaQfErShuL07PP3ezdqsdMcdB52L
7Y5AZ56zGMnCuLo7tzFZ08uAo/BMqE+n3j9v6odcGzsn90kEsS4IwflGccuDqKlS35oWTa1NwrpA
881EaZYHtgPNKUCKt1EnU0dxjXH+BfwEWUuRQWk1FLKSQWtey3NqtWRL0AVxr1ZqlRtUSVd0idCp
iI3cxmWrAPjINFNCBULXfvMDS36K7qoUUaZ1gvT7wNi349bzzvgN9Lm8Cb9pYCPmf/Pt6/mU5gQT
8w4JbtbPGMPQubr9mNvXO8eIKLuaqCJoOq4cDCXFLM75DKs9W0PG4mIELqXoQujrMFl90t6HPB6d
0IfsKkGKZcIkN9aU23h+mhz4Ux1+qMdl326nzoxCkkO8TS2ePQJeiEBYQOzqatA6SMDODTX2MGvk
T+YFfh2DQf3XxKR3xjP3AUBawiIYBh/c7+FEc5oe6pDQnSQdu3002LwrL8JNBGdu4QqodI4lN7Np
7vlsgxWfmg7yYStBXnvXKjnzFhTvtAiAw/9/7YEA0hMfxfNdwmRSe/2609n0psK0H1Gxujptqbh5
4MPGuYMXYGEOhqPt+dF5Sc/f6x3lbkGZL9qB/ydyp3SxfCl3HfwTHlDjhv4DNPYizsaJ/m/0wUr8
eZpdl5mfeq/l4ZY36ETkJ9m6t15AFXYf5cq0kxmBQ6jUgsK3ayUG8Vtp9C4nkLNNsqMJCqqGNpLV
eFtlLNiGMgprK3mcKCjklBDCVFankN7ofCVwggZF8m7EdzJVhdHiwloOMFAipi0iAzVFKxbx3Hlw
dBEK+hD9ME4aCk7FngMbsOf8duvaDaMmt2ooOoNo7SfPfKbKY2m23kOsgGUyoMkVb/ut/kCLrrzz
WLc0Qg+41Z3JE1VP+LY5c/Lex+CJkZSQWNPFa4MrMCJJPGx5wvB4iZIQBPnMMav7xJAOeCIAJ/uN
2AXG7Ejw1WYI3jqDf7XhBzQ5lyERwjCK/WdMrxgBv/XFvmOx1P5nKuMyA76OAKH/PovWa4F4iQ29
yWZDYB3kNOz7b6gsPOIbcTPLqVsKYXfyxDqL8/0Yb2GKkEq5IitUZ37gHd79X2FWrZXieyRrgr6h
DzLS0ybi+W7HY92obCFs1QSnkySSgXIN3Dz8cSVHZ58CZb4Qn5UBBhC3ovxaUuTmEqEy0dhGLfCr
alWV20puT0RJyfNNDE+ACULC0gsearo/WsS9BQN6wKzR2HSb7XZQ29eips4iy9aG/AF5G2Pvra3X
5NoAekQTuO0+TRUQ2/lKrIrXamyEO5GlvOltD8djOOoHWNAnHV7VTJMFnD5+1wwM8yQq/TzG+Zoz
K8Eo5GvS+9P3lj+8U1QzQUqdM5nn+kWMe54EUTkRWchVIFZo0NWZO3/cQEGiWbpt/f+EXymb3sX8
zfEFc+b2JXLqKdS00JxGCLcwYuxwiwe9JCjGF6ABOZ/qxoG3vFgZSFOSoNNRPCooDA/6LpLwzD/H
sSpNjXzYH72+5UWr4vP0ghK5BEUtaKQuIgEjbU7uhUl/8fq9qkYS8NquC4DUTi8Nbf4RR83oKOVn
jzDDbnyVk8pxckHoUZ+EdaB3t5Yn+CQJcagcBkasxBenpxRuz8p1FqBFRWpo85nDkx8eOMenM3Eu
ijjcFLm7VyQc/TNq5tk5WJ/aYuT4OYtSprqtva7ntyLZy+AsA4sBUCuWAVeerEHH7QFAX3WxYZ6T
mlCFwB2Gv3KJ0FxPhhCKD2xS2VyVqfdxRthAb/tsOFkWBXp9vxidqpnFHyN14uHRzuLDXj/AKcsQ
HOtPdHfasllG4gh1eCE/WkfxVuIBxHMP10pTQ/Ig26pc2PYUhQ/aW6zRhEmgQifBxwQ5AbCuaDLN
8AFcjORbL+8XDAc/vhqLhx0lT06azrj9AIM6K2NKyqcXem3o+3/kBkFRuhgPxOvYwlfg4Eb4dKWb
2CaeU02GSQS5HsDzlc2RFTOvXgwU1EiBroUDD3x9XgqffL5QnvdCA2+Ks9Wjs/ts5Jm/sQ9XYrNS
S98SwOdx0gbWqv5xVujCseH5Ax7xlRcCqg+IHwFYzu3IvXlnAjO7xxGat1RUeAksa8OBwH43es9C
lQTRrgntVLtWReTrw2Nsqh3NEG8xYBSelYI9+vmwTobbru1GI8RakVZMZ/mHPf0cC31t9JPFve7P
KvzjClxlqcCyY98BcfJWmiEUyPfBR/cDqUQ2gakbsJig49/0414Hn6utk/SEdJi74tJKY1J7CM49
/8QC5kP+DpsYFi+sV7F2v+7ttUQ1D2o613Pk4SnVEdcodS0hvXY18p1hX9K0ooMamARstOcIvn4k
J6mCR0YmisL1ff2M/dDNkA18ciwfWaHJupeHLVgQU0GlJqeQ9Fj1OB9EAL0MuHVpwOZbUMm3S05y
M617DvYEwj2ucqc6giIuMXuXG1ATPp47SOKxs0zfYjehGudlxtXejekdj8FYaB5mKgKg5EJmS1Py
OO7I6Ze0T0c+j/vDcpaZy/ffu+XAD3xaNZ6HAA8ow0Zkuqft7zG6VdTsNDY7qsLZdSVpZjU7OTuy
+iTW/Nl4irOkpXR7ft78JTyhG4CJ2K2/Dw6zxulcnoZMujRZGO1ZcYg17IfAKBBNsi4pMYnIViBm
DKHvOiq3F34x4X9cKupJFnjWQfNKFg3Njb4BGpQEXBXE/0dogpWA0m4zFRTbJDo1EWUVU4JKSyFQ
9407SHLezV1m4QK2XPBiA7D10eNImvRcObV1Wr0lIFRNcJazKgag8PMbt8w3jhuhUDYZXjK/ewAR
03taPr2aFmVl4kluKELwsH0sWbnaPMpS7s87xTmzSaDdXmnzx0QiNCX1xrZK1nMoi22zJWKrrMn0
qu71MNoH+Rd3KpfUJj7+wJNozs0wIlwm/GnYzEH30FiFRLdmJ0NC6Mds6d1W4UvGVKEaW/2IncW5
j7m065rDgW6xVJvaeeilnNbrJvCRqBZQWIhtyAqlwTsOq4jaTQD3yPxtux8+ASK4Lst9V/ya0JyW
P9PiLdRvdZGc9E+/dpmGSzM84I+xuo9M4Occ2le1qG6KDVZgF5219ehyibpPyjszOIdTHpxpMht+
RdNpypj6ncXoW5ntOpcXUkDQiRQcNL2iLouzvwLcs2AXDdL5n2ZBih9xzodwALsxAvWhzwXRC6Nu
psIT3DRii0zIithvd8xTFd3gLg5NG2h2ORgzSMP65UP0vXHsG4KRv8kTgwq/2NeAnTgcm3LdG8vW
/qkw9fn/ktJbk5TV8tQ3sZWPltG6uBln9QR78d+wyUKiy2fB4KbXDMDuAZJN02tsWe6moTYdYpnS
z5JZJCOt8nIBt87jtW9rOHzYDysElcWA3EgQhF7tdZWDQTOOrTtQqMCx4aMJsGGTg1xjDUbllIHQ
8E2i2rp7dWP+rhPFv/5W0ZBNx++qPqIrZEBxT8uvDW8DQF4zEZ0rkaNI8b8gVNx4rx9MhQi39TDi
F9QKOdmOKOeLjDnK//ljlYcj2zi2/Z6CJn7jweYjkMV9LChesTZGPygHAcRbZWCe8a+ipxl+m88Y
M5WnjPtqgwcTDyIa4R7b3LQR41RGQqR+i6UbZUaM1+QsizCy0z3rBE6AUEqS17u/gmHtHi9KGNrB
6Q13ngTIN+Wqo2hje8AxG5lQCagmReE5xCxRsJoJ+tzyjJTHahEuYFsIBKOwwznWIUBiXIGf1a0v
FGG7cwKPlr3DPBYWCw0WnMYJmIJof7T5FBAZbOJAItoVLxTs0/MGu1ip7hM4ovLZWvSdM/YuZIBE
mYQV6Wd8QsorEVnUMBeuQs4eLFBMoUaOFkS2bSlfb17iC/YPxQt5z240dK3jIE6bdRSrhflijDPq
ljIo1cMcMDkSGNvpb8idQG72wvlvaYPK65SRnprUPCb+nn25Ra2mYmf4ygVDsb01Uo0XOPZXSogE
b3Uz2JLx/Gf/vGgYs0RRDtC1Y9/uXpqfSZHZ5AceUZLvhDqXSDoO6X1RH8pJ8qUAJ6VEf3Xv5PSY
hrs1zVYRTtfMrddulCzNj4CExuiV45BLOLerH4CzrNwXhfcPad8j7zGKDH8XaZgfM6h3ec68i5gJ
4BCtpG6rVi2d9N4D4aBwHTKU3PDw1ofYebqXHbyzfWEjxyAwpjLo/EWyQ4HmPPPGcpcGXBiReelm
G/CPdX0B0c+XUnfRwJujIKOfP+OEBU1BLE2cwtA2KJx5HMaTxbcJshEKwNvnpz5SXKmWpnYewGII
CRCnrVUBmkQYzSMZiDU+Q2vXny+S5M5SjOqWURVe1YgdZN2zeX/pZInUrNWmuIBv51n7xtEscn6D
1uFhL3S2EBTPOpyoK3kEJnNbmKLQKWoW/1kbrUBwMflCTfCP0WyihbK/PHF6AW5kw1TgOZ7B68jf
VqUmagrogy5I/5nqYBJTMfCua7240RctqAVTEpYYy7NmhUemEQKf2NIy2HGXJadEO4NRRrAfvTWh
rfVihmiOcP9PAd4VlIrXE3mJMVDtfk1uod7RKOvVvrrRFsp/aL+fr0stF1Gq990Bxgtz/jLScZ6q
Z5yXudyaDkKBxTvIiwwqG08Ka6bZzCcoZHyR8ka2nojbGfB3gcWLp53CwIaCakftfNB2UAnfib1A
BaPitLJN67xQK+56mKzlcu8/EeV9w2y6OCbg+YyuReHDEb1hET/dSBZShgsxG2lhKF/w+ESOUmnX
4M3NpxjnYR88apdURjf1kbVrd6xNkYzHwBiMvxfoveOTVwOAj/DYwJurb8gWxu92wYpCdhQHgWsl
HG4POJxWHSbiD6DrszCxMhNVaPsGpiqH5tDP5OiEg7os1FrsKL023cpL1EWaqvHyurjCmbbP1GzI
eonoZ+CP0wyRDVwG+VGUf+EP6/Gjxzk1FAe7ddh5x5M95iZslnn3+Cv31uVs05r+NZ4XpqZ4tcZB
up/DUjBX3fOCo9M9jTM1BgdvMNNWT8DRlGI+Rgv4cKzRxvi3gOjgctI1qiBbIHFwbjlXUfjhDYf9
RzRpN6x8JT2BDnnhpGzeiSN+PMWIUgpavNZx08QQTDRpPHLbeB7A+N3yK0bsjsnrHEDa7g4rvpea
74e2BajPByq3RiDm02ilIKuQYV/zz0+7SuiZ4ZUObj+85hJV//DfN9ko5GtOw0QTRoxBc3JOrVrg
eO+VQqDFBix5WxEbflSUY3ciqYM4KfdB7bWLnKjeWseQoLZc7T5U+WrMC0twUWpDlDU4eMI6T7CY
bEaMiPmTw9KjGTXC/ljhd5UErJMuMbTQMFBKN5Dx3chQpbfT4YVU2KhBtmejqU+i2yECT1sDERan
zIwUHDfXAxEwIJEGDxmlTim2jg74KMtvY4z6RzBL5GGqCrUwNz+2UaO/1kDbx80QU+DY9uX0Upw9
6F9W7XpNHVD9WDigdFJrTGPDL4vC5IAk/pnlasyF1hXSUolgH5aoOvQemXhNmth1cJrIzeB1hUM9
hTXh6LBo4GH7hwD5Vae3N87zEMwitusIOTinsMa5PlhL4coQqiTGFrrmEfjZBvtm2TW8xEb2JoPe
/kdcaUjUFbXUGYGLwQO4sk5wnQLhsKtt5ie3fyl6vok+wADLsmj2nsQeO1eQ7NhNYOZ57jJCUrFD
jBkukFNufhZltjKR+T46RqNbTd7/yjNSGrCbJz0nE8hXicbQJx2vsvJEWFK4sRJD5VVDKam0ZmjZ
Ko+UceUKRaN44ABdsa+jgYITm7LIr8A6kpQWaBnej1GjiBJuPy2nP1LLG/3/AgcnBNMUSSzTjzDU
g8epx1uBATY1ngQvV4bN4RSupNUts7p6FmPjAsZPKDBgBPRC14162ejNdaN6Ub0k15rXCctBmTrK
PjqFCfRzr4rQROS4UirVpmtbzz9Jv7R42tDr7aLpGTfx4t5vBPMD2rz3h14rSQU/nZAyBXrx2syT
cDbvMQNn/HQohLwjf0GXBW3OXsqC8g0fPRYm8IYNeHBlxoejS/3in5xlqB+usUG8c/ZxBj5KhIYe
rk7nQ6rXNixrTzAtG6oEkUbfWbBvOVEX3lklf/02W5uW7rGgVsLCHLFMbCS5JRRI4UTxbwrfk6zd
067zqT4h0aY8vlZ1MjPuOqEZGvCGiOraHpBcR3wd0E5LexL9YSI6LsxS7J7HnI3jZ2zEO6/wtVPR
kjL828Kft3i2PBhUU1D0V4xWPP8taY8WZmXEcnb0QC2U3OyrGXitgx8XwNLiTgn2BxQD4H93slle
g0un3Ku54uXOeBFIxek/yiJgKmrAYDf6+yrQh1LN5y3EGsTNIVidf9Pspx78MmBLH/9qbbbEs7b5
GUaIl2ZN5pkAHzJSjuo4Mlg/tlbpfSSBmYzhltJWaB05j1TjxNAjyl35qMZoiu5cW23OIvfidVvd
9PpBWMnjVlLvPleGaySiHS/ZVHKjjx1z3VdiNkd3Pj+kKQ43mG8siFPAeruKuOmQox4Sd0froIQm
3DzIbEwgcB3Iwgg3wanfTmLyA1rmGJ0u9lmgVyjIUATmEbnfzbXvGrGiVYszJgA4kBv5NSbWK6Cr
GrO6chWy/+epvnARmZS8uCsopMiuCbuHtg9bgWKCQt9KgIVfmhRzASeGyG7tg/LzZLWgd4F/FIGf
lSCDmtL+Tuf+OUvrzC5m5LuOYBd9pzQgapDJw4aJvIEQBeDIF3Z34f2ds1cP9TWpN2teLaFSUNvI
9A549h1HqD5waB8QvYGGFC2rcyDLSZU9ZWTJ9nELm9TYIMlQxw9Rbb3tKfCmwFbuT/Vm2DmBOjnn
mX5jr4wjsJLuUCtTdIA1yWsniOqaybEMJ9QuEN3CUAnI+5isUMjIvPfyt6lvGIXPx+iP0VsGPxfa
iA9rNt3GAWW8bpWjDnnw9gW/fvsUzX4cCMcGOgts9Q4Slnw8CV4k/PybH8peV4kKws3eL5rFcm+2
8aAQ+oi+9A7dy3Bj5LkpyNskXLHh72cX1SUfgAx9LcR4POdWqXhxp3QgxDlzID+N9UKp+A8r5Dmh
bkxlreReo1Ms24V6u7NAxjHD5avcLDPl7dggXv7fQLMPOVJ9Yf66QSQgMOOkDMhWIX3bn80RuhLn
XCW/A3lJ3ulN03OblmX+JaB42nSljF8uI5bBWTVDrsgx6WMv/CV2hhAEc0qCjZibiZysoDRsPyYv
yWAvrsAXAKAg+78iuAz28AIt0wM3KlCNEePvl0V9tyeDx3q0iDLj18yGqOXnN1DbcNCvXh1uka+N
Hs/mkpWuQaFgEpMOoxpaCdD0WsRE62rIBjf24Eo4p+xrqlI4w06Eke99IrfRFyZgf+K6SDXjC043
r5NW4AoG84DcVnv6ZO6scsGjGG4xSwPmA2u2fEg+XE9frmaHImSqDrKdvH1K2dWEyeMH4nM/+EIe
vUvwiprQZzAw28GNrbuhiXABovOPGR68/eXVNBMrbAj0oqiG06JFpmUcFulqHVq/x+wDKI1qMUCi
ICMGvBihg/xf8/PjV32aNBU23Q4RFdxtashNzG+brmg7Q0LSEhV16mDcH6RRrszwl3bS24TLXBLt
hughhB2OAxq80Y33hUuRtvLxk6qEeu//b19oWIumq1r5Mt/ip19q1u9EeposI0/DU5FTZkJ+vyZu
azudss1zMd7K4DGDunAOrKimoKRoWboGmQb/N1sUgFbODI+n/kK4LJSgoVL+1EA4/JFKKn3TwDS+
lf8/zoJAB2mXroAL8NYJ+C56av6ORdtdUw29xU4iionLUll80V6UW/MMmj+J5v1NsMAAnhmGrdMq
UWzi/5yhlpSXEM1mu8ewfvve7ZuIqAPTaAI3kw2kItk7l5U4nhWsEtPmYkyoTeJ3xXTcv5Vf7N2V
YjqCC9imCcrxE2svSuY8AI55bh/O4HVRZ91UyZy9iwJt5hiIiqRZAuaNi1TQiGS/AVrfnDtTJZME
eNG1ZH0ZSOArF40neOkjuUvdlcGHE05Ac34BAcvY9LcaQ0vSMbc7EhCNtkz7jhJyQJWP1uMWXqV0
/wDxXzhEle/MJ9o/bk/slH0VTsaOjhOprbS2BLn0E+/xwBFd4oXmy5X7a1XWc5g8YHXV0C/yYzLg
/Dw+vhJ8WI4n0Ew4egakTyyYYGnkgIB/yjKIzCRAwrOCmYYtS2jk8heY9KMyEfAI+sRQ8kZF53qD
kiq1GLxmGNCd/NvIrghmtinJEaTGh6KuKN1qxEfaq9ce4YoPyOrS6Ajyv4tUIetxXHX5h+9PT3qH
WB9IWyC5aEgu3+kJfMldkr4HrqnBoPKvSCEJD3P6Cqh9HJmW4CTnAOObfsh+TfHs1f5l1mANPmPa
QYgKm7T4KqdPUHocoTn9EB2Xt6gsp7s87f7CHFNgMEevB1/vNV16bIfdxtFwKco2E9GqZovTZp3H
v6+Ia1bYz9sO+iJ12Q6Vt7gywnJG06pV3uN9lDDH6gkOSDQjlrHED+5Bg78t+6SiULOsrDysQGRV
AklMtYyZuOIfhr72iWT0w7RSVShXEQPPAm1TE0YVB+0ywhoUjM2ThYkGCwoGSyqPjlk4/7xMFP0r
AU49aRo+7DZWs91GBMfbBcGfzFywE8dhd6nMfsqZbXmwiVzhy67UdNgxxRPuUQGh821DVvcB9vjg
M6wnOL3EOyMZsgJuvFpSEu8WkYWfy5vNMhGDIm+7i6x+D+g8pgfxfGWIYhoBZALtQdD+G+R6JMxT
sy9sOVL1i2XzLj1Xv7EcFkX51HMlZFXZBmk+IietRclJMrEupsKs+ykZnpZgno/V/s24O7OuG1Ow
f5pH3yNHgMctI/KjOdP4f5Po6n8DrpLpUYuxlnAeYbs69uyN4/awWTvvRULNfVidzOKk+h891JSD
L79oAECFOfXcJ4glUhV2CH7MSUCO9Li0pic7v1vqISf6LgSrZQNobKgVBo0+6O1Xs32u1oQDua3s
6BwT306sT1ayIWThZ0shEk+5BVgWnWoCYoovW8UPFKdztcwUycBFjSx/wIPyeR4IJbKJAOfu28GY
fIPUoZ+NB6lFh/2pGGMOZE0CAJGd0Q7iKHowZLj1kjsMyM5luww5qVp60YrdLCa2wS0IKh54qRAt
aSRH2GQsdyhPoOI3RXgwp+AnYxMFA/oX+UPprjm5aFv7w1hjCwbq6Cs/Mjt4PACEeBP4btqU2m66
SieALD/SfYlzydl0AhNcq+1gRdWw8D4Y8m/9wVfdlQaKdZcuuo5ZY+Y6XA5k1DDKSSv4J8KNezx1
NBpdkKYgwpAv2qx5U1NHUquG09dkJVMImSzUjGSvOqAVVB9wnOzobp9X6yL/IiOUOIJwzYLDl5pM
tSsB5faD62Sm0kONZ3haqO7YnqyfAjfaXIVq0HwvPp7vUgBAtBSLK5csVPdPpxsQp3n5oMHCGsBx
9KaQ3RJcpvhuxpb66/75EwnbrLlkjiTGsBuauVyWdS+1kjB9AvRHjdIbxmu1CfmYs2PwUa1H59q8
m+uJXqUsXAT1Vxd+6qH5KVsUIJgUNOTO6BJz6ji4TaBqKgpDlzOAUcoYPfEIJpzvbfT4CtUNE+L0
nNn8khpzeK+C8VU6adH+oLEGwW+1ippRiaHbr3ujbdYKunP5IrlnoTHuH2GzMHuBKJzTllaz0lX6
jptBHyCfQpONysxlX4mJMRkSIcNryS9aHOk0nNZBvvT2CiMLk4+uryO1zbZos4Sb7mf8QABCAu+P
P/Avxf5utGeS94WdcaaYvguoofow1MG+hbA4vgPh19YYdt+gRSM0mTbTpgRD512X8UbB8u//q6k6
FC1IwcD2aS0Ez2CuH027KEL2IMBIHnVyeKKn+7wbTuPEmzx556LJaInHs3RhLhjzpsCXDf52N5Dm
1vaU9n2uav0T2JZIW0Mn693YaR655hfe5Uqj2PYHsP4SU6/LO/ihwZlX8s3dkbXExGJykJIkqDar
FyBcgd94MfEqDBqUJ21BHSlxM2xBE6s6mpL+AJO7aoIfWLlYFuPEkVlftr+MIQ5hw3yPrOwkWyZ2
s/+r19YMuljP+S+riAhDkpfCDK2fLsF4GNIS5zs7EsKD/BrAEFsPAMZIuOImWsdIU30bSfmp5Rw0
V2o4J5mqQvtBzY5N5t/aLqKLhLzZ11IaSaK4vogcXOotWyO9vJ5st8UA0VSy0+1RBRHOW40jelm2
ej6EYFJfJXxGosOjArbOaaIepuzPYpLvMmoNNpSzP/6EwwamiLUyjMRpNRjZ8dUq/8TcYfiE+itz
qM0TAO5U4hqir5zms2hU8wtmtXC+K4wxkN7MMxYVc7I/DmRaFGqV173Ti7Zt0hJcmsXsoRuDsjcn
wOFcFxU6zEQGopfCAbBvpcKGP7WIvHM/RoJn1QxZ3LzvGsuQRLzwyL1P7WTUH76d2YhHN7SMnZul
I2Wv+dlxK7VC82X1RHDN8hRqCgIM+v6roGoMpDAlMERat0uOg6a+XFyh+CKh5ZeyeQxEvyLLofAc
5TCO6vxuUw7JsNs0DxA//mPB+62BdX5lRi97vJWSlMEN5RlcebAL02RUFa9WLFU82d2xCNdO31se
mOCI8bH+zXtRrtBpExCIor/Rp2W+Zci499sOmkUR/+jtIy30x0GRA8XX8Ke7Od6L/bHU5KiLg/QP
MNFObO2yq6kaeBdc23+qxEBo97H4T1e37x78iBlu1yMFKE2P94FyWLkTRfacO1LZxRebjtSPqFy1
1YFTNuIIPEwUul68PT7sMOjp4yhpFANKqBjQMAVvzxR4AQ0B5QgsJ/XEw3Uaawt715qENc0D7CbI
ftim0WAEWlY3s/DLxDT29+n41PD4J5xRfCC3VIAJJ6A0LN0/XGUllwkWvKesAu75+cTGMKnf/6NJ
bM8MH5jKGCvuFEvQYPc7JptQmGxgFRdlTLstLFc7VK7WoaJOmGAEfKphmlsCcH7IiM0W9UtPe3IL
2xd1Fn0OoLTySgaheRVagdEh+9U/TV9CMnkgsewXuLUtlbAKlbzH3tN4xkJg8QX8as60N0j4Mwuw
0QDqNiV3WNxTqxVPLfkBQrkHy0SPchakXaWDEzYUPKbheQ+me+bmL2xqRTh+Z/W1qHPWJJXxRWTv
e6VFW1/lpO7Bx06cbuEOgZVImY04p07pi6Gl367/IDk8Vo3nXqaKZ3EC1UD8JQYHQBZrMA82wZhu
AH3bRaLxwLQFzHDUnXT2naFiwZ8K4dcyfJldw2nhbsGEvpjjP/vIC9C5pEf9FdV7ZJ3DdAhRdAN7
TBuZ0FCBxjR5po7JGyKPHkqEZjP1eF1R8Uk54am/8R5PJ67xhOYCoeV41q7t6KJ0ZufUPFfimcyi
jkovEnoAOAsIoNHIwA5SArw3605y/JguXzUrotnVUu+NUX21GDUbgesY/8suNKrXFq2cYr9Sw9LX
WP2P56iy3Q5Kg3wGLb/YV1XU9lrNcPpcZtrx6bU55TXDSLbjjkH5GGCH0+5UHRWGxRiFvnFou3px
GdnsxdycsrlOXToaOyD+7/ESUZjggKNEM1C6uIxA3bNRPc7KeArIuGqbk7QKR1FRyTegdxg9BKs/
IuQAGxW2a3bcIbiKYrhZwiw1Lm4oOqvU9RzPKKtoOr9DzfLOx7DzHcXADS0kkWXVxPqSaCPYKYVw
rTYOwIaAovpBb9ex5ic2eFq+LXFGxDxwW9aN2mucpCXAR4FtiuxBY6SbIAwhZZ4YdNmVNojMgTah
6/lpCmzsGijseF6R62ipRvUEt0fLB0rYq+Nf/QbSnbsqtxz4udX8wUZWe4Im9OpXIrg6+ESh4AjK
4IILOlBzKZLBFsQ9D2dCqFf8YPqXhOlNiLicrfe2xsTZmao3L/WhleEkBG/HNyQiyEoOgElYF+m1
R4A4/0mgR7DhxqBcjHXhRTLTdbLooBN0Zi5j4a8yAIlBYPlN9SDIWKFfqKBY4QcdT9aAMoORyaLw
OF0VzXrKszcMvUy2988a7F06TmJsQ7nOS1u8KIq3JxGPqFWifPpEXnfVcoezo1OhvMl8UFdvNR35
W6xQ2/rG0ndR9T62R5Sgg47e1dHJ9z380o6NhM52TbSpMssAH5uI1ZS8PKDWfKD7kYz5a+nlrbuK
wWPFoLbIf/72ytVCdTqz8LV5QJkH5Pt5MOquktsi4etc4AMFMSHzLWh1rNVUFDq+g40foW/dVQ+A
u/Agx8q4NKktm8Ig8c30RevhIpdLctVG3V0lxlY6c9rT6YC2pBOd28V6HKR5c7NTdj820rJPh/5/
wqlnrnCv7NIVuCB4J/PVHwsE+cZkMTf8V2Oo25GDLQfakreCZ4QzajMcto4/AMcukFLvWxQNdM5e
gAlGpX4QjJ2BKUO9v9XMEavFkT5Tu34lHp9EhGULCVM2Fa+QchmkGeg8b66vfwBIrcJ0BgjXeikO
TNiO82GiQGlx+hzK90O8NaSwMaECqZFUcKJxmwujIoFywPpjrAswuoNyVbCT+thlFsz5u+pjHI1B
L3IA0SiiZi085HZKcrSH5Nzi68UkGXga13MM3RDmK7rmuyi4N5FNdsdCY+rt7ze2WPbXaqWIu7g0
TTDIlvw0RXW9qlmH5m+Ah9C6kkJ62MCETxHlMF073Xw/R9T/YPk1aETr3MNwAhhH7PPpAW1Y5nwZ
5kMjaF6V7A5fWrUr8I1HggyaQJodd5YKuJdjtoekEx6UsTBVC/FINsJJXm1n8fV1pdPJQxHKQsaV
9X1BZ9TgONe1q05awAxzmT3jhSo1nVGNgiRlip42uI9zMSIU2qsTVOUU4hYpiAJ9ayGCkwDVy+nh
uEmuY6+tNHpuJOKq6S9cg61xylXCozba9R5NH8QBu/d2P4nixYnmFN0u9v+huyLL49B8FPHuNAWv
aq28fXkLNsVnXS4QIOkKWZ1/BZKvUwM79AeZx+bQ8Ta6u9V/rImIkl4qq0qDcaEvvNHw7805roIV
p6qeIQJNwmly2jWggF2v5/XtbEMamKY45/Lkd57fizMxf7lEx/VsY5z8bJghUMKduLdvtDvYP0MO
3vN/6Lz6bUdAa9mKkIu1PxdUhn4XbOmBvpVNRKC1ScIdDHkLvct8h85Ss6WCdatdGna2PU4bdDi/
NvXqlOwA4vo9dI9Er9DxZKQhwlHRtn3c8AdaWHUbYvAfpQiMcurMXeyblsanvgM+Hkk4vUS6EWtu
e3nC616RNlbBkmvo3KNCSm+B1GgWvVUn4gPuKVFrQBbXUzzS6WLV0y2LlrYFRjJwW/+osbeszmgR
D8OmW6fdXfUwXottmg2O3ApTi2y9IRQi2xjiXVceRQw+/aml8Bqdrkayobu1EfbwLkYWVTm0OdQN
wE6nW3ZpgAGdhGHVzWr8QTroViSzD924HZfNEFpP4In9NX/Ea4h2SULKqH80RZ6VJXKG55ytsWVn
a2wuJFfuGCVHZdHe1yOLz6Pui6SxNA9n93umtz4Yt/x/zWLXnqjOVvz038ZaXSxXyYh8IYAeNr1z
NfUlg6gZTE9P8DkZSqxzKTuzjMley1zStFL6kCK7Z9NYkqLeE/K0rHUseuWGwtAEHPOz6xEhCGaq
t1sYqodHsJV0OakyGRQ1pCksMqk2d/kWTIGiDsOIg5rIhrD2ORyksGAAg9EMiDSOY4tdrA75+Qfe
k5Njp6UYc+vB8Tc46gMTCK1vQ1IVNcV4RQmwNgSjP4po7BGtXuuuKhj2s45/h/+oE+X6iY8K41uX
WTycHYK/mx26mYNrdj+PapeXxlsXq55IB+cntmYZLewANflUfLUx1hhzYowIX7+yrV5Wo81r//VQ
xcHLESCc6k4lwptDwRGpJgm/vYgGL7SShKJwWQ4NjuiQ2iHqWORtmH6RkoD0sBITYh6zypg1Wy7z
kDbjG7WqI1EgCgmCX/z/m2yGJG1yBDOzgbrpWeMah0Qwwtp7ooxIMLlL3ex8h05DXgLfZquDlV/b
AN7IAH8g+ypICl67Ezbpw41OAIfEyxG7Npi8rhq4mvWU762hZxGbS3uHLNVldCuone3ixq8QdfS8
RfcN8ZLn4iXLF55bsKzK3D4WD2nQQyR1OGDPkyYO218+5IyWZnzD0z7W2xD8TcAI0JKO7cJyjqQu
dmxE/PAYspAJ36YtX9rwYkQ6oBl+V+/0LN2vl3vR7mevfLyPhTumcqVQ2Qq2VqhTIZN5CU4+rVfD
e/dV0TRdN1iJb9evyrUVRNn8baV1RYNTABVJ9duejzgxMnqtYVViEcyNmZHlBWzKTNifJunJvgNP
k391tV2/GxrDD5FTRHKFEUKWFYA86qmYM/+z3ZXVQl5eiMmVhQFn8QNYL9nLL2ZvoJD8FsASeh/0
n42Vz93ujuQoFNoXMB1DBT+JYvke59ENbq/YU0KWfRfcjWdqwF2rhpFZlLGU9Z8g4jOVFNu7ySdL
iYr5dawzRUDRVxo5YeyIc8VCqGmCzP54eGgrgN3QENriGOPX6kyV9xAn+KhNFIB5FZjpDsFg2Jos
jdkiVoaKbDZG9RKjuOPwLfQkTvfTVonqMk9lokVnCAly8Gu8YtQ+JfqLwljAUJ5qCIXlw/Y6/c50
GA1K/EunTlWdOgC6cmZsnBu3aG+u/OyhFi/RqNVlvrebyB3kpHMe2XOFrA8KH8pDd45avrc9OhMC
y0qTwYGdenWkPYsx3UL/HC/KRcTP1EZcbRe1WN97IeQndZ2eUMa3AE7qkTB3aChvF+xq3e7Jl+UX
weK8g4hbKlbKwoKfPLbtr6M0Q6ttgjVoAG0s9eefZ3o8mORoAs5F0HOVElTr9w/G5KE/6vuCKP7q
9r6CCxbj+XcUgY28rCg6Ki7cBj95tstCwE9TOkUnjntH3nsjScfG8zACoJQh9gFzDzQGkmv3/ivQ
T77abUVfX4lqXdAWXumC37+btRdJxAD2Q3zAcppfOJQdBxrsJVKYHoUDEsyr7dvDXCCFBa0WWNFj
gMww/wK/eKuj+Rn+kzZuRY/ZmRbix1VUTcKLJ4J5xWuLOXraSLChQ9qKCrqPMG85v/ASdjQPvq7R
2lfq1BJKkFIFkhE8hz6+9gUnN84C6+ThaNR4Uey02BOYfLihd3kBTGYGntmXjCNm4u9BhSBrWieS
hxTulu557ZdaTjk0X/ZYqcHB1kXcXQm7EzLvEkAG41o4W/N8PwxJ5bFmU1qrSUAhrXvmBD1V0/VR
nUTdTAHBRqIlayX7u7iPSCWy88nvsTx/uFHidsQ2prtHoXliikUXKpG8UhYquD3k8odGHF9s/Ajn
zFAYL7McYlXYyPi0F7RbZq2ehCv6RVUYnXnYczEclIRusRjZGVmUtpjhj2/NBqMnwi3iKtztRYME
tMk2Uw6ZwfWY2kjMGgR6gUWyohw8gCo8YXmTgm33GwjXp8q/eo93tHvMAxim3kouSCz04hUkGgTZ
A27zxLKynkiUP5CYqcx7PTlvkWcmHsIkdNCxylvikUupcmDheXp2UVM8wusber7DU8QdjeC7pMAe
gNNiM7t2KuM2yqSIm/+5fnyUQcEbPQr9dZI5HqX1CNhKmHY3sp1RauWsZXWB98LLch47f77jFlVc
d0dZs0rL/x3ApluPBI6FIC4FW+tw0fBCCdbVliYlbO9tVfN2KC3ZvoOguQVl5WcwvYW6bChAXljH
pz7btLh528hkk13MuZEUnN2ySTVwgZkC2LZRW97BtUZ3bDhwoayc/jtFyl+KqUxW21tlpZf+rNPV
ls5DkNAUMg+IVSQlkP+gX8SEKibLE08Mkj1bUEUd8r1z4/grCGjfztuUCZhNg9OGrnz6HgdL8P5L
0Wn9m6RhOLYWSYPCgjKKgN2TjJNr6jgqpol9w+KL91mAn86OmBtPqdS8tmn0Y/wBbzlFeFHX+I1k
QaODE6iHNll5usSjbYajmY7BJW8YW7LtSJ3mneAj2lkjfVMLrD5TGU3auUaWzXpL7Fe/1udIXJfm
HTJ76595dyN2b5Iza02TkXeLxZWEwhb5eg9aVLbYllNZIIexjxlOpyZniiebTj/V6sOMPC3W/6R0
HqYcCvxz6qAqBsbYZJ5bnER7hdX+dTuivMlGqoLggaI8wSBxd7JcWaPYwjl/1H9wrBmFgbmoCmZQ
aAOyScqNFB6PSb58f1IYtXPaK0E5vstMH7JuSCtnlqNtotLzQqIbE3ghr7Icet+FO+N4yAwPk4I0
ypJlpQb7db5lRKRkXMa0qJI9o6m7p3W4ByAhrU9DsLE/EKNJavaMeTs5dkWkEuQZhmKou2dIR1e3
K3zjz0GUN/mKtT97L6YfuFhUc9lk8qBmqM+VmNo7kNafxS3bOgbE+l0/poOTYx8uteFnXosw1QM4
wnICBEJixPWFyiQZhZpo0scdhuKvGJOXciunvNtL3gF4+Zx5sE2UPOerJ0O8h8AnqZwCgHTnR6LR
cfO0TfS3M1XZkotEyOJ949pVKzL52Z+0TyaDs9uNWHC84L6Tkyqy7L0C7yrjctIenaae59Qv3Xtn
343yM2mdoouxYERkIvhfCxHQxNOWIubXNU5JGCOIZcT4rFiMRDbftt37aAdFN6mHXBouQanJsnu9
xpYxc2+CMSIiebG9QF5iW0DyGN/XxkbWk3ipej2BkchYId0uxhnomB3O05OvPF5KtgIIy0yTiMuq
84hxV5v4Frkj5X7Cd1IhZ4oIm6YraPCJPY9VH+5BnGvtO89r0US5rdSDORYdlirl4hmIvr6qHo4x
SJdUoWoMW+2vvwM2VEWZmtEcNgnZlPdOwv+4SluclLjagQF7g2ltASXrNKNLNOJ/pH59URnQHPfw
/VOBkY76z12X1zfc35eUPmXPn3FjpEPnTQLbqt3XgyzRgb8v11vY6rQjyPMFVmrCDSjmqteLuWJi
MxxeJNDwer8vNBYPWcqngzdgCgALW3Zve0YvpP4g8wAO8eeuZuaYxUwP1GeJ/e4CLBZna1itvG9m
gmK5SczajtNgL1clntfwll+388IQCSox2CdwhqL/0K+kiAhRDtcpwTlE3HIscQzTwtx5Z64i9j/y
knrOEwUze+6+tScTQQBO5ZIvUxNmZuMaSQcz8zfOokEgmVZsDoY1CiFCHbNU54kam79nFu54Hles
8RiU8LMRGgFRP5MYlmJDEXTLcr0Q3SS9Uaj4A5Bkdd4qMfko87HmVzTip8JxqAUtMP8vdrVmnMmf
Wh1Dt6Z1Xqqt63rN3STx6gjV7aUI1zCXApcLzDasPvSp3WzcDTJvOw61ICpf/Ij/TGfWRKndhoOa
kRnQoSS2wmh/lStx8DsW3GSXKAnVKWlCPwz/emaEooIqfNTiauRD/x9YirYuBBRtPI+BGFdUyEqu
HqJbR7bE9XPc/V7V/T5aSzu16VIbtO6dSXLiXWKAJlMZqjl8GPzxWSkPeOjo/B1c9EQpgzCOfViN
0PUAnpcJWQKBKaBUIsVKWxbhyorZfczFNkMdpi5hTB/Xs6UdC2WIa6YcZYz9NNTzA6E3ExxYsbuN
sIuXUICM/msH8F5XkOTPD48vqrKlrJ3Ib3m3148/4JT5J2fZwjh3iGz886Td/EphbdUYRybbhQ5E
a4N8PI5hpvls6yq/gkfkn23vk1fHL8T8FDRHNH6KPGbxbVO7t3uGy0vQdpedBguQkq0R7kf2gEC+
xbSeflbeLF+cwpJp3kSWWShTeyHe22YEdQzP8m5XqNxkYGRWxeq63yRDe1ZwkqDRHcnX+pnDl08B
CMhCAnQYTSK0GPEgZyvMwACsMHkUIF+H9VITCuaiwfRRdDJJbD7yvHSBbgo0ykooSTnABUzZc14S
bB8hfjJlJAVAcKQvT6XLgnsXFpBLcPz7ABxbc71mko+K1ssC7PAinwdTPyeY3A0EfSrtCiBGlAu0
sO/3dworQ+aKM/kb1nSslip/4zbYKksVMo4AuQENSO4Z7XSVoKZFTP7mV/43pvkbjY9x0uZJl6hX
84lMQhEaGu02/z8TCiuFTbne8ECFOkkJStko7uU0Xq99nrg6AcgTGzqbDx6Vzj3plrD7Q6elv2L0
a5ikHOlhRgVoK4Nmus7g224mASV6/+Av1pX2SzkyVh/65S4b1Dzvpxe57PBzHlgbFJKgeeppVjbq
XLBCuWywA+CMmXVG24lcw9knoS7TY6VUtQ5c62r6HenIe+DOX3vMfLeNAF6u4l49JcnAMnmbF7dl
G4sooOemM5PPmgEBeJ6dMlDY6FIDCWNJdSNjMonGaiqYHm3dJoh2/2ItIXbvU3WDXpDqgYY+sP8T
4rEDzWnWI+irl97f/DgEY73fKbBs5QNWXXL70jz7C+ksEHcwv/KZZmre3BmHu5du0zTS/HmAbvKY
ElNmZHbd1993nCyHXryTGYaG3FSm14jAEBMhgckBCrpqSmnWgo7sD+Lls92sPjqgHMq1UJJ++yNJ
JAd+Siv+kon02ilvdQ2mnl6ZCgkfvxuJBSdsKYosJU2h+TwHWVVrlkXFmh1mgB14YeJu/4L/BLNH
hZIaiI1yD83k/65RJ6RZ7AdqYgR8KuqwFRD6JtQhOgrKnIj46V9Z6zJDL2B1vULVrKeoHJC0sFtY
Bi7DTRYfRhfTlQySmU0uLEfsvNgemhH19B8CaSV6kTAfa0fymTeXs2hqdDnHHuMvpQgbbfdVYacp
87M+NrqxhBSRLwn6BJ6oTxt6eX8cG9pHlMsmcY61lDyNf+27xZzjAWH5TSm7me82UkkSMmDUWYns
TZNcph9yXakfIjFbAR3+nz6f+tt9H6Np1H2/nbtEceo+WkYqp9Y1WaU7rPtYm871uELVf2YS0bdu
t7+MryC1EGsG5G30uUSb6K4yVUektbo7ZocNXSBzGSnrYFeGmikZr3Tb25SEzfyUXj6593fLXCYc
XDLV9wGmqcWNggdIsBX37ESnLKoHRYZauIvGdFOdcJd7uUH4PLrhnwzYKr4GW9ZUpnyF2ik4qIbU
9xj4jaMWIx+ZMqNKpdHCQSp2GC/Dkjpifnj7BAQLYHHXfnoQavMY6lXq4VvVPmfpVDZ+7dUnaxIA
mbJnRNfbBKAoOMg5mbHKzGVJ+xp3kZWhVt5JJLSNWPyQZFZBSTeYezCnWkDAOEx2PG2RbR4F9saC
VyaGVtu2vVHHiNVz+7hFCUdkCGZ4odc38LkpZn9GbzZ2r4GPegps7k5JhDXz315qzjpIzxwRmC9C
9AFYygM82Pj4MvHQ5pOAN4Er20JlXGdaIRquggckYWcUC2bkuPi0QoifwympnX/M7MR3jki+F/fa
g/ZT10KSg4fa4gViaYM4fTZGv5rz67YVPAmvnBb8Tu+XuLI+2qaMT19yLS5JlDHKN1ZS9a150Spz
GJPYAtCOe9wxSes7Pdf+NueDnGafmrkF1fwEk/5YX1LzKHohNZseSUrckq6xDr2mvGqZcsygJkS2
YuJoz1uRgeO2W2uxopPCo+BwOh3GtQtVoM6RJOgFcEfiVLfubWJ9eiQLla6CdCpFGtHCqDDL/XTy
suDw/S8JbPKx1mTSm8EQ5fmlNdp6gcTIl7TiIs6V4dmS1HeRaffFGkgMx9QRXHhFd92S/LjL/gET
YxY8ndsQN6EchZkYGELSM+hNmYDdXEZznAIus19fjHcRh7s4Nj0XsSn7T5nrEb70JqNoVWFub8VI
/xpwKC4DtUfITZYt1zDv1ya6Ldn6QPZUDBof+2dYrzAKi85Bm3YNgqRCypbVMIlOU/OQvnKnYj5u
CPmWaIYu8hAwARJxrRg+yhmoYEw09f7+0zDx8zMkSkr7pULUG554E0kY6GXEY+ocWWkkrlSUlpB0
820+qAF5ldHh8/SnRa3oK+AIo9jo4eD0nqCQJZrGfCAbfxqQboFqq/g3x/JZa++naSuREHO38f2M
gJuu4xQwBhhfTcAPb5Q+43vg1wFtbz3ITrt4vYX4kGPfTWkc1u5jCZpMF4Hqlq78MDH3WdyqVI/z
y1K9wbXWoPiYLuebkzH9qnZRpPPmv4YDT2O00/VMwU13SQgBLkP6jvU1lFSXmDOryd4O0lOAVhMu
CjvrTgCjDUMlR7Gu4VnlcFLTPA8fA0iKMgYupnRQxcNMIaLv5qyHbU2KZZbPbQm8tShiXr1PNzGi
0lYfaAdQbCWBfBvtys9PGf5jPxssnp0WV7vG4MRy7Uh078rB9k/WnfNouL5qWSV994txsGNq7Imk
QaHnSwHab6kwrINgp8zbEp1/bUtzgdXwQoiIgi2VOfSfZijM2H2853rW5EGpeTImXgUb70mEjHB/
6dF4GX4W87qHj+4t81C8frDkYaO9RFzyFXwI4oVM66j7rhHyH6PEY2YtFD1LYeYJ8F7f5a+UdlSX
lNrWoTAyoneexyPoQ74LLzKLB3Pci7pDHpSPdQQ64TBquBJpKLVxlzW+GwvWLQYttiMkleZ//EYZ
vEBeBBOZPaJuuUxICcODo3Fpq/EN3Rh4ErPYGdw+dsBA/cOqNn5e4wZYbM3oJ5WgFW1q2oEqa6wO
PG+6EY9N1eWF6d8DTMWf5aupvGqMLB3CmC9ExWnzm/cYblCtgE+BWYoCXmtD5UNmgjyu+1Mm7kAb
UraG2y3VyOceen8DOIzKt/sDAycrSS7bNJN6wXy4o2Yq7MUklZFYFhcd88EGgLHa3YrwBorB4LhI
jfSlPzA2oEg0dlxmx0rojSsp6pEV2L1f/cLM96sJyieGMW4pibjpkwzChBWJwXzU89wPrOneoJwQ
Z/M/dWOMVi7UNBzgzs9HSnYuN32lapjPco95bMuopWLMJsBUvo7rMHzM8pJRPeFlU/TxA7MAZo/2
n8baSrzAob+WgDB2KD0W2r+i883MLtB4IifKvSyP94W3XD5QAzew9Vjvu+iUrQBJFyT9GDNTsCd7
v07jF8tIHM0cpm3CrohE8Gjv+TDEPRfwBu6olqZDSHugYY0IDnnFCP/I1T0lcpzf/k8my7xfctRl
nHPAu7nK7Z7Jhe44muYv5lS10kUafVfizqsgMSN6y1KVJOhD8Hda6xS5w+gWndhp5+/dD4Rud7q4
s/l6oI5lznmWdbkvejwlDmDFhH8Wtq7fgp87WKPXAhRaMOJ8URZZ0/Se1B5F9HHLq6CI0rfrL+iP
xcrB6gGhtZ4wfRntSyyt3LUVJ/KCSovsaDONclp/OfLW/eb3O9oRbs8ZI5+OBQPZalnXxcidK8Sl
vHNQiGA6w21o72u6vLf+OAt1IdugcwcFNMJKH3zqC3inLyjz8GXkjsnuT29LaknyNMg2LKTwU3UE
7P6K2x1cV2cwEBkON9dHL8Cf92CmB5L7qLj7rSTVloLRucOodCHIlxiJlzExldRsE585qkhnSjaI
paCp1TTZq0l8WreS1h1mta1VECVnCZ41fZdAkXdembQjQ78QCYK/C5Tyfin/VVvucof+iVkRL7wC
eZ88Ogr2Rn1n84V7fXDbV+7vWTP6rsmKEpnibqYe9ye6BxChFIJvuBc++5iBSXCtB8eQxIq213XJ
NHuYsP0swBBgi3uEnMbQnisjj6ou3XrfVc/nFdlpquy379VvcOfwsgKi7f33JZ0ITvzFtdYS1KAI
fSYoGpBw/s4yedI2M2YLh5y+90nCeuaq6mIeszW+zU9KXPxUNPNFYlnrTmPcVGaEEgSIDiDxJpYc
xxKbs1f//1kZA4bfN22hcyuM9VhyC/c1Vn5vF3cH3RE9CIn6KeeRE5DU5lA7quOIi0UNnPL/zfhk
oj6XlFQFv4lu6kYvVkw4YvKz4kSJASn78P5pn0lOzMCu+Wsh5jxfP7yUxnXghkCvedPR4SBww2nQ
Ts0bgtqeX0eB0LvPhxgYASBfJVFUoOSHPonGbBvmC7hFmoz+ilZ9pwCKLjgKKEU9I+0CCTTu75pI
hrW97Ve9rZK3MDdFMWTNh9x3PZPjN+0DTAy2bcjhi++76qcyc7QrjAmhwVzdJz147eNRkkVH/lCz
MSBptZuJp3MdjB4v7GCQ1tDYLq854LgK/mQAUaPPIDOkoGgjlWXXGC78a/Ous6OT4suQsEoHdrRY
Go3Yaf1bB/2zoUYHneY142RLqqZ+MQMZriXbCLBKRPrv/0YU9XYSafMk8O1+jsxRQD0WLlVdbOSX
WDIVxdEdWOw3gpOkXLl6LPUiL1gqkohMgt9RaIwFzTRdDCi1jqm0G/Z/9qPZfdnm7hSF0ghT1LLR
6rqpJhL6CMz0cIPiDmF4jLtRedzfF4FCRs8n60kebPwcFJqb2TLWZk6p8uITt7Sh1xdEK7+lvJNg
nmFZgNTUWMdcBeCFBNi/jFy415vd/5i0/OCu8guY+t6SMfRn1cPXrUn/VYO5kZb+9l4Fj9Wg/sRn
cPGp9KSmqQDQzyawFNcO8+7ItZlsxhzg3BMPdNwdeGFTlb54vOWjlqwZuKSiVucG2p/tHtAalxTc
vfrVblI3P9ZBk9OC+iY2nWqbUWIlMFpIj8uTm1wJ4rDvkLO+gpX5Je7YGzcQsTF4MxdD3WkG9TGq
0kkLWrggXfFV3ogdTnvkhVuCjGGn9+tNNuCcKnil1jFKkVEkukL/+9vrFFZ0Yw13KQi7tZuUeyre
DU+OA7k8mNr6cZ4FTgkZsMS5q9LfCzHoVwIaHYZcjs8tQm6G9lS3FxOsczVwxZzwbEvXMmxjNgmP
NAicXQk915bOX/EzCROrzq/eIN5RZt/Ayfm0oQnbqnPXu2hgErEfyn9Xyj4kxSeteQ8SVv277OIj
plu/KRwoniSyKHriIEYYEcLmCKk3ZIfMnkRc1khJADQl6T38O8arSxxv/Yn5hbNTabbo5QWiHIHr
YYKzcNW+zcYJi+vz8PTr8UOO6xWaiz76lF1uq1Y09K08Z9z6ThywoY969SMLzSpo8oQ63OuaB3oj
05fQBuisRHbPa6kfqLI4j7E+cSRzcoXHPM6R5q5X67bWMoBB8q5NovH94LojJ+Wk2DAwTayMfxQ7
LB3Lq/JfvmwopN/sPhWxUkIT58IvTpXtjbUeHuGEh0rJXGdmo8S417mukin1rzIUlhbsn5Cw0IrM
L+IOvEfeDgevBRiu6PVgYE65cCTlb63brNpHLLh0tRh37IUMom2vP8j36M/mczhsWoC91DDCGU5A
ppATpGEOL+khUBVH19sKEuJzKjC1i/uslJbtLEwsDL5saEtROe1luEtCyO+LznSbuTzEq92bGxdT
PPPZXAglsnXO5Ir/8lIgaFi/8QBqNNUvO7X32B3sbAx3j68xIX4uUvou621R6JH5XbFS3SeOO/RP
iqrDW/jppWMgH2W7wKIOqSAiOuBrbeZyDhp+3akHfufTNVwUvTPvQCUrBECte6dXWKd1+MUlKFBR
z9w8ApFgwQeYbv9bGR0UFzW+VDHdZ6HB3D7+KieL/Oi/k5DjGyT+ex097ceKmD26d4RBPZEQ/sL1
tCObkd1p/7ZGY6uEgRVFeGz/i3x3zEfxQ7qZmex/LHHWgIvnnMsTLvTk6gfWrhpvIkDDoGHYU8ta
V1RpfrjZs/B8LOsuMqOrscCN4piLYY0PttpPqqC72SUMjTxzxLsOaaxnRUVcN6gDk0Q+gbyS1L+l
6tpPJwz4moIMbRbzfBU1zcYecpJ2tVZNfL6lXFHCkrYilO03k4txI4LxB5Fi0G/w7s9BUa+Seonf
sWorNFF0Zt4Qeiw8oEg6PFkqGtXctee0MI8peJcHeqXAXee+UcBy6OiVzMLFWJgCeSYM4JRSWSEa
I8uZ0YFtox9HFORVp8VsUQw3z7HqpOGOpDVygv/1C8GEMC2weIsM1OFnwLB1Ks35I8f9Tck95Vdx
NUBGzD4rG5xEQEp9q9goGk/IMeKvf1Okw0tFxm/plYzpDt8+k2jAAUu5rruyl6lJZtT8dqzk5gyw
/iI9KhdyeJkXignDJQyGAAN8i+mjPD3cYmTFJi/DIWneOa4Inj1x0EBkfj3xCLo7QolzW+i/UHky
NO2MlHVrH5cm3WY5Qx4k9AmurRgpFychn5P7VKWwrbhyCFUHtSEPErNfJKDU+jPid9zYwcb/y9xa
1XWnwYR/sWBvMEZ2Pf/tohtRZ8No8zv4rLlWIN0OsIHA0pwiiUtevjxoFSKqj85pyUOwV9YLhR/1
TQ7cuUfuDpdmlgCk2grw+Hjz6tr5ZbBg5M0hZCmVsyIvx5m0RPDHLLnUI6HeAe2dKpw3F8hPS+nl
MzoB6p6jS4W71kO29trD87vGGEiNAxogM4fYQVHbUTJc0g/Mgjy0ZXrA5UjeKJEo5psf2W1BoNBA
WAiUjL4lJxx819EQso4XBYBJ6uLoyIsVOn4ZNv88b3bSNVr5VlmF4diWUQqpLehlwHyzWfAzpPw+
pmmDQ53GSgymhTOrfXKDPpVNPUpn0jvZrCLzscsjfSAAhzjcHv5WIUAPiqBYXyWlJaI9MeW/JmrT
bwV9kyUWdFpEx/hnXGSSMmfk/4+qI864K91Ds1cot6LpMxA7qaVxFaqXhrWu9/OqtX+n4G0yAM6U
Az9lV0ozQZWe73pDHazGY8l/pkxYfRaY28wUMXFFphXpLL8RKv9X0USyzRi1sq7ysBApkH8gfdPL
gI/oa9ILoqu7usnGxHT/Bqhf+tSlBjxqBwa5oddsYiLqnnzUP+32/Dkm5cpnFawKLgwAOwE/+lL5
f7oVvSugHO60JA9dGQD2cTmKssU1Lr1MtaA019B7f6FPjNdbdwEh3XlGwk/T/7Jg01RWPTAPKCh8
k2rzNEZ04ttbWjdKGih9ekmYQpqtxUZYzGAIjusV9Lp26ZGQuE0ZRukgGyNPkEhl2UQ1pzPWZmDQ
VxV55CRG+pctHdg5CKb9G2zSqi7F/9BvlRkz5u/XJ5ouxNaVJYqw+y1kMWfkZjqUhuMh2zJms9zn
Qzvh3mRCqXyTWhTAsUDSIOMTXUVpnhQ9MlNPyx1oj/GNihzZcMhDgDfxS4uIwgFgFNJ5cgZfqk5J
47BreuqNgrjUaugDXZ7HhQX4na5CuDZK8/vFWE9lm9SunV/g848f5ykJCLSUDmIi5MZ8Q7v6laPs
B5vu4JAaH89oQGko1DRLd7Ij+jNwOtns3pXQqM+KqwpW2C//LlYKPTEe6wt47VFUu3fSUqZwC8bl
V0AkY402TgjTPx0K4kA2A8kPqDjiwPkhQ7UOxaiBK7LjEzgBMf0Iw1oOw3naXBbxGJ6QVal4fFlO
mFIdQq6usRV5/eqBi5+Y2eAPEbZJrJW7xgGIl3hVhEMtLgXUUVyTIgYjDkQ5W1w44y6GZa/aoJBR
RsZdnF/NHkEW83kAI2VHD8CKdLIeuZWPbGKqEkvK6BSbRJv8LhShEvrOLASlw2GWD1/B9mKADWY7
rSOXePRzLJkWsRni08Mm1KjGShFI+2BAyGhC2jcpalTcRMqvtvfr5lMNEGWwVYB6knfFXTCp97RL
iRHOsdnZDKpn+rs7kfaTL4quW8kRrP1/yQuKOnNMSuj2VIcKcksX6R9yrERMaFbQs4Wwx2gFJjFF
BiLgVh1aN3u6z2m/Y1SG2c9rVID0AQSpgtmfv9krIRgMSALSQrN/ctRCMhJoNAeXUfM74TNu+0qb
o+KxvZibm9TjRg6Ur9yO6dK8K/KfKbsTt3NwwvxsU5zHx7K5e8n42EHceopxijiGX+5i6J92lY+N
hrGMuuVHEG0/uAk6D13Axm2WN5Nc1J2qmaQeN4BoHYL7OfZn+jaIsKsqR2nYCmtJDiraS1jpIkkP
DAC4TzHhRMzo/cyotCYUB8I5fPzBjyf6DlxoNJqredb6GYNHL7/iAcsIp6EVChpqgBzmjpP/bmuh
Fk/cBbIVWxlHaxeINz1e+FMVt+blaaX5lsZZ4M1w+zTtmcUKzA++vrOX3Vmmn5sdH4c62NigT5k1
CBLi0XpP0lpThTS0wcbRG0eC2VEpUcaqX+UMikAAMuJ83kOWNUYAjKCmnVdZhFJpeUtGAtFBzS2y
is+0mG5Piw8xkQX/RAkEnzoCL9mD9C18F/oDSQZDn+glE/clcjeX5t1xA/x5MJwKmwHkVTA/e/2F
v4WDB9xFrCFOVONU1hLZU61fcOWTMXVTvQMcMUezT9dPM8Sii45sy9ddIDFDRwyzUojHeg2RFZj5
+cpHtUZjepSWRnngQGShPcfG0lvCIiiS7y9P/jKlA70Z600fwlyjVsjKGxL4+058/7TqPfpwwwDn
KN53plcVxBLZAcgjkY8IdQtrJryPuhUP2jD1mRAYR7dXijTgbFrpHoyKoJ+icYCEp0bIvpzl9rni
OA9mayy0G5aFsE1nwKQtDXi2XH8JvbtR9Kli5mKNeRq4xcGe/fTRS0gJ3tWPPrZQ93obwQIcIQ/J
Ta6Ajqc1plxEvTH6+/V9HQDrZAGleP5eAf2s0r7v7akfp4tbck5kR1fmxNr++eyXQyzwmGEvQbsS
K6a7atsbo+5oqUZuqGX9Tm+q0q8UIcc/Uc1zsDyV98BN1ro3yDpj1UCqh7m3+Tz1tRCK5Q2vHIVR
ckols3mT6vG9xB//hyPCa64nf7FfOF6hRXuIY5dIfUmFYR6yOG2wp7B+hIZLcUaSwTkvOry0K9xc
cAJF776AAYMVodkZ7gA0K9/mlDDAe+YN4HHt+9CfDZMndN3EWu5j5lFyCdLwrUhAS+pMduRX9CuA
rGe2vWQESq/jVO8cfDhALa1pKVLRMTyIoTGHZ3DiRX4MfkWN0EdxJUP+wcBLZMiWKlUCln2wpY+P
RgyswJU8cCC3g2Xl3R5UGzVWok27PqI5/ZOyMI7fE8bJre/QqfIregzgPvHU774KcArjYd+m8BZs
kMaSZrd+sEOhwF4gUvSJtv7M2HIv0BLYLFNeX1Iq3o6Ft/unHBgm+KNuXClagTv2fCnLHLwgzvx6
KbQnztXxX57Bafue8mDy3+mIxY1lDK8/S58rj6B1YkneKQFkjdbmKoGdBcJtFxpGrUeaX/ayxdcI
33lHNDqFIHqYwOrRJOvXd/7x95qOInAUps651p0C8fr5csd1Rbabgb9ngEP3h2R+hPMcuegWydni
MQAlHkNfuSjGYj8N7wRzPzTV6sbFyLdC75tIWwgMZkbOHoXO+Ioae7Z9h0yT1QbkLEN7+rWiSBOZ
+j+rpv4ANNKVHgZN6JARghTadpibb6qRo4VnON2xRTJFtVhtWfNSR/3fpYIqBJIeRi7d5MQdtpEa
mP5NtyGcrREU8P8gF19+/IFEcD2cF7lkhQbjLzQbd6288kANGioPEuuXU/KVmtPIIAbHGGSjMpoR
HAl158cyOB/vb5d+ckQ21mRnPSUEPBXrkS7k+KZ504Izab4/Enq8Ctw+CdZBG1azpX8N+lKAVace
0cxzOkGcwyYSSK1thfpvVPKYwKifDCzIy/jLFk6yyQl6xoUzXqbcVe6HYxwPc4/EEcY9jZbfgn1i
gJONy6STuPOAX1c5szQqYNCTg818HwOJYEwEw4m0LVlTShVGVRwHZxxtspNYh7MvF9KnxJUQm/+s
NIHfrTajXfL2b1ZKpA8Jk5RhbF6GsuDxnkVScKdDP1sZw5S9Ys9vqWIMCrQfVDAtcO8KyL1kjLSO
5YyuKhBNGO0a483tKXy3prEEH5Llhwpwzu4Wb5W6hscH/pgw4nJCk/2+1NIow2fSKAkKPr1zw8S3
zSpk1kdgO2cf6JdEqW9kMXaEhmAPxblcAs03oaYk0zHeWwe7a5yK9UDMXTxxORQrnrKSQKZPuFc7
uCwM99gdDLRotKDngqKvH0lf2PK+lJeo3eHVsqJ3IT8BslG1LgIoi/+NdswR84rICGCctF7hcODf
OfilqwohMC1pVjylpWV8pXgRuOWf2XKSV01PbeAjZAKtnnvs7GXyg4dqG1ThxSAIxpc0p8CA6KwI
W3xxXgs6oCQHDkFfk/gLbBcf+3EFsE79qreWRGQ9GxDhL0y6zdXnxFNujmYjUdTYutH1vO7/v3LX
cJuYkbZNNX3qHnAD1XS0zKX5eRlorPBInr85Y1gKOd4nqo2C6P8b1T3Ak1eTx0oxHB8Xw3s13vBY
usFGAdaa4NypNlEc5jgdNH/uZn6WGZUIeMeHyHoE/VkL4U69Xrw9yXkMSB8CY+0/IJgLmlyGoXKD
SGuQO5yMbXhdOy8vvENHIjJbwRvrjTfawIYiikx4X46QLVk9dJ4AcgNReSFOoH89zj4KTkPp3Bv/
78CPrOws2MVZq1oxE/jcfzONd1BrdfVnH+E9MJzxO467EGsXMJpC0ipXk1ckFt9t/DAAvrgvSb2d
4T4EmU82m1FmkNl0L6k9w/kTtEW+MUVIO15rqYW8UWUD+U3XJbAwC6TaHRloGbedq0dXaWdeTiCs
XPrPqpRiYAGbu7n9TfmhXuJP8EwDTqlZ1mow2jGjlTy/69rgfiqKEKa8WY+OcsNds5NGqfQLbXal
t6cOfn5XS7wIyeUtq20FOR9S7UrnfMtACdAHyXMWQF6XfNzDHG3M68AnJZF36gySc3Zd4XmAUvoI
eDgRKp2rvxpdTFklg2RKvtvSgT4RohojfluH9H+5bSaMTIt+bd6qQy1ewlLOD5YiNrGQ5IjcqXJP
8HyGVT6nu+lXyzS1neJV6J59iejafqgk6R37OybkE+FYAGwLQf6VvXDC3tipBCy9BXweguvKZz/G
3iJyHjjt08NGFn7Ns8Rg60nGWef5t+j1X5eSmYYaQ/Vl+aNzCK660DGvZAy9xQOsRrbxVQBAUfx1
H6NWU/t+B05gPdMHUalxrfshcO5IHPks57lt+ROlcMlURLxrPz8MtjfRuSfpzx4t+KR94ZaZkmxX
jpHhuUD8ITUBTflaSoSw7wT+GB8BpOHeWP7aQBZrvvLaVfG1OGqyiFn6CRdg/9Fd+KfDNToCRzXU
MtHT3fOJAX1vDEped9b94DfGkR/hSj4VLlxrEMrsdO3jtAc7r5YgRvblux91n2StVweBSFRw1/dg
YLykJE7GDBcJpIHatqjhV3E4Qq7g0IA9Xmj5OobxLdxdQirWmuwoghu8tlSuJZAVWDRW9+YD6NtH
d5UGcOC2raIUqRejQhx3qXt9jBa4JruGWa/sEVZd6zRmxnFC3k4pvwvY26Zr7aGT5f9bZf/ZvCuz
bLs6YwTjwfuJE4TfHHjCmM4dfXFoAPBvE6izsTOp+q83Z2dsQUPzLSlHKs9eJjYORWJCD9oxEzRY
qV0npzSt7ZmTCmpU/nXEknIRRVP3gec84tS8gF+2BkW/dXRdIvv96jSv0OSz8Sg83on4KGuZVkit
UCBKhzXp+Z/OLAx5ojBST6IBwwvBwC4BKWyNUvxMz7kFBRFci4X9hLm1XGJyZBZQmKs0ldCDggve
OCrVu+GoTug9tL00epA6ZDIe2Sk3MnNikWohyOZATvngEnIbbhuXRk+aQ/9os881Ymc0Ze1+p9xZ
UCphak1VRGRlRFBwavV/W67WUWFzhVJ+lu5iwf6vQMfa5xmHpbTSDiWrD0moSAccc248R6icvXuP
Oe1b5ymIGw6H1NMemHgFi2vicomn90YFTbUxS+Lsh0H6OvlbE8ItXiQmwRsx+Uwhj6ci07VDaIuI
NOTvonNgKjuuyLaVZuS0IBGB/VrnNWt8NWVBenbWt2WZafO3PjXY6WMoElmm1srJx5WgWQ8KAFqh
YldYQ4CYznuTmwtpDYEk+Yq5KlcMr+urN6ipv0/cqoUJxFcU2dW+TBGfITynX5qzImT4c5/qbyh3
g9x+UMuaUB0SFivXHkY05KdVHPqEGnH18HxRrJ1+sgiK7/sqEFjFHGRG8zUxctDF7AyemyATNSRh
9omTnIm0kyT5aBqtsckibKlGTDN1ofarNGTxoLdu38btP+0EvLGFWPDKtKHb+WcAETVPiETXbb5f
HQU0V+Vd4GdXgq+gLmfB/SgpdyAnX2WMX4Rs11kFij1HHa6kEy6W3QX+sozb7KL7aTH65WAWVuNF
F+eh5d3WAcC7zUkSUGxarVqXbIDMKNc+kAGJ+y0V183NRKTM/L6vYMi/1yIo2kATBkkayUeSr+3j
MYtmLHJLTDT46imISn9IkOMamaaBYVD+CJHfmUMKWVMavhyrV+j8HUfk3zcQiCJuNSbyecuDloIK
j+fEFc+1yU49qE0Z2AbNOsi+dng+057LiKDLapWHTNVmrZZJHLy669rxLiMO3omjkEb3dJj2mCKw
29YPW3m0Ak/p3D4qQhNtijUefE6YOkOUH64MWxmszuNHlAMyryQW0ljafyrW4PlpFu5EM+ty6QRt
10Ou+RQ0yA3V4XVxDQcI+mOtqnQIHUR91oLIlz2tseauRasMrGaM1uxi00EiOJRltltxjlDeKM1e
qm7lho1OpXT/KyqWgz4wcOQ+4v35fNT8/PEdKxS8DQAvxZUz+kWDpjb/wE5fpbGrsUtawiq0Jw9J
MtJW74IT3yVTOerg3BRT5v468uGFx5pi4Zs7KDNnVLFuWdy0TC3q+pX/n/ceDqtxw9ULDnfrwyxq
rkvBouKVAeTNp7HLbSvOr87yCD+78vgdNGORdWVbOzLq0KBdkXOyb2cWX+Bh1WeUtjB3SlamgSwo
Yc4PCoRpWVWVAg3pGs/ZEqm3G6p+5lGFS+PM2kACs3Q2ssevxxg56t/SdYsooSQc0/sUeoW0yXnk
UzLFzF+J/BROVilDFr9y8+wuCa9AgGCfwHX5CAy/mKn/jKY2/fgefRsYDJyLz2dtkL9HHMCl/xrE
cIbW7Kjz08VQg4A2OF1kWdDBq82XKxnmKvuU4A+NaPPdLmyk/OgviqawAA5yeAUQqgpXghYqWoS0
P9TUEythFKgWanK1ihqd+HOzZZEuwPI14WRdI7mnVqrajaGOPhJ/biffC7Z2e/sqSCQTx9PMayYy
wwR4ebeDfc5EjZseUdzBxXuKaKUcmq3Qd7GlcgXzH5PbmlSEzev5ht2hkadGd/b44VexhxwpuYXc
2vcL9rA0wETN1XU9lFPBlnHsz/cu04wORovYlvAAO7h5NvBg9LGZl5p8XHjLEje9gYuMLwjittMh
/neT/wnMGpDIIYQAvoSqR8YCHK1brMGh5v6KyMSUjvCdXLViGbsrccKbWQTRZSy6dsxCPatVFrlK
ZonfBt5szGVxxNCSh6HptO3oQ428ovb/5gYhNDNIe5UTXUp9vH3Dvfm36rGKDlzhaAtPZrRQIrlz
Qn66YLmA4dS7dHzbioK73XsfHzrnSbkXXfr8xvdVlbLxCn9n6TPrU53SGY09NyD39bMNzXuz54yR
lduc0UsQuPo1UyyIPyrj277JBpaU42HHf8FSmd+2p0pjmkT5Me/LafGKw9axTzx+Q9KsR5smLWOU
lCGyR8pUs8xvue9kQ+nzfjVB3tNtBVg8DZw5qar4IIBSlAPynX5KI/5QaBBSiLNS7Mlge/ys0Yvo
r9/XAa9LA4eIFjygwC7SEEbCH9vm/Ct025XaL18VfCJVRcmF4K+3agKAix8a6ZZnhfGErKa98/Ch
9sAd6Yt8pncbYM9NeHcD1DmyeGw+DQYB5vCPhqlZCnoSSWxJfGdraRLLyB1vhtWmPcFosCl/bzmP
RL4V8b2UGoOJpd4tFmgzlkbP64XRjOryIQPA+bVqlnBPY2xAchTl8jCE98hDBPL/jG57UxomurtA
Uaeb+1dxZ4PfXpi0fIicKiuEjUk+amNDH1u3361BtCYwPhjt5rn0l/vgjxG7X+Rq5GiRKjX0uFUC
1JW+IDYI0sxcEP5A5w6yZpnhndgBXptU3X2WLCdRlXVBRmBif0FgzODbABPS0qaquE0M/rM/iXLz
Dk4ukRLrqsx0LI+ZIpHACer+7H3mNwuFu1dMIkHrHdtqB2xh0c/3yPVIOUvgRIrWKtXcFkhkGt6G
zUFkffPwOOqs9iICdtBhn5yL4GR8jJyewUx+ftvg0c/K0C3b/jasFVmbGfHLzTn2veWkk9xLifg3
2wUyu4fVEBlZlcM7GUEmTnMMTXEp409fyB4aMvX6jqf2RKy4vGGWOq17SUI82h/n3zAyZ+k/uxkV
fG/tk56AW2aMHT6VOD0w3lr1NcKtLv+e48ExaqukF7zAuJO6VR6xwu/j11ZE+g/yAVKo5Znl1aZv
Wsmd6sBi5hcJXprEgssw3p9jFYrv6wsXGdZldzWcScLOLuMl+Y42l9CNUX2rIdiY5ks4//uRZscA
ya0HzIS40qyZdE9eLvJskZI+pIAM8YxgnvGIVZ9QprD1N3eVbQ+oiA1QqaxP/gbyK5jP1krvw4bp
eMMpQZUyiAm9aWrUy0H2Zmpe46r69p7KY1XVxC7F3U/36lsoDKEZpcRUtTFtI8fT5vl2S/V7ymL0
EmTDkztj0uWVuz5KqUR0cVMjiwqlYDYUnexepGB6qnBA2J9KHfNVnuP+rz/o/AXXiWJQn7eH+WSy
sz5pp80IO27a+26OIv85DR/LgoquyvC6HAJEEkxyb/2eoq/97Su8iDWwS9nWTteW0c/HgqaXGynb
Odx0RigEtkEnWD1SX7OiWThUQ4qFgD/XUBl5PpkABtDYL7Uh0Mn79VS7kp3lt2nlIKGHBOZ9X5oz
fct/K+8ReoxjwnDMfWY+Gc6zgr6cE06d6A5za/MysDwn4JNMK1CxqC1RGdNBVSHADE6qCA3Esyui
5oecgGtJvyWLgQSH2+Ke0H7YObA3/pFoaFOQFdcfm+1jduVgqcjAf/0PEUefX0Sx28knt4+e0m3c
1Ewk63wrBBYQfPHVBiM4xqZBUMVB/LuJPLcgTtNRD0haKiNaIxZlH6SKuIHrKrVhGtDm5cu9vZmh
K2hDY82SyUnLwWcgPL8i2AI6M9Ok3m7fqp782Ydq8Dwh5my/09iiGPU57e8hSSY9pGPouJtdM6uK
uO6uceirWaN0Bp0y4swU7hesVbQJgTSSgoUfdHdDXopasA4s7/a++k3G3LeMHmwglPG3W5Fw666r
RIasM4F/zSn1Ss55n391lIn5a+iFsBp2PEae3+/qJTPc/HuOv4LDqMRBPYHUUBJoObxRCaVKMxYC
vvsgosGu3t6bhvYJRWWIqxQW1KBnzLIc4f8YLkShOXzzzZvv1WeZJv6rBK5IV6BaHSLQ/bXQ8ZjQ
mix2vw3A+zzB8Zl9cn586seNGCr9S+1OH+Pbw/0MODhaQG21KRaMKRnLejJWsqdEeh0sJ9C2QdWW
w0pk0bBUHFMQZnrhSa2oUhMRZZjPTx/WWV9ixoyD+QArL8GpvcnvX+qlZGEH2AdSPY/nSU99ave+
TXhV2Zx3T8syk4YDbm0f8wldzaY7Drj325sumbPyJ3/9Cy7z2J3NNtucc1FgggWWuR0GUSi4+3wV
CQf3kFR98dN4vBPxwuLE7N+HLWEWKSpfTFr2udVOKjBFzEeUHx76b9MxnOF42LbTDaKPi+Xwe9em
Hn+gxHKdjH6dTiRlY8+o2GMDwU0eUv5j1P/hj138DnmBs1aP85XgmgNsSD1ryZ8WF5j9b5HfVYS2
FR2NdKuOkwnE+1x8W5dPLFvta3JhFglxjKA0aLQUAf1jmRHTaDxMDk+wuWhmg3tkVM2rD03ZOpka
6BHBPNhObkkkcOFrtDlqQ6cYPh+HQOLTUtcL6UyXc6+mEaRVtRS0yLaKyVGEE/WKE+G2ojngC61/
cBHTEktxG8eUz3/kzy46kbzFbw8R1eQUc1vMmNbQ9uRJY0m0kJAgnTvGuqrjrgaHWERu3407TiOt
1xAWcPcYyalusy/sl1s3G9zDzduoYoYU6LmdBPMXc2OrC5351dUHC51uXD1dc93PJ5+EIRfVPmZ1
1wS7F1slIvCXCBPB5/gQVy7FRBMUAIofQxtyp89UTPjHaxV3txiuNWs2a5OrUoLhfxPKrCVH8wW4
QB3jUo/poLl0azIJSgnOGSIyFi3gjaASoZIZK2iINCcV+D6RrrP5wKp8vWxGdLywIj4HsZX+3leF
t5/9bsDEGHa6SXolL4icqx833ZHjKMOVdZmc8pb0zXk57knM3V3eX01lFvFIoBdgYv4dvYmHH/U5
ZmVJinu0vjHUORmCn9zKHqkRaaVaD7N6h0zyJUluZ55TtuiPV8g+oEAx8ZYPBOmDibsry8RR/Y+2
YVmtRMP3FGbEo9S+TiqJecrmW7nbJvl4gfwlTw06waTNdGcuqOuXoseOfWOWaq+mPpjCX2hDYaSy
aHokEn/CvP5hEVe4DJtVHQhvR7k4K0ZOeuMkWbBjAfkIRnuhg31TZoI3qBHDvGsMDTAAGnve1dWW
1Nn1S/JNGkmCe301v3vMljishlbYRZVY1QvVUh0FIyJBwwa9DOe7VSbHOb+rjgRhFoWJ/RBz5GTX
RXRS4NeyelgweEFN3qwPYlC/Rs6+SKN/XwUOhUtrhVAUyxss+i5UkJ0LiQbqFaS1ZdM9ZnnG6glr
BBSqM3/Q1q0fKNU9nfU0VGQrs48JoO5jyklhatsnh4Mh75lUvPMWc4wxVwH8A5O0jX2+HINVxqGW
CFKfMHSeVPhl7rWdTto9g6O86ssUZOyDnnZxF//9XOv5FonWgK6lOhzxDO6TV3U3avg6ZLl9wGUJ
ZK+X1zPGeU436ROx44yNp++Ck+D56+Pc1abssuBTdDmYSri5ptu2P6nTmpJS50Zd1VU2TFJi3cpG
SsbgHh0zniXLO7xuVdMLND5KhYd2sgeqoRxat1+xRSQfNdIqoIis3KcMl4cb7WxgAx0LTf+Aefgr
31N3N2ElIU0PaND1qmlW6Guk7+Mf1GtlzoJTyD7X19wMzZPHO2iyWpu4Icmcjf4DqLPuTnoOJp7R
U/C88ZPPU/kjjyQSTeba8QDQ4nWQN7aO1IOEgejUOzdkcw1djtzx5DIqZUsILjlrMOgbpI5HZSyv
om24z9Et9lJ7eJ8B/lNAhOPfwgdHyo3xTevb2sy3fo+IH94fzuH3UBDrKJMjjhWPj75F/r07WXEn
2QZXttNm0VxXnsg2Ro9oiAhwPSr9ApfLVMILpM+p4nEEA23aZNCJN2y42wXrTJlgDR28muC527zS
oo0h4ObVkZwrpm8yOc2Ozu93dveAGNKTC3E0L0+OtvKhM3Z8gOEEERGSeBL57T523d0iU99p6LN2
RuWdMncKsB8x7pD5SbeH2KVBrotYkVzZ5QfHsq1qHJ2kzNx4+lgX/0nWOvzBcHb5cL28aeCcDAXM
zwjMhygotyB2rXf3EVnyswrUNcu7sbiCUR7LHrM8FdUG18QVlcvjmfcRyrAqypYGU0nyK4DR/O5Q
3KKoL4XwQ5Bsm9/BA7GsrFiUqOx3Tq7u0RlFvxJGPG+uusJMljrWmMyOnsnl7n1IelG67v8OzCKk
jyi7vQDx3a0RYY0LLy3COfeNB8Nzk403C4euTY4SM6iSOvXVd2MZljoMfkU5tmQov53xz16C3sxN
idK9o1z8bjFYusDNMN9i+1SWbl1Il9I2EG8WMXp+5KdDTO4TIPoXY0nwsLFH/bIvzMTWWzy7IoRw
yl1fxKy7tqMENrcE+rVvqbMveFfEQc6ErRgmGWNRpkQ4dBL6vR/I2ShL6FXx7Pd7vYOLi6x5oYki
3Q+sOBViuIRW84vOP8fMVHilQ82svYT1pTXFLBI5l4uoUUOIj7fm0O7bwnWGFOmACrrWNZm9Zd09
/IJ72BPYCfX3UzSBGaycv8oCo+8LmZf2e/f6RmwPfUaWw7cj9IxKNoOS9j7ajyzhk7Cst+TrGnhE
trAFiNYgV4+xlfjqSsB++2wWKii/9mEuyHwsP/vAGI4p5NJ6WEKNWTUF5N+Z0mdF24mqwuUu+A/+
xilNGwlBc7KSEaZeXEXioQU58u6Ew5mTcEvT6d25DI/msUunYIXiHDeIcCnGLLuVo4dkpyn4EW++
evq+TmXrJQLCqz3k7xUcvq3meZkCXQAdzT3qIHA3Tg29XurT5tDlQjWFbqs+lmceF/R9kNUIQWGG
g7GTZrmYkC5EviPknArvO8vTXVRn4FzCuq9sEjQJRDmjfNgqH7UTzsr/kWW3+Vvkcc9yzH91in+h
RAdUDa140oxzrRT4honWqElcYVNwAXGyZ+26TO1Ahmnjo1cSaHUCDu+vWEGrDIMaHQ+BajkFmfzd
dFBxwdgkmwy4pAqM53t3TaAj3o91gC+u3tNV8Irez7X15d7NfQWZDTUTZw1V8TzWX/RepU8Pd1ad
1XEpAoAwOwADqpgosm/QPNORPoc0WLhcvujeae3r/C1hzY2uXrX+gSBdspFALwy10eirqdwzFGKl
/kslVyHEl+T0Go8bCWRp5CVw1HnGiAi47yybxaTTqLJtlN1t2OTAIXMHd1rIDIZ9t2Jt/zIIwhLK
vj1p0tsiwd9Aov/fdLKDdwFBrQUrEvx5R6aqSsFrEGZFYtcqXiw0lgnBd8ct5VFa+Lwpwk3NW1y0
uHcjvCMCZtsP+a/fDD9OHbUG2MbpsJkZwlX+zcC6JzGasoVuRrHQTSoictuLpoYzfJkS/ywPoqNQ
qBXrcm4Od+gWlASrGgbBZHfi/EvVB1Z0SrVPwPYdkNPyi1rVurHoBT9hzDRgu8rB3r6oWfi7qVpC
UvwqM9Yv3Gb/bgwNFe4j7VcTTPbmIQ+PyE7hxcwW6kvkGX/lmvkH49DrrApEcmULpyJZm6rY6LDn
AuqBUEgmU8og6qWhvOyB9ZxrIa/0tXd+yFbAgjRPYAjiCRDBoUn48eelGKdDfT1u5VVOO7qbUznP
/Wqc0fqiKaDi0wFll+3LDM3sUHqQHd/ASU+5/LZzgOVcG3HWvawzPGUbRJbFWUnoRJkHN1PcwcUr
Oeu48vYMeD+EMEeI5w9ILBLYx1KsFE78CJ+2nFE3wdEeFsxHYWNc5xRyjaZaOAeoVxdxlqEcsSYU
FIthzrfNr4d9QzyFepzFNEmUOx0fydNRH4gu6BAcNaizNxhwEndcXegzixwuHROSqiB1Ek1oW4HU
+d4CH0MtBe1zZBOOWxvJS/Nhs5Fo92G0F9KhPK5kXtXMzLAA5WjhPJiUwHiYvz9Szrc9+coJvQYQ
biy2MkZg/5Tz5AnF1Yh76L4yud3FTB1sJN5wFv5b3FE2bA70io00kwokRl1/mxV/yjg++A2ZWt1M
bGXHQiWi7SPzuUx0LURnyA440FoJ8a6ofcyM5HlCmQ3Ua+vgbgTSZVWwjWQawE9TzQ3YCNhG/sjx
4+aenr5W9UquHkQmAKyThTh5FP8Ic8Oi8CHYjI+89/zALsCotLqQE8eM91oqpgBi6b4RaJzQvq7V
/X6pwDZQjuu44bo7NzS5ii1si0YdukwzBeSGSt8XSONIITFQc1JIi9gPo2b6C6zufdeAcuwAmvCY
OOLsbduh2SuyiuLqSdsQLO8O6n2/TU6erS4h4fCBlHS9ORwaY6UeIAK8lj76oeo1zI1S+/miaY3Y
+aA9hfC/tA1Lv9gLNibPNk+2lAvLOj2g6CqvSD2WMyXS/XJFpPJRWTr1QNdZcSx6j3ry/63egrZA
xHoSHC2WBWaraBFg48iW+Yd82+/jugLeyxTPztd4HcuNGxytICl1XkOiIg8CTOkSvlAqt4ZXPpBN
vW7xYhKFosKQ1qV4c0vyEdWC/IyodMgLHPEj7UdMd5Re6YFemvyB0bplggCUcSZ1okK7F2HfeOER
c/NGCVWmGZ0gWlXPRBnrK0n8Fn4hU/LgOOTl0rPddw75pz6ZWy3/9G3Q2wQR7zl9nzbrN1+UKM/l
POjVNaw5cXxsgfXTa3r6tg2aLuPnXxOYNTniSGq0X19S2GXMB8QVzN89qJq2Z4x+HWwi7QgX7X7r
aZFLjnRCJ4Kf7eir2ulzbOLNeIi2O+rZ5184VL8hl1CV853zBwbu241EGOt3KSd30M+EjP/dqoSh
KUDq14Hyt3KAWvu1VB601yvvYUkXEJY5KiTYOoUfMCmogaJfwsl4CF2iEts/veeJd5aGok0qYnIh
LBSECPLIdv0c9Qyph6ssRx+2QZeYJ3rNE4BZNrt/lwmoQmtThw0/N/+dMepJKAPW6/foNRvouWq8
HeuzWx6lwwqCBwyE+lzffyM2RU0pFEli5TLvCMLcli/x0s5+NX6SueDoBdX+0uwCDChvztVxLoAo
HZJ9sYvL/39CscIB8vOVZZCzzV+efrhocf6LsXshv6o6D2cQ6joL0RxUWgFjUepT4cQRWPWMwo15
7wflSQ5Dd0c4CDEyfrQZGeX325rz0EZMSOmWrVIyQ64KlAbHFsuKo6HbK+7WmdWX3SKyOS0pXq8c
WekB3KBHO4AYiCliL+vmaMosm22dhCbaVaqNaA1Me41o6QjK/Xuu/3UmM/+og8vuDeSnb6OmiylU
pIcK09tYsrIBgDn3wGQdjaW877Hj0vvgdVqcQrjGWFxMEylVwn1SIl83IRINsnW9DO0Tf5xe5GST
n32mpzRtwgBOtoHeXImKeG6iYDZkvrC1pDfOy/RXNru8QGl78q2Er/oCjfrpzQDwAqt2n42WknYC
EZLHgppZa71Z2I8xmd3lbec5vOdDASc4uT8uyJWuUiKmJD/lB55TegDXWLVW4B4pXKzD8OYRnvYD
Z16pvNQ1aeWinTxAUDvLI8cAqRS9GYlECoS2nKI8DIjbFvs563zSWdhjL5sCY5bhOhR8H5kOfoPd
zlmrUrBiDPxh/Mm2WV5pARFjLkHjTCSI474UpM1dHgM3EPEYr7zdxglGcwxc/FgzPW0Pm9EcC6GO
XD5SQlVkuC1OJvIYRZWxm+sEpLpCH51BHg0K+AziizzhmcM/qn5KpXxDqR3aSluCJAavpCp8I9BE
NwM/AvxgWdfHgtLbul9rLA0rfuBFaqs3VsWtL4xe9PeO236+hvH2W92ONgr3940utT+M2r5DXw+s
RORDLfwwrpIC43mZWDT4M2UQli0KiEBY9z1rejSb0S3/SyWZI1AEiAFg/ZMfC9XdQx3othcncrBE
6OXmHDLQvYOP35T1jCx4Hr/4ZednJ81B4UkszcHd+DkF6sLisp53bTDEMceRtxyVUHX9BDHqI2SW
q2fy3WXUxvIx3z0YU2UlKBIPz+1Wu4XjePgT80agzpSNalkN+07GLYhBg/lACBX5V0S5M9/wCicn
biu1n6nNv78tkGJfrHNNeSlYowa+bT7RdDjKEU+FgjBNnXFozXxQ3dQP5eARp1oxGB/OmjSgWuJK
7yp3pf6tStsIHtXgF00uubACdi6ZiNh1leJIfE7ll36u0b/4G3x4JkQlsxK8qXJNI9D++sudM80J
qjQLx7m/BrV2AumMOSynsEb2vil1RTRSvjn+/dLcp73vH3hke2Cr3w7dGvJE4z46HSib96sETDeH
spAUhz2MlVgO3afDSJgJe9kEekmMmsgnWEW0dz54VykPB1W6KGqZy4bF9mXbsPk/BdAW7v0mZPHj
PBnO+5G5VNmwlkV9VfEPRt9bHkgv8eOihOwAtpHRtVH1WJbxRpNytH3/KMLoqZac0g29ryQpcRLe
27kUAhxEDrAUdMyQzBW+RxKdHCq+lIDOMft6vOaKWZVyvm8D6lfYnYB3M2RhH5qeUrbNEAV0fvTS
qRizBcn1PNgniBd/BMhO0bbQxqPBdbisrYM72g3zyDKCySlKbGoH2lKP70ebIhNhyVDh8/81za+4
aZuU1M21xdOXWmQqDqUWY015hxFHnfgzFKkxpjp+sAlTtyUeluBWM8Utpody7wPm+i7VRPkWCXE5
yfy8ooNDT3V9kEKco7R7CHc6Jl0kt/xU3+L4fYZYhTWWOV+GHGEsXT0wOSuVIixzB65+0cksEjtI
RUnFX8RfhxK/CLsOU9nNJ/8Kjj2cSe8f+EH3F5s4AsmteKbIGPOd0h0YlKqjtO5rTf0AK4F362Qr
nEL8OnJzwnEaXQbTCQrLuDOX/3T8qPmeWbVFq9B0bT34w+GT2ZinHYNNoUsY1hwJfTELkOEjDe9q
eo+mCSahNp9bQCkcsqXpP1mrnpJbYkYMYz9mU1+6N8V0kf79yIM5IJDmTiSTDJRdWv9RKtoQcICn
kDTzIIITA/XXALtMyPfWoyjTSA+c4833c8aHcc9Uca6ZEdWdcslwVDW+4rM9F4RlMXaJrZxhHmcv
c531vt6V+2LchfwR4gSp+hMbu0iva5L1V0tAvMs/4gH6vi5pSP77t19MPKxgx1FdYpSvO1hGTQ/3
oid6svlQdSVUlNBX3Hptz0YbuFnzuEJffobjPogJdq6ebkNMFjxv7QEnCQtBkDkTyBrq/TYWOcmM
AxCieis3c25khtVRd2Bk6gGfz+TG61aZbp7kLPbi7Qv4gS0wq9vh/HlemwoU8djmXLfQGD4HXn2U
0IpNVy35asQrIWrLtghaAcoK2UE44v7qrZCYd2SXllsgZEfuKFHxbAqI0z8fCZ0TwZDEmOeIG1lQ
n4fMRxWyK4U7aLEiODBr6/XWyGVgqGKX2adaPV/pHiDH5MnRtM332Oef4GI/x5ffs08waRX0nGqx
GDedP23caawiPuJ8AteNt+xdQZJ1gd7IDMFm2g/KKqpkx1CcZxI9cevdYyf1eqw4mBKoWaqvkDR7
yS+hdop90AKIKch143caq4+FNs5XlfPzrvWUfZaOesAxDiKg9wpD2fc1+K+drt6yMRC7RPs/dnAk
7Wa5a3w2S7wk2a6cW6+ylJRgeeowGYIaMgjqGmyiXfzR0FVjpsQWp1AKsLZXbVu+dIouwhyeRLlQ
kDo6LO3AmRV7iz8fUVTA2BFrub4VN0TVfx5r004HQUVeG6B8R1UUNDyPLnZtsird4wCWcPDAdCl4
d6bG30SHhXFZV5sj6c9os5seqV0F+UBc8PSZ0XMo603JjWCdCMskJbiHe41ED4dU2+t14PL1Xoic
CzcLbEyc5Sa5aY1eS8Cd9i72vnTg5N6VcNIpCQ52iCecvmORFFK/bXzPKRM5xW1jzFEhDsx6EjaJ
2nTbY4WIg0AHFZzbYIjnYTGK/8zBMADciRfCmFHwc3jbZuWARNv6B65Hi3MjoLHkvPVa+JAIQ/rm
4pbMBJN6IXZ18/5jaYHnwJWJp197gYlr12NqO56+EllbvWsWs7hVqUpLoc5u55l8uDDMjq1L/iKi
4KwHddAUbeFdn7LtcEkTy+lTP5Gn6dOTuUA8djnkcihqKIukmD1DAH4AKbqP3RIM+RqfF5bGjDy6
4vc9jYNksTlkbUXyRYUThvKU314x8JEsANSXDIAXkiSNaU12aO/Di8tz6NSlEfyhD0hv8L7oQYHb
o3OQC4kOQ5V+ETgW8SPJJ1G+jmrNNanEZrNzGhj8okpjvUSL3Y1iCnbjcPCIdAsZfYNocNmB7kdF
nSttORxrNhRZnEYQmKs//fy86ES2VKP2b4pBN/gFUthm/5ZLwaalB9vgtcNdf6FSsorf/gUHIyL7
V5j/jzPhYqsJiB1HVOfz5RfMqVuyiW/BeKPa09CGrIKPnGbQvwdYRePdEm+7bXPmV8iIk58wW02/
2ZSSHDO+OzwsrCQMJF5gOeEehGcVQYBEwLwKne8AbFf/GAq95Rk9/aEXtuVCIkJPIC1xPlSndA1s
WQUMhNZITX3RMnYLP5ghWg9xHWy99DJo1aI/FwEUfhCNo7CGd0mlXcJHCw2y0U1xnZ540pQiOe70
5/kWftWqj+k13A7ABcZkwPK0RKBtDfThzpYQRbRpr9eAivjWQ5J89h+RC/O1kHm1gKbMXZm3ohD8
KMD8Os7lIKdWtg8m18xWVLYVZ7d3ndWWi2uXjSlOcACNx2jeU5IxDkzYU/lW3LwcrSuQ4qKIIrbO
vvp653WVjX2bZV/XmU6AxKmMfV0FATdYl7NuIBvnT64B2Z6BoNG6NvWXJZ+hQKJjKLvJXFOeMG9p
4znBgZ0DzLSbFcDI1dVb8nnL/6DLxOMegiUEGmvtTb3bgjVxU6tcdav2WWket2jLV9zt6TwaX9sZ
sTxv9g9c+x7QqJ0eGmQynyDF10xeWdoPjA9LYD5lt8yAREHAVSzA214lMHsKUEcIVcu7/4LysBpW
t6JO3J6/VklxPIAugSpaza64du9ayUEZJw1G9pWeeD+Eqz9zbQJwBm03AFOvaJz0NDhd2DbYfxiQ
46SjGHv1Mb76fQR8e+5PVfoD7mJxXAbbozMnSTNx6E9dYt+XOCEzeFLk1wuDRESRIfLWyVINP6RG
mpcOgJHG84hnHszS8r+jm9qLoqTA34O088pfajwIFE1+j/MFBQT7FUUJhesUF+5I1b8f0eQSJFrz
4GtWjhT6bdniJVmNJGto3TweUMYMVw2TsRQ3lNr0H3h6ht3ly0RGD1koZmND7+Ilw/LcEmYCv0+v
V13VQdqaoJpFvQnYoRqut55o5z55Z51xg50YKCdi+ezOLkz6+x464iIHPv91EESMH6+2rrpskwOb
72b4zkl3CpqED0bBjTWROZLnwh3KSafoOrNLr0c1Rl1aQigIhI+ll4nWfEU28q5ibOdtyGb10QA6
jb7A9ROmnmeKO6lbyW9gVTw9QVKqfdeUWV59cOXq8536JdEu7VbsG/aXbfdg/Gs1t4DzJHZdlWgM
z8Bjm6dyEH+e736feGBvhrC6knJXSAzK9b6AU8v71QDttX92a2gehl1v6Kjp8B8hYNk8w8NDS7RX
Hsa0lRRFXoWz69m9OKThbgDu1zGsua5hF3ry25GEWTYdfJK0bNZSIkr6gIBZAPrenbJR+jT2/eIy
hKTZgRe88aa29LxtSPGnlBDqMB4nzBM2td0Q5yvgk7hL2b0G8G54LAfek3ReNsdCz5Xnx7r+bKif
Jp8FcL5l5nfFCk5V0bysu6drukh8Xjy+vBdrjDPiJ4jBBkfmSAWbD3z4HBvjIm//S7TaJob99gZF
l8C+sCaXrM/9ICqOlpIS2wlAZDDeJG+vOhFbPrPfNh4bNGRZseC9prj8o3YX0RtrpCa36kIljWJM
D6VTNQHyDtO5gWr79bSdmUZ3ax5IMqyVdRCfescsQ99k+qSpkLhSz6TsGq0dP1yHIre/4Qsmx+6E
cb1CCkmuf7ydPhuvomdF86bg353umYZomvxJtsaU4iNIVKkzW4PvebLVW/NIR1Ycu6eO0noH99Lq
+eW/hqX8hKY4wnZ0Ay0XivhoONPL9CZnrxEy5+uPHkCKgbakDGJgoE4Q4BfLJPFgaWIlJhOxT1od
Eo8EM1HLM0beViFKgDZMQ8r2LLJiy2MUGuB1XDZQaztqiSBLG2TG2z3iJI4fZq4gSrvXlskua68w
5KmLj0RSzlxG3X6QxzhKQdsMtB1IdHN1oLvl7oOhnXhSwmE4YlBOm8nFSZWeP03yH6JUGt9bgU6w
EkbA7HFQ7fYnpJI4vZcDwCggU0fhU5w3UaDDbR2nKb7DlaKCHNAhe0q48nTH/UeTc3FoPg9LbwWK
lLmjTvbmgDUTUnh0sIrE9S9SVjgD8XJ2yjJ9JQ0KkBPohnVjHjGRNVlh9fCFtUvEVp9N5/axCN/s
+uuSRoRICDVySLF+6/NRx4hImYZQcmwnACwmUt8OkHoRNEJbk35PpcMi9A5xJV7Ap+T+k3q1GQVa
mcY3ESXnO/ll4M4P/9851C284TXeUVLWEVw9ssCYP0+YU5uGj8bIjHXjRsxtELfX92GYVUoBa1ab
MqczuAFz9Wuru0CQtNAomsbpCqs7O79rtquvqyh6PVS3kWjjTwp4/KSSsaAtRTZ1rFTQ7s62gSiL
JJ4zkmKiQn+n1ai3v2GlAMy8F/MHiACoEnwsmcmTG+xLedD07Woy6N4/2dvmdjRHLGlury4rJAkj
/oj7q/o3nk0TZF9um/7YcmVdm+tLCvT0a4um2TEuxJmY3AOR5rxv/AKeC+nzALUeJ9QjkNvSA3h4
dqGjfxfImoyvj7fS00vc8f9K9esIYdlXmb+9dpSpn2DxtsxzDO0o0xG6dIshaBef2GPqRiwoU8bP
GERD3CAFUn8dDxz7zzb6c5THyLUDxVSd5x9ZoNzAjltlyLi3yOnmcvaU/G+MdgE5h6gp6xsteNo7
KxUW4IqtKmeiUwRibhl6gytai3aHeEWwWCMcUxTIocazgi79HHPMkc920FJmw/3YwqioFRXYzRwo
JBXNfFZek0rv9m55BwRxByHPVF+fj3jXDj2sTaL37b5bcyTLdXNQK1HVt5fMbfez+5CvHxGRw3Il
8KK6mNYNwPy/Cm6vizwZgF4jM6hojIBgN9QAYNBSLb7rUGK6qoIgWd+/rHv4HAgjJAkaTi0ct3Sp
JYtQ8xLvkMV8vKQHOlFKnVrsEdxL4xP8xo7cyTPX3YEGTUDlPthegddPOTxXcP0upzS4abka3WAr
l6KWcFY1YsdFxA5YpQusJzZ8VO6vKSN7x49/o/FxS8Y8b5wiIUWfRY/MtuqcbFqI4lnaFEJPSj2X
y01B5LF+6JZJPRZdBoB0183OC+8NEaJz9eF7RKandfsq2nuRvqVe3OadMbDUl3QuONBQTAzfls40
V1CJr8h90PFZ6ZaGoG/s09xd9M6m43it8MQQu0deKriAU/Lk0CavUOCih8EiPMVclsPu90C6Rdmp
+86LEVuXNExXj03O5BRNPW/108m54g1Rrm74fPFA+C060oQWPQ/wjIjvUv3bM6BwCru/NGdSFAB7
wKWBgAfyjjMfpw6Os6XEytvyBJTXIRPpeNPZp7BJE5qc/ubG3vwOwNKHh8nDc13fX4BqbRxYsmB9
+Yzvjymyxhubx1g3VE/9+PKLQ8bZaFxc51Nyta/YkGpv8c4Ur1YMYynjuuT3Q5VqyJWYO3pxn86n
r5M0exhEahVocnNm/OXlF8walt11ilW+tOkxQU4rt3eT9NlSgbefO+t8C+o2vFwfrf2I1Pr7iu+e
llMvd07rFAFEAq94t6SIA6bMr3n5rl4kqjR1s1N8hXxrF2I9h/XpRACCgLqy/mxHWiyMvNz7AucO
RzrWm0VuH+LM5gaNYSKNWv+d+t3TwIF9NeiCqKUrZdZBCyWoWmbDtdHgkPJc7CHjk9yAcrEZw41e
ctvn9qXjCKtaaEF94AQERIvPNJMO2ogMEIyDsF0Ho3zUdTuy0lhu29MZH38NHLU5dCjf1xXM+7Ca
3vm5iS2fbn+0H2vxEBo9BURfGbTv+f0Jjhqsnye910mIsyHq8H2qgCXbd83UutbVsRR6+SzkgaYB
McGbI2OxwKxVbS0j7prPanaj3yhGxaHe6ujogSg6gNOwoOWRl43E6enK64hUiV608MvF1m96Qnn/
0ywgQrUo/5yiV4iWjn0P8tecnwWeBfEL1GbGdVLsS2O/OTqvIkTfkIo/dSF4tlxTHIRTctuCKfHz
ZZuMJF6nvU0V9xVNb7VFQQr9iQSca2j58H4mzbO47O9qiRyZRfyipqKkkwRdF1f2/pcaTaP62HrZ
+8w0fnSYznzO/OJCnqztcFPqUKKvLaRG54wCReq+o4rBbTlYTmXXN9oWpgTr/Hqt/cwSodOr13Zf
n7PPgJgEKT7RdloL+Ban3s3GLQuXivEWCoTOOjRRhTg8Vf8r92OOQeIlXehZTxhV2NQtqg4jvIHq
5Q+U+7wkXEJfHON5Rlb6d6/abG217JImcnjRUlUnEiyfonj0tRMKYmXFu8OOy8atdfNbhgwMLqIF
jbrJDFp5MlHiAfF6P6jSwWR9h2m3cQDKXCpwEmDKTrCwQV6TX3GDAJTO0nphaCamYr0aXB4k1jkQ
B5567YxGuUDlYlDTTaY/pVFiF7ipaQMzIrD/saAUbHyAfFOKN1OniMqExClnRX+kokySVrithuOW
rnicOJfdHA5XBvyw43RdIYs7U+gkCtGxHj9zuKUVJRlaiWGwb5qfh05X0nCmhx/SBT+8HUQoCfbL
c3c4zR7+DzT+MOwA0hh4TP0jJss62K0kQzX+s9vntiM5cr5/0c8goZFwLT5FT9192+qZJsgcNFgv
SQAJle6iKLSUZJGP3Wx0qrPe0O/ICi+0zXVIbQ/uE6OHfK5U5LQCXDdPJziQCs5RbEA2YxlYm0SA
djN7vFK7Rw9X3LgukmZ4nuLaSpWoK5KCBLVYQSNpyYzXSfd9QlB0DCiX49b1EMYorvsHClEa5Wxn
cyyWZoX7CqnQnqU/Yl2utK6Yv2r8HfhAN19ubJMMO7nT55zEfJpl8hMipTtGECtvhEiCvtIPhFjf
bDJXasirPjB+737+OVxlYFDEPPNkh+EFmX2GqHJMNm/p8DOybjNfx+iIO4xJPqPZJRPDR1WEAjz+
qE5LfEhUJQI7oSkJWWu/9Tkk0gUgUpC3eZYMvJ52k69nv5c1WAC9wUgQ0c1pcxk/bVkPS+gioJn5
HMfYdFbIweXARZB6fOx9Wf8oYAaqPvPUPGHV67VeIxMRzqLgWn+dc0J8Z6FyzybaPSUtffJ2iqNF
9EcwxsJR3/0C92I3zKwWB+U0/UVNGylBG6S6iGhlIiNy0/Hck/ArPJsNej93FmjudUZW4ofDWKAz
Io+W/eeOPFPClY4LBhUQn8TOX/EqwOXgsUtEY91P43kX5lks5T9xkKW54Meq7NgCI3T0IeY3YBcH
rOylBGQrNAOCC9qPyuJObyKtW6pU15/lx+Ld1YV6qvMxo8xxRjQMCR4ghnn1h0oJhq3eReqCzBSR
ouIn41h6v7Q0Ef1CBjwzILgIKXwkq7yluzsvrQnnUuydRH5fuG2oRkftMDTqWk9WyNBXYHc00M8P
Pz8z9Z3v7/B/CLv4YyQnDC2Xn1aY6CcTDa9Y3ram/ePkTxiCdhBgWLHQQcubDSyri4n0HSBpHU3+
jRI58kyKcnqoDwMAkRNHk9OfohPsYaxFKk9La49kQMxVVSPyjGV2P/l3H8BA34dV/vtqgxbmQmdM
Y5n7GyrS2GWpCrwmb6ovkCmywkrDmCOkMhFlnvsxQ/a443l8w6qPKfoL9HEndZv08yU1GMBCGCYi
ZiLyLPfYXq0lOZoLJwDe/OeXV+2V2nLk9C1fNS9ouMVyzVQNpuZC7i9o/zPEHaxcsqexhrPcM91P
2jZncW/LbDUSIcW14LtsqdthLIvCb4oGmjfPkVxmQqKGaknUuDMiC9ZIkKot+AlOVDx1Zk/OVM4u
7tNC0YjIpRN/ufBkKL0LsB/LOO5mYSsE/kzSt9CwiekD+rcX+tjCQ2Ntxn3yRSWqe5XLIxhKtupK
D1eOCFBMyljWOZEkXm3JvFZ9ZShVnp4HGQF547l7782497RbBb5z/KHzeeDMf02ymQtXH75WLrJN
y6yB6J59jj0Pq8bXIgevTLoxKFaRiyf3zapDsnz6IwmaQaD4rLrxJB/9Otc/Qdu7UgaQSnLCVCnE
FUshhKprXviA3C0lkqM1o6816y0NGG9GNYJrrmnL7M9ozbezz+wUgbrqoOleRRm8VzNblQuALZX6
SABPuPuBdhBVhXflEjsiKiWYOQYQ3SUFVGChojmZB3rCtL8Jdxbk3sfNSuvJ/vqmGDH3kAGPayP1
70tsYt1mg5DG5xu+2JcgEi1O9sndsPSP8HjNKxCy6BcFymVmTzGzNqlJV/tGFvy4VdoT5ZYqsA8l
t9ADTCoCOqnfQiozb2pXsTTjmwrYSopOJFTzhc3d1zbfiSNVsdYxXV+4GOsD+gvVSmhGCUWV5P+b
kgkl8padaQPxtm7Rp/8xggtWCuDAXHq39OiQdBEqcKhrEt3DsLBbfj23NYptGgJEsA6NPuEjtE2X
YF8AlXhwjQtItLnAwbJe6T2nASId8bUa4ex96HgtdLMfHie4e0TQp5cGJeGIMUMheLLG/wT+Wdky
jqKA96Bzuku7nVc4IyRMK+EHWW6El7KwF5NXkNQdGFQFVUvaZKj5apTHYebfooD1v6qmWNz4X04Q
RQnw4P8vbs2xgj7G7NJuRS4R497knVNbMSHkE53pjUnadoHdgc3DvAo1U/IbRUaDzVxAUWTkhnZv
UGD8aspX6+m9XFLUhJL9LZkJURcMVxi8mHlGTk+CVqPU2BeARAC9+1Fmxhb5Ciit+EeEMEK8yVeC
20kVPMCqTPNwRxws6u6sA3EDj3I8QeCw3ulm8aHHcvrm6armL5GxPNCgIW9qx7x3PklUJoX9TmOF
tmmqq7LdWpimMAgn0gZ7IBbGmf9XNhW6MimtaGVvuoI3XC7rLs6lrFbrlbFWDGh0cT9q1Jcb19Rf
05y3D9fz2K6/uihEyJ+d4fG9xoaAt6hOodkZ0LhX6T5W2Z6h2gqkg4GFc2gIShMrf/6jhG46bOz+
wKseFENTB5SL0L5vvirLkgsLFhBhJBfbYtNYVG8V39O/BCrE9ZCYnZZgUh4eTefhQbwcepRkMss4
8d23NVonAYSTVWSydEpubJ39L+W4nKH49a5R8xkhRWFMUyFuX6jw3cOdQaMl4MVF2Xpi/XEFjfn9
p+gV6fBe5rp3Ui3yfkHrO1lPp5SYrralyVqTgMLKgsPwEXLJV6Ggk5mnH+6jH6PMqLP1rBRZOZ43
O+Y/av2uisfFA+TT7NU0wYvmDmKbj2eIhkHJyls3bXUEaU1tv3RugrzmVjOKex3/FU6ug+Ul0UL6
qGjaJelwP4ByumJLlauDqKXdchST4Ni9OI1vo0gfq9i1iJf2ZXEqa3kxxLI0BqonUXNR8dxgeZK5
fMGvDm0GkTrDF/aYCExf3YWjAJuRSTZHI0Gpw20Tocer0bL8tH/rX/0f2JMeUMnFCASm4x8S+LzK
AxioDMN57zYRO/j1C8zEu4C+efNkXoptNA2w1oFqKW0MsIC/3xQ6HOFGAMZJweuNLcaFMZo3kWaD
rCgprMduZekDU/e1hPalMzHTU8rRwzG/53r130BdfLV2qw9n6hjV6GPjptH6vRHsR5NeBRkTKpyn
2vL0WrK13JjSovjglfW2ixJk6Ncc9AyTMa2Tyx1X1pcnmmhS/NUDZAyN6hiJmvtUCLO3elMB4zw2
v+fiLqRqSsJTyEl+pwuh0FEhOXxTFuvee9NkuvvJfqb8X1kF1ASvPzdQbyQ/Dq39131y2SkYIiB9
VJgbZkGp6ruc8OFewEOmwy3+7ekmMMwE1Y04VKXP1yONcERqwlB0lSBA0sM8lBSC0AxkRMT/8aXi
AiWGs9+iDMXhwoWcyU/GskJMNnxOrCiE7Pls+pq2PWqpZQDkrRddEPMEYgH9+vweBUG3S56ih4mw
6RfDh3AgW8jtC7DywryRte5E3ocDlIKvIFn+f4eHRb/6Wh6M6wDTtB3GjOJCmRc42s8N4ZSHvH/K
WWKZmE/SnCqm0IkKPVkXQbv+Xuw73PN1uoM1n1rbr5XpDAFCdXHL5ULz+FE/xlbjayn6tDicf24Q
AonxKPRzA/eXxSt/lORImpumpNMM5zW6jYOvzfbNDPbf3kKTpJHoGkTP/bRqq6Gn/lu0YM1Deun0
PCWKbp7ssM9gqkT9VKXtCmI63andkenehbyuO3UAwxfgxJVtd853UnDrS2z7wn8LKf1dLfH1/ZzS
PoMGWfzVufFj8pqXcSrxexE3/Ze/U/xIaTv59EB8idJrwEGE2h59Eh2CT14WcUvgisYeKrMsZtDh
3ktMZuR1uPeZaReJ50d46ePX7Gez5SwZp4gSmzmeUJ+vOHW6oWeM37W8nJfthGixA3E1jWeYk1yA
R5cy238nB/OOn/xhNZ2qY34E1q3fqjhWyHfyck/vxYHIfRvsBno2EbjNMp00s3+BrMxrI+gjnED/
8i7DQcG7r599dKqO9xgrIw/X1cQ/xiEwnKT73gjCD8pAKZWoNLanR7I075msaEofIXKyM6GZCPKY
iiQbIkla7ObVxDFBTsZLrhD/8lAxIzlPGlZtQO7DVUeTYlq07dxguHRvKLuJQB4W/N1k0B7obhPh
ZJWBhL5lj0BbaEaC8YGz4FrobyM/HYBkoVtXKp8QaWOR4BWvGboZGy83DgkWYqwuEhWuvnR5xs02
tFcMxdF7N6EWCL9a/wWCOtNWYRvf3Y7gTl0AGZuIGJiYlpxeBshkUl6nG23ygQ8FyTcHV4ZMbX9r
6ACO+h4yjAyUZm+uYySp9hbL0gmcN9cfByVb5N/E4uafHvwmJnmdYs5adpqVvbnVV4Jr7CUjten3
vdCn+9DlNUNvW47c0SMp6VMBM/d1DAq6AI6zOAoMuaitwuBP9/aQVVQnIXpehU2i3q/rZk04XTPH
jJi4FGQNvf0MO/YYHpUDaij0fjFdGMHAuOfu3LPwDk762w7hhkFs04Js3oVCaDtKMBl01ZM4tVaZ
/CqbdDDAXfTUuqyDp9DD+tn44yVQ3KMr6px50HJNzH/E5fvgvZ1/H/uRHAZk/WDLAIWG3WLKdmdT
0lTMiYXmCD/I8PIC+OBmInfpSPFXn9g03cNlahfvr9AAjBseOSWaOlAfkpQXRbW71UIjKi9ayDTU
vpZDi/NT5/ckQ5cr3FL9mWkRNZGRw28BTGaEG9ormZKRXhRL4/yS93InxXxahrN0cJDMxbWUDKjs
/cemxpQX2dYtE0I8Dl6dUvtDmSukDPwXyt3TTFQKRq1NJNj4hwaZFp89+FtAX8Le4MQuYuDC6bcH
aN8eVhV9Q8EHxp6fZI0cLz0z4FjHfDDhpn8VZi10JsmP3PMP1TtrdqM3PKx/wSMkvCzsZzm4+I0b
FyTFvtRfXU9yjkkaybKHlEBMXiCdAEmz8z5Cpcb7fDpm1xt4v2y6w2HMXf+S8ckvytN6UPV998kL
4BsVzNOKH5M4GWXpqyvQuJMV7guD6YEpVmF9NEpndnsNuBa5i0Bph09XyD5tslBsbO2RiqQ/HYOy
BFRkvkRk6N8J7F51rcuBYI3kg8INlwWke5Ug7PUrV79SXhqcbJNstZfjA0aLndccCLC0eZUwmT0D
+83j8yXk2xTSZm8mKzKZBj8+/lSVEuuUXjWfHmYgPp7oasF6Z6HQ2NM0HQ++ThfQITIIugwpCS6z
9k+Dv4oDx99Xb3EUweK+2GRLLj+UucqbQ2FstYEPnDbhwPT8tKaCOJxKpYqEmOyJBFC+VvUwj/Le
5yNSntaZMuE1FNL+oksXhyWbRs/CRlnzP+EJBWNuRIrT6vd/u+4gAkxwDFrij5JEQlbSar10CvYo
aVbq9IQo8Xuuet/NzfrlA5dG89goS8BnQKcwzdtt1s5zrhfU0U/Xjl2I6XvIthO+DNeKYt+RX8mc
Aat0NtNnEKOGzP5mGmKX+r1hABUz+s3RWVLdsCminTFzTad83f0jc3fVcasXpQ7JjFZuRWpxrHRT
gMmb9hj0o9Tae3SzH3oPqYXcqqEU7nxJlWl/+zvGWT5qwTdxvlPe7QXbePaVfN1923wKd+NPI2Ky
qYBltWb3ataWWrnCyZcEJggvpTXkr8Wi4p9d0zXVEiJuXc3ozZaDlLp+gNNZKWzj/edM2awTZUry
lLqjzpG3OElnU8DgYRZGA7+PAoCtWjUj9470uvbPMFX99bIubtpsXCsDzDirK0fiHtANb7yS8tyV
5zM3fwQPIDBHVQnozgP7PsfZ4r0gb97T+LABSDeU3pbEaNGx6R+tXb1skbF7vXwQijIU/pQexBqd
e0pGD3b6NUeiXmUTuHeQl3fV8e/9XOKvLhBp+YvyiMrRVrZjbexK0GiH33VeR9HqzmwNeyJus7zh
94egPliUqcfGMyORhRBpHOdnE6Q3++/oc1UqKvIVHFYDDlmS2tk70DdCexPkeSENwiL9Wf9ZfL2s
ZL4VHmmheKPF8BqXmZ+xQYD06qfNiozhl08QMFoBPIBxo3h47ujwiDhgNVeeR1OFw0NPutSRzHnP
SrPgwcoTcrjo7Og8C7sqt0lxmgb5fn0OlEbOHj4loEgYt5xfXiN4Karpm10FQ6aN2iphVvvZnrzN
38IzSOODSlMcXaFlsmEMnaZpq1BZIGir0Fxy6VaF/2ejKG5lf2ddSn9eQ0FNmYD4dTGZ2biyH+wm
XPspyywNbpk5Nh5R+/13k6faL2WJs4GAmHA8XQvfjWPDbGsEil9FBRxL8ji8QyXm6VzpjlNl4RlI
Iqcy5P2oYgh0Se1LDj+04SsI2Yaq1WA7AwTQt7n2h/bfKsIZA3c61IE8z1Rmjaf6l4358xlxwnOX
w+NabHuX+U74/XIo2IfivQ7bMrWEJS2H+sjQhLHjOXG5gUWOd/hzpseOy5nbdXXEEbWPqNt05LVG
RtAXrVqmd4Qso6+P+bTKxi32UnFiaV0hEoDGybgyMot/Sd/VMZcArs43jRh8V03fXr9+TSeaKbl2
XE/KFReV7hu7p5gWIl6GnQlq4qPwhhYRtMatYeLhdE3voOMpvZCsYKY8mQsq6Uy21muTov1/T9Zd
Z0TDUXirTOYUdH1reLigtCDr6WczVRv2eoEeB5fN6jvL/eeWqtYKaqInxrLXcpH2UuVcJmjFiEyQ
/TwhFzbj4Nynn+gor6QizIvk+KYw77IJR0qrqTi8fiktOsDZ82xaqed0WTEVT3nacD8mvWRqKjJF
TXVSSdjjbTKdoB5RvN2q84WnDdly2leGQzH6tJ/fytDVHHOv9OHexn/3HKo+0CFAmIyCEsgxrcyl
BNHSBnNPDWFWoTl12668jj40vIXdPxsOnHeNPY/cMS6TlIZbpAwg/ytzwQ4n3uRJUQ4aYVjZTSub
ymb930s3EVghZn0+9Ct2eXPzzkzCUR/LcjPjcsCQgZsqzLQPBzPe/KSjoqbzHJCLOEs6aMYUV+/D
TlppUFFXpiFgo70yJAGpkypkmT51Q3rn21JUJDz6n7oFetXdVhp2DgZQ2GCbVh/JHEGyTK8m5gnb
Lapwd5uUWDbhfZei0eWwCbTeMV4oMDLtb9jSv3WIfp6o0xA7eRPUDcMWmzzbssnQ5+O5JXAvUuZZ
5bks4M7zIZ2p73dhV+5LMR4iW/eBcjiJR0ZjVyA2bFGILyQq947bAuBn4HqWkli+r4oNQDkRLRar
fiyG1cUVxLqERnh3EKvgFaOt8GxY6OiQsVtl63D4GcpsEJqgmhlk16FeoHDkgUrrG6u4ndKW5zBS
TQUUwUD0wrjwzWbOWRYKJCEsRyr6+EEYKI0NTKNUgp1h5n3v9+zzMQNLpQJGpVm4PPb13neQyUcH
o9ISBOouZ5Q3nsyHksm7NsvQmkPLHAHPimhXFlA6vshhSVuermrdNtawRgjsRpWzfPtEWDfKfD+T
Icpg1uHrvRWHeT792QevlNZj5c64+3cVdCVFVP3f189L4PXfIg8snI+3nfW71DZNEEtdXse5J4Ht
Pl0MvMcmf303E47WQf2qDE8luAPPu1s9vBp7P9okiicdneFwIYUYpUeNvNFJQz16/rlS8Cd0OnDu
W25bd46CTuHUtcECopdum+MiFidezjSAkdGSliBYzpj1vf+3zehJMfKBaUXCME9weH12/xE6pIxA
NYboBZXr5y5Mt28TmcbraMGOyBJ0sOadBqPvr66RXwb2TD34aXVwNDWUX6HPoAmecgwEPkPn1dQs
fFuPfDXNvTJh1pp0H8mdtPvVf1vSbQLKBRKEH6t9Em7D8wkcAH5t92RnT2Y7sem04OUZuoBsl1sy
39Lul/lEjO0IcTEIsosqLrq62vNqf6L7O2abmXzgbEOmV+8IcHAWnA/OVMju2Vfaf8+dSgW7ccPF
u2iTo3DnTpjfANRvf47MZoHrpQyhgOG1C/DT5RSNGEzqByTEsB3EsuLgSUOn8N5LiR7VDOzWsTIn
PQAyj3b+muwX+WLPy4KX58sGTlNtkmUPIEUMLmCAZz4601pb9KFVP9mN1SL/FdcCg6R9IoFBnE/+
K+AzGfNUE64dLSsCgsBfCyI+wt6pawiT8Yhkv4jkHASpL09alZF+V+73hcmiUE49vgQK5AxlyIbC
eLlQJfttbJq8ul9sKp6e/J8Gof1Cr/uHqwhHZMGYUkj5qqLN5hPOWB7Z0t6QfAUaw1xx6e0Jskyb
FtBtsRvEjv6KpHWS83Em/BXt7wDgQju4NstupnpDhpiVRe8k3N5uLQF8hyrOta3vq/vGCxch8w78
oHAcAQWMmgonOdp+YR+IVtifwdsiMrIuBG9aQZoIITafAYOs8qK05m9QnpTmfps6E5B4rGBNN5pC
Lg9azyhpCSimOW8WzZHxRBX/OxpESHcZQamPRBrcIZABqLWcSt7HNE6ZQzn4C5xV1QlsUiYprwGa
7D6PqyipLxI6j2Lw1D97qdho9PT0LKLdHFzltcoGj8mwxM8yIgC/e7vEnq+zLBnOND7e1oQFdj2K
DC2Z9ijwHx2QRdGN6O1UXuUc6As806YL+S0k0Ber1c0aVMOhB0Pjc4wCU0yZ1kAEMs0oeCmNrS5i
obr8uLnawvp9n8mYunDRCLIQgAXgCJikjKiJlqgp1/929LYIhxyoVjKhI7k4VdJiynMbMTO5bKWz
oNSK0+Wwe4DLRGIdjN6s1h81si2pJX+UCjI+TZ9MV1/hy4TheK3UZu62L4gG7LLnlSUaGRKLe70Y
Lot64qLA6qJYsS4D+hCWFgEG+wu6i5aoibSNC5fvnbDPhXfU7F3o52UZqujAwp6zfeWk95mAbVfN
atgQcmpi05ug2t3rkQb1wsktX/pKz5FYtQAzszC51pJjlFWDHF0meBiQlma2+ARuq2YIdD2I1on1
xTIWYDHERcO3EsY8yWNWZ5z0fZDescAvZ21G+Ywu4rybWAr+jW3712UEeBbBFOq62w8LffFLX92F
bkR1bjbT+2k07ZxkFU6u1p5hocSEqZ9mPDxFZJdoJVJMAWCBJOm6xmOX4/hZFtKWWTly1DLdxpYi
pb4eEVbg16ocabByhC94kHESF2aXeVzEcFXLUIJf3/d1mrdxHC1GYERTnHaaOtlXWsu+Fyy9Ag0A
b+mmtqg925CUckOrqIGbtgWEWJGIAAhmczsqRSu0MJ+nJs0TVRKHsFnAvXxEUK8DDpUo4JIKFq93
ZLwCb7CDvjxqdtFBp3yAVwGfMff1SSNNqEfITyOpkncESwT8pH1/Zw0XbulPEkHxJKLKdcgjta47
fVn+TBOr+NKpYGQ5iYBttUiIRuqWge9x/QaWKaKBi6iNM8dOoTVjbq2l0EP2H1VJqUbRooHREpuE
RnwEPz0ockdh7CMWvP07M0EjSHHKWzjcpYlA8FI0S9DVgGBkkJSze+5/ztR6MqGJLjx+TmsZsl/h
Sod3HhLgXFOMjZJKxtThlD0K5zO/Kek02lJ3J6QiwjBpedlvP987BG3vCHBwlu2QY3GRNLbbhqa+
mJVcwXoZ06C3Tlwfsk5CHF1AA/2KBWYJn4OGw3CFUsCa4F6/ULd8L1Di8tRUytADFttUUV9tNSiy
AS7r7fZWOB3irSdBZA+oFGXp3bXf78bj+WP6LYO71DBC+cHHLKKkFSNSPI9DazGOyPwkAq6CF075
usMwxmrS3UDWxkDt/ZQtsh91RI3oiCPa3Tk2QFOsMr8/uTylCNWltLpWwFuCYCiXmF0i8UjdQh2m
3WoEiymqCiwQs2hNpGCJeawoIOF1g8waeH+zCkAxSuhsYigl1JCLpKhbvTsyd+of0qI73wTgLo/T
Xicqjd3Cqvpz/PCkrubfxn7JsSCZ5OqcTfcoZSf0jg6VDYRKmJyLvjcSV6huSIwWqHiuYeNcmDwa
RPJjVMPRhbhFxOVtHUDCP4i8GJQmPU4rxfzVEQj8mPUIeRlgb3uW60qeFUbV3R2OVF6ENTAJFreS
Fe8ywhPsWxbEd4yatjWE67Tx4w9N/oxy2uqwGLsl3YY6hzNWd/pt5Lb1C/JLKM2Qq7Ci0zVUYlF3
7BRnFhyw1IZXqtEqYdPojFlAHWVaBnfwuWU01ev8EobS6RPmlncAC8S6GBAgDw3bpOiwoPcnKyjn
L7xXP2IhmDZLU+Oh882RzesUUMEPGQ14KW1e+V2VBLZCapyGXCTmF/bMeFJi53hzfz3Pt2P5waox
CLI5UFMKVUQLzDO08hYF4OIsNoU5V6VoBPgjJUiCjGfuO8AuM+1IAXYakacKJgt5XP4VlExVSN7/
bLfe0KQDd2+jf3Vf/SG1ipFPrKX9Yzg4/KMZ5HcuHdN/MQi626z/xLLfvp0SVtnujBYu2ArQepCt
bzjoq+4LOA1WK/P9rb81r362EbTk8o3E6R8XKZi1Bo8n/bWk7brXZUHFSOF0y8JSSScoMmsJ3fa5
Wiez/hZzRvGSRV1gCuabCTxeJIUDtaHC2GaVMjZzzo3lcCSL6Mtn1RnRY6B33pUCW3SoW9Lc7Yr/
8bd9YWWSWde/vCDCZc+ONTiBcRE5D2QhLAKd1jX179emGYLHnSF895NBQEKjUw9ulblv0Ct7PqYm
yLarLkxUTnZbIM+hNOu5ovTRuWJfqTgJmesGHyu/LIQbjvb3ggbjitoRGSaemHgAZebPXQjq2NlM
yNVkRN2B/S1nUOIrVXmd8vc4/REa6eXBx3J0Gw97KR3OeHta8/VtUVHWIFRev/s+HWAwdHoU3fct
oZvc4OFC3f3pibpCjfxyHDjePHPqr7QnVKChURvSS5430DN9xfEvVj8Ci0dD9+xjDN/Ql1+YBq8G
v67LjgwJ7my14jNBjpHRfkW861OtJ2R6/EMdg5L6Y2TfnzW12dehrOLyURZqHG2ZfYQLBAh8n13E
AmyBGav9rSpFX87W2JdN/RF0/RZxlhpYhOWadJNDcqECqPV0gOu+Wle1DVxIZ9WsUuML/W9xh/Rh
ypu+EBd4PVZAFQ8KqSWRVTCJ+jregitioth9kNmZD6IWGE/qMiAltn67kz35wGm7qQhe9SYTNDjX
V/MO0N8q9f1lgGnrvlaYnvRZ87Kbm3+2a6WsbCGy26SF3E19y2FEmd50n3HXAMRZJ37LTmmuaGVa
XT32d4uephjjbtcizu8BBE35JZViFcmLPrwNR04N2qc9J2VHr8sWC97H9Durn9RE00kyEgvIwonn
wFTmXtWx45QXkhRh2XjLrNtFl93LqKhm96FrXrVSV5aLOeRyEE5N46ejMc/vsJSLMaHXokJJOEpN
Nos6mVmF+zoI7SJ8VnWTGEuOW6ZMWcLNaKdna/F7IjPCiKFoX1gNE9mrJcUevzoL92sIBsU5O7Nq
jB8tysbEc9pLdahNchyJTWPJW1xxSV3SV3Twuv2/8/BNYZ9DjNBAvXYkIyQZer/hRT5xYyq8aL5r
Ce/nhlcAKmsth9ESZZdYiyxHFvubsTUwaxCRJYdKACKLLY0vfLBCiroXJFbpOrzCy3vcQ97ya8DN
lyglaauJq6QII45IwmwhztrZ1KbF0Lm/vSgHGIwTisDmPjrcYRLXIxArwPcF1PqDv1R808Yhf7OF
Zlc8ws2jKG3OGNHIGx4o/b2kMcOW/X6G+YZm/WzmAlQXlWosh4I4ISYRGXroqlIKB8VhstxFx2Lc
7u36UFEPKkIVUjnSO6CaJ66iCucUGAhwJlZVpLHqnX8bRgZ4RdAWmYfEbOFdj1hXtV0HQzuQgF+V
+G2yhYL0Y9kgAm6vuhXUyno2b/M8Ud7rGVWWRfgUpfv+5GgXHrcR0CTLsaETV32xTdl2F4b8gLhM
Cf/ttxYdNog3YesNpDccuTsvPPzLaxUgd6Sut3tczUwOerxRe1NOLQF4/FOZZABurUAIMl1XJayO
kmcyVbUVmclQF91cxqoI3lZRUBEAsIndmcPXmQYliPCgxC27whogFfBlt7D2kZsIfg9Z7tWcETfJ
aWmtHFT+N34tgNSiBcSEVH+aqPReLUSoJCmu/HoasGh8kBs2aLUq2WeJktYXedsybR7L+eGGMdHb
m6D+W0b9y7+9S89Oxci6RyQGPYbnAsnl5/Hkq3eIR5qkPY+ToRFKwztmozgNO9VWoWgR7ttKjVcM
2pz1UB0yAhKYn2Efq9p3QfmMgnWljBuHyMjxcLbXeI2cGuU0JSi9hqNiLRPJk9iIN0b9LoFLHmcX
XeLykNU3/fek812I5a8qDhEyY+88nefW76LlRR4UOXwpa7YtsyANnBSyz77/z1awfvbEYLNKSzHA
oz2pAes1beDfV7FE4zaSUvGjO9D7UyOGwBnkrNjJpO/0Mlxh0VNPdxo/1RSqgmpGKjM6vpKiaKww
pE0NFGtx4OhgxH4uZkX1Ou1QpiBJWpUm/eREC8GyLyYSJu5wTceFCHG35ty6oMSkJeQAE0G85a80
uRmE+ORDTz+2YZ4qnDwizQC/GONpV/CO2948cED+WwDaXzzKsi5LvV/EST0pPB9M8Vc1sxKQ94/r
bNrUJCwCa8ljCatQt9feNS0+5gb2mWGURPazZccU+efayhPG+oyEaHmCkKpKvGYjdAFiAHr5bMfX
QKjdlLAHZx3JXiMlG7m/ERZBiO0h3/nzeGpsHyV2h9NuQbQ261vi9cAAm43c3+wwiOgrP9KjONlw
xy66Gww0YZgOK//5v0o7TDO3RzpOM5CjdroVRChSlayJHkYUw0x+fsTPaogsd1HbJ5ML4N2RaamF
Rz7eJfwPKU5Kwx//jF7n2t4kdsvPrcTmHEr8/9VeBM8KEmeKFCP275UqnG8pAZPSlyt5i6hTorTX
fWrc1aim0hsx72GJZJV/IZb4PUmumPvETjYS0hei+ObRXTcl2dBPor5cPOU49Peq0ELPUE/G8+o6
du1BS7MDmq1zBzYtclE1FEbwUCsCdDL350GY6+crLIfs3dNMKo3Qvaq4Nuw3bWNEToeovIBMmj1L
LAtAFArsc2dHNAFIrInhGHY2wzQ7ZzbSK8C++T5TVjeF92AcB25SDD0IOPFz0Phfq7rtP/3vBw6d
Z27RsyKczVd6KcV0pIvnPUNfe3/iFmvBrD6ja2CWEryMGL1GF6YF0H2tgLFB3RIE4+rBZrItzR+s
v58E/fSXR3Eu+bq2AdkLT1fvtkv8cu3wVLd+SQGZMLpuiqJCE/9d/m5yejcT3OZ7ft2AHuSSeiq5
wP9gTZIkdunCO8yGOKEXLcEiBZDYlzvz71YE+P60tnprZanjlYIjWp1zngoFQW5WpPXjqVpp9WLk
oEHY91/5rHs3Dt9qAf0YSO9IbMoRGgZ8Ij8c7ucpFZn80cdVsVn1pOoV3VbeLo3Iw5wJUWrPErwk
WhA/JYeuCYyQxSnszqUr9Az/vsQ+m2qUTGEXaPCP5C4h+OZr/6LKoxJ18mTnxekNb2++n1o6I4NP
3nI1+W8c6Hs3H7La3JijR0j7eGc6xoaFeIhcmp5FgvgqY09HULDtnIqdS7y2fDTCQ+nfZ3///Uja
qlwUB+fIWy3vVZaDlHsLxi8RxgNg0Mr/QPSQd5JoKmKIhg05LcJkDbEM004St5z2eKFUh8Zjpdhy
JT9nZFecbZS2Vmd/PdmgalX5bEHk+HVYSN1d+YiCPLEE/W3kUqHIJyDuX9vqBU4bPSYKnG2jYPBp
hWAwoCmocxZoHfvCtqLD7oeL5OnzhxE8Cv3i9DOnxnUn2CGo+UQDpY5XEWFHx9Aln4c+63o5ybQR
RtR56s2AeddkihHQaJPMgd2SPaagDh+cm3heZzYdKvMzxkGkA/H1L1ICrHSKHObv/649LX4JpAH/
tmVHKVRO6Q9xLLjj7FBVpaUkJNqwc77Lwmk5Q0OXOvCoErQ2++407b7/J8/Ceq/fwxMcxQJ9bxJ6
UYrr7EB62BdKV2UO+0MKEaKswy78gJjtjwmSFedU47Kg4gSJP3fALTrz4GZCtcsFNx0QYCv86/vr
FUaON5e6AEYJcCfYGuG9EOtghGa4Y7s6PuxuL7s/AKKPG2W3E6qo+khjFOhtv27YNJzy/W1SAR5y
nw1qDWoSKzYMHlE/W4zh5J3Ne3zv33cWdH2Tmb7r5QKWIS6vmTAno4htKR1Ny0c8f1m457htxTW9
irlX6FQ9jRBw/GD4V9QhgvOpsHH3qX+sv44sK5lJkvU++mQ1tNT5+5934zkPrLroWnf9ioCnvKrx
m3TO5qx8/sPHEf6E1+1D/dy2tlXonxape++Gxpjv4N4JEP8POHCc7dhe9vQhUwcFzjs4FP8kBjzV
VeFA4Zsi8i9kH/gjcPKc1Pq7f3J9vZdeis2nPIIw4eTFEvklnuzI4u1/PW+Eqcal2SBJsJ1lIV41
LjgRhx2nV5WYu7raEhSUeCTdusQ9jdM6HZz4YyXZVgU5q/7yqhkyDxtShqJBjY0VCqL7CjVpGIuM
7v2rF2ftwFB2nfxzolq0+YZdeaKFx8qUjOE5WctBWjpuimXqxfjAvfiK+op4rP1Eu7YgWoFhdW2c
OxMzAsfent0sY0fZZD4fcGoKuXvTbkXNVqQjBChCgDGNBg7d8eCUnqkuoQMvEFcd8vWHtvsm59bk
Q023A5STifHZF+5rjfmxsEPEGkdi18FAsE3Orv5YhbmNrE+rtZx/cI3prnxn2/Fd1LN6TeyUo6WK
VPSLBKCRbwrDr1/5hQBCCoDLDOpP7D1mtm9cBnE0JMujEbNLL18s5lu7fWzWjRLFl2kdG0YpBpwU
9TDbTKnSzdRDziwVcjlMAx09vC03BgRKEfZzh0/CS6NELOx2J9khRo1fnPWlQ2RfHyjx0FuzzH0f
YkHbPaPnlUklvEh0c59PsEDgEcMIIrnITaxEIn4BReN8YIu4T8OcxYhlyNhOLqF9DtMn64btWjWF
IpJwVnUfAPX1g4HKMx62TmR7jkfZsgBuxEEA2BFyass/95QeNAW3duYg2+gDGNX82b1TdidFZHGI
tptuS0pbDqxSLWS71cy+lintX//uUBlKLTpvynhUsOnP4dvuD6bP+x5v6rQcgbdzGr206KaW9JYd
7nQBgSCmqX3BDDT4a9H18Pr4MEGAqmeCZUkyAE7xMyv9Fb8TZaVPBRHgID+r8Xi0OVDJXgWdrrW8
UT4NogAvys1Qg8/l4UuTxsEHjPZg5ZakjE4mn0C7KOIYx2ifEj6NnkeHczAoEU4NU0h6t71yFeyd
+HosIqDlV/QYW6WcA8Y9BQ92K3luCzym8hcInqWHk9WEjmVTsoXwWLLDgGkPMMDSjXGCz4oL+amx
xEknzUS+k64OEFW9tq8nIJmM1Bi7XtMiuQsOtGrLVG/CTqaBUMNp2Z+6Adirt8BV///7VvC/tObi
USxc82LUH5QUNp4UwhYgdOm8/4jZLQ7vMltIo0gBoCDGlR7KIG4AIqZWN9Oztby+5q8DK7R4VOjx
JCHZdhIpZuD/swZdAeW8j+1a/m8z6bjRGiK1/5KLMPAYZ+0AVg4Au6N31sOjXYPhy7AnwjcFckzX
opYJ4HzGyVyU9TZ3vgXG1CjYIcggRGrWLEGKCB13EfQWT07GMLO+pOhpk7vW2SRgufKxIkVTVfJG
/EPnObL1bWtP1zMHzdjhpLQy3AvJMETmUKPw/eojybfsurnE6gU/v8Pn052ZYy0T1SgNQzWcMC5y
l4xFd82m4OOS8WQv5OThsY/lPhRC7ukIoUGjQ/hXJeVJEolsSO+4vw1PbO1h33T5kIcIRQRYj0R0
A/T+HxOFMiO9+EFOWWESO0Rg16tf5lMA12GJ2nYkEXrrHmfgpifoO18IXjCU+QsHSMCP8G3HtN7c
54HHI+JpCirBR8tHDOjGgZ2SG0cXO3U273THH/V1TNrkgmfcMnW+H/bkroIfXapfa0OuJnrcKgEn
8RYuWJDvX+MNkZo85AoAT2sMjPmuYzWLJXbSVvy90Ri78OkRuj2w0TODGBRutq9dlLswJMD9cFXa
f6wjdJfPY665D7X0ThovE3Re3D3x1afllUZF+VRlP5zulcUDQJOTfxwoXXa/Fq2WSnK26YCme8j5
ZnQM0EdZOyGf4E8tYovElQU6/XsByi8QrxuHY/HrObCPQ4dnS7E6XVlEgiYp2Du4YVvLkrmDxQbR
CYhaOJffrkBoHx3rfB5FeTXqdDcN6u1GWW7Jo9uvpdqUvXUqmNTvIK1kT+VPIaIPPszbVh7SKqIO
mHb2FXd9C1he7eCWHpe+BjashmKvj7gHFd5r9h0ISs3UE53mhUnX4RP1nj/O7rxvDGrgnX0K1uP0
LrecmltIpWa29QrPrJAvfiCjGlTa2d3NM/bj/O1jM7GaiFQGDTAL9oerMuX9Kgosz40KILcrj3NU
nTv3a9taDsFeElN7FrGa2TpFaZtL7HOG5x/KXXiE/ffphx0kIgLVe2I+6zh5BjlEPGZcFRXN51Di
uJIp46aCUkkJJfrLh4wJDrQf+xdtLPVyT70KFio1tbm4OjajUiYttaybCAyBRI0LDzPfzEKIGQRF
Yt9radXPRVOBB7opgl5vPc1xWuvs5CDmDGvR2abpnd+wARnPjQ+r0MyuMcGh5fstW83rU3FEGaEa
MwwzoHZMTdbCscwzaY+O6CD7f0u0+WibmROaIJuTgJDihPEa4cUwduKs8Ct5G2akGGiI4rZuuZ1M
FFyjM6qFspldQnclvWrd6IEkCHzuZ1rEtdI/hg2oSrkx416hoCJ886LwT+JQm/gFyFLxqfc3no2M
dkukQnwsplNLyvZKe4j7G7K6UMUUdj+z4tfj+1K+YeT1pb7Bqif4vtVJ6IMszxRl330aLU9OXRGS
0b2jrGa2nV+iDlwgYMeCSfyDD0CKOGvQKnZaNDrQ56o6qkU7hPdUCiels3FR0HbGeBelX8Dx7lfy
nUbmx2IThJL82O8d5Uy/tZAHdHu4qt84xkbAXQmuJGWxZ7jCpC7lmm0Q/bu1O5/o6+2SG5rYMcCd
DQOfRu1Lqcd2u9arpzWa9arOf2MET0BEbsdcxq2FJ1JdgLqZoQ+TEizHYOoHo5a2NFoXuwaWfiAQ
M5zq2hCg3a6qpuvFp0ZOMfoy4jB8I03dNfGrEL6+kRIW1HWHvGW7p1rvkCqvXPmXK1ZI9nHDjr7R
uMyNBOSIgpeb9BMipZKjvkBioLtoEllcLPKEo6wm39cVIeYVz8vCvttvJ+v7A9FbvW1kuKFwsbsL
Mg00Za9r4dswQIqjZsXlNraVJECom4CGymgEZd4CxrKFyMk1Yf2asU5ZSGq0MSiIGo8xe8UdarxJ
ARv1mIxHh+oi+t2spRLENNzcrmdu3ohAb64UAKrXRtA8+zjr/ZL4xkqUQxsZNd+HlldwZ01OkGqE
Kr+A2yRoEpmstXEZCnxHhAuo7tlrrpIAHlTcI1KoGzvd51qw4g4QsAQOeGosS9G+wARCbrEBEZ6n
PUz+yDapOWsHPglp5vgafU2l0z1qREoraIbZD387nMz6qb0spfF1ExG++EO72grEH9ISq+4hmX04
8WJTCXqyMU8Q2QjZPUmXSuBRbzOQPoAqCwP7VaY39MIVZUbhDdBkRYect7lclEW7xRlS71HUDVHM
V7VxNj8vs9klQh8Ov0JC/fAyd5n7GApoU3Sjtka1zfka02Cl/m9z4tbDhvOAqqWA13A5dW4PzhWj
WFsGM3PxmESARnlSeGXdi4t26ST74hB9zgetKdvupjwSCU0KRN36ye2XkjxE41T8DuVarbWOy5YO
Y4BUY2m0Ptwb4YPu5OrYVvet6z5C8CoRnakz1NSjFlRsLd88GjWho8o2eJj9npFTUm14tRqtj7np
EXtd5NCeud0pshk7CLizwo4AYwoeZYqA1UPdWW2DFomuByl49gcMb/Jds6BQ0VqmUrcnQgQhLXQl
QNcxhyqJGe3LWQumzMerskQZ03BTPiVfzFXu8Ysff9Rz71byqNo5ZyI2BhPmTVZrX19KolWtRUuA
9WcuVcbMGSS3lZjM4V6h2eLDkloto4Eqsr/sV3DfPMuQ+/GU1XNimuzFUrEf0FUxWRkW4OhWjjF8
/MRAQubKuxZyDRBNJ4bNqymcfwjJPrK1+mBUuhwgi+cQpdvhX8iZLYyg5CeguymeUTB0fjPPGYlU
wBwacf/ZR9V9d7cl2TkcSj0PW+LOV6hSaX8803CgWLIyX0jAdWjxe7+GOlC19R9hIJYo8AO6Ynp+
b9BMymTvwhPfgxp5BukcfAUqc+bQoPJyI2f+UoAQG23+gs4b8hk3FlJq5x6FkmemyeZsA/FytePR
mKnxrYsHbvAJVBKq2CX5mMwYpAVyEHli2t1ELJ7T7fjHIWN3gUV+WIuCgn4L9y5FzAN6CWSic2QH
MYC5KyWtyW9KzXuAqCLg8jMGYlk9hbXZj62K4bxucFpjO1ltY0iSNqq0qrdsr7NtDnoIt91eoAfH
e+ta5sAbl5l4DX3oGc8NJYwiJHANxFokYEmf+/tg4SHeYE7ncDpfKaoPMWz/ZgxJBHl9fDeZMBJJ
/RroAbLMvPLWrhPgcK+zsRws1DDTrcG358KAWfPvnEa+hfA6DC56fSoXAYb4AZ+i4kvfe6za+H3Z
1rkVDN7RFPyOiQUb3CCex9rF5CP/aeeR31ef7GWAu0978HEsXCb9sLakVtKdC5lxzn5vbdjK45Wj
uhw+c5DApr9C4mx1YjKc1z2g29qUdIpn8xi0cBG5+oVZpm4jM21GkDk0r020uxi5/SxCdCim8Q24
rUgyoY05OEb5xSjqz+cWPIPLnfLckBiiRyjysOxL0ihGSB0dI7Gc6kwjaiIEUHsQMV86nI+ztq6z
HFhe+gFqBp+b09gIsb+KVZw0aGc8+WXVxT6u6eAUn+AhJtda/p813JQNm4tVB5w4d8l27FKhyzoA
lHm48Th0GZS5BOKpzNnLQfyDJiyHIEnlaLUMu0h01lbrKfJIaRx56HuGHd2tpHIZx7yrC1afmvXo
hWZgXVtNR74oKnjc2OAocYiBaQPZf+udGLYP2owUSnSqZ2Xr8RYLpQlb6p6H7rtfY7JXPD9aPt8K
Z7H9XtaLxh1ti9oWStK9ytr0qOEJVgxEACV5uu8XFTaA5XSrZ8O8UK207iaydRmuQQJF42ZPdOTR
6JY94bBvhAekDwC5dSJyLAQicF5d1WGfUujRmITD39JrXd+x1i3D37C2mWvN/sqPMKmaMiL6M7cF
JFzsJt+nJBuIWaxK0PWxlvKbtSsJ7zPIcK/JNLKCbvWoQ7jdUB3vxlpZ4S/Kj/e1OtxIJGC9gm0e
epnvyS0zw+Wx0mUZXoGaNDdwRdvrPQaUkJw7T2UZyfjCbynOViZ+reUMGsCirgDB2SJqrlBPZjex
7v3R/1hBbhAA0xxv4dg3vWjvmFS6ZgSxbHxyct1r9e2ytdnWDITsehHU+jgBNXK6uBgxsOB0xBSO
kNhGI07/j28XwSM5EYsjoLgYBlF4RDuIXCH9ev656UeEYYZg2OQf0QZGNJaoRN1NFzXTP3NyHRn1
NrsdV68RCCFl9rABaQ/cxnfLulwKVF6r6G04RKTN8O0vbwwbIj/LbbXOacsPaD/Ebso6JeSmfxNJ
1wYqY9v2VmttATGapckyW2qh2uR/9Rv3RjCB7I9rhMMx0BmXqMdUWaUJwkU7bIdSSjQWk3PwIkLI
WisvnveSEobrNJMK+3PVQrc1Lixmhm3k5Xu0XEsqomU3w6IK48w+YbaA7xNz7mGw6nRo1fdMAkin
5h3Y3gty658waPeFqMTqdugPIHkAH3//tgulVCHcQCTH6Hh4Jqv35uCwoyaEWjnlY3Sy6q9FSnTl
MzC0L5kUkRkOPv1MOC3gGYS14fbEZdKp13w6MH+BrQNzgGAXhQXJz7lHRWVzU+v/sE0cDEPOnz2r
jZXAb8gSXxwgx1R3vZGMpggGF+vZ0wLMA+HRVhwvi321DwdDLwn96IX3ceXo722Y3tePfF2W/PIg
Hmg4qyC/6u3ULHMkR9ABY+IJSzA8IkO4ub+kmc15pSNQikR0s3+Z5Lvd23Wm6OWeQI8lfiWWuMmO
oCbs/jcvjR1cxuggy602poGlPj+k27Ebt/6xaXj62YR7wiql+OFV/jiOP4lFhN/5Lg9jXV6MWA+L
qLV4+xwFE3VbxNhLUeYBt2wkrb39za4/Vt9VqnaxMcb8gr27Fvo1sd29GQNUetR9ZTywkiP8gkXA
bRL/TgFBa7rUMNAC4QBVX9AQdDDS5mG8FioweIhsWLaa9ADwt1wDXM293D24axUNDWeQFF0zM9H9
Vcc+YSxhWwZvn4K666ELCcUUbmFxgrKjA6EcsXn8lAAdlPssvXcbIuPNJJuOn7btDbe9mjmvyAkG
yLl2o55XsWJ/dduCuz4U/lFQAYEwvN6Q8pSSHIlE1YN8QJFJkVSbSEawj43Ts3OOq9bpGPkBu1Gq
4OpcbXgmksTIicBW7bbY9p69J37s8jOZkOh6un8kI+GIMqwgYtjQsDidqM6QgZlI9cvn2K9J39zV
huIbcmoMbByJvRfQfXWA46aowgeuVtQIphOAMjCob0fQUgAuSQoJ8Y3X+ZYt62czR83swTmJ9RxP
6QfGHxmmY/O6NueC120QMU/lpGtX+oQWwFoIJFscowu+ebm2m/vpMUVZNxTyqZsKrRTKpNzN6L44
7DQTIO/ds38xtTIonCUPA8tUrzlCYpeb3/5nI24uu/nwANzdWwHg6D2mKB1+W3WOKW/VWHIa0M+W
oIng9kXVrNmxELIi44XBta17KdH/u4ThmAXbZnQv4v7TJYUs7zMJxdg72LgyL01oLyD2qnZWdWeZ
mDgDo92QuL4CW5TkbQvLhAvFlh+yv/xvQDcaUrlb6h9jXNcfLhhhX6CmWb19z09iKhN7DYhYmb8y
kjAMeYh6vE3sqM+cWjHwYTeB60DYFjwndiRV2+s9uAYVbdSGfeHVKw6NjAU44qGTwpD9Zh5gFlC/
bFvRtrqvmONzBTI4c+Mb8IMutQvOWIzSRGDnJjsCDmKIGhdy40ZnyamKOZWT410uDQsIY08A+tL3
TcqcyyEnV4oWj+77LYfknbRJ5AJmA1VZcVUxMzOf+VOdz5k/5jVLjC58pUfjbUkrI/QbAQ5o0lER
jWhWZbj3zoEGmIzbPWTLtpw98hhofYRmnOyYSVlqoy+5zL30JO4AaxFfwqMNmuUnJryDNoiXydjU
ouL7o0Dz1qgc5cgVg97h+0goDjea8tEAqZkMpCMmhJi6h95uW144kChiXvoF1zu7RJiCh184UV+H
kBLqJ7CLLmj2gYig3Slz5ETNErj6MxM9K4TFSq6XT7Mvnb9JjOtrHjRyk0erEcOHAvhRxTG9aEBq
8KdiczfGEUD4ykBZoNrm3jM0QJRI5AdhG0NkPAqNPXRWirN6S3WTaisLnPqzEnh2zC9/cZovgrnW
6aXPB07cMocSwPr1MIgC93PzcdVGXORXpJzHXPWgCPQ1j0MjSBAWM9Liu+9FWJnEgj50+W4S0U4v
UmRhZRYnlH7KAuU8WvcbBrMMR9wEXKBUcX6EVjUSQ8L3BB9ZnIgGCBVI4Y7GcuNHYWLLZorXqstg
IFTqNhdH8z4Issx+VxyRLcNV8K3acYDUFWwd4ShfvpTURCDcruGL1ltQRKM0iTk7e/xcCNHs9kX7
lYQ8y/GROBfCKjAli90VqNutC37lUGZ6j+08/yFD+Jv6l8/I87jA/U+jugAvFp06heiDtx2uzOdk
kgshkM53TldTODbAc4R9HIaTbt3IDu2G9cHTwuSwiECiIzKO/p8MEj17CzhxK0lze/23sD0KxR1I
Qh+StSakkZypUvSFBOq8cNO9eB0aImgIEW+oXejYFUyXL+zVJLYo1w7kaMiVL9u1L2yue5Pwc7OP
5DTP1Skx4u6oTkyIw2MnbKTGwgiCckup5J0wBYSuyZ5scmNkgoncCOkmyG92OBG2AeS6LNNfqlUc
f37URq5j6S8XapILT/2iPK/iZTigTjz6QWMiDTFPErQGan2fArFJVKcHM+97JBY3K9SdPzPhPpP2
WkxMkDglM/r6i35Gqd+h/D8vBWnwRFZwh0aJmwM3K21W/Xl+eEMmBIip/f3Nv+DmPmRL6eH3ZJ4P
22ztyAng2ifMuEPG1F2eOIr19ehP7dUY+sEbhebrFf+ymtqIG8PL+LQtL1Bq7MmlHhDSr8FKq5Wp
gjtlnv1FDkuSJuFUanN1VU2wZDEhuwykuTeb88gO5GBjX1f7BGXz2M+UMhWyCGskAqmSJf5dOnfb
aJmV3IH3K8U8uwnt7Ztgf2KkS/kPBRsir6zbaDpoEf9/i/KZ2994tJiJmFcpTdHjrmISv/tb9qIu
H0Jbc49KigZmbUuy6CzHIOWhwtc6PzC6TmIddrKpxih2ZqQZ5ZNSrdI2epyQuaHmNBCqOu3wwc1E
FCzPjdBtn+uocUKV9HqeGQef7TtrCMLiYFt/TRwST9D1M/DJiCIQTNZSD4Ql0hHw82b8SwrKekZd
vcM9qjjnko51aGhkr5ZRKRVt+uuxy3zO7JKEH+eGKkJCVr3YUGTRPFfVlSlFSmoZxAxY8dkAgI5+
c7yI0caawfIOI9+Sw1g/NckQ16i+decN5UFdlXeOXp0SqOJC4gEksPNKegoZqYKOMrzTdL26E5TT
1AtGh/S3/B2b5OWN5BsBo/+HDP23Xu+ZOCKdPsycAgepIXZ1KGM6tGBtDPGLNpMYwnndHqcIIK4R
MBkOiqOs0tKgXl++HQ+uLaYGT9oFgYSim32ES5cvuklyMbGs8BBsFNF5zFsetC8oUKmXfKLPDVqO
wgsEK/JL7zrv8NC9hvUDerUYIJ7WRh9rq3C4m3nyfU2UNc88fmrSPLNbPlDiN1cy/QEUHj5pvyKB
BL2dBacURhGHKCwOFQtWKB/q/cgU4Mz9kLgya6TpYtleF9P4DJnu7YbZMjCJHwpwQhpF227p+vdx
IA+xZrSchhkG3Bur4UTrxA7p1yaTLASXDvVEBWB9rJC/GMHSJLzPBy/sh1hW/zkletp1amYJwJkc
+SDjeagGl5zmx2AjCg4co4iYH957AMx0jq4mrV7yqy3GKkctcOu6rWjhFUjiEs7qxkWxAWL2QiXm
a01Ppa/bEelVLW/NQvBPAEBTsLGa/5TE9LXCYUhBo6p5hybEw2gNX5d/de+42nxFWa3sBuaPII4P
GyQaOp5IDY0E8rzfG95YTmZdOJ6leBQMAfo5eUi4GaHaS5s8WQham/bhgE2/Esy5l7+F+KmoL/c1
1ncm0bq1L3oEO9DRwTk4Snj4SMKUfvNBwz09s+CmEb9Vu6mr4uxDk4FkskGwQ2AKMYWZYfILs1L+
3asmsn2Dm5Dh2jRqY9IMPh27e8Llt7e9mez1rgeN+0crgk5PFaSeYUIHqF/qYAaTfM86NCMZ2J0h
HWsxJVWehrn+cHrS49r5TwMMSszop6DbFaQ4B4wSzUoHbuYOBU1sF0kGBSmChruXlvuWcIVvtwB6
vaHoVyvKrCbJmnYeRkT/hVpSyOZMrhgGJBz36cGL1uLeRMI25VIhUXkCGwF27tj6QMDeP2dPWfp0
GLFPu6W4X5HFBzgQ7aDclfmz/5Pr1DTLFplcpTDHfu4CN+RIx443+ALaQ2jObF3mTKCah/kZF6UK
5F6LuzkS4ZO8PwcdQVJXqRERKqTWBV2NinkFPAE/6Xjfsu7cnA7/7SPlnPIMK6Zhns71/W6K2gv9
PffrOl3jYfihenBBmaiuoltKhIFcP0/C3FQcVZIdUBG2XAv88kTHbAejF8OeE6acpnhCSrDRsBJE
Poq55MHzK4x1VRuLN432Q8o+pWKFzrs3gRY6rpP7NTy4lhy2zDEqo3Otbvrn3zbpLcVKlrtuuIpH
Is+Vf2nzIDuKGq6YHlylaNE+sdKBdayb14pH2DPQsVUzYO7K658CiDZpdH02eh3/YGHJ0tLfYgum
ywbOE713q7pq1fGfIbY/Fg+6IEa25qKJo5xPq2Hyfv0nK1+gPNCf4sQbKpoF97qJpUieIUOyPn7h
eDELcCY1NiDDiTaRqVu6WqAQL9vpK6w33L/4/fYLzhh2vbrBopu+mTUWGp252yOpz9gpOHRfM8KD
gI6N0e9XYS7YpCHTXwWZEApchIRPtkxQlXEAp2jRMRqdhH4RjEHve14mvis4matsmGeswWHgKRo5
Wzwe7j92/j4FgvpOmTLTYfPVpgtxdEBmDdQe53oP3Naw3rmtiwDJixQpboOOk+vfAzOWs3gHQp0t
YsUXpIHC7SFLKBzX+nhy7ikg+I5VazjitTlvNaPmgeojlJRlNylAh48ao2JIWIGjAIgXBrYjc0m4
23f/y6/q2paWbQMTC7TRzKGNIYGueA69IkZ27qDCILx4EVwW9mQLsEIA3ffBofFR9xQTUor7ZUYA
2LmwDQAyRubViVjq6WGg7gpu1cHtx7eeUQgyrpsS9znbDMIa3ghuOKwrqaadjL5LpPe04TE9xMjI
0Q7RT8YMtCCbeqzEgse18Fr3QPOARxcPXpXcRJkfVNFGn+96k38y3Ywxwa9gTnezVzMA5wDxsfqJ
FyArVXjgqotGEJ8IzNymL1Lk2Nf/UvtvgXMQLJmGbqGaHwTl9w+Fm9duVELEAyrroT2IhNBN4nLT
IrQuwmdy8YzHuzibErsQQRsTXpBvAG6ygZ3iO3rTuM99cfHjjfFjmMmHIFc2Bs10+kT8qJ3W23w6
9fLekd4RPzq65HVJhm2GwhZPdAZtAnbW+GppFny8Jc/jrTkJEX2togOyMIzY0o5gPXjA9di/ZZox
cInJbgVkObVj7Icrg3dka/2a08JsBP0TwMf4MpW0yaDCnJV6Y4CMNmkLY4nu6xi6+rnhXY1U1PxZ
+FBFAXCPhjF8driCB9JUW42ORT0Gi8vrdis0VTdQw/j7qm59HNX8CR3tfnLbxVJm4Vq/FGw/Tm+r
FyJuejkKH8JRpDZj/1IhVkTF1Gv5kgpiRaqYaazKK4/zv3Zg31t85a3/MSoTq/NO07yDU6qPXR79
Bv7yjsm4NJ94hHAiVpnOK1YKMDljxdaxK/Wgb9B2SG/X35Hg+1z3t4XorfvqThmtCK4C27PWu/t8
Rz/Z4N2pl2BtCJtySDn0JhadAAMG3pTus/DdKKS4zif/wPYxdnKq3m0QfFDPjpS4EkchQJlBPfMg
UgoEKuLNPs6sbWxelDb8KsC7Tolh5fKzoiA5uFzx/xaObSsKdEOQsmcbkmdOqdOB5D7hA71kmTPe
u0OmrW0unTRnA5EX3VhHDYalsuYdoHKg9mvaBsZU90ox5n2s48CDvbGV1pA2DtYpmQxzDas9sjx4
IurMIJb7ndDMUt/enU7m0+nKFMUEKSmAJX2OCubSwxA3RqrIIGtASBl31sVkkZDizRzl0kIim7D6
2tkb7ln3i4MmTLwqr9Cjw0H6kW4KaE78aX2D8ErTDU3sNq7OiE350DOw94hCxhPtj6OHUP0iTx+9
gUAtc7W0ulssdMlEE09nYmG/E6p/ukI9KQgv6XsGTcrSFbodF/0KZhpMHarHAzZKOTL4wa6G8NtF
jTf3AAXQyg9Ao5/13J5aUWYP3gP7MMtvVO5crX98NWMNeO8bYUE2Fvvrsczv6pYTyQze0/zrp+kI
Bcp+rajVqmnmrab4ZC069xYzTjjUdW6xjt8VNRSdYZMWGhiTuhlcT8dCE8ztonuiQzUjVRlHp943
3VbdjjiT8gb9mMqNflwLPMiSYKCb8G9YoyBZV75yvP/I38gfBjjBuuXythCcCgmaOaSTsliSzWiL
pNzRkr+87JGoWi6jyBlOL7lxqZuQVZi2t6Y00NhTL4ECoyBshYwX/1QatYUUtfjzPiNG/bWIRS/3
25EM6S8C9tY6E12zPt9liCqp+LWFfLdjAhJMkGnuibKu5bQHftHMr10kGlAHGA+Qt1xGxbv8400K
8q/y28+m705EgBcWnG2otyrLKBll8CATvYP0a+HCBVeBdIzre1o919tTK+vUvnopbEqGF8tHhriz
0d2an1iAzhwyePtQmLt6hpu7JWGkgwZYAy2Q6AAS62P9a89uaNSM8TiynuaA6hqrRM1cMmAIwiq+
CtDV9mgY5RO0hAX46idUyHRPG3gou+680pvMHPOOxLVls/uqM/piZ8QY0h5dfLZoUeH98vuEaJ3W
oS63kTx1zYKdX5xDj2nsAHjVNQI35CdR2JcE4hm/7823TXXZ8iGEI+iTPN95pzuRRgm4vzrSp77D
uOdRDpEiNNVp3VjbEuQiTRXmBrvcuXvTB2x20maCYaxQeEVDrR0YLEEM64m/jkTe9thjuRNGdOsF
3Pq/3MZF1Dbclm7VxopmYVOKqJQgc3I/DR+dTKD4yhcZZBQtWMrY3+qQMA2v2GbnqW5/DvZAfrim
/8lK4k8K5Ug6EQv8HEAF2ZPAEJ1s7XaI1J1unLMnrtHXz4cfOxUf6EF6f1qcCnFPDR+5pcbzv+/P
/E/yQui/6sdZn6we/JAhSYCHiLjpwqRSX8cqMwgvx7XhwRqPgdpVe3/TUNJ6TOlNgRQpm+/sJDr0
f8A1bjEwZqZzvUZSv2Dk1DQS3d9fYrCO/OVRR9Hu3OA9A7nFgdVYcfKOJxMaFyy2p7vvlljWfzpg
v0qvWX2ZfLBsZxXoUCyuXcRVtd7NYALeyTb0hu0Up7chAkpcY2Rj6/N8RIaAbfwJcBVqLo+kwVXG
syeN8iiPd/ghuuTaBh9fdQiXsyDhNyuo1OZ43U7DCMofB84sWRQsW3+7KKwp271nkPsisunyWlh2
7WFn71xGMECGXVbpBUGkQ9T2G6RqI+cn7DsKHI0y0ILiAAAstQeqy61Om5gyRu2t7OiYx2Es8zDW
OSKTlKc5Z7WiMeWo5diHxfKOPlQCeUdBAHk7YJ8ADS1i2le9Euo086XfS6ndT9HZbNe8sLfyyQ92
Wmxyi0TtS3fsSegT81rQskaD9rEfPjhJMcDsOF5z1jC/264rw24S0YKge5hLP0c+XNFm7xCR7QIw
9Ito4w/41et34Bxw/QXiB49Eoeo8yv3uBidqmneZ91e5VPOWrp6g3g8RCKxl9kn6UsATBsCmK9fr
Jihmwrd/ycNwlDr3AO/aRknbZNYWK3QT+rPykh8si/k7TlC1hnp2WuOIYM3L0/ci22XK3avYCkoQ
LvGF6P+lCmegRbCIq5nI1yqAbtpSAyRrIQJtMyUTGZxdNJyWgQVg184VpXc36pUdkBa6zAlJGsEt
bA6x0PTGUo7CPPx71LyO9tHngMMjm6Ajn5bERa/xlTtnkj/Q6KNMdlBgav40ASBTBt66u64RxsqI
83/2Kq2ejgGsAacvFqFwXwLmZldTFbCcfoElgmG7YpErUQ9H8y+vMA3Drr0CXsD+cOPu5W81M9cc
M34y6f245h2UdEnh6L22cvCSMWCnaCtt/JspIxBu4urUwrn2LtsDejXUasXdi9yy0s402/TbDA0j
IG/9wxGI35JCT4RYHnw5sHNdd5MlMNqsst2jRQSTtk1DH8odZFocWQigYd57CWIloOVLHuFZnuY2
9AEo3xECctEv/BKXoDrMQL2Ym8GtRI+V2DPaykb9MZgD/D6acuYFUN9XUOaP/jdLl8iOGCR3hinj
7K27NwmBBdJI3l4qL5xVPB6PccMdacTu0OI/9/C13Ia1zbF5fLPu5mbkB4A0C4Ety4vR5Qm7Xcoa
Ih2E+eP9uJtTCyFXmEjHcyulIqs1/W+Vp0UUxCjSvfUo6SCFEcv+2MCU6pEH5+pY9zau020XcLQ0
NSjHsAn6vZLIBpba6IYF8Kp0dAraW1VJePk6J4104F7JFvp5JwIOzBxIZYIX/FDg6dP6Y76mp5hh
MJCJ5tH84pbpkvdUifHDYWFmq0+WA2pjYn8oQ+tEKAG90Tu1SqC7XhzMDuJr8br91l4EHAG8NHXO
9MFUTLNg+W3VglxOxkaSA9k4+Dvgu2I98fyF7pZBBp8CLN/mZABm8ilCnQN9rhXN/Uqv2sdXGH6J
pP3QfYKP+1XuxfcZmgjaghKq0LCveMX6WCeceNV8PgwxlYHGpFRo8W9LBiNazbHQecPODQV/OpMs
CFmow3CFQG8kuIJOMsO4P7petZAXy1O1Qy/iee/xXBAFrA83vE04wl6lSpQsgoW6GIgWwA+rlgI2
90GcLl/769ZYswWNoh/cv4Z38A+bl/YntU8m4mSCFAYP1banj5ecFkm+RwM2ZmVXXislwAgZWuUX
E7VtEqsHnxvh6wNMUsSQcn8xHri7Wn50zbkSXRFKHM8lbY7g1evx0Z/Cvz/qY22XAaWAqHtoI2U6
Lzf4dhk1CFn6STFqpTudf4IVSAytdomAqzrXu/yzioix1esx4wTcszQqjywUteOrRUyDQpwQ3CUt
UzvZMOBFMXNvGq1joeXzKmXEclSXwo3j40F8KwMIiYYGNn6ipCLYj6m84m0NMKjj48OAzUjiaRB2
aDFhX0zJkf7aY6bJ5muZclYRaEaa8sbHet42AwkuaKTHwp4Sf7OplB2c70afqdeSUlH/Y/STvf79
8oZjxcHrnQvKcWoE1tBzw7Part272+FFQ+BLhLy8F9jjYbfm7rCHZzzpm+qYn2NKsXEsXlOxQjk6
22Owyk1NYgf0e094n7lfMbR0xqVUmlyE/UaQ5/QTesjZGhpkWcX8HjKIo3TqxR+e+YPsFHQC71yD
gSkXKBxD38eT3K9Jjy7SWs2N1dafJJyQMRj6wOuKT5Csvg1pR7C+B3cANLNKD6Pvybky7CyO+jq6
cEXBlK+O/K9qXYadEcOy54JdeGdXEh5312TEu5teHrSkpXDayoHahGHrWndenAaY10pTrbl5rfLt
PG6DK9Hx6nkaRFy7yvkB04X6LcboktNMnLofpYhqpaADl/pq3Fpl2RwItZM3h9UWEn32YuX+CNGJ
CLdgJoDptAgbnw2Zsq4cNhggXiDsMNYMjbTqSvJw+P9FdZ1aGH8e1Ye9jPzhyLON7OUMBdpsRRgH
ccIgmznLQcCr995sTDDsBi8/4DRV3fETAX8u5Nwk1pyQmMSuX1zm2VnPo3UmNSDbSZfL2QJhv0oc
hIN39KaN/u8UlF+gLbbsqHimOUdiuY77afbz+rA3qymKtNgRvU49fib2EB/Rjucyj1wrtxdMmCc4
GGlOdQLvCIp4mWLGKGeSHM/KrpWyju8TCc51mFmCf7KJ/DdTeYzkM2ht9f951NjsBjn2u6C99uBC
xsKbl2T9hsEvB8rZKRY75ArHZTnYIig2tj95U0xWQQ8lrZKZ5mWd3jxMySJJtDKr277fQa9ZXUSx
77lT5Cs3OAXlfPi4y5AArRtfTzslU4HYi84isy8Ij84crsW1qEawoav+xQKLCyy3zOACNgMx9C4r
rn7AYegPusQzknKvBCF4w9NHubmLBoTuFmPn66BMbjK5tO8ISi6ugvwGayaeFRF49Z+kpmtF7GUM
DyZ5EY5J+DBucp0e3HTa3X60gUjMueXSVe0fU8myBxe3Ynjv+f3HuI94LSbFUNcBcHFIYCdM06+D
niRecl/PFT5A8QcMtfQuUwSB2y3Hq0YNUCUksdaGrUciT8FYe3m8UeG/N81HPQCalOGGpHOLzcwq
0g74nm1e8apqAbV1azzj6V100kWqQmVjkOuLgEdOPARV5SjfvObLV0P6HaOXPdvvO+1Ggo6rIoBm
411HcrCGfzt/NA2mvYi60bvkG6Moy+9n1F9X/ccLtiDhk363pDZea2DA2p1WGEBE5wQoIHfHGAZW
bIj/+B0yt7H9uhOgsKiTXUcP0sEo/trDM4N0FYE0Cghh7jvmKUqonbJlGLFMV+h6/Z9mkmUegFv4
sjyPIRf1CRfhuAm0e6GC9UEaVnLETRTZhpfoKAyCU1NwMd1tsE3O53AcMyJX0YYRArC9z/cfoypH
9XG/vA1joCAohc2Qw219qn4/eV2VFJHRMBq6QrTB5kDaRqj4HBzouFPH1myFZwhO92ELitmXn7L4
iaMdbrbFK0uDvunHG9R/btbMbpPEAOF3SMVzjfjIGzaK7igabuu3onJfzSnPfwu3LJb/DbnsW4Nq
WEaUdcUI42kuHZUjiCzKPYfIrrKevg5JYq27QlOJRVw3w4v2FYVXj2/WyGR44LAlVcqOiIOQFlTc
sbVEIW1svXSmKwYRHClZKhijPHmNsl/R+4UwNv2onNYksHEptS26G24QrReNLWtlr6cZLGWbVxc4
qKPJ4bcjWiuOmWcQR30j3Ec0qg4M8CXbTlm3110U1Z+oNPDa+F6z8qdPt26lPIfJmhXJJ3/Cp0go
D5LCOFzpRllz7AthAuYHQI3L40qQ08LC2A3C/80sI9NSsHHTMKm2QlyZJIjb7oOKAinZhjuqMwjU
lkZTd8nB3pwBWYwmVRSmgZwr0Udg84vrJ5VF55p7ghIS/6IfrhW33hq/r+GM6MxToMB4CwqTBTS3
SORmBmnMsbgRzWcg5fuz//Mag829waO6qrvEg0Fc/LLe9duM47Ar12auB33VNiR2J75LuAYtFp3P
rqwyO8Nhl4Vtu2/lt7eSQ6GPS7Agtrg/icBe5UBj2JCuaYiTimr7T3NgqSjx6lL3VPyEbgcUppDI
zTkUrUrzPUN5ScEJ4W2ClO2XkISvN59THbDcZgYgfWGE3vblNI8sCU5p3pw4I5ab+/zq8SRuH5TO
O8gvGhrYHwq760Cczt5oDqkGApcoZ3Ws/dH+XLF1dX6FMgFWci7FjYDebDVOxCw4JKSgXZ7Jpinm
HzYLDnOQQ2V8+y15I8SBhbCfpJGH3xB5EdJv9uJVUmmtYmCT+BceWuVkCu2QVfJFhPRM0T8hLIzi
Hv4yIUuig7QV8CPnPSa7UuGPZ/YvlYrDwXN8ERROKo1tUtzh7HDJn+5CApdkQR/2CoKKC7nPNpb1
WUcZyoSSm71AWsw7XrHIjHnTmAa9seNdVFPCoXJZWpupJ9tmlx+/JXYqXluFfWmUlUHMRyb17ZPU
jBWP/di500LofHr5jlUkJIoAHoAObWZlMvT4BYAJpou7VGLMP4dW3wgP/EJLlh767RBRc+J/s4RO
bY8SS6lFI65laE0f9NzrfRqftW95TSUVpdsm4Hq/jM5fTR2cgXhBPsxRWmg9HCSyT6oNAjBlPxMU
kwnn9cIEnossrbSw5Qns1ND0trA+HAfiEwkeBZnYMS7bFS4q1EJ4JrzxiWqpqFu0kccp1LrBOws7
QaYDHUn8yIi7YFDFbPi3qIHuj2nVSuBflWJSyQBUMwCRAMwOC5mD0LD64xT1PfyoHCbHrnW5OmL4
wYCEHWj9UbgSvEyDTP7fA9mvcUn1evNt8+XY7qIL6gSzD9Z9+hbgskFcGIgJkS4xV8j4WdjYOPKd
cXsuqtNRroULLh9ZRMBARdLg51UdNUwZwbjArgAsMO1T5ttCCgti/YCMcC+cnarsNN4+oAsJ/9I7
tQzXA6WfabL8+cI+iegk6vRBj/AlM0wcQ3zOCcbZ2go114yD9pw8Em9DM+xeTzmYNKtcO23i8WEH
8ArnV47qwopNgCiseC4EL8I+6GKqCgQQnBGgEL38oEwEGfBiGH3V5adpbixLaE9yLdFnCtAeA2/o
EL5APXkCdV4nimOVZS7vRS9RD3ANHDEgAA5wsXgRXZggujy+Dyz5heSe3P3FviS6KMxgLnQABhWP
1O6n5E3EQELFFucdWDw6e2cWr/RQftocFW9/tAizUwRaSJWU+hanS1/N8sxbsSGCOJx81GilGJnW
sFt0bMdSaDL6+3ADl7qSeVozqsfl5esEjMabgqxkX3MnsAPMk9hRfdEYjOieSo03svdzzvSFwpKv
bU8BgCRFP7EYqoSHF1dnbu2XysRwwHz9NOPwmCOlqC+P/Sudr0LjzvUOyDgqZ5k4sZMiDPdRWqJC
4O2VL/UatDVRGz8cYsjb545mcy024fE8HGFYEdPWXMdQUvsvVW4C+G00c0AfDB2FccjfeOTpY1VW
geadcuCBvoAX1SCeo2lM91zXdzBrQUCQNrYqPvwPglYqWod+c8NSyJDO6pvxgTZDbEJZgyG6s765
atlOPO75wC2ZTZxdC7IWE7DEUaS0BXWKywGdNQDnGhuwEwi9KqFqLCsJrCjVO+Aica3JyLZcSsz2
UoaU9Z8Bu5VA5jRo0O9RTLuxbtdRiyzIeTPRP0p/SFg7r9w47gHUV6xSCzASp6ky8p1kB1sYU+Nu
Q3ZwZVI7pMPmZWJA/tPu0XUOy/WlsfyhTcBorwTMoBuANLFYF7If0Wry2kI1qC70Rr2lCS1mffi9
olZWAV52UkaH3dW/DZvxYZp8VHZifzRJjzBU0smHTVv9Rki5ADKfPPqWjZyivUZ2z40Iv7X+SFNp
4nfCUrnyVlAZUCyHd3E1q+LdwHjBftBi1YJ6FKMnc6EnlMxHwlN48PF+ObcN/oo8H3qqaOVI/+x3
MMQaGAKvI55Ke13mT/qId7wBVqiczQADfdZXrJQ2AhYJyGkAjIKtNIL+ZH0V9jvpfL/+XPNRS4UQ
mn/uSBauD1JyyJJO+m/jPkWpI404ZAR4LBz/IOOR1gVfUH+eYlXwmt9tOnlKMk+qdZqeZIkBmE15
Z7K+oBb8g8sFe4gUTPPGPZFZbQdQQ/Ixr59C8uGToD9vCH5+eumyvQAqQmvAKLrL8NDGWNKvuYHe
L6YmIDE9Nrgmlu73oCN6v8c04NFMUEurkXuh3VCtOxndqrAK5LESO2MzQEXPtkbH8KPoyKPdxuBa
NLfKDrldB8TSlVwhJs7JSCr63KKkBeRmoOMXzBtpzp/me7X3gLxDsh5vlji7GSRnLCYRGxHqeSbx
4EKRuZ1CEu8YYUW/AOfiL+cW8JwHru6M8uxO1sxODXSFMi4qd4zq++5C3pcJasWYZIC2VozZGqdy
V47WQkQnXrKJUlTGUbtfmT/AvzGwzCOU2uMFPXKOHP2QkfXkJqEsu84kPMusedl7hsnvj1qH5kXF
izaP1uDYF+k9s+oPxZYkpUwBsce7USk8EO3+EFqrdkTKVVXq6etlmGhjJegdpob2crmkIweK069t
1J5RwUbcGo5DxfKOULf0AYCdEl548RE1BEKOyj94utbeN1peAWWS5pofo/PSfIeguXoseMP36oPV
CmDYoc/upMGWkH/fPWxOnH6grmBIo44Y89uaHHsFng7do+upqUbfPxHGz3P1jLt2ZD7ppgoriMpa
F3JxswyNPaT2vy4KI3ygU/cKrVaJGUQJKbYCzUW7WOpnlL706p5ZdKqBaFxnrjBmukpfzyasEe1N
1Nr4Ew/78ZDY0/6bSMcCKM5itI4zOAnNgB+gzsXwKV1YbbKk6i8i7q0tj0so9Ljf4GrJgOqeD0dx
gX/gVnYje9cr7L+9UDmqHhp3RhoELuFtihr2G+j41Vl78kYc8BPPd1X6x4TYWbhDAJLxCAYtIeEC
+rtUhr6D3uoF7bfsRb82f9XRGUgnysq2HgvCHKQYGrs6ePsd97J/xXwMPNs4nCKkqaY5y5sWKWZw
IdBmB+0n7Ti2wrk0ekls9NPpcms8KrgypQemEEND+vbRqFej+6I1dC5/L+06uEyEQjuKNuZcaXpt
TYoE3fbawBEoO42SbVS7NnV/F+OP6Vg1J6Y8WlyaGCldVL9I4QauRimN+FmBd1S/IesxO+fBloWy
xG5tIR75mpESPyXphye54oDzzrs0aor+lb18xfiuPxY3jzpShq8ZDHmHENJ9r/6ZeVUUZMVBhxt1
6hvD1Bh9rPg6n9PKEvZbpl8ofw4Q3MJG8QPTiawBCfBgDZLqzwJK34R4IT3ZAWlop6OtCpmxDJtO
kwMIGShF0cKlj8i+y3vgCyJiNR+6poFhPSdC/QCSstsYvrbOoafzxK8RxfXvDGdCvZGcwAngEtTt
Uwljfx3bmWyuX3ArExfT22Ne0NMgturXIa2xzK9/G9hQtp+8ZOx/gHZ7cLftjs1jAZAWJgqQhdD0
mahzXyRxqXhGv++WKRiGrc5i1bctts8eg0iX0ZgujLWUmKtpKVqi3xQvtJJ4g/RFQNMUG1xN92ZD
vrb6IWxHIYwngh3JQfHlJJeXm2Um6Yc9RXkrO/qjLQP/I1bEQeeCFR49vGoaMS/a1uZ+5uouyQwX
o5BAkpHUDqxSrLfG6zuDrvhTXLXW4/ZGeq+NjGfENmndZHPDsRqUVz4WULa2xVgitGVSG9HXvHtK
hulUcW7myA2gUdpYkWcDtePHrz/Yo8ChFBE8p0dtqwYFSjZN0uWaDNXLr8HbFMCMzFpaIvg72/++
5FT07DM5gAFXnWYYCddKDp4XPtznjF/QYi2qNX2GY1Vw0YN4f3MdeHweHb5RKtAIPwv8+39n/vvQ
IV4CX1Ju1Dk5Xb4Mpxi/vJgZ3MWjH2UmhxFr7o+qINuZbt9sbjp5eG6wBDSWzY3qE4Dhvx1eWpra
oTisNOcDzGZGXyn2RkYB12GmunVfSg9YugGflpBzk9pISQfie0pvmGM3MM0kEfw8lQ5ws09FpXHm
/6EfxU950wetVvqV8VQkuyob6mxJTyC0bYWq1ID8DH8sIHV88Rz2TcRQSTQfd8kKQKaWwWJVwh6T
m2dgVWTPOuJNEd0xFvBPk88E/D514ylTq8/y7VTHNIX5mpUGul0SKa8118oTU9DUPdeFvdyOVVsw
zk1kl2Y2GMLYjFkvvjUjxFDJqhu+MjWQ8yqDYIqK8jR9ssOtLE7Kz0k8BnXdtS0ojDtyXxAjwjX6
y3i8cN7tiKqlo4BzOUsArKN8zzge4tZGtaIU4C7Yi7ElAZSvu+4xb3VyiZruDNQWEw0A84dDTFhq
Lu4CcAtGpycpv1qxzvmp5hJQddtSlftu6EF2ySmbOnPMWAdh9PxnasuB7QCVd1KQWXij7a3O/QwH
17fvuaCOO25+fDhHfw5k2+2tHE5Xk3IJh5pm2/sZLQ4XG1suy64bihtdMLQTEYC47E9Wh9He4KJK
gvfuqM6h4yN8uwFFcWHsB2X/QKEIQ05vAD0AhDX9d8LMOVz8UJ/4lj8tU7mek+30fXIygsyRy1V/
Son6LWA2/NdbixlZNRFku8AUKVyrl6GmqUfSaOh4iNGRnLfkCnMLfjaugU42l0FCJtIcbXETG3XK
DpSfkrQXkxsEfxh7LDdOqfgC7dka46Rb4V78WzSXD1DCoUrPtwQ2SIrJRxLOZjIKXgmRYGH5ilcb
+ui9HjJ0IrCohVIlAgKeSziFtjUaE+WiPsZKEuqcysokzsfDDJ48YUiqPYoVgJiReIK149ub/fpI
V9V7C2xNFeOylqfwwNJomtlo9A1/V7ZYHFxmL3vDnMoO0XpKGm8nohQZUXtj3EdToBmPQQgwlsdt
Jfi28GUWPpck8jMeK1U9kP+Txn+J5UgNvHC2cCAVFA4kGg05bV0ywixUTm7p+aWipFEGiPIhuXwS
+fuGTPtxkgmqNCI2Hz5IXAP4v/ot3hiRXieJgUC9PF51HvMuizb2AFARTtVpQQ8Zau0TSLYsin0e
FiYjGcNluAIadJzlbzUk6m1O0rtE9dnF9ljSmpYkx25wPiPWkdmf9qFDdXc7dTZ4LBvn7zAosNYn
8PTzDoLOvoLET0OAfnahfNZPwIBl8A3EViNP01A5UHLZJONCSxQCFh5jJz+yQznAKMZOFQQf3MXq
/tZvZ8l7igNEGlp/YPe5gF2kXK7SdcHuvKo53hAd61XD5v3OTDXhVPeq6xSEK9nxdh/B07HCaJtk
n5XMwOeOLOdj/NS/Rb9gUDUCJqA3r15BH0o3kcRM5QxAdjRld2fJaHaHBT0HIr43Ooko72diPGaF
hOkglD2mUcqYyb1w0BJrGecGUMlSsQvy8VjgDMgIEl/9X4QRYPhkB8MMcYJbtTfMGVqe2n4RquTy
KL3Awkx7xth4ub9HfI225jag8d6yRSciPWub2nzL4qizcu2lFC40CImlTBFLZzToMAXLOOi2DSSZ
lOM9a8GjhDBTh7PpNO4XereI9qdwIe8fyKNDszYXpiefq0YBuLPEowPUNV/RAj3u5kzOYivQLYsn
LJQE91fHbnd0/TMJBJliuvBNP5PEwuQvXn7OkaYRfwiF2Q9Xbd0M2jJJ3eyQaJgHMLZoF53yTyW/
4Sa+kVmSuB0Q7C9Kca2KjZA17lgRyodgl9jcEm1l6aNop8G1i9ZpNTuPbk0lRWG7Rdi4nLBCJG55
y+kLysd1FQDf00TMV5b7uRQ/IS54yCcZznBm+OAsRfomcF6oYJsjk0tbJzLNDYWOtAUnRJFWjluc
gRan0Q6gMRJuzAhp59KXA46ZwUVT5/ql+duIXNEkLn5ExYWn5aQ9avgxVrqNBVKt+fTMomXzd8nj
bZhrk2gj2w99tV5RggbOuz7aZvHWo3c+Rf2NOoyr6hb1nXVjH030EBITDU4szAuutqJrmFZu1TPF
4lCuTTWNCf7Jldhs5fHpb/fgTZNm2jsGuIIAWzTvCiHJf9U4JT6SPCFGKNRBddQeRNr95XiptouE
tcwg4dtdU0zH5DJ5gjATlBYnocoTAxnDfnzb6LD7RQVRI1e/Fyvl7eXE+ee3AbMk07STodh/tzm7
xiBWyri8B8gZqZCVCo3xDojbQOXAjPIgLE44uJHjr55n48hxOXPM+3UrOw1zIylY5gOeI0oQkGoN
aTAyT/Ed4CkZfiMKeFAZh7Qhh+fjFre1Z1NHt3SUx+cpNND326yiKE5Oz5B32KPFzGuNyTfbFbAk
xkxuMwdnjYGer9/OwvpJrSMN1RiTeSU0EUvflUFa9XL7nQtmYw+hi6nH1TFdszLHMZm0EMvWQNIj
VqJqiY2wM0nv+dkVijsaumiwxJoCDFmf+aP3bUg3Es57GzBCPuyrdSkMDUiAoSn/83jjIlatM28x
cdPKJiMKUiJUGjiS+OjDwxJFj4g0Zqw9bvjr0Iy6z4jQDKygJFpjlFFPXROUMF4hiZMbuxmEhF6m
I+xKbr6jbANfI7FofEaIzxS2x/4rhVzAFxi9ErmSk5IbJ9SVxfFsR6+5Rn0D77tAwobcA2tYjWwd
yROU/hCicRRAQ1Jz6vmjNCAdiyxUgE8I/fbWbvEiyPNFogJYL7nR/+7i2IQY4NP9HTFuo7aNwH7N
SRTX5VPPoGlCjSIk95IRISU3FUXDJXVV97iCBPW1HtDmjDym3pv8Xa3hADZYmuNAc67BqnFHuENX
IS4Ny6hD7fYpMyqoTBfc1N+6FW/7mqmOLXnHHdO433OwenOLJeZHTPcnEwwrvzmat/fQE7xL6nz/
4lpqb9k/0OWQvUhXYEadWsaRsJKrrv/WBVVr/W28Nf8gfaGyn9GQ1ILYrfcrlNlVx+JGodWU71q+
goSX/LOoJA30qGPat8x3/D2kjQCgceScbZX7rlZmXoKSs8kvqTnRYn1mqz5z9MGybfw8xsnst6rl
t5tHLyi2e89nJOdfi1xXKLhjtz/7uwzSqcR0H/42vsTW1HMaYtXLkXQ+NaCDKTazIG4XBEkiW1EY
AuWPBgg52CnCqdEvJwCetid9lUPcn6PUsUUvvu1I3AePbW9D5ZQkfoRxexJhTFwEaQeCi4q354e2
KCU6yla8oslqip3705qnbWMsmq8WjlrlDxsul1ddgxvKTmTbgMPEexmxwZLzhabA28Gsh2xoukP2
0sUazvo56QPoU1jWIi2PJ7sF98mMHQINau7Gp8LflU8+KfYSJz9ZxUarhxfrtnT3l+rj4zpfkpqi
LGr3VL2OC+r9QOqFaUZy5xk3+BiOBcWCnxwJQ8yVHxqeoK3cRak3UtYeDhQWTC4f2mNxbpbH05tN
fgeE2OG5V6Bso/me1yYntCcisg6jRV1m7G7BmepNbicQLLkVV+VrPriA15oqL8Jzi7RqTFpTK0XQ
jHWJffuxP5uTBEVKxItNJ1TIGyt/czNLHYHoCXXGrQ+3900sHQwSjst3+oucfa+7NIfiUKHNIlJ+
Wuy4NAuowiwAjZKksjz1OAR0u4UtujsqA7KsF0QMEFBY58tQZb1I+CWaX7QuFmJ46mZAARByuVHF
PMHbRGgPbY/FdkZPtgU+FdYeuohB8MmOerapAaTqsLXqBZDGnYjWpe20T9fYdPV3mwGl5PlRyH9T
JegoiRnBdeGbr99zJLNca95f3s6aEbljTcweieo//b2LD73LzbrXI3miQmLZVaFL2WvezrkZ18QM
dCl/cYNikp4XyOlc9RCtDccPK06Ctw8/IXJKWPJ5Xb4oLoX0HRM3ANSAr3/dCUeDu9HKbPYnbY/D
xB7hyBUTT+jbv3jZXY5ysIqwvkhcYZFlbBkkkrTSGMYBOjMmEEJTGkWrdaLLkQqdXmkQfKi2ePTV
JynWIuoSuhQocaKdQI6fotj87wlU3m/1nUkrTXDP/+YqJ2RLh/IrPyFxxwtq4tEWk6gex3oig2Pf
XbDdgJyJi1Jx8OBI9Sm7CFMrk6dOq548C+X6u7oIkwLG72LGiIIQZDd5XN25bZpYDLTWI3meNT/4
d+IxEexLLLCk7MIbgpAiXfzBOcEP6Bs/SU50bqdozQv+6zV1a8ZXMj8GcJDmnAVItQ6d68fp/Rjs
NEaXrQXJoQB6wggY/iEz0jhdQtIMwxkkZAAF5a3ZiQ/apYZWknnZ6+j5cF0B7rTylLHcN1GswjHc
3lTZNG3yorUP2b1xYbGQ0Py4dTWZsmxc68F5eyjm95oppIQvZG2KPojbKaCJGLfp67sTBNbDrKVp
h02I9f0C8YD4VTk9CrV3aspX/phn7w2GiUcnerRGpUbDOpWj1asrzZ1Sypu3MltUKM1CdwZkQJXY
Sx8+OiJvAc1d6/yh7f43/hliDCA37Rp6A8VBF8Uuf0fXozWRVEzaqkPmW46zh+Jnhv8bOd7HN/bg
EFBb6qkXLjWGm5NBKVK9FQGV/DPFgyrLN9j6CUnj3MS6+DLzzYFiXlnSwEg51dWzQrMgZx/aU7w+
XqjfimS6p0TUPlHRx14438xcYB8u0tOtbIDQ75XhnzEC7fhbo8IiAiDJuuNXosGXvLp7uoPouy+7
RxVsUxdB7QmV3xTUcSCWLUGPOgw7dSUp4bK5Ys53dQHqjjf3rHpPGDAUX6lC1icy/ZN7tU2Jnrz3
iou67mvZimUeR7QjoDRI+X9F0P4LsgJtp+wjral/h+RgvfhZht0A1/SVR6IqBhjbO8i2wpDmUbyz
uJr+1CDFd2+xQRlIgioc9bG2UF+TAoqoVh42n7yvsN4qU4BbK4SQJl184SQBX2zv6u+RozM4y5zN
Nx7HItRIH3I1gvPAVV5BvQPSCioHEjRuMF9wyW2cyUM204qHgOKTlVi/2r3BmZbW483k1qgrybpM
m/MrnciAwCXw62EfREHcntDUnuL/SH72vjkcLWSfRIKm3ytDw5sBMt2i3tvRi79Zv9Tx+B7pngK0
BXELGov6P0SZoXJSW8F8VrFZMV76u2Ewz4qyCVgxQ9FISf+E3dEDXBy650JfpaprydTSFSp0HpHP
dn9LGXDi/8DErd2BL1VhSGUQ42YqX8SiImETSsVeRGSQhky3lI3IISLaOKrQW68f7HHYR7UtD111
wFpoo3MkRpEufuShVBlH21zNY31OAgaBxpIhAWj9O4JnGXv2kUfYZcLs7KHIoZKULzy66greDusb
VMOyq+H1DGV20LWQXDZuaiS5iwqLisqn6cNPpKj4BU15CIA5+kaIkZZOkiwvsKmZUsSAjQKHYYff
LS5Eu9bL+R+Quof34KLCWavl5Lig1yl9cURAay/7fY8MPbipyuN17HX43ry/s7nADqO4T6A+vbrO
CFBKIFJ+2jvWZbydIFzqldw3IkLZcsQ3Ly69O7/uwhUf0UnkyPfmFOh7jNEEtZpmRf3tcua9yw6+
sPCnRH3m7sFpl+BjCWiAgNP0kgx7P8qbp1NdjI7XD7760SfeSy9Euum70Bja06ipImWMe67irRgZ
UPC76byFwQI8DluzxiCrTthX8OTtS3KjuoaP8SsYI4tNCJe9ry3/EfZmMCmaP21jhlr8hGB3ZBhI
PrlIaofIt029Jf/gz7ZAygOfsrofaPIhoThc4+9xh4RXBOIFnqHnMbdTRDqkYLtzqvdEoi+rcKcL
HEWJp6ErETAdD+oaMiOvqH10SYYWF8tOJwjX7DwCpPygbYF5dl0KSO9l6Ll3UxpciqQOqrfvOEQs
XPUXutnFfqF8lHgJEeVnP36Iie5YwrBdr4Fs6owGEhCHhBMnmcHYp55AtlXb6iIBLsjVwH/Dsxxy
X2bvZ+nNZ8s8fX4k/FMCKqjbF3CO/ut29UGkDCz9qLKVjvHtdtAvjRrxcmQms/BDfAfEMWIBezd1
ox8bAeJdn+GbL5IaxBimwSu0uJAnRmOa8FZ+TgyjL7yUGC6GdXswV64aL1zaBLhLsENTnnNwdQ1w
TxRH3Sa9DZhIcGglpUPFKQUxGzFY++LwMWPID/crQx2gGJRJdLF+hNCbUORq2lmOAoR5ZSiHZN+z
/Vx7nGxwnHtsQzYON+jUTkMQJhn/wyoKUqzOj1TDJkD2hz7a/Px+FkXiPttL2vlH25/kPx/ICaMh
D4A90F+1cFJ83xkY9PiAlJ9IgUzyXAhZcVohRlTNxe/UXZ4HPQpekJ3LIcyeDpm/Ud8k0+bUV6t3
/zGk2fz0XklkMZgajMQ2nhtODbjLuccpdXnyFtV1dKK6pXnoWOPguVlMWjDZkhm4jg+qnGBI0BXJ
UqM3xZXOFq5kdHFzr9TCh/r6qFNaYfRvCyR0atptIQlkDjAjqRif+WyU2GqLvKDmY6z08e3U/kil
W2a/fdL0/9KHF9Ni4ZYMMVaLPO5KxezCdheKk6AgYoKcaE8xP2vdvTBFTjj9OR0Y213eL/XQV7Ob
4+tyLT1sxmVXHNplMTMRzHM6jnS8Qs1K4w77cDCgvZhTNkL2yNPFbUrcjCy760pfdJl+jGadSIS9
51Ed13SCeFyvb/13L/I2FMqxzWZk3srvf0mY7FiOYnJ96c/4E1pEJZb6ByUQySJzkHt7fTc6BT41
BXbLiMCYHtbDCRVHS+uDHHwClk7JNjuAt/HsYgtQoyEaAQYcGOjy9v+poOKRt82sbM23F8jZj3JH
vsbPOPCGcb6Nhzat/uqLrqHjtgcRZjR42hAosxPfQ9VX/tUqI+cOy0QLA5y+ncSwQnoopr006zr1
88+2f7e0dscp/ZR7kYV3R/dcMwvLJvAu7OiR0QSBGKR2FJEgg04v7j3EUFGWsSuhRQOssx1fgIM2
JSbibxyDilqe9p2BWK+0RZ13/rgGuUmZUaw7jiBugx/f4UDHbZYHCOYtp09TILW6BQamwVBadS0V
n1OPjTR1PX36RwANbvdA6ZE515poU4fWDHYGV2X4TN0+r+BU6DqRjJXABymTQ4oYpsdjH6j8+UaP
e9J80PjvRbX2wnkBTzLaKiTQSxVz94jhoAqDZIugUXXrgc4HYH04Xnimh3emvhJ6JOjzMDs2w/aq
/kpYAE9DYvSrf+a06YhodguyWmcWN/4fskAEN+la3YMAhaXkJv7RHApIPfYB79z9osPUo4m6lUPP
4XVgKtbk/7NLkBqZdx4/lqJ/EXxYrtm1d4QGt4r71B4QSXUkg6wJukYEAv516HzKrbJ7VLgsH0S0
gzyiZC8//fOrt4qBhXdvUMaOewOEJmRNDkG6a0aezmh1c3X6v6dsac9B8ldJPyZINcXK1tI12Z9a
d7ryVzjM0nhRDz7GnwWEB5QchOkp/PA3kVaOK2o1BhEdcDhc4Lp6Ch9JPGrg/PLZoH9OU4u5ITS/
eRkqgQ6Tc/5kLFiebei5sabTg+MetsliHUL/8piqEY7T5ClPqrDLCs77eM+rhBO8CFKv9arnz9vV
iardXjSzrbMQ/1KlbYrfahdjLL5e0Ha0CCHga8D6NIa6OPfdZNOoJMfzCSz+yHfFuSDo47mU0TxX
AAM0kOAh6fMGUy3GlAMJJSnp0lGezys9cVPuQwedav7hmHHypvTmLOronT7NFVC+ZVEE0dxQWA+K
RBpyzFhfQ0ImBEcMYmjuWCyxUCsLXkb6gSjyp0+1Uar8Vx9CdYzLbeAwbMD0A1jvxVRJnANvxZYK
M/2vkkzr1gsVF+Y5dTKYfbDdjc5cdp4ZQxZ8vSQ+9OzOq4HBt1LTrlDyl6xAlUk09VxNqudS0oIk
dekHdgBKnbwM4SKwTbaJI+8Qwi31xhRiyCMJMfhpmuKOKt63NjinudToz0XKhiImryLwpPstn8Jm
CXcUo6Cza7tqduUpMnOpW8U1UWwfZglBcrWpTc5s0kQqzQnsLTCfgSBEdSxrdowGECBXo22wF2Bf
re6PMQlPgZ2rLO62W8b7Eqh0ZLmUUredwiRa6wpA/NkadKxB3cOJp8+gqJoWujlwMbLQvlkyE6hn
OJMcFyBN6LDPp3/3ByuEmU8jYE5tdAODGBdLT3bD3haUWUaGRKZqYrhkGGey/cgTRAEyfTrlILVr
EiCQtVTrKkFzm7TCAswbB68EqiWOULpnu1WSdrZaSjnnh9bEl8Vdn8WjOULv4JkSomVSy1pKEM6q
f3k+p8BE/EOonEX97sseLXnl3bIO7TU+7Zwi+iTIzbsFnUWNdSfGNWb1DSSI+P31GrrN80PoMtH+
qPQwR8dgMgWIxBOiax/VXq1gL4UcndQb9XMiWVrOSePUoDGssne0VhrLG2cgasv/P12GejyHIVGr
BxWz5PQtAlnKK1D74bg/ihn4oGzR36j98OUser1jEfTzq32o9atl1VBNb9kIYuBpYaQDgSv31B9e
AQNM3ufoKetFE4UYghHwi5Y7h1yYhP5jADYKwejR3SPPBIbjVm3cqEGoh5ftSoNwFmTn9VSYt3Nv
ZEUQ84Dk2YPmrk9Gf+HBizyV9rGkJT+78Sum39SL1y15Cda/+43EbeI5yxVjzR+q/PfX+6m3bDg3
QQagOh/OwrpHaXGI0ZkU+jGIbM5s0wpGgVARnSFYkjLnk/ScWZFnoFQs3ILzK7kxHswe+2Km3i0w
ahcalBa+Rjnlfq0SZFzhQsUBozQlBQDYxPPr1pqfugUwugv+1J7xwcKLOjbS3AG1BVBZpMiZDkWi
iFQu8r/R5WOYKivLazMU34iOMbqnjxFi0IJP7wfdxCrX1K3UaZO83rawbLUPDJDwmnhsXMtp3kcS
k+htBvOv0P8fzJVhqPpOsDlfDxM1VuI91SJOUBLY59u2+ZDO31b8QHUFHlvsMAs4SsKsu+h3zO6Y
eXFdnkTFTXgqsP4U5NUMnZbO82w/6w/ExHLHLcRt8hmBEIUWn8N/Ysf2aUuQCyOgRB3sMiEpKZu2
ysIM/KvHkAxx4YZMxB1gvARfUrvJbJEu/+zGidWYdFC46fBTD/UQCGEIwN12shyVWzB/ryuYjERM
mQVl/oiHDKzuQI6cOK9QtigfEVipkjYPGD8LK0h3IHCA+rNXgfTLU0EF5erWKuhg9IOtw8kopOwD
ycScW6I29l+9+/6bNK0rEyQtMvzZRB2aJdEgAVLp3kI7VKDVDImPxmVNJUdjOkzoCL2/y1KyoTbm
0O2wNL2KS0keJUvfveqFmDYUlFTdSMM1wDGemZXMGAU+SW2g2bQH2WpHSHmPXb82G+Y0bDdAkCak
lyg9lsgCMg+QQCqEO6ViR0ELppEfBYFyu+P/x2MRsMCLUwD2R/WkpMX4D3u4fSKslD/Lzw6FlI0t
RkaeuNPlJt/+ULtJODmgpgo1XV7BNYmIjRO3M10RxKbddbqxbnmmxeeNtd4cC0RIjesWH6T8MgBf
HBRHDo5EY6NgSzvLCKnYAraA0yf4It11iMa+kEZ23ISKIUM9K3l2ubizdJysupPoAxFB8shL09TV
sV6F566LNSznM6uEaJ18f8B/dnwEbtnzKy+coJEzxaGz4TZftg7o/9LovHLLRuueJsb+KayN7v+9
xlm+oo9sw0EVCTGj3Dsn/BSsl4PcdHIS6LYGDTs1dMLAIIsYs2U8rEI3urTAQt4TcGiEc0Z7mqrY
KQv3/JwigHs2ADeoLCfsQAj4LW8ogC6QAAMGpwrRfn7CRVgjfzxOqI2soBdBJjaz/fV7GytvefTc
GRlfwZbmHa4oh3vaUGRp1vcgfv+AmFpfzNIXfQk38j1UMx67/mk0lCIkmG765aQduq+v1HDESA4i
38BITh9tl9ywfksOVACBbAhX9nhR0e44okuDhOmpoO5h8nTEcEHiJ/jOFKhnK3cSJB9chRkG5grK
Mfcxhoea+u3fsg36Rr2/v0qBKdA32Fsdu6d+KeNrcSkOQXTYgRDR4Cxtbj8GMheHZo1w93EY8pu6
A89hHdyaTg3S8DxGET77lYul54KWx0zHplNk7OSgbsmh3tA69W2sdfz8cPVwwVHZjd+0QImuSy2u
/ws6d/99D+Fjego0AbhXcd8L9cEmZd/eBmgJE9GzCa6DdYQue/qL9rKHDhOkTaCiyw0d7QZM652Z
y+wcaU7Vl3CGbydx+Gb3DSuB+I7WxPx2rOOrYYk39HMC2g18ys+HGj7EpX9CE2GrDxcEgb0Pgt6a
muqZUb3S+wp/ZqmdjZti7VhE24w/e2NQTtkh6pLaRH14amHLwFwu4/8mpfOdtR8CYBHXJbHDxyY/
UCXNRNiY5Ufbq5GbuuNrmFBg55Jfh+a2KFAk6f/qD/7nERv0pVU3UQQz88szXQ+EIBolLwJwIFUm
7VTle7j8obsvDlKnUBHN4Q9JTOvX4N3NX+HigAt15AVGl0JODVv2GjVlPDkgKm3Lvt4RPJ1wqfFj
JiJhMOF/Yu2bDKQ9eGs2FpAkj3cYU6UrkZFgxgw7dB4xZm8xckpDMhA1s30me4nX/F2jDzmOrtcD
B3FaiONndZ5KZfdAgBZV1APirNLUOERYSfHBn7dyeeskELGEZyWeueNo9V/ZaBqTCaVbCk6vKjKQ
YcAlmfA+VC4AOtyaWTCdx/Nsle12LnPijp1PaimPX1GsZF327COzu8elkAH8LdEir5rW5HYM7Jft
Rf+cSp9n/x8AJbY3N0OL4AE/E95nI8OICi6vHBUPmojpwwLBo9TE/obyNF798R3yWFxVdvzrUjMT
d3B8LtziX1icXxv01BL3Sgsqi8aIeRA9MuJySYlj1kOr1f/xxB9bK82jqZM+lsfbd/iNpua+UYRG
6uvyAxXHXcie72UI+aAZ1VkwE27N+R7jhMfAOz2hOSdyRnsEtYjFio/OSEmbcZNEfd17UxUxeo4F
DLaOXO5v8eRi4iCWiWxaDvOdXyhvZN5E9bOszE21TIDQMr8nDIo6DR69Hi4vL44iTWMgkJofhTB0
eZcSg93EAZej991f7PPYyyqHc8SmnCmRJHriTRv1Sue1ETu5NmRcm4N3YnHZpeItPcz2zAv3hfIg
T55ZvyvyN14m/o2kdCHRdpnXz4ZdwfMRU2/UVgIQrBPZ6GqDbnFSuPT2cJvoP9CKuR9vWEoVm5Fs
ruUE3rn6PwQyoUyrVq63//i/4r69EbV6PLzZXION75FwfxanjI5m8oaAviABz4kO3xuxX+1S0rXn
qAJCrIdmX9cNvoQInJVGf7QL9DAccZsrB4x9XPP2l8kizZ5w8M5aQw1A5Xc7V3RvTOmfcjDNtlDq
50a4aCUHaPfHVz1wf/Xb9WJQbnh3kWp9TXzl46dUdLCrMMLw0AnK9Y/hqMZ11o8xg6P6/FHGsIiT
043IhPkzhicDWJTjy7MyNJRhTnnMOTSljfe475hpsAfJ+q20nstwlvC5q8X3nYqrvvAdv6qiHTxT
9P16zy8nsYinSm+6qS3gxRqdP4uYNz09c+/IJifaRVif8uVLeTifsycgOda0IwWvurGKund/11EO
BfFZNMugrRYZGRP6Xyl3F73b77jr/HtpiPI8o0IwrCZ5pomnk/EgouThog+p+9qkKH3+05W7Jc4S
8HukOZI+ZcfJDslUZbNibfU/uirdpYVs8F2ViP7oOP+WeueDmhws1mPTN4nYnw5Uv5l3aMNZjVHQ
ErFCJUzmaUxIabwnO/aH8Y3wW3NWI6T77MT0PVg6dAWoaJ9YkzXnHbzw02YYznRkhTMK7ZHPhXD/
VrE/9qtXMlQGBsKHXilegcCGafI6idIvDvYd1VjxcnVkhlDoMlLI1pNzLTLzgI5xUyJPgWQRCoyC
Pxo3nG71wiU4vuhJkDrRUdTrMgBg14rB6FwQ+wmJcgsWoMjVcMgZ9jSC19l9sNrA9fYMqXFoAJvQ
zjm6MEnRi4i0ZXWUchVP14ZaFofYGjjUop1ZUzjTJp2CE1lK14bSIoJcR/tAv37PHPaSdEMDLrNI
f5bwJMlkop8d7MY90UkYmDBWrtxN4P+W8US+COAANaDHPMULUeeyzzZN6jhy/wgff5Ed0xKtqKRG
/bkLaw+crCNj36utio7qMFxbNR1yBQUFF5WTVY7g+je3gc4XkwfHEyVwIT92Xgp8XAnr0NPXp+yR
vqeRmRx/yHN5pJHn96DKASw1dyvNJUmx2CCiARe72k3mtUr8f9O0GkZ8B4qdDAPnBwVQrfAQZXCF
X3UMyeu7hFTVGj4bXRkcIghfs5wxd/TEC3YgFBOWmnmaVtWkV374z6fPPH0iud1l0hDYs8GmBeaL
E1fNw1zYq9UXGhhe6AofEEAE2CYJf0NX79LigQ7nhxS3g1rO+oWQh3XUk+ilyb3XmGg8m972Lo1M
2daGlPuuUavlmi6gisft6MNREScirQiIE891DXtWVGNu/I0piqVBXdxQ/cISNZqAjGS3qeFQLyVa
sf+wR9eA/1+rW9tPySKRRpp5IBWP8QGhDzpEGxzB9fCkIyJj9Swq6mFxkVZasP8PENNIkgHTT8eO
ylXv63UPIpQ/x9hPPlSInN2xkAqVQD5hgiYaRvzc+vTN1oAJiIbgV9J7E0S97Hp18aZP6t39z5GV
JrLfmm6TUDrV9tIzoLnVp5iX6iQvFKNdvAGdNPg19zjn/jwd7+PC7yz/J5GAO7NZmzxj1VZe+T4e
1PbdK1KivbzKa+mrpmSeadTRnLHhj1N5D3MA6HLzS6DJoCbbFpeKVjB5O3GRNPpNfI265IfV1WvF
9XZNacxj/kFPwo50sutzzTdQce/2+OP+dA7c35bU+S57699yWJpYdjgviSdxmXARPZTrD5ouQRC0
TKz2we7qI/e9RkxpgkjCIh2sMhh/4CIB7K2f+GbMiFp/3J0zWn6lc/mO0xuXBB2/WxPgnHGkHFq8
LP3Y77Mu34f4NEC1cV7zpR674n4eqE+2hCfSdkxWqVDumsJk20Ax/2uHSIPNuLgXWoZVmZA81y1a
9PlfDupU/1QzvgGDuoQeP4W06clnK2axng4TcOdG2Spg6DJaf1/hAEiT4805gDpFf8MZ3BUam4dh
YtUmqMGKcQPXxU0aJ6N6Gan07fXBJmtHPGYemGcExVWMW9wk8vT4kONG+asYgKVv5qB7hA/ibwyY
YJeq62uZprMdejKVRzAQmDXeTMyAAq0AdY2BWl9Gxv8t/9s6VrqoDqPFCNkFu4dOHLNAFuk2GQJU
Ii52f8hpm/KG26QfOtjbItcHwY6ubR7K8/YE3PGNFtb4h+bkkKBr5tPwkJKgdX81gUrPVY3AfmGz
KapT7rJniFrPZi2HDD2Y3Z8L7XFiltXRfr18rnWAhPXZcBWQAlqRlXxU4iXPNjesJKITc+zORuvH
gbtYiU8H8oxIorPyaqVoiteecHGFEliGqoWahI0cObJDSOcBhwk1zxcYB6VtH6f9s61jes6wEhcZ
3OzH24nq5+hVZfWqXvHEaXzlHruEj7542RWfNT9C7BbsJ4Dl2uwm/iogwgqYa/1U06CMq3iPTnuR
v0MUqh6cctQArcF2E/BXYAokTn+KfZa25d15qNivtn63y6v4WuGQ93cGc1xsvtZFeHQAGmRdYy0Y
Q4eQUylKITm4WkBbKEQpTRGobQVWP+iS769+7noMPfZHvQvIIyyLAXqfUFE9i2svdcuepVBtDSUS
yC4msZXjS5WIopafVEbv8mnodYWRPAa1CuJejsysuq7MJfEvl+LNoZDMf4GQJ9m2IdatBW06DpBZ
DdzGqt1YPuQXflv71Ihl6vKjGuQBXtARzkSAi9iUt5h7nyMPlOwgO+LpEDFYCim3Y3W+c92yUfny
cYCoGQQ2tlDPSUXmRWQpkvuk6JaSI+ZyLyVzsrE3ANUpqNoMgzAgXZ418PXcm6sNG1wCNySnWVRo
oshxXaE68ffyawc58eJNAUE+t+mM6HfpX4ZRKT0kQiucWlHKJ7EyuugkcfxZtpeB9usGRPPkzR3p
W6xszUz9JaufMyFJcYNaFVTwVbxRqaSAFegpZWeDpdcJ4U1aaLAua9racetReO/vF3GjR5Lkf2C1
daA2y89IiIpNUfSyY9VJ5kS6/EU6ffPezrQzO2R3jOMr6NaeD5MR/rwoTiG+alaGgtjc3E9KXCZT
PVdYypG4OimBBjTpvMTzMREeYXri3M6ajem2Av75TlO4UHP0+cnxyeYk+GmNpNZfjge7BVxEZBcB
2YDYeSzVhIoQoa1SLakorNkWDKRmZUa+7hZDWefz7dzgOTUoKo3zgMx0gjRQXbBMRdEIldg2DyA7
xpTbCYyznS+bXkqNMcuzMH31G6xOH2BCugxrBk8k2Q1QQvgdR7QXPEayV9mIBnOFtvToApJODyJX
pTa6OH6CNfrwDgVx93Q9NknG2kQ0NZrhYbFrW2ahWb5Svh+wY5iJkaZ0IJAY/18M5RBOqOZ5Y4cO
DkhOsd4dz4SZsgcM6MljN5VqTqbnxWAGUnY+hcGQUQmPOGtGwBFxkmv0TvqoIYucSwKA4qj4pOdM
j4T4iy0lTW5+p6m1x9WS3MOoIKteedfvBS/GonrG7T2+4QY2hG1EFSXgSmd9PEagr5kLD6Zxo+Ly
I0DEZH64M+MWJM+1JNJWnSKInTo/7zWtBUEX3hWGKIXFwz4Cu55ejeJF3dxVWftGezaD3PuKav71
z781SHC1R5lvo52blB5hdX4a8fCxDjDpg2ZasgYalgnVnnktxSrPG8La8CXApPlMwZzjmCa964U2
Lglho+qBbDYAm4Q4jGssX0oS2wbCbvTT1J4lhb2eQSq6B1KkqIFLZ5rZV3cnRqetrZVFY6/0+s6G
vJlNlksiiSufWo2HKi4KoQmFTh/w7WjJ0REGzq58fiIvirOdMP/hiTzjsdmOJpYZZM6Rvc3fUzCg
zvXrd4Cyh1IEWJrSBWw5Fm1nSL8w6Y6q6aVLs/Ytlibl2u2EP22CdcrUqdThCnbVXKiDG5iPkJqQ
hbP2qaB6cmkWTRtjJjZY68OuTb/90cwe0bIGV9ePrvOij8gLSZ6Zf4337gyWSRwCVF6qMIpJwIuj
LtjUHfUuMKDCzQz9eHzUmtimlBzwN8CPUGF+MDbTbX/G2Q45CVRjABTDaXMLKyjLzak+ArXqkoFk
Pp1LXQEXMCfD/MZKw7Q0EkP1PUZJ6DXNwv+L3VKpxnQNJOIxITp093GjVtDL6A5WG0ey09nqa7fs
29lxVedxCvrOlT+ouISQk27b8W+c0cjbG5G4SYKdkfYXZ5ZAfz1YvayvwSiTX4LOBgKowmCdcsMH
vF7jAmMiPeXRTdK3l+QIOQzKV6FQu7dhZkk0xyQqAsv2znK8CWmHukvRiycRS/MWwX/ic+pHySBy
VEKj1zz9Bo3VTGD9JSyXdNHeR3VITA9+hon7yAsvBr+UcChrJawP3nUhkuEwoATQESLkXh7jCMoS
+pSJVQBtMeIbzi9I40jgvJVPmxyAvik0GNOvEt5xwZ6V7ur1SVLeyacjvwzG20oY7EKh1hJg9Rga
8OPC7miYDxD2KvLhsAMj4hSRNFGR60hF4XojDxADtJIt0W/IU8IxkqGQ2Y1eBry7BJuSWnUYOnZS
DZdKPuAmfxlIRQyQtrQbosx2Qu4GlhHaLKg37IR7JEuyj0cGEa2vccjhwwFbyHE0Yjf40lhtBd+C
4crZO43Vx6xl0cYTb7vUHPVLn68gZ8BwgtEetUV1HuMkwo8vcDim6LsMegiFAZct28vOAUFpxMNF
EBcblVYVkfYWhbLt/pQYbmODfqcv1zZEXYG71ej8ji/hL+lVeX3+pyZePJP1pYJrqNP+AGhJU9yU
NLJiO4ykIPt4p06pXlrt7qLcQRlPKDm4ZLEOHORXcrcDU+Q18qy157E7jSaogriouM3sp0yalZF9
Wc/SiPCmfuLa/5OK7y0ueF1UtWmrlO6FTziP+wzPqJ86TjRMwQPQXFbf8V0yPoz07tljVC3fQZFV
MRqMySw6fHpxo7HtvSi8R583Ahf0CjNP8ZIqQQ2Mrq3qiKgLlWDTo58n5PcMF5Wc8yzs/P/RGw47
pbPpfmVbNvS/4GPsI4HgRItO2GQAwKoyzOPgpCm9jI0vcLjvBW9FaEZl//Cxi0dNYM1HCc8+fCr2
Hh59plGW0pcfhM+ogJDN4iteUO43ic8XJHpQ7apfx53lnp1tsa+F3iTvTrAr894v9BykHzE36r5O
s1fQLjSZIvTWCIZzjDON9dNvJ1I8j1Sdm1dGOgXpJR5b7DkUEGs/K2NY2W80SQqdZfTSbr/wepte
RB3dZ85pPnvSDEQlpwMOuAbS6n2H4bUmg1AdoYxOLJPT8/CWObbU6ddywbsC83giblH6w9VV2STs
qVpPZDb3dUoR9gH3VrDMMd2azliA56Do1cVadndQMO/5c3XI8ZIVuyLhrwoffjzz6I9X3Pa6nbpS
QJ8sfKrFdhFXswBsiSRXiC8H+2E2uhFdGJlFb7KzEQUDDPphFeOtYTcheRlGNmIfdEUfr9aCXgQQ
KFoXBvSTGcL/9A4/zGxp7+1z1va8o6oLFHV+9HuzmRYnewa4w/FRLeHtLgN6WpVAHWFeeNo8LkmS
YA/K6WocxiW6QH24O4PVkNzrgFU3xDFhJU0UYeElDtb4XZcadt3mytov/7vClhp8qHnHjJGrK7si
VFNhTWVJRWBz6mTKon6yMzUUYQvWO9h03Vq9TPu6AlMzey/u6JLBB0plku76wJ1I/YMu0eexh8bP
cifeyERYP+2girCTl4KT50IX8oGW7cD3QfNB9ss6uREnEz8DdrhoLUXD1MDz2Ki9nSBpYZOQpTn4
b9EsXsWEHzTJ/hq+P3tYzB8qaqL5oAGpY1TunSG9rOdwaLSExp66SUXdvBtxuJmuYGZU6nar3wnE
ysIFyQxS4p3m42KEB1o+2dPTuRjMZ9wnc5E0Sh7JGTyawsi4g6bfTCeAbqBGsgzRJ0g6DzEiwPtM
W6cz+AwQUD7n2kXy0iyj0vLWVDks9SmU+EWqxtpROmJtJlq/r9bCOB+xFhqd1PAj3yreQyW+89FC
B2AoJ441M26fVROn7UZoai3kdtZ276tNB3wkC9VwLAmKfpsx+kZS5UkeK4pLhoSxrBi3FT4frYXB
WqfZCIL+/GmToQAPU6bjJI9qZ4DMiDtj2Z9S43luFlS0GW4GHjRO5tx0AbsW797Us3pMTW42bi7R
2X0cvPMXe5K5clpftZ9N9yOWEfcvQixIwVzmyO7084XP/Z1KlWCDTuGEXGPZRT+cgoDkWGcOzbnI
r6zrVyQg4uV1md0w0yRHlgxCFbAUlaz+hgDuVnXheSjK8AdvW23NSlbRLMEQRM21cdRyoEz9jjmo
Wx0D2j5AUFPKMsR+ixyymln08+hjEw8lDd3r2h35rZf0ecq3wNp3aHOMDbCqIXbT0nFLRO6JWjJ3
diGM0AUE0CIzo+dySlHzrQUeRRQIZkUw9oPm2emItmdcxVPyJt+jgebB8ZBoUusnPFOYBG2jG8DN
Enb0eMZNfKuvK+Y+PmKrDl4aaOCPVGRmr/Sw9tjvb59G/pMJ+yew3GPH1tFIijTIErogh79Xls+W
1xOlX2mPHjxQhJ8RGVyCXaLmG6/kDde601MAsR8hyiR4T3CQgqtrRtvi5MJDHhZhaw3EIxmt8mvb
JvFLypBihW49JrWZXaZGGsZcwIpv+Zk+ttNvXg48VyLNcQNkL9oYq6SAfky9tWk2F1Dt4lQNoB7K
BrM3zCDwOyo6jAGCPi5o7ygCZECl2tAL7IWwAhMajp2d+KkrxEEQ08rIbwLV19P+xAlQGETAYR6I
UQd/fd0CZhsEdgn7Hf+f4MHuvg5+x4fw8DIC/4lgBnd6BFITZlVMHltjoHEtYnYRpHnVhvoQOaND
ZXBgtGqMr+I8ENlQF0Qv32U/N9kps6Yzj6bCNDi7zmjpdYud18ZcQGj5U5gRmWkWtI1HCxmjAwh5
gM5rUEdSINpjZqLdH1ZGx19zYJhyOGTZQdZFP45IledI9foj/8fqbCBSejwXBh+vMRePP7e92Ioa
1AZqWbePFJ94OBLkXVxyU8GvKPBJFf60WjeLYpNuUH9SxBzxRmj8ug9aGt43b8W1WwJRhyUSwzsj
Q8pkqxLy+q4cEpirvxFMI2OI9/Ic8occI27sQFh8Oy2NWsZZ4MBkezdx6c+rVCN91DOIG/OzTXQb
9veBpuXV5diIhVqyFW2IFBWdT/R++FMVluh+S00D5E4m7jDoVyB2Ms32W4t70GGzQcWaUdYrpAZK
1UrOVdeeyX5oLQLGT83Xjpf0nigMIaZxIu0WZHVVVHDEUxbgmJBdQjz7wSxanDyz0mEH4v77ByKv
k0RChuQV+ZdfCJY6ASC7VjGWAlO+I/zea8mrQiZHKEtzO8yzSq/WKLStwelVHM/IXHZL+tLzpMbq
gS4D1p3SN8myeInRD6I8fpfwj89uAOeuEV3moZIu3etxftNy7DlPNGVkcZesF1FblWur/514b0tS
RJCj8EBXYaiRGLUR4Ei+BkCqYP2WBb/JssQL1T+E2kfJEtm2hlFvMI+G+PeQqpOdNygmPWFLRdWq
j0NSVidfAtgQ/TRVNToonCv04IUUgzSOLSfzm9D8jJgwAFyEsTFARzqdNGUOGo6L39QOpogVVGqF
7V35WfZKZdO0Bk85EikBSiPSUwCk0wRfaZunQ/KJEamXuWKYnp43u5qZpdUZueS8i+1PwCZVLcVX
XWjAlDprk18VCWM7QZ+nz0blICdJ20H0zFnAvuNajfGQlaqqeqAaEud7TWILe72v+2R8cc+R79wq
1ozR5/7y3/t1f8wBcbrolaBboihD3l9FRaE/76GpDMuphLWWrIE+RzFDRIrTXEVpEUXaQ5Gkjo4h
yORBtZkEC7eyWI44ru49VY2xCY99cTVIgNVZ1GTvGZqsETjeC2FLyqF+eF9bzEH9vSHMWuVr7vo1
DtSA2TZ7jZpZyAAiHu6BU2oOoraCRM2K/z31Vop37oiJqBuy3x3ncoCUUP8HisAddTSjMKkylIo3
DTIq9LEEuSgUA8sSXtSOsXUZyb1yf3l3aG6XJDaizZ8VLbwIfsSIz7TCEmIEbBNtD60tfugkivTu
VoEqFYes9dh1VV2kzf4Rk2yWzj9Xsfpz7Q+gkwnPiBtNyQo19OflcbIw+9n5ImDF5J3154Hh6624
bq4uWhy4yX8hcueOctSzIjhAyEboTtyNKoGlWD8PUfKpji7vzmM5h8zGuxzM5FdpYRYdBUPklTkN
r8eBEwEKxvCv94tCYrvFWh4Wu/rcv5vsZ9DfKBXjxoMOEFU4XMhXAME/Zl/UJ2AkVXrm80ymV8yI
3kC/9ahHIWtnFOm/MpOTJ9MmCr33G31i6L78t6QEbICNUbaYovhkicdvOY2o0vguqoGW72zMCsrK
snRgsU08j9402Oo3lV1AsN8xFQxV0IacNacpkT/UnzrcHVOfmuHbtQdKSihIWeWMdZJYc73tzAQY
QY300vEyiNI/yw1yZMUezsKDzb8O4HDtKbu3IYCaZvG52YimImiCNmilgsMIHqRNhknW3d0U3Qtm
TnED6ouCsBX3qAKAf6lukYSKcAX5YDa3qScIjQza0AtFs0kJfwHCmGMnkVC1sgG07y3JJLSWTs7q
jxIjZLgXBdNIiP/xB0Xcx6F/rFL14IRWblqYIxzQRH6ZB4poCw83sXFu3wMFDU95KWjvZOA6yRMT
egu/Wr7O7xFRWGbQ5Bc/fSwYcq+PJA8HSVNXATf54UmqMfEw1+8t2O9Ngcb4wwifxYR+eNIv1f4W
IcqQxJxqaPUP0S2joAN/sFt+THnen0BWDaZUhaKLMqOOj+HAEHscQH9OH0Pe8s/PK3FLhftaiFmo
9gmSiTmGsFEyeneBPwKf4MXUNu/quN2mOhEdHWpTC7lfxRDXjjJJZP4aA0iHIO6OF8UYnz68Wd/e
YVNt+lN1gZKm9z5zbXSLndLJWbbT7mIaXvp5taTGT3Zx4J+roLw6x+Dgb6eHbC7fxzJl5Hg9Co0c
pkdpc2VcRo4h4Y7TjxIkNWMwMseA7qpeaKJYRjpL1jlrXyPgFsSyRR7ZhdWPSr6RSQ815YhO2m14
1bKf4Onmtvdek7pDpsr/6C6z9HPjvavuMz8bo8t5C8I9q3xZyqMM+8eyGEfUG2MFgmsY0kmpRps9
SirThAnnaRGvx89ohPbB+HGcpKLCn50TOAUblL05dw6SiAN3G5b+IbEUjccsW2Pn9gmYeUgZDiB2
Jukz2pX9pCbKnQ31C9/9X4kZMErU90UZu2EGQhhv1OPLFRHwTbFEC4d5aTmtmMCH9Dy4JQpqkJS9
8eTHxpEEPLu2jmn15EoxuKP+Mk94RE6xgj+fQxDBJHLU76JeHhIxtOEbL7H1zxQu53tqrx0mrf0b
V8oM/bp5gotOrHwv8Gz7NfiH9c7LbzO5U4W2tv1MjMPsX5kc0kP6edk45LlAwQiRJtnTmKwsbUYK
f0yI3E8jjvTLQdh55/c4js2U/1WkO9Xsj2YKauWEidHkX6WYz5pqhzFtPZu7FrEm728c+ADxKBVK
HBIAVAbK22fh0jeD0uPRh+pXYtc8aXBOdZR9m9BeBxDX/d92Q8poM5KVeqZcQUOwJQf3ib8oFD/p
d3wMSCA4FEhCErwiw0jm61UHgnc0KD66idcinuFVMg/A4kCIZ1VB0AaSGmMbgdHCfCjyYRzMoC9i
bYuU8fQjETU08YrkuNwiZ8B8qQJsPyUQoCa9crfzZUVnm/kLhxz5ggmiiU4vdqUuI7Xw/ENiG2SO
cynrLPqO5qD42MtWSBOUUy1lYLUf1YbM7/kSk3Kir+eAyizUnvqrz5zvSU4SIb5agpg8WOL514NN
0bF9vqYVuIeplUXTBPQ9A+o7+ApSPTiw1SOXTsCKJTfa9jTcpHTOG0SZcn6nxlmTBEPe/z91PIZf
/K5vbCQa160zqvEOtg01zn3Hef9lZXd4ivuxYebiI5eHvAguSpLozk47qpqxHICnRXb8DO0qrkiS
AF/mOsoOkLvUqr9KbXIT/P1MDScgvy7LmdTy+bG8H8Q43CxcpKLXtp5Iqm4MPlFGFjpQi/rx/n4k
rWWMYYoG9pUb3CxQVqZ1IYxaNRotpLard5G9BMNIe5dhgBp7FiZbajbJ1VZ2fJaER+OsDNLkoKGy
wlQvUz4xciOnyQRzIHYeXytxgcHec9l9rbRcWdrlV4mfoGg/LhhHiSI7ZmPzlhmfg6TlCv0ah01X
rA3ISYTFQxMz41Wv0hLuGPiSiVws5fBn7IYtdzRBkMRGb4ul8VfRAEVbhyx9X/19muXwLJeFJh99
95H0AKQkYBEb3Ml2zR8edTIzeInvRb0lxk2/xmwDlLCj4bL/aalHBFwlnDnxA4k2DBge9kpZivID
VY4GeW9aU3/AN9Qypzq/scjQZCVCoPMX/NrsCv9l4/QxG4eCzC07sOTzG8To2/Z39VJS2NYhyF/z
Peok0ZTa06gGR/J4Q6QV8W6jINhiUEzncmk5hz8vCuRKmsCVg09cPFb75ow+IIiG9cr8aB/Ior44
15H5kIijJfzfXYgb29WYxaRP+O68pK9uHaFCOh0oraRUtVNGO51ZvpOvmmEqq2xZYF+NobH8mGpv
0fBOWKjhHrdnfaAq0TXQqkcuweRjmZxqbP5zMS7cY+AZ5xWvYvks3ACaQixuY8v7C46Mo1Afq6+P
mx/OGnXitgzV28wUMXJJkHkLeDQUUHNJuSTG6+MrU99qu62jMMub9y5v6VxbCc8Rzy3CZ9ilphiL
7ttg4bPi7AnQ4fcCyL0VbwmLfb5/laTAHElkq/9gT1LJFTjVtBh4x1LjFYAi1QGOBspG1SWt0OLI
FrDjzSzyNDRnygCLgBkGzH7CuSPk7PyB+EGPAyrNOV0dDQtM0sFhH0Yiw7hIa8tAZvuxEnZdoNae
zDsy7jpbODDKj4OvAk2GHwUPF70dnfzPcEOr/+jDRzMLHGibFzZrLdikRbpKJHxAisCDg0mCeK10
BtY7PUt89Bgi6t/G+DlgL9QYyXAC1LzVumIHJ0ZO+jwdbDU8Vk3SoV+0PaA2lDWk8T3JDeFA7wgC
F+Ue4GsHQIVnhB+9Geib14ykrsgNkk5ujaLpMZGH8vx77KHEK4U9jf32PF5Yz8tFNINeoEG/txky
vsfCPFkXZpIbdqydF1A/hoptLegd2+TC0CqD03yhpFZZ3jhSEITZFTR9biu9cTZN3EmaidL0jUiw
mVTN2hoe4yiaLzj4zI55jmEit4duu6KiYrNzmTeUbq7WwAYh8wVjxJG3Ud+bpvjJMwSYEviJ42ST
Y0M7elIy72J2kLkcXX/ugYqIainMzPKBK17yoQnZUydKNbneSExtrjfVfuMOFSeDDqiqGc0QG1gv
pXpkmEDLN9kPW2xUAoJxq83uX8pkKJfg5nyM85Uslvje0FShYlB0E2xGkfpz6YGDSlsD1LpAA/DH
p2mr6obbh5MwkqCXqfiSkxipyvRGuUd9Educ2IxzPudTWFrsIV6zK6dftNgRpJp4DtMgNpkTx/sG
QMiACsCaUvlTarf9C3jpU6NcARGSTF+9ShRXqbKc1xkjZry77PQRXXpwqHQ2SPBmAyViuVF8aWN+
h1FXHsKTy+4fgmXk0AlLKykMQtl0CFLe6UG/koAoUu0Tpx341VCRdQKfyJiblTXjZ8l9MFuCQSOO
pYntVgQOvrVJLTHHmMl5OB+Dk9zr2Icw10vsjwe3RTpXVdrzBAt8VgWfMupOVZLufWMl+ALmvnTp
KXFWgDPo3toXvdEdKMq/MpwMLVFBc0JjToYJoM5iIy3e8qdIOOaa+2m73KxIu7lrhSLLG7qiqvK6
Pq7YCVMd365ZW34Z84J9brHBQQsitxbZh8M2r3LN7SqDTUBD8ulMHsKfkaoDyyAwBMhRQhdWELGj
eiku0nhVGkLPiVGyr3Zel4QBJUoi0Bpqq3VGiKrzvHuVPGYWn1HsClwZyyGvXSIu5TedflFFNQzV
Zqkr3IRRtVef7zC3BGnBvcquQkOfRuNtoBNxBBEgFd2HsUgaH4FRpp8NhvkAbLq+53eaK3TRQP7G
POjU/yCoEHS9a2tJaruXxvSb2BMttLMjGgDbEP92yRLIz9vrCq7X/RkInV0bhMMWbk9V+dOpRInA
AnxxK4buAklB3ALe7MIirA3LHTchyBpv4ChLfm+BfRLXKJNTPE4/kT14+AwVQDdz7jI0/T31vZTi
o3mFBBLegMwwet0mC+v5V4m5cfLHLQo1DXyqtOMF2H22oWF13okhCwnxSki1oKwYqOXvo9vRTqf2
PGSxG+wTHo1aDKpelCpl/CmGUYeBTtNqfP0opIY1rutCaNKY8PW95tGNoL5vMPuq08lQUztMEdKj
ZKBnTvwqcsdzm+iYn11GeRTq8/Sqm3nhaMz69XRx0lUte6Um6db7J1IXpzhH5AKV/Z/vhuJnRCYC
8lhAGvXSTUc48V7p1JwcSmFH8tnKa0oqEuAjsATFYmuH5GbCaBbnZw9Nmxxc1wZQUdDGUCNYIfcX
k8F69n4d2SqIhjXQ+tLB4XLaCoBBBzzxgM2vqxO5Dg+umGJX8Zx2+s+cE4rmRJtM4HqTB2/0KW1E
+sFBLqWePi3a0VSnuh1axrEO/PvGRjEwH+Ut6V1eQIXnLmxWm64zCTRi5MDq66x5lsF4LjgPk9eK
ZtPNcNSkJMtoUJM92clJvgpCBahY0mkEyDf/zZf3nT7n3MqklcMclrUssGRpp/e9XJ/WLf8lVhSU
99CH7d3Bd64CLffO+jFLKVEnc4Ilqmlq9znzo4Zo6IQuaLwf85wOd/iaYFdSWB9WVeNZ6YeUNK7G
Jf7bkePRb4CyB5y6u72gk9XAYHmLhAUqknowoTpz2I5OgsZ2FelIn7dcTEvH4HPfgcc0C+nACa+E
5HwQAXgaegLavYzlEGbjn0exbMaKSNeGFCVcn+KLZbUnyHlPfbTUh0qTMM0n99MSMOOvvmFPV1Oo
AUGHDq0e63voeNTa63JB+HYkzBS9f+ZlMMVuZz8+IhAcPL9LVKcYgeUQvbuGX/mVtwJeKW8bKYJO
+ALz0G5CIQdNYKNj/VPuSatGt9aJOQznGp8asSkPaP6xRuTUPqUBYXUZZtV+hFkyUhRvMN/3iZh9
zNSM8cdAAmL2V3qquqPrlwpm703kv7JVqf7t+GXuAg29jt9ZR05753ITwaeUjkgQFp3CptEoaFI4
1ieFLMRzjQCLiQ0LE7ynxxDSRqHVOm280D4PDzWYwDipwhTrXzLanLNg6kGc26NFf4RfJVpWKG9D
Fg+0QQZvQw/wyT6MDW0zO4SLmJ203KfyXVRdT/Ku4CHXuKQQI6si5bdlOalFwnRfcBF6IF+0EV+X
76+9fjPGt+JOqyYwNpJBtnAdZ0kgZx7tFI02+/UGysD35/vBc5UrIVgpibevBVbh0jsRryD4iMcZ
H7r1GbNkiB9rGsAFAYzEZg0x9dH7dcQWj50H1Qz8PGTL394EnAcbusNjiCd4aXUFaaJwsokgQUJL
pSppjB99gechHZesvjr3ZV4L0U53kzALbga23/gyW5ys8cX+Enii4tYEXutBC1zoVBJxxSB1tdrK
1kpkz2MPoVu4dQAFNn0QjyKnRsv6ca56BltCzp8z3LLS4F9BP3UZCCCX3N4tBeVwwsPa0YGtLlV2
rmZSJVD7exhWxtkv1JUs9/Tc17RmOmbKa9rTGuH354bhO4t0uSkzXBZnWfq1pvaApYRZxd1Pgnwp
fyM//Y8cm/VndRSV8wNhzynbFvgqDmK4C4dbxBWK4TEdmwOatRn87qVqRDxwWijjZ033pxXoCgVf
7/IjP9x8Xr/ZlNF031lxE7YgBHWy0EdlqTe01+GuOIZG4fTuGHqF6Nw65nXD7Cu2oCNxtGHEQp2p
BX/YrIEXj2ho0zvN7EMsjaU48DbBIVFZCzB3/BCnBJysRh5UzdyLuHq81xWGnM2pu+9mYQpFwM0D
CjSC1stGsw7LFXC6nSY9ZbAAXlDNgTWn+4BgnskMsU6ZEzOdPdWXwHLuK1rr2BemfwOK2GhOuEQc
B5YjDCK2bAovB5gL2tghA0mkwpeUdHBS9dopnvhQ9x6A+WuItIhsd5pwddfs0uqCTIe6DhMh0vB/
SaJvs5KfyZ4PzRU5kP5L7+eyVVddCI9mJNCNNfQDhInNizScp/Qe13zIlzTAuPeMcfP7o5zxtT3c
4X0M+LCdYfASNS8mzptwU9evNAQnEUhTmCaE33+eUR2NV0THokqIxLK7AdQGWPCVD0Xf17FDKmtF
XlmrKyt50Fl53FBt7OUqgiMf3oCJQ6yZZliYE8DvEurDYOb0xGrBlSeZ2RM3gALc8oaeqAuqggiQ
wtXGmzP3W9JDxhKJJQhHvOWfvzpz9+FOdJ2ztFYPvUMqDxDdLpjG44jjgqGxex6hx51x/s7zvbG4
kVNnwkg3muRlsB/QELvGHcXtECCi1Kn50/iiwlBJY9JY/tsf80VT0Q5TMA3dq8GTfNU8HoPpCm05
aS9nppDFCrn8aJ/cs/ClcUw+qM72dbHaQrJmhdHZ75yJwAz2ntdQYDjkOhnbx/0WMIcR5AscoGlc
d07AYUUp1T2zm2HCmod0fCuwL9orutFDEGd1bTXzfmOO45JFFB9WW1KH9wo3UjPFNCn2P0oohKAE
xJmWOs32KSIGhn6c+8svlhtTybIMJlTOEFEtRNLl0aU8skeTIGH4dh59Szu2MsXYZ7qLF1eY7UAm
l5dVws9jVo1U8geGf0+ESLYJZJiYISPCRhPA3P/Z/FFAWzszT3qaq4tT332MeCz70RxOjORcqgaL
L/UnxbBe8b5bwXKBCOM+27UCU7705CEELgUbTarUsIqgWQpGYZ075FVSL98kzUNmA0L9/GyRIXM7
KdUO+cj9DlzIwGKwfc6bLznuWmpx4EJKr82w1D4TkfoVCMI0WakXE+HEeku6t3N8FaculkuLMYxM
888g4nsXN2BKmEM6jqvZHCuMl4EOfy/asWqEt/AUn7wHNBlGheAsaV0fNuurvtmkqnxvKEpY0Pz5
aTA5qMH/kPVEGMpqXP9LlRoLROq0qy4aXPjpkGnxkhXxoaPJvjJpzllK/jbUgUGqOXRfG9NCY8of
3aqAbtLsoy8dctcpb/EBcF27uMoWkH+Kq511DUSXCsmWj4GQKfvEeEsMky+0qoQAy8NRGGxkCoY+
Ncb3mJ5NPannBl9lL2/YR1KmR9CMa7bT0dNCJqHIifPU6oMrUwsGWrcnJqRCi8QAONl0s+L0BWtX
OGnMevhP9Ox0d5nUL8RJDVjNrhusGu8Riz0DOsk9qRHp86u3GKXbJfYQuppjPm73al0sVjjOCuN4
duYvUy+RwgwP+5nsEyVydjamWxyLyiMFOQGmu9PniJEKRZ3BmfqlYn++UVWFlm7aO6Mpv58kAAbX
apHjlLJZcBpWV567fT6WWsvUyP3NqaPONKsu3kkGvVhY/K2ejVU2WQzdk4OcZ45ll8naweg3H06E
Rcdh8N0iX8KUylhCmBuxXJEMEDmeHtiM5NwXN0KrSTEUCf3nUtfxGtNl4+CL/YeskDGAgEHdC3g2
GIcQgMIJCo8l9S8coYJc8hSJWOHuIYazieOH/81r3dQM75htYyS7j46WHEcLbsxu8z5WGCFIoV/f
cYO0v1AwndCPNiWM7HsDqIv3fZ/AN+frO2bL2UVB/tvFTLY24u2egdCZZF6tMyhwTvzRkZxy1KcQ
M4uyIFR/OWxo29pw7vuvr60cGaq5KZzbLF3IQeX9U1+E+zs5t0STkwZ1WR2/aGzu/uwhlzqB50XD
NnVek3UpIM4NdoPDgcIBX1c2ZaAu7WoRFugjYJR9AgAKWYwdmtdDjmSM9yxT73naxVAptDvAUjoI
fn+2WD+mwy5kaIR2oeiD6rT89PpUqzHEJgeLKUvbRcGdSzJw8/WYzElgw2YUfFeHh1VN1au2iBXA
kl9W0YaPaMc0lt4gjYlc7WjJJI9uAnSIyECI/HV6HM63XxUaJ6inUyQNnFPFgTax/qZTygmlCgMy
QsQzXrTic/4zsbxMGnQa7sWSkR8WBj56OIYFGCI7MHWJ955znZHybZJ1Kf1uMumqkzAeBsSwLzSD
GHvoTv14BWosZivnTj/Mi5G+OjyvZNlC3z2X+NFToY21b+jOhDagRi7xjHsKICuH0WRIv8m1YTda
24rE5UaG7/KeDOKdHALdiFpsZS3ozPUx5IB6JcMIaT60PXmZrp16ppSuP0GKA2+x4Xr/WH65RKfk
xDpwlShPbm9mjP4PXKKXpNlaDZSPqCji1k0c8Er4H4nDnSk72IgKhEw9DNLLvyiXjabwD+WT4Ba0
XjwTawrGGTuAHGtTG+ix7l7NTIokZt9O71HfaFINZMoZeIz20mVciVYFebrqk357Y1wMwVxS5KWS
d8WXRqgvsDzc8qcJiA2lrOf8Ccc1D3LRNKzsY2S8fcUP6A5R5uXVf1Hr9adsVGQXn9Kh6neMiQPB
Hf6EZz2xsuHSoHfzlciYrBIvvHSsklIjAFdWB/A4aPOIegELP+L3c0dZzzA4ruo37P7cvPhgEJdA
KpDFx+soFVdByXRoqjluGEH69PCYazVL5Jy0GurzFJe4fNIy9THqSvUWYl4cIJRU6leJcQCJmVh8
Ih0T2Z4LGQG0OI+9TF0ZyYzAa6uT8u3dorgYrgVcKp7LhY5MPZ4nFFN7Xsn5Hnm3rr2YXNikEdXm
3AMIetjQY4WHLcXMoCzxGi7v11GI1AO5YaMOfhlJaASDTNhb8rFAtMnv/DOv7ZmMwOINlKVjqjcJ
DMtKgdjPxGVtyJ2h7b12G8SoQ2Au8xUBhznarCS/fYM5A5WrN0GGYtEc9amg7ivLnV7+ikdTWJfi
UGHQY11jy26dhsmZMTIPBW0MhVzTB++lUmiFveND2KcALKIjPsVNS5ZPqo2+ffTku9UMsVhoYAU+
cW1oP+17He2PFHJlnMVk/Li4o9Xp01DJKDAieRy7Jf5VHzIKnSk/tk8V9k5zdivsYQDx/L8gyeER
vCYe7YyiiyaiLyM1HOFzcH7i7IPk803thY6kCL1OcMXy2jBOm8MJQLkcNccVQoqjpArrF/ASnkKV
7xF0hQ7oEYBe17xKoodznGozHwBAA0IiHWQCJD3GnMADOeg+X9yAioh5LYsh8XcDcLcr8OLB0nZO
nkhHQsQBkq1N+9eyeqNCqOg+nFu1QGz9cyPNbdg2fLXLtDmmpm3jLZKrgpSutg6ggaEj/FLjuSeo
qOlH9DamyeqZ9XG98YnwwCpl910vkRLWUGS3BU8kHUITt2++Fvw9PESYa01lHwFVkj7qcFLJUj8B
snLtTUCGdqEbdQGu5Wj1mld5lIOaBGQGR8ra80mg2T0+oRrxVHpWz2hEswgc/mFTT0dtfnXYaYDI
fc3huflyPz6BDq/tfrxnDrEcIrKxVdyIrhev3QFTqkqxNzNp06A2WbreF7WkCA8i+fzZVJhnlqlR
uCxgFwwFQhyn3rH4A4zm3gJclTchs1cCYqUDLUFGx/x6kGSgrUqS+Sz8d7Die+crjU1nUv3catmu
eQ0hJQB9r2K9P/I0KYSQw/OCaQZnHj7DDCP9d8GbrEE+aSjLkYaq7lL4io0iK+d6ZG2z76mQPyDF
ViM/g2Hm3/XUUwJqn/lJWq3Q5Mps6wOvhrj9lBSY2/Iw5WZd4j/Nydbk6KDF8RZnr8nGlttF5sxv
eM8DIw82tKU6ASXj5yb3Zg0I6DEVGrfTncR5hTiiXV5XP/otHfGuYcSpNy5wNkreMr26WBY6YHrT
063eYCcd8h12hQTegB8Wp+Mj33L2Pp3q2MZ9lGrZGJXiCewOwX0ftaKUiCIgJcQozyNRzkjRCNWs
CZpHGJN2+EXvPbIvY1qSAG1yYamBtFmNN02IFjxpVodVXhnLEr6DC3bQmGIWx/cJZlH7KtJ97U2z
MHk55ojQmJFQVBA+ahiUueZBBGq7drOFJLfJZ0dHSr5N+ElShePqh8mK4O6jNXs6knoBvo5KWEx+
8Kg+QOS+Ma6QBjssM1j2YoL5EdK9Mb1i/yJBHrk2hN0+QdmnxHP94BqHKMIZye3K569jHc9k5xrg
QAvXQytfl+8W3Tvc0Qkw2LfTjmbAwCa4OOvBwveCNUOnDBPQcFEJjPw3LSEUeWXvQ/v+2oZYTBpo
krCPQ/ksYhtpjMbZBTfxTDGh0D3206DMYCZ80uiLqrz5SZUPvrGCD4UKcz5KaJ94T/X3TmYVhojj
PM0CojkaigdzCRnU7jydVlmMSHouXh5+lrLXzYP9+CagedgmrQDviZwSEUcD4NA74KWUanBlZA4s
VqeWP+NW3ve3cjsTARyJbotTElmMrJT3prGCWSAMVM0SidoBNDayPPToLWVvWMGo+W8OcSOKJppr
I7WuwAT+E6QnkSG5aS8dyGnR8rSJsDAPAcLMCIKq3VzfwzwgxDCE2T3p1Y9h79wNl8r4ZRxO4wuG
49WfBg3lFzNWRhFA29mMfvvHWxv7ErLAXB7wrFeqeno79q5he7/EFBobDJbZpNT5pJjpyDrhTwom
EvhKoeBUYJfBTOHobcDFEZjcbCn8xmNRnfpJn/Lr+SGmr0fngOC1LsIbrj92A4WzMU8iDt77VBNG
p7WuQce4X+JU0w8U2+DavKs1aQhIZTjlY/IcBgrYbSDnJuhn0J4ZuDmjpw7BPifShMAn0gjEy6si
M7bT0jNSFVQDFWtUnJmRy4Cgyo1PN9XXWtNEhELKDWSWmOyvDJAZ107eHCcs00QVNZbOV4ytlpVD
w9/Wb6DJhmwHa5cXVw4c7JF9Ei/XRjvurvClGVIXRlwUbgKXMKVAnyE5A376J+z5Fhe3fMBdhA0M
BCg4BatmbWtaZWLsfhNY3g2xpOimJ0L7lILjfL7svYb6RbYec4OwyjrxOEtB5cNYqAxjhC3zHw+G
2FuQ57VklcrwQNyCliR5Q/DDg0y5ZhXFUydabdTrxrcfP1nmLVwEXkr3/2p6Dxo59+sd0wE0UVWs
9tNuAMGJ+tmPyjWtzU76sSLJXTLyl1AK3Jvktcc8/JVnltNTn67OQjVi8kFDqOlWR2KxHYJ3vY2z
MNl08CSoqBTcGpk8aRCTnoR16iwFHsl1ZMOqpUHhCQbHgBw67SOwUva49ox1XvQe97/Ak1H+/ce/
jRzRtU/0vTq5Et/HmvBD/3yfhnaxseerwhgT8HOgKRUpl87+3MtAbycqMUzCsq/4FKeEItEvVnfK
Ip+zwlm+mkWudv4wnJU0cF9g+Wz2hxIRu5jVWCI8fX43TdZrYkQuoV3U9anrEDexiUEv7Llf351m
1P9UZZxtnW1uM9houY0zUkvyPwRgvIbItGhsBRH1U62XacVGKq8R3bbIdD9esIgh7k5EI99a6KXn
yNUDyGp7aDICqzvwzpgX8TJNgUlesU3BiTsrmvFnyglPcpF5qSEFCQ559EK0TnhxosWQTgsGQ1Nk
BezK2aocznU2vBqMgpEziESoUPvHAK8KIE5el7gDu7vEre6a3WzpodeUD6asZLSOYdF0UTHaxY+7
wKtKNjDsNjXq9x4zPzq//WXNEM7M7DrvG7q1AQq/8wQ/yUDN19AbI+S7Xdt4G1aflMq58me7/Mae
2DONCELULz0d97RiFThvBTLum0/BVIhzaSyI9jXGCkfV/Dr3ezCDdMTxAhkW4bYVlg+ftfl6J7/r
K1IqAL2R66KD5FoVfpaZA0J4WxOpGk9sWs14qEk2FZ6jGt33BNTph8Pr87v4hCWzf+KMlPLHA0Q3
Q2dMVXTPT4Ce+z/BfL/ieUFlS38TlQbTOTlV2QH4SBu5MC0IDACH3YYnwCGhITdRu0cWZHI4bxTi
fD64YpOaXiiLBYvvuX76Yx7/89Yn4abopOyHDtD70aevOmTuHhva4dBMwkHJHQ2J/fDa29X9HV+s
RF6qh8B9LRJUiwTAnnVkZdICfx0e79D0oW4qM0NaNT/2E/qiY1bxIf7Hb+FMc0j0a7oNWj15DWTi
RcnA0QcgT7H1l2nB7WAWwnR4A2zxU6j7t8QNhXXgGKcpt4frDKf9K/fKWuhR3GT7ftZagmqfyO0Z
UXEQYT4BoMisW3zziwyQByk4dlmmiT+HM/fYoqT6vrewqdjf6GTlmR2EzbMbjNXxoSFVOBxG4qgP
s2o9zfMGxPzFohNAJctFL/icVOfTwgC0sFrOgtoQLG5XnLEmqSKV68lvrV7YVM0EplQ7vRo8c2HB
JjpH2Con1rEXXGeOA6gHLDUeXgMxv8lZdiAlotFS37j9puXfRDsCInXQ7xjp2hUHw+iIZ+rolXu/
HhnnL55tPw6SnIe+QrY2GxeebmWBs+tgAA6g3JdnKxC2UnHipooquKqP4oFAinYXUyU4TKZmss/e
X10s0hnOjoevx19lOwsltRMTliRJDyTd1lJP8k9X7SBud+NFHDIVZDPhhqGjRKsNRdFMu+oEL9CQ
ipyZCe5bPyE53AEGC99WqWrpyL67knX12M/i1RHaDDNbCGB2a/jyR7jDAjgS2tx1fwITic9C/p0/
sS9vYRMotvMLXs+IjF+qF82m3QyuXktKDS0zzN66fUjNb0fjaOGSNUXKxQVYNqvKqZvF35Hfydx1
yoOrKTllI2iFQtszC1TUfGlVBZ1dGBo6H+yEaAaP4aXabqJA9+Pi68mjk7yneBEvvSJP8Fe5DqSD
X5XvUXthUF0vgGylTXmvi1CO5U2HXmXdZNQrym879wi7fcQ63H5/E/8Limdxs2Zm3mVcmNCWw6j7
0C3aCNFAt+DgD7IjQ3M4rsGqohtKwSG8SsgnRM7k1kn6UoCQcPAIDrgGMfI89l/8aDlmWAqX760d
xOH07SrbKt5RA/IR2KXFWnRPgo5/K6k8Y0W4UY0PsGUoFQIHQUND0HExtuSMwbxhpxHYiW9VBLtv
gLyupg6hTnmJh5BkyS2aQK5DHx9+if+k6ll/tHq4UVrM1og8WGasLD/G/gBn7kBkO5XWdsOkNiFg
Uzc/qMAFCowclioa4F4bmirkG19KJq8EKy+EOZEYB/wPE2aarT5uRVTg1KuUqFgxgybmwCpXvWCK
niHz7LfxBtsdjQ3sj5L/QquAsxFfHDcG+ibZ0WFHqkfXwKgdn82wuAdg31qT9rTkqHcLeLrLL20q
BGFyuigvFu6Ep/fXzeW/JmYBym+pk+Y+w28n+wj4v881V1xB69QrG3baTigazzkPyAwPOfFEBMSw
5tJoJ0D2dV1nj15Qt8CgRc73nwGG2/bQ0NdtabSgZCm6v1nHSykg30Z2N02I/nRW1QPbTRSB8zow
WD8PH7AcRLWulp75Jjdlzuk+Qnfqz5GgDUqAPypYbU5gb8oGYe2mPOIOpEZFkoaabbvDTCwc5LSw
ms93nbQ+Qa/xcWDKNnBlTwT3h0BRCbLgSkwDFKuCl/+L1zXYUlPbNh5IW7n3BE3a9o98Fvb5y6vQ
DQ0UTn2eCMqTgmshHTf3TWDa0JHN8OeRlkSbFNdtlaXWXg0Has9arRT8i0SQMptSO1rJC7PCdc2X
GU6GXub8lXhcdGdOzXaaSuExxmll17r5PLMPymG5GIlSp9QCM2XTFKIR9uSazRvL9EX/Wuxvn1g6
CtRdxRwVzLCDU5L1hVgrWSL2XIbtikrCs2FFizXGz+yx4DazaVjqX72fBI6Eq3/iIIIjzA6y5TIm
hjYDs0NVNsYrzGhSjqycZqmcuhhDx0mwE3gNdpnv27Axpt/MCFZW+dKx4td0Y+CryfR9xAPe7whZ
wowzdAjtHfaANluE0k29fcZIIVbQ+nBcK9fAHU3Yq9U//rBHFBAs936XZfPX131zTBNQE6LYaYUp
wMKoJ8j3Ztyh9MCOhNJA1zIeNhIF5ykFnENsFdnkud41Zr/HLeKElAb7lCLYaSf5FYhg6rrXr9LK
Hp7qCl0pC/4dtW8rNdg5NYla/g//YQRPMymH45ksH1/mPHxsRoP2P9deipCArEBauGr4ovWeMYFy
x4Vw4cl8LkU+qypktz+t+V6GG//Ojycr8n5eL7rrsotumCC/WXgiNoen3rS0OJX6X8xEJoq2QMzl
bZ1PrtLmdHWtT9nk80uUVSoC+ScohIpQqr3N8/TmuO57ckA8ev97rJzi1lKWYWkocCe9DOgQ6Ajy
pDb9EMxnhtGYYdD3zhtwDzf49jJvPc7AiSQoWT866bxMZRgc4KE6wzS9cx1gSxzQ0LeXAGKRI05p
OwJhnGNsfr+kAfkqEa4ng+HnBJVxVuMmFbpzJK0yMrhFj3WiZSzCEwhEpcwFYdvG4mhkMYLqxzIg
OsB93GmKme3IcvZa2TAlX3Ib8pKkmQIBOzPmOwaPan6roHy5gNchMSQz9C4Sanp/ytoe/bsturNW
65JBTFU3dv5l0Y5Dcu1QJBprl//hv68fWkXCCVzJvXQazqrqM6UvZtyg0wyym0tRnWQLe3CRr3IC
MojfmM6k/CgErGsE6QAkF/j+n3fYjvF6BsvdfFlFcNDIPcO3cPMdJON+XaFWe2zXjwOxTuBVpQLd
xZ+SiTBEbcc+gxkHt+UoGhekfh3n6gSxUg3EgXmR6L6W7hhJaeW6Pf5NHao7Al67MECG0SI9jiTT
Z0F2zBnFYjrwCM/dkEGxxlfI5TMWbn1H21+WcyG4Dqqux0ZiQoYj88GwZ18djELYa6kIQg6J4Rg9
68d8p5k9+AEZp9/1QrQFNfrDOyaHqI7kQpXn6GJz61T6/TkPBgJMsmNHwrK4Og9O868LXUow0uYn
ucH0Pfy+qiR08CzTY98e7cvD26mCXFYfd9QP2rXr0GcdXJNGQZydzK+mCgsd9w+cG+QP0o45gmOB
Yyqdcc9ZcnoixIcGdJ1o73B3eWmgRjMNO/n8KH0nEx4r45Es3lGsn277NF1eiRbOYVxcSxuC5tb4
t811hAwVuNV6vAV0d6F9nA+lpR1gCsUCsh3S/rVut50fTIRMIfTFD3WeJAuUpngCHNgzxGoe1V+C
yAHSjWXU1Odfufp3ok0S0jQxyUDSBHIeY3Gjr4Mg9AWH20a+NxmeiGlYchsFPU4t32EH00icBk6M
LKQpXww72awPn0FcWB+iqgkMo53CQcKBmmCUzt/Oa724T8vPNnBEzbSDMhNfZLty1uk478VPPng8
2LCb9qdS2Zceas34vT+mdXsHxVzyWRlMPz+guqZDvyMlOmmljPJuG9unzT268OawJfbRHwtK2Pqo
n9LIyY5J712y0R6H1SBuRDDtnVkeBtXLLwJBYRqJ69r/CIXqPFuBkiwWTM9kp+hyU4dfKtvflJKy
JfZxQWIg0OBV1pc10yHDUb58ZYwVxNNGMU3fD/gaCwS5BK0FCLcCflB27HwE1Dtz8ZKPQX5ArqwW
6GoeTeMYXm8q9AxVFACTdPOefSTrIznyxGVc/MsTBnEjvCReaHHXcn183vd6uxInNmsMdbtVcHSh
jM9EaKU416vZwgsqI7hgRXpMwuWibyVrxpVyRjF0wrM5HTKZZozevTex8h2OWV4jNQ8qVX0JCpDT
srjcMd2iF06sSW7zxWOaUsHpI1IkOXu4L19acVq3+IDRABwhKRxW3NK3SLq7cS/BCauwofMMr/nw
HWcGhfavgbhwAQBeguB4RvViHYzlAuQOOHcKTm3FxssDHaSQyxP/NVuZH5a3s6R/rXdGw4UlEQYk
F6g7iYdAECJfNDSLTBPnIquj9Ljy2Q9WH08fMe9U8bviPCkKqh3P0AN8O0U0ZepB+PBete9yTJRX
dSdSy7EXQOgdfSL8W+aZk+erDxPvN4CINcn9RVBlmoIEXfYI5Bmpa7bYIbTRFuC+2TmTSkeegqBN
/FgyFm99k5sTn4kDNaMUJRGhkiXw8AGDbJ+ks7fShBnySuM4bASs1T/QNWWl91WtEamznI+cFvVG
PUIzWk/0+XxW1xi1Cps2OAmMl1j85dkSiDIZQMfhzxTdW0t85yG/ooP5R3sa0QB4sypaGq12m6e+
0rVdU4mixglg1uHlzrZ2+uSt/nRZaPb08LgP56R4fpbai2qYWGvrelNY4opTXBKdXyTOUj6LumcN
AISkkTP1M/v34/YzD4j4WPSJAFL+XqiZmskHPmB7WcLC5bZ24UqlxbEYj0xEc9uQAELS/WFJ6/Rx
5bSe9lg4WpaEw7ClSQDzYMWqsV+e6h+IX7sw8CUQVrRUlcDQWrdP5m0Yk1JA3RGtBIbjESICfetd
dfyi2PW9NuLvHti1ylOcJxF+bbO42Juh5Ud6uYFuuZ7JFfIvm6HrXz85LAojzg0prfC6jwRa0JNa
r0cGwdscxXvnU9kiefk83ElPo6yoD9CJiDLkmeUXA1RFyZvt74aIda3uB3ALy1h1Xi/S/cpULxfP
Loh7DGACs6/fZUV0/n+CkOF/qyATGNr5o+F4ytIDQMj6HImHev4cWbJrI2SaO5Vj0r0+W+/7VTVQ
TrowMRq/qozxHJKa5iiVeUDawBXiGodOX3qypyvO+vasbfURJgcmt0JYLgawFFcJ/v6c1Pdl6erF
zd/OUuwL5Q/arbqqySVpGGBF4enu88Yckt9fekiBEbPpv1t+PTaHpOZTHexe00gwFZcV0eMffx5b
rM3rPxwMxx2Y/VmCnU+c6jKCM88arn/APC6i158NxTyUhAMBoUPYCDDEezBjEvLr6ryckmj2Kg3K
Z/XRxpvoenez9PHRh0HWox8Dh0KiV/zmdiYx4DU1qJoAVc0INv7vg4+oii19qmPN3UxAw8X9MSsg
kKVdlRW5ki7isa2O5mqiY3OyipMpouEfp3+IxaaeXMwZeaY1Yw/GtBvAvfYXf2vE4zEAMSH4keMh
S+nXOsbDd3nvXw7nKAxr5BN4hKlFso35drgar25uTzSKu/nQ7alKcPgtFfz1lUOkB8Kt7aiFvpun
mlgN3XrABgCpykQcP/IVmsazdx4Tr+efkbyHRAe48Nri+CohEEFa6Y2rMyMVuU/3/UsTA2ndE4gz
SbVUvhM9nlpiZbMhNjohUrOYO5QvKCIFBb0ZvRk3kIdK4giFI3evftVB+wacNrYTij584yXDD5Un
4AN9SqQKTwkmm+WwCfs4rlZJu6wwvhXRN7vZ6ccZ62MjS7+pS4rhGOSrA8YS040TZ42o0jWmaCUv
n+KM4ikeTo8rHnw6ctAMEI824OZ5t7vrS6ZpLGfVt/WeI4YdXj3cZSsVsPnozJh/u5Zg5xKj13MF
X8Vq3TBeH7Z68p5Qi80Jt+SaLY1tZ60vLac6a0XpIJr5249MY/ahCTHhwSgzECvMMR3NDwx5pfc8
WOwYJc5iLnh8W3/wDo/fMwqWuzim1kIb8w7YpknVpWCpy9rlheJAwdyZ4NXvSp3tVxxjJecCObbM
rPJUqUpQDylLeT/ZPZOf9oW7Gu8RgjFe/sG79PPMX4NoTcq4DZlPMAPfpanhnU1IhPclYaTvIe+f
v97omTc0HxPqipn+q2aflKmfPy/gtrkquCnz7/vkPrAW+8ss7GKRY6DA+Y1rIGs2tARMGkUd0xCQ
clkY1LVCNwBBMgnaIXG0Yd7QR805+32l392Q64ATNlvu/FSBsE6Q4E8kuQl+Fa49u5Umcu7woXy+
0OUyL7eOsK68xpxIV2tvfX6tIZPmZubWiCKziVmu95xusSImsB8jyHxrAsFzFUJEmfZM9iDVAGWg
gP9L4Gum5ZFfIpkRL4c53+PgR5BPbAhEUoNryzNLNgrjgExFQrgP88gGfwy2+VEayLIx/2GgvrAM
Xm24Yfgqpi2qBwnMQNLDDAlg7lnZ5V/MtYCRIFI67Ie/EU1xvyiYsf+Of4pUF0WXBYPx+IIzMlr7
X6ONHxyYnLFq8MGUDdAMupvZDi50F5pcPXIULMje3Wu/0RQnxNo044cWP27O8cmh4I01sHjRbk7H
SFH3mnYKYQuZcfRqGie1Be020t8pXlSk6ajojzQgfx7COlYvh0LpuvvPuzHvGd5tEKFw7TH6pMdq
uQ4kt2SpItMVcncfcxY+06Rq7i68htR3G+NQMUhTbIo0XBhdBUmRLRQ98ZI40GKY3LGEWWItcVWC
YEdqJGJQGSq7ijfwZlLn8PEeQHvZlVCayoEkV85JtaZk8uduHgbKiMMmwi0H2tloZHbAB2YBLkfT
4YgD8A5tv2+snQkmjGb3xtYpDSYzilhwMuKf0ALIub+QBQpqKLu6irf5HzObmEdu+eBY14/D0Lzn
YHtxaqbLTABXCXpqNI+bzH6K7ADFLtYY2nbzyalcGRXT/sFRPzIgeQxd+kX+lJbd5XHZOodL6gI4
UixbmPTVb6dUZoah6WZztnyjza3uafvVJGZB1Cz+9jIIwfdJ85eyScVq8HVWbEhYalNJhjkawn+b
uR4k7mUfGbxwByR0hvmEXnjY4wbR6euhIo5GYmiVHNhaN/zYRHCNofyrwEaffaIges95BmLaXACy
gRbt0bUJ12k4LNoWyqGsCgpGwSmmbTj2GESDebeULblCI3bgihuhfDLNP3Z4hNofySlWIoaBKkMa
G21AtpeemZMlalHHT9D5gFMJKVaj8gOa5OfjAImOylMAOEUnaxz1l0PpFs7Ot4IOC6HbjJLlxGN1
bIxmp97CbWVj7UegfBdYr1SExNyiVcPf5G6gLJcPvn2MKAWrfd8PrEcmxqLNq8bun0Z1/aNZYVfB
Zq7pfGZbjbcXCggfi60ZDyKZLnbKO7g366ZHQkrEpfZAPK/CuG1/DS5PZK/+a9rwYDdU43i/RChG
hzPLy5gQK6z6Z79ouxykOewaRp7Hj0OYntGmnRqOX5wWW8swDtuVH6FoBYetVZrBRxeFOzNYGWqz
In4+rwvD5s4opTm0Ro1lLrbClfp15Lv/Zaze50wYaAvRP59Q0oICWKf6rxSWUSguaihRNxMaO2cs
f42tutoMK+lq2O5aSCTl7Amkf9Fy76kGg1WFzhjTPjhH/TPlNKDzKMbHSDBoNgFxD5GCNrymZFO3
+0ae/Rp1Va9BdaMOC2NT5L1ygetZ3IbAykHet1kyRiS89FHgtLQ+sBV0dgbQdbUX8KW3ZUTE+0YK
XR2PfTv/PCaLK5zpiFmoFUVSOQrKmvOUhd1SrdYE4LUPICpvcFjBGpkXxG63Tht3DGpomEpTIBi9
kbbwPnUv+tX6vu8s71c7Urv+m3uI8YsjtsRB1r5ul8oomXuxo1p1A+Iwx9FpJLXazJEmgxoOi+HF
cc/mNDopFD8JRg3GLcHm/BSBBgWzLLIL3t/bE5JLLz1DGGBWBBXjfMB+4L6Gwm8VkxxIAkxZDtRV
sMuJdPnGtFEcCJoS9Ff4bMbW5JYWaZc4U1nrZsf3n0bvi8hJliBc/tqQ9RDLSC883qcoRpE09t/0
1mEpQBPFNxdCVBNuY4VAkXPLeKHgJHFrRjpc94f9WWRhqBH9v33PfnrCb0/MyEtLc7nux+NOqebz
9FUzy9sx4utAmwT9Lid3OoaHNOAUD+OtkRb+vou/MQpfGmTOc0hTsJF+yHGfK/MIhqiLU1B+9Ajz
97EeFGPj6ThBNgyN82oHP1k5ON+l18oN7KwqbPmMJYEoX8SRFmklwwYvvUT+2JQ2YkZScRn+fziU
SAmUR7ZNNFrnjzPYTNu0c20u2kT+v3Hciozgchxiq+0DjXfkKCvNLcZTcwZ9W5MZe8T/ZRYSEB/m
2p+ZI20k9wQcuoxyvkJF7qdbgxEhWEqcm2NKMxgGPlHxgW8Q3cirlU76hEOtPamFO+h8LKEijo+m
NA1M4FWpODsV7nldeMcF+QttHj+vh+QN3FVEAfM7x60cBp9Jm4Nv4z80lSIGMFUJ2/MQw5g/g47g
UzWLhWN9Qa6HqpeLdQj2IS86LkBvhWnNyTu2mUf4+QzJpmT45cnc7ovPKQoNWzm3OvNodsFyP2eg
keJ3D+wT0z573vdyVKTFs8cwuXa6iuLP/yI6C2u1I+rdAude9TipV2mwjxXWP2E2dKNZcfxXl8EC
L6P7RT3C1U1qguzyUdlX7NPbwBKLSvrcyiQ4fktmDlS125L3RpeVZv1K5ulThjZjAJzn2V3jQ1xz
prkPrGxzgAxfG/PvZ6X2+C8Lspd+Lkkyz0WRgb754pM01vCAjL637Rj+GTf6NABWGywGT/OUEl6C
x9MEzwztWqwm4paERb44zGAxqvzwlThFpgGd9j3Vp/T8c71fN+yMDmSEpC811J0QtdV07K83U0Gh
tdLTykkf2xZ2zyrCzK0TdtIrSG3zEHizolfbncUADBoefe0c96ePjKp4Lvr99T0Ptj0z2rVi+YDb
gBJ8WfvdUxk5a8X0PUfyuf7xugtjMI6hmDABD/D+TJF2gKWcQAzS1uz12fEZIn2no2rA/2f9WISt
YqmuWz1bLq9VPJm0lqSlX+HCqvyPLNZX0nHTDAcGEUgqLXWtASjbOKGtk33HxtRWj56Hf6ot+v4u
op2eAcYAf7zFd9S4AY0XxC4IfGYdNwwJm//lvldLx08C103123z3qIiJrp4IyXgVauRIrvCvYyGB
E7shRxw0yCMKi7EGLUcypNpzsn/5Yu4feSXJetYlpk1MfAhB6F6uCvZPnq1COOI/g71Dg9xPON/L
wC8YTrLUIKvM82mEGgx9Qygj1bIF+FgQvFoLLuFyM64D4OGtS7JjlPuSCzdaa/E3OY3+IdTbhD55
uAcvQwbzMVRWGvVaCXM74nGoaBi4snWS0Vb+cxG18FrjK5UcWw9NkH6CtzGQ0qwS9X/kutIlvrsc
DnVGYq+iyKQRLtdxZ2HgQcd502yM+GOYzy71mQMluLwlom48QdvYxmGeE7ih5pvqj2mGLD+mcQFj
+qcm4Uxm/L4P8cHUIsP9ImUC3FSeJyXCP2Ul+EjySSyNxDAwZQYcXEQSwSZ5ggNQQe8BWue0DSnH
1c52mf7TDVS7qnBcMs7FwIJii08AZaMoFYxl81yELlmyZtSByn22qOYK73F0t1ahJe7rKzK/HtUY
VV5geeWwvp6CW0i+KfIjghfDaCwp9S13XHl/apcBrQqDH/eLBNlFn1T6VPrJPUETwpsypvFmLB66
0OJVYP6lPo9lWhY9zNjbCnKUjeWq0oqGZ/eEQydp3HBh005cfbxE/6OSzeDYsIrKv/A/P/yGG7Z1
Gc7ddFWxVyWEclmGANzPJ4zIr/3lMwapn8g047PBeK99aWwsglo/gHTbNC7Gpn99lpj+UtHaQtpM
cQY/W0pJfI1Zw6IKaTAeDGfsRUH/vnGwJYohe90DLM6qB9NyVIceO57lB9fpPVnX4YH5lzImJkpK
4tYJ5mRDbF+1tifdfIQyteFqKhG/8FB1KW+CJVdidaYg3XbelFmdau5TKF9lXIkN8CoOJXJ0fUho
JZuuRkJ0fKgdWWlz/5ZXdI7+hkC7zXLz8QzfkL+xsnhkg+RDYybjPNQZgzVmlo3Hz22XxTJ2VHCh
A7J08jWCykLza49H80OTdyUJbDfOcF46SlFNBtU4wZ1vGhlEa3n2OdNCv1OGYcHYfu1UzywYPzSK
dGkNRBk3kyy2EsdaJzynXW6RDEjCwU6YeQsFogxM9rlvYHFoveV/KOHrenMcYNvaacM0/ra7npLY
W/FIYkrDA1iSND7vQmyvUEG62ZYZBoOeDF2peDKeWXILrIsPssBIhGQaHdSCvJDjB9KboNKCXA6a
qCzq+xCITk45j9LX9wYacvc7eOOiV0l28kzM3kTCT7NBeCVlhYNLR1+VaVZK4iNK9m4G7k/fNP3v
K9k7G6Dm1KAtofs8tJP2ol9k+AVx+1izID91HWsY5f0e58/YjJYSLBnOxAd5aimtuMYl9kiysuyW
Y/9AGyGlIIvJPDMjh7xt3nbi6UnQmBQEs9p3x5RbThCUuSEORxXBoc0VWo/evnzCmCK5H1yC5+c6
gS5ijKZCMeYu+PtMU/OaqG7oh5Jl9MEF8m343ssAcFC4UXdWkArOH5q0EOKPT3N2giYdR4M0qUsk
gg62I3mzBXH3Pj6aaSelWAbHC4hGhpRuftQvANVATfMcgnPWekDJWc/nN1hQFnuf2KmMjz3BXMW1
3X9V2lDGK1pOMyYhMbHAhFfkyD44SXP5ds22uZBuYzypT/2tSBuKKik+aE5oWJPhP1NlytyB3Pw1
PsAD4vIfC9lI8fG0XzsurFr+ojt1Pn6NnOZyevv6fqpCaniGkmwkNR6xy7AO7O6JvXfprtZUZecq
wTU2DhVT4cxdAzsUx6NG+JBADUG2HFlV0eUM/oBeNqDFZgbT+8gOcAIc0tyL++aPZUKcS4yw0+cN
839cQkvnwGjaS+w2dDXkHw9tK+/OfLmoYK563vIapZBSWf64sgiofq7iEMHH3cjegpi0nrXkWF0x
sMPjxjfomwthAN3ApoDphVsW7qQhq62Dq6MF/yXqE9hBQLdNLFxzwZ5r+biiJmjeRmj6PRb2BS1a
GNksCBgUBkdWNCKzDSHUhDmM9RihncYMxCtzOj11PTyv0bn9ZsfUSbnS7AlpwNrgUchU7/2F255m
Io1XKjnom2jLde98Nm6orE3Ai0JBllv5C92UKAW1YSJYzgZWic0FqPfCPiwEAqtdN03bmBptyuya
wR3ZidCyihgKNIcd78e6fV1S/d4hHmU4dOdsww0rmTIDvJkBQoWwYH3PkEnyYcWhhUujN6Zvt+U8
cAAPks9vWoTMEvQgETGPrXQtQoEYCWCjpwYNNaV8wrZRFVlncT739dZSMkQHv+GvQmcgOtKQ0E8P
YsYI2trVeuFvZBa3hppaChPAVHCEIn+jd9anGnQibIu5JOROkjpVQitG6lAK7jNQfsQQYl3Fd/Sa
k8dv47lMEeeciHIAhJV/8KPHG8sIr+co+p2FA2b0ThioCdefolqm/U1hsxH9UMTFqtHPv3824R0e
Oox6MYqZvaTP1uSXImRVUtnKVJxXcZRAcnB5yLTDpFb4C247+6Uu6DOY2NQ9snAcySwsDxVqUt92
SYfpjxpDCQPpefuROBFIobX7YuXJG5wYoTlu6a+t7Ispk6yZjQZOfKqQR7KlVOcOPthWETRGjnMS
H1NqysoWi+rKge73jtU5y991W1GhiVDWfySj4aUgdX/ujrDzY5U0gdSzRcXaLSubAfZNMyIYPB0k
yB9ena0cgtaKBcd/Q2jGYLj9ErKsfGB/E1PzptzGwEKDxjmqEUWTTRsQ0X7hk91cJnDivw5piI69
/St7Qm1EGXPO6paa4gapabxMq/mSSFJp03MIHPTIa17S+RSjZDIkmePBzmtZWFdoBwCUsO7VVWOC
A2xDrLxaexgwOVsGyKJlm0ndxUF2VDyQbYCZgPd5ni2GOuwSngKsuGwC230yo+DVF5OyjVbng14F
VP5UQV67B5VulBg5qMstZmF5DPFiB1LrO0QgCB8Bn/svoeseG0H9Mt7Y9GXoW6t+KOvOIYpJGOvC
BszlfUoD5JUlWPlJnCU5eEZYvFR2jFoecukka/qVUDwxxB0OqGw9gpacvkjWLM9SGzWijZL5AOX2
JuFT0ccyPYFfThbkMl8GqNrgpST633Uzv/yjkaG2ZZ6mgPs+4TkmSo963lA73me0qXB8rACyQpRz
TprkJJERos97ZjmoTJAJTNg6dUvJA+B5aBIYuOz8NtNL5ObfdofVQfmtzdgarzfI1LkonhUsFJM3
w33mkrLS7w7JCgjOVhVhMnc/g93FiXR4+EQS40sFGNUuTfVAP/9X82o+HCyMEH6HjhasQBtDWbpj
XU/E8IQ0jF41NobUtE0C+FrZpbFrCnl1ZlKSezzCKTEVWTmxx5R0BekE9qu8jQNW+Ma17Vgy0mPP
Wu0AH0/zEDpmgsd1WLekgfNM4zwsiwpE7OSBz0gjFDhD7t6NTP63UyhvamM0Bv7FcGwkwZta4pym
A0UvEVANNR9x1SPIcEGDdRkpRnjdKCbgWwsVP2w8M2rkYRNqUqO1otYLGeL/2M7k4btqUuxe2qDL
EAJpviMTwmdACnxO4Xfa+e9WLdskeWRMl+PTBplB+ugmJeSkkDr1teocUy8KBuV1BAJ2JoLumDwh
boaDP5Yyn4tXuuM1FbncpwsUPewwWCgxzrZ0Qr0OsQYEObR74oXhXFLWV6YkFi5EcipD0fywMssC
NYNkpheItOWbDYHFWmYehmE0UNkUANKUWZ4Gnm99oori03YGInwVuvmrMb4YP3Dam7lvjGz5Ljk3
PPTflIZe/KpPn2EmTWPSjT6SeGX9gUorG3cP6j/lMtPN6ywYh2yZfgcyb7xvhlGIfTMSBmFqH6Lg
iy1AJXxkuqtkIVy3njs0F8fBHSq4iU2f4d0IjjVQnTW2IH4BEBcQTe04AXa6hIZsuf1hdNP4b8ms
e+h4qQ6bFI68bUS13JfdPDRwcqRBdvH5UpxMIsVt+/YT9FAdYE6uV/9ft13yU8ueOZRGpcrI8c6i
MaHXvT+frFsJ7nj/4JJu7IJoq8bu6bBFf18y1Ga1rn9Y56ftJDmlsK5xYvrPTzhCD+wNBBHtiM5D
rW5QktdECpjCqopSZvgwRINS/SXMXmNiugcOmYCwdQSKKaeof52F1xH+R/T1/haY6K4/1YdGdvsn
qet0syf9z8yx7mK0O8GIOjDIh7pkmXPfzBfosPPIi+xCED9TUqwX0zr92DI49dxod62xkMUGaAUb
BQIu7dIFmwFno757bzTwc9vih51Y/vQxliNTYcG3JoVwHSzGozDIvczHj1syGxmK6ZAKHJMOG1ca
G3qCLynD1xDNDw32NTMZ0EM7E4dmQDhRdCO/RNMZ6m5FajBm8z2jRXHJa8fpIQvKyD5gp520/3Ae
KDthh6g+XuGTP2lyLFmCzbyH65ckSWiY0uQduvQmahnDoW6e/21G/At5SdEyhrYHNgie6lFrNuL+
lVlIH4DYGqoePz9Y0kg/ddLOC4EmZ3UOjVA25M5CmqBZZGGjaJCtGC50JPkvh1hFCuFuRRjsvaTb
fCVtgvTAu5Ot4bkjauYMJu7j5Y+hkTI72HytLetok+UGIvEyRRXSOs3sUckPs6g4xlPy8mU8piBV
pItXuDk6ULE6jB6KGXR92KDHFAM2mx7m12ctRuwSkdT3tu65edZvk0hO0aDG5P8/9vF70G/fWb6b
bOdu5I0JN19BgRGtyUGkjBbgQ63hLraM/7QJ4MLvoQJv6czKAGAIuxrgG047WY7P7Tvws6XPgUmH
4hSWKIOMcxNW2GZuM51YjgZ+sRLD21xEnQXhLIMX6dRIHRtTHTZOHXTOyzM6BiuKQzxZFZ7Roh6I
gwYXpT2kg5h4E58LCq1veVz2xhjkSC2UZ84C4gDaWVrFmXrE8Bch+wtB7Q6aggtbAtEsfCHuKUHc
a+Ra2qJ6AArU5vyBSYrh8m/SKSSSih6WihQ5ZFZH3aL6tcnI4bwJxKoSWYKal+7lAKCn9O3fJ/2q
1i67GXRjDgBCmlKLP6uVdOhQ9xN4mOE1y+n+FLPKpv4DRYVBk8WLoIIQtijkyxMJ4k/E+OmRSoXk
CTGmcpAnOuGt33ZJ1kCHhjTHG88eDwx2wefFl6nwgNlNRQPUMsOrYGYv+oBxDP3jPPMToVx+z4u0
wjB068ymnQwJBPDumulS/S+47fKulrFLZPnGGmQj7aDfNNCkuLjYzYolFMQIncsac1yfoEe3nYi+
8dTDwpR7qCBHdZZ3PdqvRRgb81r7j3j+3ktr8KKlEszLbtgxYgoT8M6GIvhl0BAMVKV+4bXoSm/j
rMH/X90qMCspP7b72cwNin8nfklXy7xJyJ4Iuacejao/Id/C2eX7TjpbKSpdzJokqGxuRy0gMgmf
lfehM9Grb+8Ga48xAH6D22wymAMOCX36vq/nSrIskvWP43eanl33gOD+fDaU/K655lZs8obCQcmB
Msd+23FsUT+dscbXaCPBjvlwS3eLxELe/mK4PV9BrarPFWVWo/lGJRmXZfIm8ohmAaHbLeGhZPlv
rNzHN+p4Ez3EXoRxgZQaFb8K6zxkszbz8yarp1Le0a//CzPeyGKGDDTv03aHZhpYLKir4mEvWVx9
Z++CkccuhJWPq/xXypVQsACjO9dgjm5K63cjkNyWm4u/2RCpGNMcoKKBz8wGRTZ03wKmd4DgcUxP
rQu/RN2ULUQ84Y6R/o/oF2a94hNFgixQ5Uj6SJOouX4uBtjBXCJVG6kizt4ablvosKjBwZ8F4+Tb
GReZNoc6TiTq1IuHVZZ1uyAWRzdj1WxxxSj+FAjJg09Zh0FNqyo4MmEgaU+Cpu349av96MQZsXAH
SYLGI2lPpuPqeN+dSDLKucPaX3EzzgGVCMgsgyPmwjWKuz1eQB1pSETNhNALNpFRb7J0Se6ApK5M
Ys9o8ioen/YutN7NvvoO40fRwX2kmAL9RIFsoCduB51kMdzCFPO5PdtdEbxQn2wFbSsq8aHH/7g0
+1+MonRaBKs+/JdndRM6ST0sO5IXKzlJGELSyM8v23u3z/5zqkGr12/VeIJO0SxGRMc2Pqg1uKqx
v3bVugHSvY9Xn0IYbaAs4s3AFJulj97gK4g5mfpWIv43rWtF0FDcqdSjq8lTJfkECmAcnxKw3IZk
guJb/ifS5uMUh6i5UpqRv0zKwTBsh2AwZr7a9ulF7PNLJOVed5/pV8d77LPpmP9fRFhlNY2SIqq3
N06Mqwn9jFdeZeDXTSJggkQCSiTviq+fyVpMheHfKzyjQPA+9ZpexLjrzQxoYbs/jb33R1OG6inR
YSPK2n9b41cZ8pdWS5SIWgZz9nsK+48F/iHzg9xbEDUt72MgnuMBJNMvAmYXILdvD/C0/fsGO6Zn
tbaKRfh3H1DXPsA7KwQpuosbaKdNo2kocpYyB5B4D6mw8RTXFo0Pi16cbxeSQlSCz/TcwHWuCCf4
142yoEovgRCDPFPu5DpSh7SAUSqGuHSfH+RjRl4CbvgUV/3uA7MluzoM7ZhO9qdMhlfxWKxj9Itr
Oi54fSoEpF3jRxAy+qfo9jwvVmNTjOOOROUezlR41O/XOSfFiHsks4B0TNv6nOpEHnracyWFawn+
mlmZDbmKvbA/hKS4fRELMkZV45KW++osg8+Yqp65EJetWe/Od4+MaCCPi97E1/xgVezq6Bo9wFtQ
ZCrABfJPJwTfYoxxajnZNWdhvWzhopmPhsY+JubFIYy3ZvtmOQrW5VdQBskXxL8hFWGMmHRAgRU7
evlG/ahahfW/o9raU2YTr8jumfRuAIyzIiGtRxvYeKvbjek7c0e6peT1CmRNr5v/rIHqo6WmxLAL
kwTz6jxtD9U+cL8B9Ycpqzv2vNyEPPrzqKOh/TMn7qDEYI5FwgBk7Z4Q6LukqxNh+8EAGMXlk+MH
LcDF1lAWEQcCrc28TgC6QDQZRKFYIE51dOLS4UKe/OzXH/wIUjg+35jvAGwCVw+zgAj0MShO1Gtj
ZHivFwmyZ+Sx62qBL/WJ1o+NlZdWqqq+sjdZdfvPpbYOs8BZ01kK1A/13d5PVKLno7m3PVqdGUvI
TMapw12vNauOVLxxFMQSMMoOfwhO7S2/hB7vKAyb+apSpSuQTV4DGstVcYVYwFLFUXBk9yUqjKxo
QhegHQmZKcXEtmlXBHFcEXjKC6R9MhfUuooEDTdD+YP2/Ur1wFdoNw98+trJ2GhqGwINXIiBbxy5
K55299brEvQdX0gw5g2VX7q7+Lv7o9WUzCXihcusmO+QCpM1rjRywSq4PnmCKBYLeFW1/Cqad0Od
+W9gJ07IHkDjPVoNf/+GK0NkhF+hp2jVX1JvmHVVDKgeFSe0y3M9pxHHEc9nGoaxCUOf/jsNDMdE
8zyFfFDNa733gqw4qwZshYirzmIgNepbUljHuegvkAmd1GuQsAOCotgBt0Oqr1f6zjkxi+hFv97q
rrK/8q6Q9TPqqU9tDnK7vXuW2uQDWsFgur+5XDn0ucUblezYVHI1kBENEpi+2MuKHAtAQK8jPqV9
KSSRug9iN9pwHQ92zPQuVRGBPBEIkGirJBWLB1KWF1doPdYTaS728KdGyVgvWEpT3mD3AyVAF9/I
7afSUM5pkfnDmusiWoira5F8K2Jq0QqwBu+MPAsv+S4xQT4HWb/Moln/Nb7A9ubKPiVxJPXsMbsV
hNb0b6DJjQgfSofR5SmC4yoAsIWY4e5Mnsmf7d/e4GLb/J/3mKkxnWuwspTZLqP7o8+34HsCdpJm
X2+k8fXC692YEfIgSA9IUSoEh4gVTRdzRSHoMNwmzSbjFQlHXLumpNZ0Rx85nByG1QMlqEksBrDh
FAjZ8XJi2cEupGYG8GmV7ZEDYOYOtTsuMBJff/vYsx6NdV08kDP7qjNdFdyoS5vCY/ax12lLoXPf
xAG4WKVpg4rJBgTWYIpLlqozEHmPLPfgxIqsEBtFoYBJDm+0Xllzk/f1hhNlaztKL37v+a9e1TsN
vrU+FmzLTdTy8WdSxSX320v4mzkjEoDfvD4d6PyBGr+FXRECdp4ny4+WICZYmuxPmiJPLQtHiZzn
9qxXqdtkGVr+XYPqh57T+lLJzo8gS6hwWI8queoU+C/i7qt/WbMnLSfeDb9J5dHyMNR5Y2tA5HVL
S1P4RmvW5i9WnXweivLD8PajQpNcIPVZkvbXwbdEPYJ0az9QFZgIgU3jOi68snLwDw2KGauOpcua
qT3Jx7TzXf1pnfyA1OoCqJthIDX6ez3ufe/i2Fy6TFMAgR0AoxRr+UXS+CRCksYB+0XuuZbQRSbF
NJ81e+xla7Oyjq9ON3x36dDKQLeP39hbxEjdUjJl/0AnhDfI/SI7gjMGZZQ++HOpBI4anJZThM/C
RI6ekpDVFKxK/at5v2LbZlF/WKVkTOvz8C3WMcErEJy9nWY65XLoc6zCpxsZ7CTfEkEZKwQY260j
axeXYNx/r3zUKHOtgM8TCu8bPR0gSVxRxg2iWzFFj10Ee1cvD1eL45rSbxRg0D+11GQajebBnhKx
7PRmIWkEbb5wHmBGvSl2jyfwh4oreuHIXM5Aqw48EKfFMaZwCouin4dQukPwyZxtszYJ6QQbDN2O
HpafEcBqdhfnBDxDB7Kic+nWyh7X9q1Hy6ZtPAaqmazQySoFGI2PT257kEWFwOjj5EUf7duLMHOa
YMr1KvFDv8gpP3+kKsTJprJjncKOdM5mAC2AGmHm+nNvScXLb6aJsvXxgwfNhrOu6ZY7726p0kFY
lollWodvX6mIbkrtZCx4UNmGGCjjSoCAthKEZ3cX/rzl/0i5vHcD0UM8HpWvIiAV6BP19y+glyO/
wcaRTKLemaNzZzjV6tGtgTtKB/pzoj4AG7Y3OASxU3lNHWc6TqXakxzZm75brTXBN7HapnlSiwHm
U56bhOH/0eB9W8AbrLcSbpXKesC1ITMcZwm0shzRbzqlEciFu3c/nArlbi9wSOIxuwaaAr1TuQ89
6mrrnQzbiYjOufMsG0aI8TQd8tdGIp3kdYEZGzxGzhr4Kb1bck90pbUjy8i5EW4OMau89Oii/GGE
eYzDBdtNV2R04XCI2+16o77Gl65V0TNl2bvv1Qq2ZZBOhuzdtE0Gq+KzDN0cYVFxVuPg7AenRO4Y
LRlsBh67K3HS8gj6bOoY3jrk3UTV8tOO9il3+9uU+6uqvzB66DO1Ib38a35sRKVIYbFClVTti24P
F7Ob2dMFJgWM/Xy/i+fIwOkj7ABob6X8o9DLHq8/OFx+icX1KLZgXTH2gv3AWrRJTLWG+HsLWpu9
hwzC/MYpyKB7HrYtkyNeFAZ2mi6fk8EyAQmhPP+5ThOKkRCyk0jek0pgsRlKnBKDuKkzFiNI1Vcu
ft/MNhjDnfy7GUBsIirWD7jnpAFVxXCberqILpAIuIXdM2/gLZlG61OdHe8takgrqaMVZv2bDjzz
1RuC2s6ry7si6FkAifw+cTeJ3Nq7tosyLq+priNUugoeqzopmcjPrNBDOnyxQEjVYDEPNQ+eHRAD
pEy5xOvqvjeoKv6dExYgptuhJ3eDxqCVv5YYGECSgDOSVdyFsyQxj83/+dNRV878hcsAAowYlq/o
mJyCUu7xpxVE/h/Gl6m0moaZPWX5I+9mvrgivRpctveV5rK3oVwsqLP879Xye1x9xFlcx7OxEJ4y
FY8y0650j22K+UDEgBejQyYwUMVUYkdAoLVJsoZnmXQmJ+X8L+BxSdrI/I2uzvHHNEgjrPNDgMrA
WkqRcPNYmjs/QZS8G+xMUI51VLGX9AsUu9TCMZHm0mKr28jMku+yCqOXWsrJcvE1PSy6DfuWqC6k
wvE5Ko0XNO72zUR+y8gOf+5u8e19HCf+oZa7qb4noMRkEnhwvcENLamRVcZnLkC+0qHHJFnnJr9b
J4bT/z/6hVHVOiMmvIsv7Wycz/JMTUCoOA85iXjwXD3l3cy9NAzJWHvSbe3vkAeD0eMHQ4lvqGdD
NcRxyoxmSIqpNb2M45PqaiPJAI1ikQVJGPosovUUPvSun0rG1MQZK/17nmhH2MH2yGVEMeanpWIm
3ITawloIQNAg8e08RI8Vahmh6FCI38EkV8GDZCRXdeSVBiIpeu657VLKFcfwowt5t+13CsD0aEkI
W2WRUkygNpmtkprh/7qsyvLQiUk12INWR+BKSJTVk6eZPFiHuO01CZcXi/LUQ8dHvz5vFtqFWfHR
O9RM6H639MRiHHWmCv0LNUjIw3rDq7uj2Fo8T6UfwEMmTjJin5aiPwnNZtEkSJi6rsJoeMjcoWs+
JMWTnjCmusJGC0rskmk/ne3nJrtH9rbbOqAZGaDkCbmNZ9s2UGg13lVJDeV37nFpzJVjdrId5Qzx
qkjdMzO23lml8Pzmro0vllK8jXJxLCEbaCwrCzG13/z8Xfg2k/ITt+kwG55zSOLKR8/JpGguWKiq
POr8ciOOkFCagpymr52SbEmRPX38QrCAjkK4LYD4z0Dlx9uJ/NvSnoZsj8CMgq5qWoC2HW5DZ1TQ
ei3wwgUr7mehCl5rHyC4UsPwx8AGDBAvpGmu1xLSnvsAVKz2Y2OHtalKVj6gJSAgmvfDVwo3rore
zWGOUTfwRy7SRn/vhcPH8TxD2S5NkU8vvCxJ0myjiVP/NjdnqAkdqygQQwc1pYHRyQ/LYe+ocXsQ
/vixISytL68cbstE4rPpZZuC3GcQnQNNXyxNCaRZ0JSTgmufafmbJ69rcHLJI9eelAIuKvrB4xU2
unxo7l+wbKSlzVCF6F7JwlwFlVMMGkWdZLOqpCNiJDiffZaqnjBTNiQVgea23aAvsowgZgS3QWkj
fh9QHK7kycscZWywmp6g1UWRRsnTmQCl7D3rT4YNE/H4NkKkQzI7lYhZ5Bpu04aLiKLm0iwTU0SK
dAoHsr6xBajW/hbnAat/qLFNIuTxMvv9eeIoFQnU2H6CcnuZPxceQAJ71oKoNCrRoVx1ZUJTh0uC
icutW0cxelykUddTADBMwhAO04Dp47frEDGtx/nZMYdkOrHkkD7Lj051Ne3Bp1t0jfIFD62PnQwo
V+3cHudcwraKp/tSNaSYmySJS0R7iRiFeyyIo2zfR2aFED+ANjPYGUm5C6D3enelYWelHb13NGVR
cpT7gFM2XG86K95svU0GT7TfdVlNXU0i9eVrgL/bxbf2T09Z+tjkAvQIULb2W7T52pLiMTBDJvnZ
Ca5eOmE1B47eFu4QnRwrUAQH6alg1kqLo+sM8IpU/ANHfxcBI/kbJjjd9hDA6wu/EnE+Se3I3mIg
2FtF6dAVt/bqI4bJEZQF0iLJVQ9wpwMlex2o+QVt8Q/Mxmjtz7PDc302s4HyWnP9LAgCoJ7VMh3N
mJCT/A3OjJfOHur/2/91GV/qI8miPa2mJ4SUvABalLpsbQWx59TEBNoaT2dGU2H5331PYS/jHRWC
B0A47E5FPD3Z7vsVPHcPZtdPQFZ9KKZ9UDtdTfOQJcmOnIi6AyJepvfgHBCN12yKRXnbipHJj+Ts
nyHf4H2YVkUBWB72QbhHsndVtHRb26YTh4Dzs99lPH9MScs1MEp9Glp8dlAa/4Rz0AalfCXgbPf+
Czd3W3UabOBMK1jjF6Bc3P/Y8LHWp+QLo1MTmLL8vtFB5DtdaLzpDsOsfCUmEDXXoxijoo6cSRur
uTM9zJxnUn1BUE3G9/R8Om7v3gilxhOiaS7bubdcVBQtvd/v9AanfnUNCv6B0HBYTqY+ean0PpTY
JVYaMOPWJekwPyptz95MMWKKuQck4pMgmlxZXPp9NDvk3M1QfRqJGGrUf2XLZbrL4GXIXkG8ncSK
bfRhtGCqD4Fmh3Q8kzgt2mwgNL6pUKSgEYIPkJv7upYVDUNZOKhsiF8d3hEL7DQEhkCTHcc17Rh7
uTmK6DV4P0BnpxVrbv6bjskwTD3msn/5KnpSiCdpDcGUN1c83SsvHM/HhJaSXs6/thVwBQfH9RtM
4SO8YZxOncpKuePkUfaBGh6uNsvjtJXjDmW9R1iSTypJlXC2XDDoKEkao5WvkQPXRUIaZU71P7cT
airbxuMIeNyS2FYS5OpvBnVGP95vC2VQuB63eR100FgVkclDplp5quobsqAQ3wHnpXbWwUXeOQgt
IDpcgx3c1xd2uJKGh+U3qJWJ68ihV7jHc7rPKNciVWMb07ocqi03orRNTXkl2+Z/7abQQ+PCC0Qp
1gEYzOQLtHsMkjQSdtrxo60NT+hcb+snoLCv/3pJ7RculGcsjhGcG/9PiSira4scJfH3mbxhELHI
FxGyugcV2MgF2zSV5SiP2e8J1ABwrjeYdv06xZSGtfJvP8sow3A3cGb5WiKon06FqILu2GVkd2hN
BMQY8XFwB81PILq8Z9Z2heomOZ/EHOiGy+tqP4tr8mIX+UczT+f7HTE7bYq9O6YUagej7BiPzOlu
FaLed/vprJ+AxyzcMja6zSch/KqODS1QvAIo0qxbcVj20ZjsUvQ3oCLksDhpK1n/XL14gnFLwtIy
k0uUnuoGbi+IuwpMnrQl3LtICaW8jFzv43/9sneJCCRDAvzUvwy04zVEZ5um/o08DFFdhaYLjPqt
vtrDBUPdwZN1qWTv4U1e8hJP5yQmdoZ/LbwkTFkexWiumXyRGv7MuexOCe6hTtRYZm+wVFz+iHLj
zqoKjk0cVpjJWEttDCFRGK7DJBoLT7XWN3f/CaG7QgiFB9RoPu/e3DW85VOLGR9NX+8jG8a2aiKF
6z8ibltdTDB6Fn2oUq8KuVXd+syXQznqHFC6ZYbhKAKpgxKOwSx48+ZTAZfDznBGVu3zb58GFe5F
KD/h0WccksIMPXBuATcDlR5GNdqtyK0zih3c2qT8X4mYReSeKv+qE8XTnh9Di2+3LlqnkaCvzJts
5mLRXnpvBPk/sIgIB5rPi1FgqcOyNDQu+EMyAdDfaPIDUz+I2rCBcRMBaBblWGgsGieYP2R27pSj
ZiIwP5oqfi/bELXlazwpGpPxJZwgFpWrrFsrK/Mz0cFfl8wnNH4QtB4wS7MZ/pTayOzbZZwqyhEG
47zQQTLg0u2Ysif4yRlM6stroA8sxSeoVpq3YiTeo2HfClPWOLYZuvQotyoCTSOhXPCpGWo0nKRB
DKwBIsfOmFdHy3TFtpTk3i1rqpioCoVSYaC7ZkRs9inqFrkKLXtFulrfGSWeKtBpyFqEQBAjAIzj
1LQwzmCy1jTSyGxlKpYhIQxjHF0MSoYMn6sWmuMulr8SuhjMJZZypv9AJ9iJulzfgsmEBDFMX876
2LrrrGe98q+yDrne5y9Oz87A8sHM3rwziSKqsP+kWoKSS8ETmmzl3DD3iL8Auxa3v2ETNRwrSWA5
bQ97yk3kLUFmfk0kqSyCbVRvUeSyMCSK7XSm4ileaiN50Y6GyqHqKadW1YoJOkuNAnNBrulLfvbR
Kz5jxeObVlnAf6KK7OoK76SNeuiRMlzt32aFMCjsVqL3VwaY4tuIUM17AClgYScO50nFHqXGAHOz
0PQtQ8/UQZbBKpqCohVcbZJeDdg8iYFrIH2PGDxJmYP+zgoq/KmW/OvuFQ67f93vzK5mpi/a7OyO
XUJH3DILC10drhunxv0qVgZ/1SW6/eD15ah4vPqvlEr7G4KakltlWr3uZW/u2fCv4owZJK4UXiOF
h2/NPbdF6PV+8gc06BOHQ91qsOyT7SIIAYMyNZttp1FyTTPBx55/DtfI5GaKcFGQgA7nrVY2zw2B
a68brFPjLSIRAvQGXw9WDEk2doSTUbDL5U8XLV2fQJxu7Qch2wUw3O90Qmy/t9ZGmDij04DFGFP/
QY0u1Y2rTq0F/3wwYbYDsotyraQZOOpb88KSLcRHd8t0CaldR5/hdReQeYK9H5vYeS2H8b7bP1PM
L3EZqma7K9R6L52BkPBofOxZqSTal0WfjAa3m6OwflYhqjCVzJAU63pNR7XqXRCc3suvfcRbK4ml
m4jd0Drs+IoyNwO0nK3uVA9rwz/Ao0ijGn99s17Oo1UlkcDSNajFT332nVyFc+pPY8FzgV3Xo5ft
WIgEOS9deNm8q831tacAFQKfoR2eW/kQFZILczMjR998ENxfgkGCX/dpSmVUrLBy/aOBOT28QJMf
DR25o74z37FHJ+cv3CJCJKAKe8C0fzU93tn4r3MC7z986BFlfxt5UFcHTJoZkMdDTq9DNYVox3lJ
8hHslQ6jycdBwqt0FLAelqaNsDwljPrvuAvvDVER3c4jz+3HGEyOc4UHAc/yBQnJqnwFkCsHQww4
Vpsx5GnpoxofPjocyME/D4pqS2Hg1zQnzyx5rOiERWmZFHi1N3UpFjSBAU7E+iOfPeeREThQGW/R
LTsFz1ZUcpj2L5kNWfcOqKnf8KYlZnP5kTOPk5h+A2m1HdhlxcA1iDLaVMyShZr8/DqLjaUdxSTT
ZW57nszaxF+xknsi+9iCMX+Z1e9VhVt2vBB+HAl7HaJ80JBKM1b71npYpULCbE9VIYW/tBprLCFZ
k6kCT00jXdjBbxmdGUZ+UqQBSUqLvqHbKG8hCYU6SgrXLBEbZRpITwh44n+lWFmNfb0xhTY4ngzm
mkTdcwUbKGZySNJEAVGVffIbxCDp6bcN9S9CuNefVoA9bKNVdvww10YSW5Gj0YBgM7XN0aqCmFM8
mWt+NMKyOcqPhvboO17o/mNSOHq7ezQxRaiJkuuUQfsO50G8km1TXKFoFW4ZmKgy2CfRh5bhz5dG
lyQFVLytyoNX0YyKlO4r/AlPSTtpu7ZtLM8jK8fQpQ0qj8flR8vPEgmm0SAFca3n1sJGr0xvuW9T
xCyTJwswFiC6QZxeLDwZ/mUIOv9rPBepWpc5go6PaQr0xv2KqeNbsCsNKtQHBMLBjZeWftefWreI
4Y/uTdn3MtrVQFe1ZU2NzAgRPpv5LnHxuLA8EZuukHF2bHZJcHgMJUExVTvwQ0a+eH3+34LACKBN
RxPgh46TiXp8UxwY2q4hC8IQyv6x1CJDTl4D6EnxANrnByRPR7C6+SGz9ecgRvf8xDS/hhdqV+D/
FQ/KOhJg/AUTaSu9/Dy5U4047b+I1cW5eILAEcs740nbPqjineez1l47/qUvMmQqkpM5ZioQamiD
126fc0FvbcFOITpekCw32el5ktH7R76CE8fTiGT30QGTWoK9rRrNpeJmGEK4svmtQMPSFQtrRNfc
ENTptUnN89fYTi95NyETtp+AfxLhzIJdFdjN0lDvBxo1uOMXAueqQjO0S9XU20WWCWFaP0kus6se
BCGs0sTxbdhpSSI4BDrgvSgbscj9FTYOLoBKH/yT3gknVr7XqWWqM8ABa6c9OlnT5TJ16QozHN/J
Y7NP2JSbxgIcLVy6QxFST3xjLicYnHjF/nytX7eF4uMk5WMezA/LRVqKpQn8q5G/YN96h0dY3DkF
rrJIjDuhYVIv9iEeipAenQZnujESoQdCNIAL4RnpNjeWNxF7cV3JFrXT4JMAyJIZg0Mg7L1LIT0b
MWWJ/rBJw6HJJU6scWYWRGWDoVcuf40S79crp6VuBGUoo6m5eKZPTe1UiaxS6zz5uN/v0AzUipQ8
D/t5073Lu5Wk2cWTtDZWq+YQds8SBA1RDgIl5cvlVTDLZsNC1FrQLOrVsEzWDVD27TqYe/fnDKce
QXTdjt7kflkYuDv3ruOB8dzEEeXwjvPaD8pLqHF+WNf69wlDMX8EUqMCdNYY3iir8gEvg8JjZ12x
mHzApwGviAeVFPA09LHXoOmmr2WVZZzBKgtk7cm8dvcLu2eAEBWB8WsTrr73U8wfe99YXtMRlxYY
1i1iq8/cAdqKP4PjFMoFCGe9qkGie1PbSG2axoMEvRqSAGStiATBRZ6B3cemb29i/iA2JmmcRBc2
HkxT96z+kurk4sKmJmMG7in2HIMaOjyVAWPlhlfuk60kxNquAuXfzFqIf1kJKBrJvQ+cKvCVB+I9
NoKQr420j8LeAW8mkKbCbZS3rx9Dn+q9gTusOcZwdzgNhkTRVcB8+xrwwOl1T3qf7i0F1OvmPBz1
vg7/StTJAj9kv61zDnVPj+oodMMAlReaSd/Y9GDNJRcnW7RqjUKMIddKvlPwUkb7gY9mB1ot3zPq
0EFljRfGEP9jnKIAa38v0hKRoDiV0DpfFIBeq9Z+Th1kpAss/yBNcI4bfw4o3Ga5LPV3NAE/9c++
UBkecqrb3GtOv4H6a6G4UIVnc3vvOUZC7rnwQ8nCIh9wzuX4Uk5Tl5Hjal92vAeKF+8ffsTWimBC
aNOrWBzUCEXlBeP6v+N4675b7lqI5aaAJNRK2sI43bYt0+DDZOsUsniaR9JBF54stwVd1Vx7W+FM
PSuF/aY6wA5oRa6/lNLEoBY84AbfsIX7d8C0S5yOX3Cec43SlpeygDY/hHjTFahLapfarQjP6aFq
Lj/IFFHwBYSTW8n9IFtdVnxazpUEgofmcdJP65uhbf64IAKk1M7bZ/LEHWlnqRabiSn4EsuY97ur
b8GRdQQX6Bg6U7/WB+mygEcOXKZOOIYjxaiFP4FRbYPOws9olS2dWLwaALSDJRGBPFyOKILMG+dj
FJ9xVZB2hxcOmY2k22A4b9JiRVdwZVzQM88iFbuGDRQ+M7HXAmb/47YAj0wvekeorrtls2BSG9vQ
l3VLY0Y8xrFVQK0jsenQXXANC9mN8Cqfegy80oA2aCp8j5ZDpqGZO2e8ZILnx7PcMHd7UpBbiyfe
omk3HK2t7KLPBfdrZkXJZo5HCCBlu0Y4GzPf9UUa837JkriOMg2vVa6p9pJa61nDAC+68OxUFy5I
TcpcTf4uY3eNuZLMcAjL47fRo10Fb51azMizfCCUIbfrYMUBwYdNh7DpTdz7xNekfA7XwYPwZkjc
3VhlDRWsrqxfTwnaV0mcVOTHpXlTG4uPwQxu+mrL8Y5K3X1LBJr1T6WogvSiNqtgpgiqByT0aYNR
U1s/J4dkw31Vyt8vjbwefkjw49cSGAuEvhlUBGKtx+RrELQUS5E13DTxiUSCvyEMfAZWeXJSKOB5
MLR5ro9meotS5LffK7exgNtGXkmMyaOG/+567k9BTSt6mVkXMw0cE+dIJlCqlvSzHkWfCicyOXiY
rnr+Sm8B0GbWiNN0TNTS5U7FTleTpGiHs4suuH4hemuHiMYDYBWwpDMZ0w7uJjJM8uFjwC3udlHa
O0WcYNZbFwBNYLRcp145q+7lXQd7k4pJbSiTs3ZfzFh2YAFfohDCgU9CaLL92QasQD9M/Z1GJ18p
N7iRXN4QVMivhtQN3ZiZ4Pn6405IU2gy1lG+RzRHMS0JSL8XSLPWI/ASQWCdEc9Tv8OqXYHQ6DFx
iKQFMgDboudsrOooV2SEKaXVMA9T0j0X2sCQyb5vl4y+LhBbjEKYRCpc3xp9OOwSCvHJzFSsgBzE
obHY8m+2QB+GMwaZJQLXwJy90HgN088auqq9Q20fxbzuA6xTrHHFMKdIQaJR2OR4hIDybJwx463l
NCDVKzLwMczn7XDHoXkyAZLZx6s+VRC0rAmFD4jsFhKVXZuDjI4ipaBweE+r4IhrnERI0xR042Rg
OUwj5WTFJMYTfxWqL8h8oEXfIXUUSphkXoLJsaRIw2YlrTe7Rcxf44EuBOyqhoend6U3TGfXWzXp
7gLd3U72jIHxGK6w2mBifHv7SHIVweisyqqA7Xz7yNL3kbvK5eG9WJTqXKaRr/Q20s9Sfmp/4nOv
ax+O00/ZlpMqv8j2v28Cqs2j2LhZUBKH5VyQ/oWuDIfQsd1immsaxDnYn78k4f+L1YHUgyYY1SCq
NR1ccQ1r2g/GM5tMD+LzgmVEfcggl6Fk90wEekLXsi6eFu7BkjtDUrrY83G+/lDcLwDX/3pW92eU
SI9JnjveK5Y7tA6ZGYugAEijyuVb1DWpadKzJ/Y01HDX2xTkGB1zTBwSzoWKL31pywo8PqgY078F
bqxgxfRhXnNZYcvVtZRuoT9LAGeBqJn8itjpGt16SGpMJ+NmzMZb/w9cpOLLj2BGzt5XmR3IJYXj
FlOlzMdBHbiC/wz9IpazjOZVOC7SbPgI6lzFFPD8ScwEJfZ/vY33ZEZd4yu+Er70jXTxhUz0igiW
qX9f9Fed0E7IWpLTm8THt1tIgfbmmPd6q1SWA42hc0QjYEKDdf4jeIgrZQWDor1RkHrbZ1f6x3U/
mbn6g3YfQJk/YKeUBJbhZf5QOaMYm/wVtUInS9nhZlu22rzsjZerGd+f4GFCOAy1sV62QneUsNDY
Fbohpn0CXCpWVZVsovDzfopoX/ywQTsPhZlFfw3ukYprZJV2GBLSH9odfvaInP860f1FmfWMTOBG
XiwBBHgwjWkHEZexA+bmKdkZcLkNXO3luLLmbd8vraxFcA85bPNtIWTOwqPV4Wlrf/L1TwviCFlT
vnYj1sASFA7HalzLdArTzeEu/05W9va4Be8ercgRB8vGD0amVqksybLJWR4Y4QmGLrZd8m+QJxaG
cWuhd+k2VV6HShaavNUkeHc22kiPU4RPUsWFD+LtnDPy4dl69KDVLs6/shlZgm/qQdHR4Ckb0VSk
F3sTYS5dT6LDCaWD+grEwndpAx3pNrv5ah3nTa4Q2KY/V1Q+VEQYOzjTjymwEK8cve98dzL9jYHR
3toVdKH6OCT1If8fLq9o5ek1xc3NWF1fmoOxdyMUqyy2tYjbFldU5udX+MHemYygX2rTZky/CXRO
CJpST/wFVZwV60vmAWeqfeo/yxKLaz0s7NIpCKlqPLpotHhQtVxNBLXhYh/gQ1phi71fiW/omIBp
9avk3fWZLBUiI9DV6VIMZDi2/T5wjq73ba9sZ+3/QQOqlAx+slUqLaSnB4bvhwuXt3MxKvoAWR9E
yX2rPwVkbczgJB8k2Tfg+oklWyUPuPIvg3n0sZvEkoajO61eIlUeRQLM1sgFFS6RxDF7VLk/VzGW
kmPxGWnpIjdhaLnU03vFFUUF/Q+xLtNfnRFBlM6sRHXxQgNhUEItzrErqCrjuwO49P2iBjKoA5Px
TyzeKJ3FoZda6i1J26taDqiazvYpKc+8vpwryOJcASntQJZqSgtrsD5A9inPjUFjPdxumus0SA+q
7blv4/SdR/RpeJmF24OS3LhYDPWbfa9eye7btXL+96/6moj3fSUnttNlzdkPweM/3Bv7a2DqT9B3
gWBUf58NdlXxSiBYfBj2esN7lxxDrcLueh1wZabhTBXo+Ly5LFN07XRzMYn8PZTa6qU/ojs62YdJ
heFeFJmUM325XKU8R8+eByzjjMdl4IXb8Hc8CBKUvIU35RwIqq3vc8CcZE0L/i/hZVrCeP8mPIam
pnaT2qy1Os7ddOKrQc5OAiuoGEHbrstRh1IamYwAIyHl4Tks8MwsH2TKmkA27iLWon6Vfm6QRA9C
yqWQ3WAg/kqFy8YxMhaOtXWc8uHAOX9FUfKBvnYMDM0nnP9BDT7gGLypE1Ze44/5vJwUZjc6eoZJ
r2qqansaAWebvb9Xv2YWYC+oEVFTTSrIFyvSpli86OfToqENiOHPzBq96feliKxxJqiZp8M/VV0e
qjmIXYDG+23q1Bqo469GAzc5U5NQxNu0FJh8YZqSYSWUZ6j7Vej3TJbAgWLs7UzRGe0aXnEEeqSp
a29lpw0EZa8u5rQGbvW7MAA1jI4EeLPm/78peeLsa+cd4c+fIavu7Lw4WiawcDQIqXWqeoURsTGo
2ZMA/A8HevoVehXbbH0lMtqq17lZ9tJzxVfTTGBxJqAl8ATV+UXKpRvumtWEWtJzjMo/Se2qb0/2
qVUKxkFYMr9mKjck40qaxuOWRTQ7JHcf4qfPEm/xuZ/dloEy0mXdeOPFwYbM7rBJiC0xWy/DK7md
IvivS6AernsFm6kUz36zKFRknM3NNVaYCuNHoMOSaE9KvrNwO3JpFEv4PXjaomDJzkgcGypKZABr
i2IpDLXoEvvFgwnBIQQL9zomwd4dQ5qwO3bc494c85bAeIgNf/Reja930PQ4MfdN0ZhOlys3hh9+
aPhkJW40WBCXxPDSF66Ecqk8BdM8/vTWt52HP+4hCatH6+Qc4mH4/ziiANKo5rZ9dYIdtZQQ2by9
9L6y2e3ebLLUf+OIDjAuTuSXCLVQLpJDaDLKIhBGDu2MZXjyn2kJr22/h74d6u1KGmulF4X631tR
43m48+8sb6mKNVj7nd8/6NL6++6BC+OAVAnCnCOWGdH4ILQb3p98VTq1UcI9zGAPTvu4eqH3oG5D
hbrk14Yx1M8sxnbrsZy6nLNt6z2dG1wlJPaQV8RQkbbcItqiRxW9jpPuUZsBXkWryYoZJs0PfyFd
8kpMRzxILff7zyHIXRMC6drHQ9S2PcFg7k5kCsbS4plvWm7Dt7qsh25g3ediA1BdZIm7fj4gkhKb
aA1eTXMs2JbdjWL8DDSNSb7b99cneUexl905d6wJiGjfVWY8asNqeE3LmDT1fk05236Kfa2dEoIe
I8Gdhe1uOJpQBSpx01NNKAA1ZNPA1dScjYWj3khc6C3ZOxeHQ7vWzzTalliVeIYoRze6D0a84veq
FhNCD6Z2amwgYjT7CGvWE/UaAG6UPj16e36DRY4IogviMcAvEg5ypStMsBovXyrQLn4GborgL7T7
tmLBQ09SrU5hBxSBt8MAEG2W/wvFwXflQBiNP2l4r/iANqwB2T+7xkcYtk6kXo7pm54n3w8isaxv
bl+IJtbgsr4XOP139WUfsEa/EU/D6ehweylfTmSRBlIqyA6VxsLIDDFd1zYbpA46zfc/5cmR32sd
WEmr9xyXeRv6DQRLUjj2J/gk/ZugdKlWHl2MI8+Mv2FAwXQVfcUDGmNpWjuxvgBmbeiVTsII2F6H
lmCXY2nKe/FHU9ccipMIVPl/0Mx0EQv+ScxvjZbw6Ors4cCquUGhgUHfHgnMBZN53pThpK+CMMEB
bKg+fMcV+35SGdicbc1CA6tuT520RDAbS8cBQE/QaayEpk1xVgijyJVsiW8aJ6jBQp/CPrQgG9yp
TKdGRToGu0O7ia6FH9BQd1DKyj+UsjJl04un+LpgppofqitBUoWtjbUhPIkfdoYabWoNr0PJa52l
i3M/6VOtbdEW/UlKxp4eQr/uJ8/RfwrRKPY+iDLeFZiqGUNgzxb9X+uv3sL4VWxbp0fxKuO9jixu
g7qaVhxInREUtkWp2wrJNvQQcwG4yBu7z7qbrQRO4iMwckzjI38Nmr1JSNoU71TsXWy32OGN5BAN
9fxprO6OS19kTy3qNYvs81MgFDsH0G8t7WUEkOUJHLG8lUunj2svvbhLuHutQEvmojGXxYBNHN52
Whhu1pfGVlBZidf1USpd9Gx0V9ngYac/uroR8N7kYaQmfpUYQ1yzvlLsfjXCVJrgDGI+Fao30vCT
yTn31oXX1igp3Hq4nXTM1uaZh/cHzGZqz2lsixh75GKTiQ6zsp4wjEg3NPZP/0F8IP7Ca0QG2132
ViOTTYjh+4dXebs3BWB5B+zcNdD2Ra55Y3l8ZWbu+1VAv8FX6wV8+0V8rhj1g2FZqGbUcsZyoM3R
sUYCd4CtddjnfWMypBF30cOayQOjqjrMG+Xgee0mgBi/07RqEbQeqqJTaTYlyYTBUHm0bULQf14J
Xw5xYHXerOoMM3kbkPLyUmBG6fNQBY5z5V7r1JBNpGu5v4f1T1gNHpFDxd8LmefUluJYEs0SUZwy
Nj5jw3e3xpYQQqvU2fnpO01ze4ghwKVTogOagwcA979rNrVsB5ltYAP+STd7C5V1TWSMGCpjP6l4
6VPVXIWT+tN26I1BJg7UYTzM4AHHtoJz5aCPUFwj9j48XpekjOOwGA/F5QHguGKUM6oblJj3kF2p
hh6XubdhACHBGpzyA/pfIBr2vnoTVWsoReDq9/8tXFa1/LpLM9t/eIMdpwq0IlsqV5EANNX0TR5X
kowyz4WtebTP4eeR+RoMsqO8LogNeTK/OomFv9uZoGPfd1tj3zN0VfQ7RmkQUa43SQXGlo6GEKSS
jfjyjWt0h/HkJHmBE9tul5O3EfN+ZhzyUNHz9WAuy8Z2v+BHKQejz4rRWZnYlTlTx/ZUgZiZr0X6
2YShzTOPyNmyhRZUiDO0XVgh7NHNfkQ4IMfkHEx6K5MVK/hHlN7Bz2wRFqUQkDQMj0r/nkLognsG
99VFheXiB6FjStFWDdSBa4pvgy0z72YCWteS8//rFOlpXPpDMkkg5beLGnHIWZZvvHW4Cxt2XJY4
0Yq/Lg9lG0YpbpFXvkNAFQYER2LHIrBsjGeC30d7PkpZ/3e5utlteDVGWmTdAsSFghHPA1+eoh22
qop9UF0ZKGkU8IqD21jV8YMnA4J4flfxuBnakBkZE8C/xFXNEeijP/eJ/kAt5ZeBG1RpYyTY3giL
P4KCg3MSBv4p/Nb/iLZ1LkGNZJWhNcTtrHEj9QhLAfpFtEeXhg3i7i/kI8v5HModtOhrCuCl/W/d
8JVTAl5yVNe2Gv5kQOD4xdIOGBSy4n618VY4DyiekFe9RsJ2vEh7qUTaGCcLaEaEbSOyNPMpOh3I
lavCTJnpom8H6yC1HRoW936eOXIgIqeni6de68xAUt3MEEgw3j6FbMfszNYY/4FMy9HORLrtyPPy
DHuddPsY5Bqfub28xKkGCXbzcmbc+NEoAnJUwkzn8p4I4MA+3BctUrS71h0bujB92YqfCvqXwqDH
UJZQJVmuGh/AR2cRUYWJbNCbFoDtPPLwpFp8YkM+MmgpDt4bwTGTXHKooYufC3v4mu37+0iO6R8v
JfUT6M8tdBjyPJ4mbIsTyxfYVuJhPkCbwWYBmlQdI9pvchfhrkSDoBy2Zejev2cyUp0o66/KkIkU
J0fi/l4Yye+o7siClK8+IJzvROGYwQ9F6BaZlV7xXIPb4rzW3q4euEmWLZ7nQ8LsSFYqhByFtdHX
ENs5MoEb70VjVkiTjXzIMzftIJmFC8i5DpbCay3gmPyAMSoIsW/QwMnpsHF9KB/n2BbcLxc4Y7j6
w0RN4pnac3+7R6xQ0y4QDyE32mASAyBdQiZP0uOqisJlL5YjfRHwG24+2wVwVnoUOET0Ki5GBvCc
zErKEmUrcHbBdUVHdRMduPAYBQTyPDwEzOqK2tmSpTDynOv5x2YKXF9rGxtvhtJ4TRNif7QWeYTa
CWSbf2sRKInSWKM2Uqa74ZzhlEaZ20wOOjUkeXlnJKA1RGm4oIEKsNQg7AJT1Fl/0EHWwva0R+8K
MCobfVRwAIE64Ndpv991Cag2hePdsicGfFC6Q8YB7nkdgBMoZpylfBmpDxBGLmcYnyctDeqwY4Qj
IVP9DnkTtEhVDmdJKropKvsBBZkV2HY2Aq/XRPSIXWmJpcFJeoEif9YrXOLkpDYd4C/u9djPJ+Ux
QJu0vJh/X5hAW8SR/KD2BoT2rAC530XqhDIy+AYQJRD/J/LP7ZH3NCHHtQUL15EmZj9LR8iN5tQ2
ahULyliYg/sG1TEOKPgvNBMNfcEuuTncBBDPKfHGkZPjLA/qq1xsZOOoQal12OKbj2vismzWflSK
wNtU+/lWlz/lE9M/Zl1JclEG67PyD7F+1LYTkHeVGqeIbMlUSjWj9Zm4/CmED2NiWN16wZrOw+or
3g0CdCHFFdPqApgo3FUG9JTr3Dk+hInzVc/ediOPeN5nQfHUxADupMuyXCmVOwr9+cyoM1W/S46m
a+4ubYQYYBw/AlncO04WkYQp9FQAK4ALDl4oNmOrgagEe4yLkgUADxQ8+Kyrr84VW2Qxa6WA8X/f
7BlPXPxkSFfKyBay0jEpAagsXBw8YTNB81mKRoC7IMmU0RMsKDB3yiZL5J1tBblwHxcHCY7dqkTo
AJTg76KKp4uPRsc7tMT+y2QkCmNtsEiuGD+gtowfi9OEA+wqitL+ocLae/JnUPNGrJvBDR8Bd/Gr
d+gTuo23ctyZFLwy4Y4JBjE9mpiyGbjG9H1REWoZYrl0VK7S2d8z3qtI0Aff5gR6/cnGnMqfdxpl
EIijGaqzQd0RFBzLPpgzhWQvD2BUvz3phu/YzqZNMFkvLn88N75gm+dadCPQYJ6dfQr+MkNvkmWZ
mu73cNT2VSX9huP4FjnkoMUo2OrDTcBq5JtkU0V/u8JKL+uJ40m1S1+j2Kw2xXoQ9Xm/51Z/CWbM
2BM8CFhMGjQR6IB/ra7gDc0fwKCJArxx4o62XE9cVyCgkNgF+NqZ8l/SMJ0dgsZUHr7z+VrO+VBb
sfc2xgxW/XvWnwtnQRKHMttargHltNlBY3OA+/cHz6t4ls5MH51hr+x+yWqYnF+M1oRusjKb69oP
1QUD/V8oRRdHUVNaUCA+KhzsTkRGbfui2hRkffX5A406sJm+e8Xpb6I16Kw2uYoh5xaxvgeW6bAQ
O0qnvcc/IRthaleo8Lf4BCMOsPJ/ily3KhG0enZSJ3VHO27cJM5pPclwawbn6WQgineEiGPL8J3U
dcAswWb+CaPzVLD4lHWPtqdo2Sz0JO9ubzALrspz8Ty0IAx7XIeq561kEEEBs1fGM4xYW3Hq2Fsd
LFmjGL90d4bdHZHVKZJ9FkmfNwlvsTJEyx8Yz+CxbcSSzzG2feuK6k1ZeQxbmxMIc2DtL+KYKI+i
uRprgMHybZ5oD1yOf6AkQhKyUmOs+OV6IVIHxqs1LOUNZkefT+ZQrHcF3R7EE/DXXbCnehjz5JGE
wUyEgfLBEIxX7gIJSDJ8QVTvpDDn37JUd+6sIEGivWacs97F1vOileklXd2jL7LI8uWeRm4THtbM
GEtLI6B6GdrFba0LXuV3V+Ko0GU4KVY1kOjopLSG4DTfR+aeVVzUsMdJK9l0hVrDXUHBIuqv51oj
muopS1b2411j+nIVLkoa5W+UJSmTU+BNkQpKd4DkY9zEnLqE0riqYd+e1if+Qf0sc4iUV0exY5jO
iC2sQCc9tI2Xx+IOwBJispBf9EgVgtbnH5/m7edH5pwbdOnyvFDKuJeW884akmgNfJkj2ExLqriU
CHuwJiYo30BaMTB8TR871A6ee3oT6YqhJJrNUteYp3NPmeLQPlyFLsPxylehwsGrblSa0ksH+lm1
zDgcydRABSem2Zmcj0rFz4xZQdRQ8e7oAAmwQN6SWL2//hnvEIR8j4rkEGGFsmqTscDOIWDtnTxU
lIqEqht88jmDsf0VXOIONKInJlZT3ddCldakeYIqSmFo3PCRdrQx9f7JAQh+4jh2xco0ZlbA25fN
w7R8xien6FvGhdglAtXuQs8XRdZjdjtVHdTENI7qzZeJgAeGY1+w7EDxmchnw6KZIlxZRWTIgQkf
wLXTicYPIauKXbtR31l1+JzS187R1UhlbbvC78jfrZncOvfg4siJvXre14HXvVF+TxHXJQqDosSv
JtFPhu234IfzzXzr1foBWzOmLXm6AhtecIvS6g95XVLzHoxuHLqcDYgrEVwA1Ntpqq8ZJMD5UTuE
T0t5GVZlilbEqkpUwqMyzhwz8GA4XzKIYplAl4PPjYzFuKYwnXDER5jsRnEVgxF6ttcP6M/nR2QT
FtOXc8N1uMV90fvlBpd9rW18ho0iijS9iIJSMZvL4L8pDcacgrbH6hYjj5PcpF3k0404Fqk+MNSg
uL5Uk5nvy62kuu6jhe+uGo9a9YmFgnVZ03S05WmYnjt6/KMV3QG5gVUp9ex5gsIVuOXMNP+xhM5A
92qRTJRdzvq/wf4sQEP2wHr5zxMr3po4tLN/wWazBb8/E08vVEiH8qki5KZwAr12zV3OcG951c6F
CDUSN6uRsTzKIEzSPP9WOZ1BZ+1JJ/Uwlxn2UvN9SYbSmQqUVasOhIZZ1JjuZikJdoUh1I882rY0
YavW3BHhkzXQRvT6CWwQFV9axVTy2aDefNWU5LPTYzwPd+O2nQvh0vH4yURbNMHfVGwrY1oBevcU
wufH5rYjTstDsWyAFbrAQjjO3nYknoBg66RmPLZ/6ru4uEnw8kGHSR+VmVstYlpBqCGojaY0jV+V
cg4KpFngIogoys7BzeGbov4TdnyccQHuqBWtdNjPGNMwfpENc0zi0ymXKdKy030pi79QvU7pT6kH
m2eKniKVbCY5jfWfVM7KVVLuSTTyNp3oSO+4hhGFftOoLNKoQeJiEK939ButewTEdTruwQPDOEaS
NfrFCTPXEPzYCe/BrmZ8s3cO/WG6VYlVyQ2TVdVCP/AdnTevdasdCO0XVluh6nGoLlU3vHomWUVc
hyq1GnygtPoTNFM2Yw2TF/T+nN/8IQ2f0QcTc+6SM2b+99hmis4CEG+tbzykblpj+/ucQ4pNAptI
8FUgIZDYw+5mEwcPdxwA8qYnQgIBUjrHgU8rlu0wPNeT9yAvr70pqVf1DFZ7qpGvkgJ8UzuyD9Lk
o7o2ro0ARbYhMeTktC3aK6uC3vi5+GK8TM27D5up1KxSxmczEmK+0Ca0hHyzZRtwnFqpRW8IplXJ
CCQeRH+PAw/cCfLgjMLeZ9wXgsAri8Xp42PUvvj/QbBMDuLuSXhgqv1wXwpdYt/kqtnge/cf31gR
9RNhs+bmZcAtsBSoy5NTQIjvxnwfyltEaX8t0uuLHS+ByZT+HXuMBCaZswmDoYsx1E7hqfZ1EZee
j+NPka64ohsWM1RIF4/8dGf9yq7Q2NCQjE3S+SB9JOjhTuhoUDFidu8BG7MuBP1ZIo9S56mErQ31
u8T4TOuBu8kUS31QLBG4RHoi9dYO7wlmcRFeecTs4D6RE+xPc0S/830aRm3RGv9IP9jJehfPYEtY
/qUb52JZCabDBuSZghhZo+eO2chW6fDNWoYWVvktu+e1vLkBv4z8anf3hPpxnSxYHvWAsfmiImTw
8E95Qxd9SN2EX6xDyvfLIuLAxDDZzudjivaYVeZdsXMyGjG//4hakDm1dj22FeS3asSk8QG+Okyf
VQLJYEtvf2/7aIHjSoPf+P5zoaqKQfpsmGekbgVaxjoQ3/GvvOlKBfNqVlMu+G3R4TAB2Cgr/hOt
QiG+RmaznsGrOqqw4mybR4vIjzmbElfnpssehbgpTfAQz7roXLzDMo3mQn6X5SSVF5NGxmAKW0ZT
NxesfmRWXAPi4v5wavJJ/QL7LL21SvscjN0LM4t6dXZyLh7j1ac8+9JsXbwKx9s/aLtr4VjKuxZ3
6tVX/giZgTE6WGlGOGEiyrbA5gnBjGeN+AELcMY5T9fAxaK7s9WzvCqTw8tZs9YEyYBKatSH73HZ
j/V6Yh7RviLPueULxLGjki87M1oQFiUlaASTR2VwnRpGHMsZE/ZdmxzzEZ2e28yvLAMgIqw6Ksyt
103iGaFhibZvVo3cTfvps4uYIYJBHLu6P8sKJoc/iNQ+nMhgKYkyQzG+K1dy0Eyto93jzzyLj+HB
hXbGUp70fh0vabBHoD2ji3haRzDdTvuS2exO/PBhvtj1bZOV+MXSFTFO/ZpL68qs0vjcgGBpL3y1
lrUMiuJJ6UVUtUmfjGGUk6fDLwWAM1BRS3OGSld38uWjAxEVLyfFORIMHRlwoYnaGQ+hrNF2PjCw
+S8pvpw5kQ1hAFn8B1cmiN0aNTrHzDBiYItBbBKyTrGt66TPPjoSHhmXYguCYL7vAsBc2mFAgPty
6IQCvvXQaLo1XeDNgd5+Yg53ViYkcnwm2uaZkzw5WcV/WPTKeR98eNHGroQHxvWpZuVdE/yZX+nc
W4bHfIXkcjg5QqPBjdSOIw6/DKGaV3YPdwiuT1jZKFUQzxrKaFZv0taGc2SirTbuJQftDicY1Mo0
Pj/n68OLYNepVx7D5dxTnMLG1Ij+YNYOqbCj+QDzNaereWYX2ubmlxknPHog7OjFJhQtSxhOanRs
61WWeMmYy5rNOaYdDPcx4nQ74x0enISPKCZ0QB0GI1B+9SlnHvFXTZDLlHPh17xjnTU8sT35OZIE
tLg5k1XIk1JEKyKY7L6uKdP5YtmeGux+3n/QsVyvBCn9NFfyDtsgH2RZF10vQgDe2jgoTL+LgBn8
awFoxURFRkPg1zPMd0lSi88gq/0sgDSjkt2RVNvh0OQ9r2ZlzYlnfqBvpLxluZ+KvK4NQsfgv+qo
29UcNVPgaKLFsCu+4p/i+x76TovRTdOGplhGGAqeyB4FkRRw0UUkvK8frAELpsDCKlhEaq/q2tsw
eihZFDnlwm4eqcDb7NAa6oMTIqKdB+8wWYxEWs8Upc0xuQjw04kLAejWwKOK1HpXWvx4mrUbhkOE
HVang7zMxHf56ONbZ9bDvU76xiRD2oj3RujRUcdCxMsCbJU3ClPKeWSRSXGToYXfP6dJ+ai1keBD
GKGfweXlvAET3ThHEtC4i83tKuqENngncfw08FUFx2V1kR8s7agA2oVWfRJ5bG5cQepVazBql57+
l28a5Da/HvxBOrzV5+Y63mY+QBTyrEYBm09VouoPe+MDihOkOfHhUSRdQWORbTM1vFJCiT3z8Ro2
UPf2NeBx6uUub97Ag44fjlXWZzy/LTu3D/0HjpscIbqfKyBTRNXp3Av50/r8K0SpwTvLE9MOj/YN
wDpwW78hETSGo1lOILbuabzzz9hExJzPH1NlPtnTOmjsBF6glwgpi7LPMzQjRMlnNs7LSGFsZ6PZ
Nw9fWu2rz8k/bi140E2DHNGpr6X5OWlRFk4cGMKwbTB2S6JA0W6k3GVhMSe8ZPbVwcwVqH1iKQ0x
Ycns5zkxCTEv/9fpjxdhVADkGwkr2PoFb99Mrj+hRya6BFNX0bk8Ljh15v6UNzql5Gg+1FyWGYdP
hEf9YZPH0dfeJqI4bB67FOi1mHuyVR0RSVEfyFcYPPSE37QngnQop1ecuWgn0e+YYkA1dQZnHQQn
Idans88qWhe0z/Q9rsYBAeCbYE+L2cDuWqLxYQi6evy1gayB2TNn9WAwZp0D0Yl8ZwuEv7wo97ag
xf/582hAwc8A21FtsSVcIs6urQm1r96TGYK8cfDV/lBqz1Sl9xkIOiHcgOUXyefK2uPVPgWVEh78
9/vtuw4nPXQKeOy1B8RgQq3RlnSG9UhNvdvm0jyLAJe/YWy2iZd+mw8lGpPl57FF+tpC8P0qeRsS
pF5l32q0wfrEE47LiJ8F1t2jNn74+U+xKxePlWWVfiFbAaCraU3uj3kZBSqnvgfriYHice5YFbDf
Ft0qjaH3RlGIZRVKNYpwi+NDxWowlcAqVOYqZsGsQZDsBmUp1g70BLJkCMLzo2QaYuPGk8WmUuSW
FC8c1jBV35rVxNBosrauW6lHpI3PDuoV+jM48dTl+cMVA07Qk7YDeDTrIbQSj/fMBTC93rrnDTFG
GJbx/MlJle+zc6TillqNWrZ0lPpaJ6skK1hWLUI5A70XupVZVCpA9cI1fc4/+bIDNbF5UPMnFvXV
XNZQZxWgbd4maAqpbvZefvxFYh0KQHymRfPkSxm8CYyNFwxFyI/JoO7Hvrb4xB7W6+nLQwnecycW
OL7o6amojeG6rFmb01G8l6vV1eEEkkwLQktD41kVn6BvQiNOQH9kX7nFC+Hg+o+f2KK1MWkJBfbj
nqIYbT0TdwhwnVfw9IMrRYUHQ8OFtn0EjwghT4zKMz4a79TbljIenC7qE7s4nmAwBw9XiXloreTl
nayBLB8kLX9y9c1XziMqcAcxZ/I97/norJqfw/rt5FRrm5I8/3j6u7PV5jqSd5Hc9TL+Xjxmwx94
ooVTsuPDqyCWfFToFX5s1ZPKp0Owx7kZHbpsZD1x7zuOXa1kdZc8tFCMBDunyhYUnSN6deMhpY5l
iDjz/cSTrExe7Y5bWfHr4BeT+Z9N59GaCkDSzcfbbR55DMhVmpUfQVaSCW8HugCCo68bVbmdaKj+
mo69JlJoeUHdy7Y+8qqF9vPW4/hd2KWMbgmy/myMI87mdImjjvd2Bb803Hz4iM4WJ7QU650oT3+j
mV/jfwuhAoqHIIuzKY95VMCMDx8HEPwidqfW0uNedqD/RZ4QMLE7cXD1TN4GQ/czYgjHybXDfXJ7
6/kL8Xt5rPchm0bfZTeExCRyTdfnmKKrWFVdn4VDySRj3MA8t8Wg5KTpn8AT1mRDN8KAvmNCYrx1
k8LZwNmhy6Usd/VhBiJLQBwqHbQdl7PUtDa+32OO9VHdic7repGGA57tNrJBvez3DkuoRIMeJ0y7
oWkMHQSs+DJuvHsbKPRD9XUSctwoeK+tCq79XRTuaq4zn/4ckXiKSWYaiVWOjVhwtysG6tkmloIU
u0Is/Ym7ioNM2/pBumxeNol9hXKH9u/uuYlwLowMLD+8fWwum5Aw16ZSeJbv9OtsktN7m0E8PiJJ
cgJD18ufZNJhINuGOsKxKaR07bZP1BFe1lcrgP2+gPaq1IAPqs1X6ylFJEwg9GZ2AWKvFlzWRvAd
QMASt30oexbEvaFsNDKW4uMbap/GuDubwBgA1AUdDwoLsfquNXauK3daWQ0uOme7OWKFA9kxPlW8
+wzai669PlZMVurNabogMejuUxNZgOZeZNVZp77FuVLHQ07MBW3ZJuJ9IdB7sttOtgff6wtrzppZ
j4aA3A2DkxeLgZohuTy3llBeRUGGb5/WsyYjfDG7w0N77rBXZF2mD9YfiI/uy4IQrpDEdDvYWoZq
KHGmvE4kriq+wLcr7l2bK75c9QqOPPEMoRPlt6HC7Oo9niRrR9WTrPOsQG/t5zul0ApDuSN+jf1g
AUKG/F7Rak+Hxjs3SIKiGXyJn13g4BAoJUvMA7kkEqWmjxLBTFc4f2Ri10lnqZfbdhWGfNlPQ/4z
7uYZpP9u4DL/u/I6+Kx8u9FYlgDVEib5ehfEfGg+mK7BqatrrY2/ild2rG3leKeXytDKAVLQIC5q
lz3jTE+RmVFXn5LahkdYIyDIWldMDopeh5TzNuF68CxMVUF8cDp0IKZiOjZpfRp5TOawkGOhl7zn
utYFubxwrAgE0w+AhnB/FFNQ9Jm82RALVMLKqJw7fTLyLXYNNrR7ZwOlwR8BCLnFwlBWJmpeDD+p
xzudYieYKQXOLT3F0eDb0QWW/LrnwbgooR5dSVy8kKtpupYrwwv+fnsjcDpCqE3WOih6uLROdyp2
dutEhuwze+/t53sAkG8AXKeDENej7Sl3/JP71qVGFfYwy5nAuiKiqTv3sWE7cDmOCU0R5yadSHBC
yR7AyXaNKmC5ZCvVyP3izIlLZfC31jXTJd+i0naKcf2/HfrfnSxLCMp/+jdnYSmoE0t4nCkXjXcR
F3I1ijV0gJ4HBbsNpzrTgaofRAMtRD2UuFz7c6qSduA3eqcgRkeKu2ueyQxTWi/M7eRo917Jz14R
fEIL6eI42Ez/6bBZqGvNzs9NXZudyDGmUpMV99F5IO2j6g6xlFtJgclffteGlr8dCu3TfD9f7pUT
yKofBxQgzdpWS64v724OnMUtd2mgOEJNpFEKX4eG7CkszqsriPEetxglSeUJWlpd1d4hYMK+F7PL
OncLCc8lC+rogoThC2A+MN+3MqLY+JeJCTFZbDkSGynm757/IohjlAmvoOLANfvG2mthzHXyo3bF
VYOCHy6f1D3iHmhpff42QHQwrKKL819hLM9fGqBFqrx3Pd1+OMGdotO0L95pmSc7cETSNnPvQCNF
pqZS1rBE7jnAEXElUp+HnmIAsm19G601hu+lE+rp9wdxyaHjUiwiYiNfhH4idYUCLqH1ZgZ7REo/
6GPMNb5YreHQWscWku2UeUW/TK3nTyqlJ7X15lS2X5pKcBpyBBPdzZjpJk18M7SjbBA24CE8XDFV
kaE+mrPPeJCj6qAgpIpwcxJbEPXrs+eJIz4A8h/HJ8pcFwRtZ++hlp9YlaXOYsJZmeFQ/D7OB1F+
7rD1flkrP/5xiFjKQNbUg+JTeiXUu8FZSg9/+38+8kvdlB8FrpaTY2cY3S3Vh31n/qMovyVOGvEE
TIGl/0Ddwr+hy+8W12wv5pnn+PTKwPYSNloYSJWH9COHtMkKE14ozU7iSQ1OfUTbeKeR92dU+V8p
WR/nYTVpG+dcF0U+4SV5UP1JyOUtAJan8DKOcccJNmlf3EwTNfVZb/de7CedEsCmANgDOpIsxpkP
o6QAGhLBApRVlehP5FMffHoo7uFDggpAlqrwRBe/Eb0KWxue6yCI6InGbSdpySG0oSsJK7UaJrQW
ir4B+3vLFFbn25x92tea3lxBWX84IdsVULCU8l0uSssAZ2bQGHpbR8Gjrtj2ABD9juK7jKco7kPp
+tArrk9L9brsqMGRkj85gkV9aPD/bFt2kHWdLgnxBZEc45ohYQfpnzYC0tMd2yAPXV8NNkvtxg+3
8QUGIXHg0Aaqlw3IoIE0U9xZ/ZvkmUgAvsb0GwWEAR8+EA4vVEflYLyjoMfclUAgfrWmp0qMJQrL
LZNitUbPPchERYXw9PiRuUgvWcaRHENdVwYN4AjMu29kjLV0T9O4TCkj5sK9hQ86uTPsBsi6gmyH
C+afjiEQEfOAmjJipe9FdtNYXH5/6Rz9NXu9aYrsOSkzHkGAodF89/YTCHJrm9VoicCqDzHqTRbD
1DJ19gFDZirLicWgNf65z8XnKE9xNJv75idJ8g89ISlXAuekFoSsqLd1CyYC+YaaIcJbN1MNBWpH
KRtxG0KZaNfBsjtvgj5Ay7Lw9NA8n4W3Rio1lyzwHBwAK8dm0hg3dM4iyRjdllME447tIhmqnVWf
Hc8+PPu1Z7P79VX+liceuXQIinBH5GNfq7z2qzbfyTStfnSai4LE1KIzLTBLsWG1wkS7Rh3nuL8y
KVeMHwTC7vTFlgJOqvwezA6X39C51k3ivpZ+f+/d9xF24J0pX1K2o53Y9v9iaiQ/hNtGhl6ozYDZ
7oPEjhZuv+gBuxEYG8rw9E+C5x4KNxhw8iqEbbwtuL0aF95SW980/MFFzA/WnuzD8q6VDkoF+1dh
ypbgRS/WDk6LIzRv8RNLRljKQZj6q7f0z+0spMIwhb/hmU5+kFIDPb+azVB0q2YoPRsEDs2f28jU
N8cnhQPhawsG9JRMOZO8r0fvWt+Mwvgu1cewPGhsYXAqSn+0hqsiGxG8ygcp+9GnbKTBv3XY94iI
RYzAeUVAhOxFm3bL2UnDb4F6UXupTYZVTIYb0mT7ArdXXrI/gYXItN++VmgPdM1lI86Ta+EbBW0z
+PaCsaV3SUCjR/zMqrSzE5iUGymjzQymuaTrS5bJYCx9bM4/IKPT2JW30lmuTOJ9GZ00ZufhNej8
Sm1fxOy98RPCv1SlSmjAJszq2mXhlHzYvBXeHTciNxOGHkvNXZN8DPq5HHvvXHx6lP78EnyZhBbv
QCcMU7n17A0+r9I2pgY2/upnTUUDV8zC5iebdv74Gi0GQPpZCtVtjnJSc5j9r7OGjOSpT1oPTH5G
lByUn2h4hlid+pHedKUqaSX1/JDH+aVOAKWgTD6f1xNNzHQ9CXrTyPt6xgqJXJxAPwKUm+wzIs3Z
60atwWU57820Ehu4sIufWqDFulI+IDzKPIGHEqi0R2skz8+c16BvU3ePYLR0obdlaOqr0JHaINbo
aGw8mfxrrg6UX3O5KWJ+WdVfeJJFLW7jUh9h8mZUNZFNF5drPlbniqK+36F7b3HgVP2F7PzEQaOQ
b3SLfAeY+EhPgl1a84Qu8H6slxDp3I04muGGHhNqZP5YZbM172U0x3ymmJEYHHuziXFOU9Vcfcy6
u6Smy6c4+h7h/aDS6uIhiTejfAetUIOb3wbDwXvOj0snxnmGhZhS2vv+ufyWuKTn65AwsDPSGeIp
brILvj2/lPWpkldUN3pdNq1my5/GXlStOMhsC6UOvDFlZkJLhuXsT7ghVfrbsu2juFMs1eAMoAWD
WZ0BU17QgQ/8cEhhGiUOASz1nXJ17BytwriIDqirRganzwdoaQ93xN1uLIiUUClFhsUqqoFgrs1+
CvzAZmvsejKDOREL9T+uFXQW9hSZ5rBTf5WFA3146J5L0IggYnHb3ZxGb+bGOJTZIxFVUZ7ngBaf
DtAGw7QlAJIlopGyVWGbwaZcbxvPDHUzJ9B4q27bfeXPAbM6Z74NG2ePgu42TYHzX/I8XtxArjzx
umtGJ2HlB+KbSR9dz/FYeAG6w3BSxFQZRp0abPrwh71DTqmvmHw/umVMJf3snsmu7fAPdU6sseD2
8CUy1S9mo7+c5qdMoqkqNJvnNqjbwZ6tBWiAoECxIIZBt7AgnM8KTwKXF2W5paaSHqqOWU+23y4I
lpPsKma7VKdfV6ul89kCXnVX5wb89LayxFzfLH6RgR3h0kUqaN07ARuUQvSAl/XeDtN9WpbRQM1N
Xq8HbkIvqNNG8oaXM9nrQ6ttqG+ENNrDNojHnZ0Ho4iECp4yVcO6hYJ07tIOaBnEyM8s5g4JNcjx
O/gGwEKapgfc45egy2ykNybFmr9F9v0h8dvzg7G+UskEzmLjtF8PCVG9haL6VpG9ky9CZC+4BO4w
pQXgdm5ZmbNK4Syz7edH1kUpMnlFAy+k1NrFTp0ZAz3IYF0IGmUiWsRXAGBscZo71m4mbTw7GyLo
RD8U8rWu+BUv7S6Jga4OgGIP4QXH9yG+5FX5SyURbZL7Akdvb16H9fKNFJVvUb2/tglo7BjLQ2qc
pTQ8/7d3KMTTvQDGpU2P0fX6OcfVJyDoKX0FJSveOGA+pP9h0F9FGv6FeDjxuQtpx9CpaljxUefE
nxSc1JYwfMZL79kl3Vs1wHAEjo5qkf1RRMlyQVcxsgmXMQjjEXwQ8sX9cUoLBAHOVl03EryDUcxE
hwLIcF3gE84Sl69UKIYdYylSMChh+WIivRdLD7Teu0+kxJjyAL+YTEqsn/vih13mDhwnFHZJOzNl
EcrQljZ2jUI66Q7YXddjUp1Kk6bxmyeo4a6CijZ8959+k6Jw86Y+Onem7OTr4sKZCO9KNzf7an23
CbjF4Xb8HtjshdEYWwMPmdFuC5i3bTwUw6SiStxeEptGCut9OJNrmaYImbYFOCYgrSMljW3GZNvd
Va/WoZPjVsA0flTHG4UYHMSMKohjjuEUJ0SAG6ZS2EvKdx+3rZ0xJWs1HKfHwM/fhxXOomMAg3a1
A5h9CJA24QDyoFKycmxXF0MtcwjkGpQBceIbgFSNtnm6Noo++Hi13jtgj6/rJsi/Zbe4B6fXwqxY
2IOrKcaMgkPcTGsg6kNrJCIluTGmj1UG9UQokZotuSZDKRCaF83lcu3lV9XF+Autf/bx7BB5MNEc
S7WsUV3F1F5W7a7NsLcljZGu3TGRdV9Jf0wcpiZtF6d3gjj/E1bhtqgm1etxPiauhzDi0ZfMdFcO
lm4uUWNQcSPCe5WZINw5YjNJd+gGXQI5UFOFhMYtfQhX5mGiWdvMXc3AlQqIV8jWZcRnMzsKxM/j
DR9Ww5m75oy4TyonutyJkMRwQpQD9HUpPGKGEGgew3z75kTXYMbKUvRHwmWGcSpuOx+dTtmPtscD
Nj3IHqp0TokeiUguwq/wWmCaOaVS34raHBmbCYKcrFxrRMgn65DgG1QedKBehUORTZ5PPXByvzp2
8T3JFkr/yV3JRt4rIbpw/VbozaHjdhXtmAe9jWtt6SCoGRNrRo0h8fB53ZG4TV4bSbQRDPiAGu5D
nGXWhEmHcn8sl58qiDwE554yyOQYHPWq0LRp/eOiJ6kLTUVD7n8lTfSKdwfpC4eNKOZznH9F/dcG
khT36uYda/te6wPkAsvhiwDCyFblklpn5KauwgKgc2xFqlixj4ZeBcYJpea1KVgBRtwqaGnJD40N
YNlaKN3JumDQWZmF2R4L9qNNDycFoyMauP1NAZUkQvF4eOjWlQNrQscr9kzYBzcGtYbW0fx/yv3n
HwbzYMRAQ80Cl/N+NueW1WoS6batTM0psSeSZjG5zSYEp0HR+JpJ9HKcut7g4+VHC9m3auTVc1Up
6c59chwCaT3K2ZTGH50PPrV2E40iXtd7JdUxGIrxbEUDW3Vaa2BQFn+rJ6ZANIMbK1roHvm09BuU
9oPNmTeJP7C+4N3MRd07OCVyqheYaqOmgfm+a+3CHb9SPG9M33U7QKSMr6aw/72q73RNruHBH0jW
/bjBrl3xvP4PaonL2mdfmiNM4c+R3xOfB9F+itbFQGGCbGOveckOgB2SN8YXscTCcfFheDmcprOX
39hSGyFUwOPdhLtaRHHIbfGzBhJfs/a1X5u9EPRa+Okd/F4RY2UB0n1zDq652Smxh6TsIbuW9mjU
KlkTLmR/ErfUvFkli/FAOkg6y87OAqT2OwzAquOJWho50TARdurXUo+OGIl+WVwv+m0DeCBR7RKD
hExG48uurBaQ7dptIcM3fthGkDveQsIycKFUieI7hxtFxwEkfUllUNuTyyxIJbbeKimkXk3P5oRS
KrG39NsYHnHQ91iRtJsKdu3qtRp171Ek89cJ7pvL7zIFq7QciZsSm6EYZVU2ixLh634l+djx3QB9
WbZ/Z/uDN2JZNMNyEU04BH0FKX8/T5TEbqdncz9xekc0F8x/6Jk9SIQQirHgd7XEqA9KPrQy8/Bi
un2uJyPqNytzx3cC7QavpfqSICcaoGWh6VGRjZvWSR64iNYbpEBTTI3s5s5Rxu7UV5iKzUrRzg6D
siYqeTjfYrhEXb6wdll0meEMCmP4+Tmlz/mWnrXCyvIHBXPnWhbW9+feTGFJjGWVJYLs7mdP+67x
Wr7Mjrah8u+L86M78LTnGI3fa+dvwg+Qv1tWNAI0uNjphw9DAQIAm0UTLkO4FaF13Db6yOptYM/o
cAp59LghKz2kNhq7P0KlJ9nhB37odzSKM8aEt7orfELX7T9ZqcfhOYt0kWgoZKfp6ukRDuJvfPJ3
6cF3chmXs7oDJi1cdr84ap4mEm2eb+F1V8cEBcpr+dx+EAIkmWvvvblKIvhPFZN3liOnC+Ug8Xek
03sdohNsfcNbzChB1qSbQVVJikTm4INrYpJw/eKqTLHhPlmeYW9CB5yAXBY9NmSxDhu3z61/sBPM
FlPRYWdtVdxA2bgR00anhjfaDoxby33vCGV500TRuJMtPIBanS+3csb35cb+s8PPCqbZwHZ1cEbg
WGPgqOjC2P4J3FjLrC6tG/0o91eMObx4wHMyEAfWAjKCt8QVPw2nusl0rxO48+vcBk3t5OeMKJym
CvWhOH//EL/f3SKwknjmboAUwFct05vqU/BCxA5Sf/UTaMYYReI8BVg0EKTMNk0E0d8O5XNz89JK
MVoM14OdmVZ77XdteSUxEY6eR3PUFnsskP+BQ/aWt9043rae5JJm5OR76n8KfWg1+hrXT7H3q8J6
qjvNO6lFFZ0m9mnW/+E3RM8jb/QAvlqlyOHddtbFHE44vbRNvIPHusnzJLicQHpLPbXXfFLaL+5w
sc/M3bkufj3YTVB3Y09OiLjBpViIEJ+OScm6bZKUR2Y23VjuSTGlXIAXYzi3F3rNRP64RlO9ZHrh
evW2IYXBUeKUhNGYGvmmM4hSICIxbSBz5Bd33PJGoBwiqXtpi5g+5MI8sdhJu4+26+iQi3RSYobk
n+Ytb/974rEFBDcp+QwCDPVXcEesdbxjqp3jeDuiigpK+hRkjnMZne3QZPHH6z1TG3LQs9Mfp0xu
gkdsc1VHNFulWu7gS0vsUXkjWIVlXTvtJNKJPdC9/tVX2Zqi30hbbxmt5gocgpdsEXHqf7YM2VC5
ugRH/N36gw4ISfRIGtfl7/wdEdHauLbdzdF55qC/di/XujVCWaP+MHmEOpTwbJQD2wNAl770EFWY
Cb27cXR844oiyCyHWz1Gzo8JKW8dY2uR0N4mSVhcWRxCyTogPJWzF+RY4a6R9fS0vEJpuD1dlHg4
UMSBOYpDjSRT3YzK7RIPNo1YhGCXPLDGLvsor02AhBGnWxNNeZ2gBX6D75/D21OA8QQEEVC6oA7m
TVO63xpHTTo+mSnAJkkzRkLe/YRdbg5KUjKxqqaP7JZH3GAjI9EDmOY8VzMtJX1g+e59jVhLBMJW
fAj+ti5JHYiLxbdw5jP7hB+g9Ihqmu9zODVxHKLBJVcjuWHFOeWSkFrCC/twBsijIIoTSWZO0AH3
r1NMjUl7QUqviA4k8DpwpcUZPW0bflV+tZRVacFEyCd+P56qIPSnEcm/Di2oILnYJTJHL2rWKwBu
gKy0eaD9KUEuWHg1EpVyKgK3PsXoqgdlTqOOVxeLNBpzQ/D+U7/TNwXztr/CP4dC7XTyKhSIXE4i
V3GuD8TB3V0pdUohu54YLNAi2MH33CthoRjSDUV1MCKPBhUVE15b6aLCJbjNFA999Y+uybVaRqTU
TA2XUOl+ptCi+cOmS5FQOmIJxTZZhj2FhJV0dqoWqkHLjS3aC+oqO3SVrEan7itiqPwBM/IS0Y5+
ewHs0qu/FSaZyP0LNzMXLhmUMBOs6Yu68hZbrw8us1Zkq5rcqV0I6r7hq+3suc0h5BselZQ3XCb3
wdFEnT6f0WTQfajUwohlbvhfFZabOrb/3T0DTheyBM9InS0f38izZYEHozQ+ra+BhH2PeUCyiu4U
lHBLKRVUvdHu7Xx8P3fSUYOnXJfTElv77kXmn3PTTeSHEX5j10TMIxvBBzrRxAmf+WRVsXHMzuUo
G2mmtfu/UICq2yCTU7ZDn+2ZjdhlzllyABQmBlen//RvH/zLqz9QmrLFST098qkh2SBtjK8i9bX4
hgGgr4eEgz9ATnAhoYJE0/769ZLTFcTPoRGbPB+5oc2IlUQgwYJFuZ9Uz9VcwF/M4Bygi7B76o/z
WWZyV5DtYvYysVhY0aXratfWmkzahjU67EoMet46rlRr67PMDRkImkazT2FMTp4BHZffXv+MW82V
uXSWzTSjHFo611fmpjJT11kCvuZLgGay6n9Xh7WZoraAExuYq4fkOgfocjaO3m/v2VkiNOXlxwcr
OElVhTBmzmw6TADeIfSkln8+Mm3rjIN7RJExBZyWEosBadKZwR5kjZj+8XMmDHF7t5Cozh3PD6/C
i15HOh+wFHnqVvbnW1ZWgcA6h3MsCWBzzHfSUSs4Oemw/AvJ1K4rmYstUYDizh1MxRvbpA/KLJuG
yMQu+23ekHMbGU2xZ2+7TSiFpfhvsGEJKvzim/uJmHgLZi+Lr60Zo1PUuJsDXBn5pEhrPyDI+tvA
Oi3YFzp9R661jV02UxSyW+4LObyDO6eDGzOy2YKrq2eiJoS4ZS9w5ySR3of/X6noOTtdlCwzR1iu
e/BvISAvx8xdxLsBQc81weKrC6550x39KkuBI3AUxfXaUP9bsIXAEk+lGmzUC772KxHihhI8EWBj
TjCRWu4O0U82WJKiTS2AiaiC6PU50I6ljdVMp+awufHglNVF9jUqhwhcoyfy0yayMMpSX9vZSzc9
jm+qidq6iWU0wXhoARk/qRzv4ApGS4Yv6IUcDylrq3YJvtVOiJyk43a+/1xDODoeXqNIdG0Fbqki
kOytxME0AWOGJggj5VaDW9v4S6+WjvxSmWgOGk064E0Qvqsuy4xq3hqo0cJgK0I4VcQ0gjoQijXi
wRX4jGEIl7JNPnE8WdqRuM7Dgx2LVVC77gl1V7UMBn33DPH90UONmUVqLT807xSBAVUjNcB11G+Q
y3OZnARpT4zAsp5r7Hnuf+N9kDKxi101iX1cdVlt2mzJMhHpvSlMLgvzMP9mE0cA88YnM+6O2VeD
gDytqmJ5Fv3DW7bkIEamm7oDcnUZLJ2T34vPuFsfCCxjEPQwbiPtoTlJUuBznQNI9EmRPFSJew9O
YsWTQulrydaiC6WmokdfzEdBNDisBAfLEx8/x9sKYHwTSY390PsjBAjHAznzjyxWgyCACCPvaCaD
L/UdUlPDNiwucpk8jel8ibEtZAgnSP1wbwW/JvnmG7MMrx+78kpPukQD0SKRjhetwA1LXqL1xPYw
oCVZjSK7P9wFG9ro27YF5/mQ+W/8H1wq9VlRi0osCFG3i4RdLu3IG9jg/ouAVfQ2ccPqJ+g9hmkY
GFw/TK/1LtoDI76MjryZrPLJzFppWQeE+YHrpcmunB8fQ9jFzPrvHbg9nXapF/RHUcBV3360yt6T
1FRR2k/LaMrIqm1YAUN9E0Igjeiy+TmwouoSN4B47a4gvbjqaZqV23HyLgZiWRPcz1prWNKLLMAn
CwjCw80t1QFqv9xP6Z8tPS1x55OFaHL1e+XrJBis2bujc10CuoyZ+ZL9ap8nIl1VMRaENqEBW+FH
fYm4Q9gL11YFUa4Y5aAuBnfZLkPXd/1ffxiF+8oyD6S4YBnOoGMNMnnK+2hR4TNd6AlvGgNDW1b8
QUE3e+z20J67qyASe5uqCYXvYPpKtMkwAvMubaRArqmrnWyTw9x/7c5AmQHP7X8fzU9luo4VLUtS
vHktd9YXmW6RvWTPbMQw3YOMNNyBNAhWiflhHmc+LUs4q8ISDa+tKcUnYCiGbzK3w6G8+Nb4dIWD
mk1A8qP7EieHVceT++UcjGDn9OluTXcs30XBCB4Bq+j4Ab0G/3RyQDhJjMPi8w0PR8fwcmkxw9pR
vg1OnhUGkYhuDcbVZ9epkPM6G8vuZ3+ikQj445oJ9E+S3WTra3GB4QKTwSPvKUk8tPtE32cyWcOr
9OUkKUlQGNKNN+OqQefbTIOMlkUzuGb/cGP/h8BeYQhu5gJlgVkYq3ihqr1gCPzDx2JAx13V0bKp
dgxT59kNe78TzGX2zxnOnNlF0uLHCoBGmTyfjPz4tq/0TJtVbKWYZ3LjKOh9y3V3VK4c25i1weWJ
oAyA28EnzMmgSGd9x3Ab8MlYmxvoTEoeTvMF7lA5NteEbYfJN059RaFY9BaYTOFTJyAh7HithE/w
aCJGaJKJv5t6IoO8ThVD4FttAlx5ODQGzKxXe7eGaDSDkKaswRDxvd2bzRR053ostd3eyXRYTsuQ
VynRnjCfsWi0ERxvE0NkbNEGndBOWSIGJKTZQ4UOmDt7gp4nnLhnoNKnUxLLR/9vmI4gpnnVZBjl
D6ZLC8emRCJt7F6DpxsDXPuf740u6QSGkVCKS/HxaoAG3ecKUoimmQcOLg13YuLtWxDvnx1/yPCw
5GMuu4yQO7nNIdTlbDhUn3q/RmikeZssg71EiYZHIahyriKg+Sy/iiYDRzMTyImCWPFHkRFFJu5w
0YEcwjsZY8a3YSNvlkC6ZCwOxJdoOlpCqBK4MTuTFgy/LmWwl19a9H7Fd73Jr8MEyD1q/WwxAT3E
N4b2NzBrtu8FgYsXTVyiEMcCHw+BRZdO5Z7BdCOjDKucy5dn6kq5sNLodtJ3wYkzdu0ZgDXRsTtu
U0E/4wHy46quMUv/QONNeSnB+lI6OkxLcuWkIqAQbczmE7AZyPz5rkDdpKw1Ec6GhuPt+bR5vPrM
+Bj+FUKmZ3GfML9SnKt7tfiVUN2/20CHQvD3SPzfPSI5JSBgxGJQ2o3HQRohqcyQhZ+tq325xbDi
93WFxN3r3hQhpv0M1jUe3+YCAhofPIqxu5/c36Mh9YM/Zj7eEqVXHG87GBcZIx82qz1G7nqIQp+z
wFWh+GoY78gzU25u4v/kHiA0Mf6z+hSt6ciB+ydGkeyQQhvu7xhPTfZ0vzrq1lEQwVKPMemGkI0n
7YebCRpZUz5+bpYx88ULBShHsTuJ0j3xKne0MGi+mI/28j7HUv8lJYpnJiUtrI7EsyexegN0MM68
FdJP0scQfPxniRRuyqsoGmjMbbSO6L3vXOIFjaB1B8Z8/JHWgKD7kpjS6rmtvTZJMLk1gJNqtQGz
0Eht83LUIaLj/WDzWTTVKOQ+h9GsC23eapG+3wkBeZRsZjzgxggKPDLuvIfzIFJGupvu+OAlapSx
Jw/EyeoAO396lWKE+4kNg96IIwe3yhBaC8nbm+WKV405H2KwD///7+F0zpzuDnh8YAajmvzBglc3
LNg+/2d6EqXpTraRgA+Nc3pHfnjZnScqnNSBv4VRB/JBdsrEDMyRPjGEjyOcPkV5Y9EaPwb/sa4x
R3A9XsDkqYUaag34vc4KbjdC9HYCqB0p4x2mOrrnUYJezmWx970uBOQHixuT+gI7SIXhMyCIYRNz
8Y/cEtSmDr8KZtyqfc3Yju5xDnp+mjZhHI/9BVLBfYldRuae+/+dm6AOh8h+nEuZv3XOKRfghzyO
KSg7QEWeIDT8rSqNJVfaAmnoaQF6KiM8Syek/YkYpaIU36e9XApbxt0Sl6qF+t7c/h1Dvb0TVdw6
OSCxFqbB1DT+mgePbofDmtw0MI2dHwfweBw33gWz2GiJLmnL5Vhum91wO/oUrLTO2f2CbdWw7CL7
rjtoMAT0ttsV2MqNmkznF+GLGvoZE+iaqHDZ7HaJJHDz7tgdS7J9mzrZqUTKm4ql7Bb+0Cvo+fES
hedMfsanMejVrg1GdqhGThjSaOravAskA8IYZgV2IKXQ0YDrKNAfie9SYn0ru5q7kUTNjlnWU22D
IJNvWHS1d6+aj8Hqg4SCDF0My/9Sc1mf0ynk+Lnb2kRAdx7xqPDarJmYUknlqFpSo/UFWKgexl1G
mLWDIyb0zkVLRuSz0Mvz/yi4chzWx7lG0eIhaV26aW8DpOgeU433W2KDaqip0dyA3VXZ4dns3NKs
5WMzC3kRcvYGx8aXJ8wjqDLgwOx5b0OoNzXKoalELDzV3Kg9V5GEmWNI8bWkWgukxbnDaH0jLuLT
f5/hchRcoNb+Z2gbPz/W/RVX2OGfX/tLWwnjC8/lQKesAjd+S7t7AYO9sSScBQIKmxr56LSvIY08
DY/9X/Vvktd+y3liYdZfDz6uZzmwakk/EgOWhezrhkRZUyUFEppmZsmxoZiRG2mRPXall8zb6CO5
K1TiWbsW9WFGHH1mUn0dfcfv1uMkB1c3JIbvuXKBic0CI2KKna3EHEMwzVoOTgp81UTiHcu28Yog
kXbP+c4yM0Ha4ZJymqFLyIYJffxRBmn6rhG1LDuTX2Z9BjQSJRbbQLqBLF2nes01eNMv/PvbLHfl
DfwhpfjyDre83WSj+0k+XSx1zofjjVGUNPPsyjbF92b1WTgbJv9WFaVnQ9R8HMRfXn0tjQzCqWfC
tkH7K3qWM5TOD3mwz1aCY7Zv1EfqyGRqSk9+8XBLnL4xivLn2MIxv4ULVlCmlSsHtqu+X0sKtAdB
jXSEXnk23XvAOrnfsnT6BXJzt+Nl19fgUtDOfPfVTAUTFun64nmhM8ZBIIyk508ptOAiufH9L8Zh
ucWW6A9gzXYaC78hzqtURU2qWySbKW0KOQki+krFVweXZptOPmZNI7NNM+vd9f/htuadSJ6x5AgY
FycxDVtIZ4oeZcvRhc5cnDV39RZ3OfqU6Ol+InefozCOZi3hpbtc/mii29+DVLhPae/7nGFnsIs2
M/skNv7ew9zWu1Xp8VHOp9uaUI7YR647XX+fHliFWRT1at4Hxf3Ldh5sqrsFw/HadXHVGmHhuEfj
Z4IrSuTaYRa4bj62I1S+tJNTHxgKgqRwUXlEBK7wijmum0pEWvpvoxpLJKsHXR/AjCTTVGD0PI8B
FQTMaUMtYVhqWLlHcq80FRbRd+zp1m/fXYQ9GwNo7scb5eVpHM29iOiauWnFirG1h4u9XEqUKt0M
K1mICM/HZChD9uz11pEpmU7bP8LljZAeElDnI5RaYLDw+WOZ4iVm22yyfzRxv5aaJo18DB2lyPOg
5sVRaoSUpDod4WfMoH/XQDhXp8EpJftVvBLF9TKJBdTUWDsNwGQhi6cbUkQmcWJWVKU1u5yJVPdt
O6fnGM6G+rm1c8kwI6hbODniYmtjCoMzXSkPO+yE68fJCJ/543ES+62b2HDS146CwXAdw22vMG1U
dmVXteUJpWjpvx+4KjuWpbinfHUaPYXulkIPcQC8NCq7f5f8roY7KjZ0kMOdLXslSPWLaGr9uM7x
ysxiJxK/DROWY35zAzVsZF0kzn7zUn5ITbAm0FUB0JD8BjayugEsy3r8VnPtJfQULnLSO/Nh9ken
nfJwhsyoFZ5ShoAQ334SaQrkDKbQID6LVL4KH1yRZqertbYvDZOLucCWUU65XLfbcVoXRffu2hbP
SwGDJ+4ZYKowFKaaI02wdXn1DPaVcR7fP2FdkQv01WreFfjN/ipybeoh7nMKOo+DPL0ax+xRKv5V
LpNQewlFORBvnkJ1jcGoxdA8YMKYox43BwD9b+MY7WBy3+27u8mD2BV4e78PI9IhgPP1c6cRF3kB
9JFKHlrsRS52cBX9ggVvaETDmKfk3cpmuyA1+/KYrZg7BY+BjsiSiCoY7npv1F+dpPK99N0fxAHI
yUgXpN1/d+YGyLqYqj06hluoFavp+/VH5qDYXMnBK1aUGmdX9Lqt0y/clhREiegzUQwX4TRZTOFW
7b0dn0fGFkkYWW0OaeFuPfSL52TS488T8gnIUSdC/kbhlo0bl0yECuIMMfOLPpt6aS/7XoSNSlXC
pP8og0iVAOs8X+il8uVBbTqYEPKg5s7b/JTV/OA/Y6pTXuxZz2acGm2Bn8Bne3EN7+YB1Y7VjT96
JJpDf9OzinRIJHBvLvVlnsiYP7REbTAr5FbORVTWIyyyqMMeKShy0Kl9jScVECAIyetMhbtnQGql
Hfp2fjmc3UWbJb/z+szTb8c6D1n+3x+2fiA6+g24NQzOqb02wDe0vBiCA/mjTkFVMM59xuPCe3EJ
tWdO39pMqclPmouArHFDsINpQNzhsf+zy6PLjvNKKh2/5D947EM3fVpP27kIhciguZRZqUZpze+o
uJc4zct4xEQVPiMfkXfiaJAfofEWzyejnNU82JOSEB9A7WXka/o3EBi9KCb7ijxTfRiWpdBSyGVf
7Z145TQTJMgvvriXeBRnXohoD3fsrh4gTjyE5mgdpeobi3wwBDWxUGBZWsx/ZuOJrNkMrcVOcwtz
Vx5/pLduQl/KrNa+4MVq8qCX1Qaby1Wdbvsc1zQqj8rO3Bl3qe8ZPkzOyUGEl0dolj/5to1e0R47
2QJ5CCzC50g37l0mgpELHBHTqwbzq+MbbvY59NuGycDJW6Gkb2TtSQX1UW4RY8MHbwV7EB2sZX6+
iIolTTOizEywWEz+7xV/aspKHoxbrX5Dso4gYRVOzCCun3/p9JWC8/Y+7JTfHHFk1Lnh7WURE2cM
DB2hd4XtS81a68624iocBtL9sezVuazLF+bS1XGUuKMU9anKaPNB380IRFoawge0MT+TVpw0cer1
KFUkECIWdn8t8Hr5RyrrdIHiolQg51qf6ZJZ/KLtZK/JHOdQSxq4SHbYtzsFvMJgTnBbYAIiFCRK
2/Ucp+hV9lWmCwSNQrkyhklLWq7QeCV4b/6t7fPMC6hZmerVVPJIcXF+iuPMXBgB/VAq0a6VyrDs
YJPAOPLEeDG9YmNsw9fMBO2dC8ivfk64kqEOFW0gdNITvCfQcltLXz0s0pcDJPxCekSiFRBfhWdY
Qc/z16WtqcEbRfUtXR/a4pqK9X4p3KQT2T3aMlMwtQAoqytN/+4usFisahTHlWBnreHTul2DvfnE
CUFje0C5AAzjE9pk7hXficIaAU7sOjaiGZQlFd8tFv/uXe3C+RYTUNwBKHut6CIsDB5QtZ+F+u9p
nzJh2CzfxQhQiPlar+sTuhlCacwaezXc1paqISwN4YW18V/bIScUAVZuSlHf7G+yJ0forSWLrdZo
mPQCoEo0fg6Rn+M869Y1Mqlno20+WSxHbiuhtds/YzYX47Q44IH2h5rB/FuMuoRS5EUU6+iWaS6g
RzgyRkWcx/B3W3fsdaswLhOxdMGczS2Vb0VnPBdSX/QX3YKyDmVILAW7/KVVllq/v5qXaU0O0nJc
p2WpLOzSIFFUqYiJBgkBZLImtElKa6qPjTOu7yi7NjTrVQlyASiXXcv6RXPsnN0PM9XdtGe9E2y1
hJt2CwIZYHxCe+UbrZBe63MsNn8dxyOlCGs35CTyf5mcwPkQTnal8za6V+ij8/O0Lo+WYdEKrUjA
quEmpXdFDIB7lRdbzqIipJz5XPejLWaHgTKFfwZzgKpeVQjSWOg4a8HU2oRU4Pf2G/JX5ukuBf8R
lvJ45QfjV3MWBUKXMaV6DiXRgqJEWITnXjcSTYSQINRjdk5o66+8929WCFECHToBX8DSwxhJB80c
aqu3Yp8Sjwpab1lQwC4ofoHAJ7S7iuyksbP+h/quBGKPh6ZsHadyEngBWNStlHrgB76Q+9uxKAuw
ed6TdFGA3YZTS4d8AZOZBoeM9AumgL0k75r+/P5H27nRChzBqjrpSZcR9w8YA7icwyElenm8Ki0g
LoGtwrJIFoNIl+p+gKnZvbCNIt28ouQi/lro48zSPziIXh4bKHJe3FmaxYkR/OzClzi/qytSdNKl
O3vh1zVhgd0jSdeMPPU0BPVcBCktzlzvFfcLRNHOId4nyah9k+fGOQLvTgX459CZD5kDrOEU1fMl
khKK8NC9/WCwj/QkwD2oMA6fNc26TNG4tcdC/G4zSVjSJTjASMP2v0gWnJNzWtEU5APDJT02Nlpf
TntIzsAHJ9oB7mkwH89+HFWpZODVhi+B7D9sIRefY54ka1eF8QGgpso1JGu4/1KphTAOadXjYOVi
EH+MBcDdk8TDqQATpgvfHs0T1/cYn2gRHoTTkoiJY2rtYuwrq4pj7khYMC9kKm6Z1FvPokEuIRO0
Fn7rn552LNz+2WchqwBTw7EKvhD6BVmd5dWPR2/+QpH7tPbL+1PbLtGG8bmjIK0dbmpul9QzAgGA
Bo5WEMZ3AyBAB1mzdNkuU0++l1WOe2Nvvy1ch/2vocpk36ahGVNrVSH0ghnElewOTyUGcSr3Ftwg
Yqtacovid0JN2hfBkOk4vLGtASGOc9SyOc+X745FnqKxB6wSjAmDSuOJ9H5gyqEJYNroS1mBV53+
e+q34jeYGqrtLt5HOSYozv/Fpkhmea/Kamgmn5CKzrzjpQkmvNmYzcW/4RKql8LDCQW7RKxqptu0
QBMapWFMW7O8Zflc1vP8XM7HBkWJVsgiQ4DVj+jtuDs+m6117lSU7seGC9pw4lJ5URO8YZGIJ6T6
8H+yla6W3SkDWCoomdYL3/fzCb/H/wVAIpONM4UaqpjbYvMAWGHs2hv5ZN9GUYLJMZ5xr06yf22y
misYA+6YzhlR/wnWzynz8GTTCDZ2e7XSB5eTeEg3xcCr7/KMONFg92R2bJcOzQ56xjXbs2yIr3d+
kydbrwQ/L2oahNl/PfKobruotwv0nBcS6jqNh0bYYRVvjMvU2cffB6xLIbTzhFPpSWD+Lrj7sZJm
mdJ2z4sEXfeD/k8BrRO7qtFsd9mGcn32w6+dcjc6i2i/45ECFOpuntrFeK3gDc1fGZrGHJ3/NmC9
GIUuXIWe12os23OLVI7vzKjW8XtgZhVf+RWYljXOAV72UnhJCtR4sIrhC196lHXzK3x7eGe36bp7
Q2qgSZwjSnisQhIigk+ueCwbzzJY4QwxI4e5nMDEMTbAq2NUHev2ZFJO8Yagxiv5Fzsduwi6rtmh
92mC/REp4b7yNKWGogtYnFB9Gw9+NEnOPnC32IXhlPyLHD0AU3Q8HbncjQTJY30+EznSK1EDcocJ
2mJrVmDbdaII7QDeKPE5WVNIGyVklGE4YsJumYr7zbQmfT0avagaO1M4Mtb3tYZYsoPCzoWNLQrI
oyrqkVkk/Dgf5604aGvu89nEGcN87d6o92nL5aiuBo4Euf4jmatP3NTTHk5jlj1cb9qeFnD0Fr1q
XWrbFc2NvrLmXkoIOHmJ3JJO07uVP2ARsqL5T35Zq8ftpd6F9ou+lGq0IwCY8P23+YUHOQtLXavR
5a2AldGCnggwVr48AQ7K4+DeOboUu/lQsnApVfrB/0uf0EgejCp0nzxyHPx1EZkC3nk05o/jNX9a
mYwZs0oo7R9AtRTTGjSWAjcKDbBQ+KD6CTfGBtw2DIKT0HdRJlAHnQTL9X0n+iLQ6NvmjJAm+z2T
ViDm8AyjmaEShq3OC/Te58eK2/LblOImEK0SG6OusjCqeqG0nM++LRirjQssS3q3cmPd0gXf+1Bb
vrndzOfzQdrHFocs6dH8v90cHPneivZHXSqxeB41KrcXitRpwVxKSxrmsWzJlcHYosU9Rej+qtnY
op+/e8pLLzc/sb2ffo6OprUKhfSSHjXhMNnKLiIa5GHbjdDfapoL+Ny0LVXOlhric/TnobM8d/Yk
PCGej27CnIL4f+3XblUu46lFsYhKmujbhz28DZU7zOPrMOOCVVXvTCYm95Z1kCudi3K6eK9grFxD
G6140CSygn3SmEdBGdy/pqRBiceaCiq3IZz8qyNRrOutkE/HJkg8I/h5VdOFDfVQWuGUCRqLmu0j
1UGcUzrqDBrSg+VekK+eRbyrlfMKJqOCdrf22e3oDdkttvMdPAVWV6ij6vC7A00Pc/zjLXXn5Oa5
fO/otmmNB8er3EdSe/3+MyFN86sL6ofy2q7SLT3Ailk1UhRpbdyaDGbNBNHN3rJLU4haPbVQiniq
tg39W2XzwkYI1QYks8phf7oO1kdxmBvxd1QcS0tF/9CiwzhzuzjTYMioxWjEZY0HI1BlnAAU6LmD
Gld+LwzlCgY4GW71TWhwgfcCrGyR/T4oeHPcurMn/i1aCsMuD6FBIXTy9xjrjFNk9HUYH3OP10n2
Q0N7U9YymCGA2NhNuO8jGF/sgjndr++tSXmin/0qiGC979CjaX60IgS/uxT81weNMO0HjSgPtsB5
EbdOw8BdN8YUlF0Pt4oYZyYPh0L94D9whj2wTFZ7xH8BgcXoU+haMKk+5T+Xq8yGmtQiwLVqfYSP
/uzuvUasK1VfQksxg6yyxBH3Vpxv9PnDvAnRj2yb26nis0IFv6K5lldFBFoFquJKCuesjBXw3yrj
aeu3R/7Y9Cl1KbcECs5Z6vCXoaFn6jL2kMlziUKTeDntBPhkBqnN0CM9dXFDEEHmgPPAKJx51VGM
YUOZUcr/n59dS57moQseHjktfP1BvA12U0ie8xpG9deZYBvc8DBnBCJPW4vFb1f+58BBEeE0OBik
+JJpnp0Dp/8MpXB0ncH6f3CWTQY8zV/OfreeJhfKkptYSoP+k+N8osivWEUNMgHCZajWv53vUCA6
kTT77x/Jo3bD+gARVLfiXvd2llw9bKQGIV65fjqgqotxafMirRaoUmj3t2XrH1jlfILn3qGDP7Mk
wttYuDM/1lMMXiAl1VH6XDIAswBH+07ElpI06RTGpXVPCnU8ACpJdFw0y5xssM8p350rH6V14j9D
8cEH00XsdXrmveqI7lHiemdlcxntfHgMvAdxi8gA32gThIWt0r/RGpm7qR7qP6rFpGR4cjfS27sZ
tF7Qt2i0QiIslpuorYjRoCRyPV3oXrI00XkyFqqDpdmT0wau7QuKbt//Zc+OSaXdvPHN8fYOpX4b
mjm+IzZo6JEBTzwvr1PhmZKvRDgj80DSFYzvoPZ+Th7dgka4l6Lo2BKZaZ6qmcDPrMaoiVIsAw/l
Ri5CiVVmuVv80NHmmsUN2aPMdUHeFZJS/kcY7NLFwQKYo57k3aPbMs98EI/VaGFzqXBfgZUnFEia
fEsGWPw6/Zf0YjpCWZouy5xMhlifYSNdxEkU1X0zsVUd+KECK/jr0evTxhjynE/Kmfzkwgs66H4b
HAODL2z97TYG/T7m8iw69dApFcjkA0CKX3eeLTmsYBcfUnOll/XLIeWVXKpMEhcWkx9KUtxOymBq
kXAdMM8TE7+R6f234aAXBlgXockASBk31xg40qopw77KDyM32CSpPudvzot0hfnwbStsKZCZ7y2x
g0fGpBMDcDR2SxRIf6PL3Vr8SKBMzkemU4shJvb24HE6q8DdJ3WIWfrniaYDsxdEUzPAj2oVnJBj
UUbeFCDa1k6kfZwE54RuNolWW3Z99FVZcI/YDpaUoyTQqWQ0i7mWuo7bw6kHFF0WDWKdEUUa9r5e
TmeBSm6VI9/7VLPUp4HN/mtXNLBC14KkJphIOQz+XyproYrn5U82+c4X1s7Eo9c0noSn6HWp3CDg
IMA2rpPbpgoqxKj4xUjO6o/2cnUqhNbZSNEu38muhdsUhcPSgrCm9L0efuh8MveiQxQZHc/7SVTk
PiuRblqpoe4N8VuFwYieiQjwTsyHL/CZUV5BPu25Lr/G4TBvVu05Lutc1nNzsy+jBmewJus9MyXT
yn9o4ARdww4sJlH+Amb4AkqeSZd7SuwBo08xDpVPhfN7C8KXFSsll3JrHeopSWWxyLYvFCJvjOjh
RgZteH5YAioX2qvNkh0P4jcimEjWkj4GysjppZtvxOs4qytNC4pZUsW97Y+F3NyjvigqCUXf6cb8
Vn34d+WOIEOtG0qYRiMbgcmiSoBqZyJNtOU1WQF31NIhj3102iLHeDIdf8Tpl7h+ChjlcXKgkPDd
MxBq4s3yHTkUd5DdCSj0o7ZHAiLmjXi0gr/maYsOToJiqw61SqSFSBRDv2NSDSsSdmgTqJPNTsbV
51kTXNhS9tTqJxRVT4i0/z17JFNUe/3cZuo+4xW1pLRQbM1AwVHejvzqzG/6IKE/S9TmtNAGtNdg
OSz46YNxsRcvs1NfdSNYX2/sPYfKtbPn4hnIE93olsrLo1jLA6gpTy8XJ31m07eB5PVLWSWGfNdE
y3OgfOByFUG5VaRxwaHZUCm3d737//C0xYpbz1atmD51l9n8QZCVMd4/4NnQrb1GZeeEuVoy+ir6
GPF3jns6witYKrjqzWd0xygsBpnjLB9KLBnxTfvg68MNGmQreJlyss8i45jZvzpqPFgPIW1Zzav8
OZg3ZvtGK/FqU+jQ/QTzzl6x32AbnhsT3UBPE41KyquK3PjWQH4IUgjkNPAP+mba8pfR3vE5aGLq
HVU/85XyXOOiNh0oT5dFjcNS6XaXdTEyz8N8fgP5zk7w+pjsgztrSSfvAdaLj0tIKRe7p/dmHzBe
lSKHlA90dE0MDQLzMoQ37nnQwdA74jK9p9NIS3oEd7DMH5ylRh487La+2JmkVthdm9qmO7BApyuZ
o/fknvOiySbURN09peQE9akRddb3FwsJUZ8H8dXDfwo7oQqfOorbpdosCawd6tpFXDb7KicfY8PE
uVLt4vXYyq4h53w2q8t/suSGgjvuu4oljeQEDJgLAr4PWiBavYmE44zEjyrfKXQRp2jJEvxXLG+/
VOm7nsAZLyc12S7gmJsLINbUORyBc/vEC4pS4meUtmDtbOSn6nSRchRJodr8QtaTzDsEduJsWVsQ
INhC8iatZ1g7wQ2+MxOXykti3wd3hhEEpvfLDwYXMPxJjtrEd2QM9guHyt1f85cbSlIl0nj0flsg
eASUUVB4JqXe8Vz4i7LRmFMki1rlaLvfReI1Hn+eINMlSdb640pIZySnUS6rQk1zYeG3G7hyociq
oZHga8rwRD4uzG6ZePxx8FjDlIvJXLNui6TWil/fQzttkJ/ZwUfKs6KArfqUgZXLKzrW19VEEMMx
SKDXYfgVxGMop2dW/Qn/WyT4La/Gs9OJsXoR+ejWN0Ps/XxLKLA6aUvD9RfG5CCMuzEZkxkKlg62
WGCsRwOFcwIVHQBBEsdWzu+xTon8rswuc1MRPy6cpSbhY3w+87/mepmWrTCQc7eif/MGKZJ1LP2i
xWgkvftdBGSzUj2dAgJpTEltLx341gEghGoSPq8iFyRlLE+xy0KGCNVISHvIktyIprVCVMytyRdY
j2OePQt4OrjZMaeEmaucxZN2qblZ84YWHgys84HHMaFFdxBWUxHghGetdn0BdXDY8o8azO9PV8DJ
WZzbBTmpBw+UXBYa04jkriMQF1HONSeuIaj2L8x/ZytEkIpHzAMl4hRifYvvd3yMKjzauSsVSSzS
DNSAUYREPY+gHbjZb7M/N4dUeTKooLZEfLU3hKL+rKGHkHbHr4pXzS41/fYAs4ndDcqEGyXsIEuj
vR6141OLrEM69R/OVmpK4QA64o/br181wnBNEOtKKiwSpU4RnP3Q0VekD/Eexg0ZV9EUnZwFfTO2
UyCNX1OQRo/MY4+N8IpXMHQI/Chf7i+bj8ukyOwUo99FwCFydzbTsDgoEA4ipJc21YTAkR4XXvf2
Nqf1dW/v2a2FoCPpJ+VOW+7rnE2cS03V+R/dpX132Ef5IYQAjJ2tBW9SDiDy6LOc1FeRbEwqrgBT
NTtuA0+fu0cMGUOue9M1nO3UDRNrWJuHbs8ZVSn7Kl0NOX+UnH2BbaJ19X78p7to7JLY9RTrYykr
vBk3ibwq9ttBdBmAJtoQYwQqNwfM7qluQedp1wB9d39g4CbEq/dM3j7jW23Uy3IuRUeFTMQjeHJz
rk239619u9gQQZk55NalBfbjTj8j8DTPMBXHPx09/hfkg3fQvBT/hQSHzbIOOaz39M+gq+YauBQW
0SyPQ2S2Y4LE191PcxPp7WXx7O4PbtvI2QammFa+rP3aoeyPLYtkSDyUjhniZU2524oSEn+IcLUZ
EOSVHI4iDQjsGXvg5r8xzJLwApz69vl7bWJ7fvnhuTh/RPur8H10BkucSp0DYdOe0lQqusDSh9Oj
1O/rCQwjsDtjg351NhaR+RySgjbCWMOUd8v2/kFWWa/a0Hu6rnBHKKZ2yYnYdQFDcR9vvobr5UsG
F0ZA6078ONbnLeoHm7+Bsrlyo3ApGBHVLzUZAfbTrjY9gULdianP1J3h+mePH6I/04Rxj74aRy44
t+G0K5QDyzKZF33gHg1K4WB4pY+XJBO9x3X6d9+wtkNAc/8qJIIyE8LETQCBnSAc0IkJ/hO4gB7q
DsunOoO33RBS7ZwBZ5rmT8ybt/WBx6E02+JIoF10ledA+PKq0SgXu0leC9tJFAs80GHqvLDxhLEc
5hOUkk7EEkxxRhg0cIDVynrbBrNriXrggqgSZ5kPnvA0ACPCUAh6yWTAWzAmBgpuv3MyKf8JYqCG
3l4whQ8XrWL9ekHjpJQy4t16Wm7igeyu4OJS9ieJtB8/lbyl79k0/pbaYmPUX0hQT9U23t6bE5K2
mqvIBE0vJOCyfwVJmSYi7QFrobb/de/M/BqisJ5ShvInoUitxancvE45ZGYPv6BDmKAC6HsbElfi
DJ1giL5PCJWWh8VYFfLr5cxDTVZndkLhpdt3eSzqUIfdRSNIEQDUhdfJ1C0uDc3bDdYCtyYcMlGS
ElhZlJWo8Pr2C36/F01zrOryS4OAWqrxKrHAbP1MyrLAKmgrpEtr0FxZHKyKxaMdo3ld3SfjcNW1
akvGuBDax0LdG6MMWz/qVKfxnUbtqaKCk11NG1ecdGy0AFQb/gNpFkjBlK7Iu70luNTSA9ANgU5m
4lyacP6mJ5A/B83f8Tw0Y2kCfUr34rD3txmswWN8FeRG4s/jOmGAVE23Nh8Mynjt9SqmIefJSzEB
bE49eO3pa8ZmfVZ73Xe8KkTGImo7KujNucjUReEKnoIPc2Y0z0UBjpgTV6xBDVQUQffaoVYJ8oAx
A6twYKitT0fnOExIXfiCLfB/bRWqhZtZ0Qz9gwdSXMYB6iB18/AVfJr+7pQO0STlMLsUVt718h0i
Jv5LxRFQU+GjvnrKZRkgJWIY0aiZHj6j1BJ/rzW6nY/P74A5Y5tl58UU2pmCS+LxdnJ200XKhnow
lURrdjlreTUuD/NYAjVHU2bHfRE3613RPO/beg2PgbRhVR+3LQzBzwi80+tG4AnoTdcdTAZckd1i
kILow4Q3vjKffZY+sLzQpG94Fn8WmDdHdsAJhfUKHIUaqUoqp2u40JQx5Pd7RwGR5/XU71BdTDBx
AjZy2wFFrk38mDzp3x2qq/25bx8qazvtPobnge28bIQTnYeFq+j/gbjhcVhQo/7Wv3wKHlvMJ58q
BcS6z3Wt5YPzzDwAoxWuhNylpvmhgWeg50UEiHe5vSr/AoG1DCm243omA8fEx/72jlxx3m8x49F+
zMwNnLLO3OUxHQBZSGBTfJ5xu2cZqt0ESAx7Hh8Amc6fHyZ+f+4cuWYXsJzV0o9TJ1RJs5UxAhpc
ZOBdO3IYXVJbV8imnkO1zTm0q2qV+HEG28svOG1K8rv7Tt4CEsqhjx4bXfKu9M8e1criJzyRWmal
by3+G6guD/iPnAKJaFTTLjjYOqZK1MHk+4+IRVpuB25qWTwT0YxYK4XAynpuWIf39B5hMIQP4DTF
3nthmy5Bu2cC64BLLhX/Qg+wcBE98q3Jbi+ECyGGy5gHHi39Vks2vWieqcveytjalEJf7GFU4XA/
K5DzVSlW/Kmiob7wQtAhMQh18d4vvsXfKL9vU4bM7cUxDTfADHX6BjN3nOOtmJnvIF5Irl9cCDfO
RIdZJ5GnwishjBpFXdzq5Kpul2nG3lgtWDvN85m3ogz20I7ap8mQh/S2h5P6LgwPRvd5GBa5io42
v0Hflj/i2HaWfXy/Fq2dpCyrAH8i1+UazQSPg8Zs9KT6bsuIvpmwO7/d4whbyeUzv4VQgB8KRLkm
rq1yAkKFePxv8PRbBIEpNtHlPlmgVE5ztKtq4BBmPvRLnk7pf9a6CXVPpqNEky1pQABr9yQvlOt8
Sv69HbjG3BfJmYhkFAtxdwXykTrp49QWp71kuekzuXJoytL2XmxF5ArkWUo1EKM31A3faD8FiXi+
ci3XM4Tyz68sBQ3dvofO9UNr98NcFFtBolzfEJZa0pchqC6+jhgYI7TENe2NMo0uV1/Mgd9Z6pS0
ptk9j0Hx5OFKSHoeldDPM5nr7KVrdQT38a0qjDvahpncWLKwny+yi2BapSAc6DfTB4d73EyO51GG
uUn97sej9FkXV219CrJWBXeRiOjipf1c48iSAfIOkPnbOPUUzUfqOE4h4CiLxf2oQ5rsndwL5OYn
f3n9F0MGuL4gTlg30Le7Q+6PFu1yFognU4hX75vZu8ImkhOEYr8CT5mhaHTfBONH9aLt4ocbk1tw
aO/kAM7laiZxC+g9dBn2/rEYQF8/1r3FpJ5hKurA1Ep88UxX7vFp2aJ9fndm8YFiyL3fP+eEVZDx
/l2ME58sFKz3VX7gtPC+RmLeVQLfOsN0vuQN3NjmNRflnEJva3sKP/uq+xhc7ESaLYMmAYLjffnG
3nSIs1f3TRDLSUia6/Kq6PYaYAPzLk9ZVuleswhZU6QSIzY6U7HZJMK2EhINXClVWTN7Y1Hqm+Hu
Zst6lL4Gn4sc9s0bV/bRH+8d1wZNkg9B2wmNHBk1JOC9IRbUiQC9Mz18fqF2a2rNBG+s2SecAny0
31anoWMA6xhGetrEo7cgJYF4SjPFr9NWH4SO0Lg2k8KVeROLsHwwunANSiBXH2hfWAbq5jJcfJA+
Mo+uQotseCUMpJczrUAqe2Z56DcpjghruPVS6KR8wd3tlKUy0VuLmXDnxpOuPtcXbk7+yH5DW7oi
YJ75hffeHVvK6E7ZiIX1GE+D1GDEJICIUwao4+BekanPl6vYYYNbsV/lhkxFbrHwQWoGqHB4fBcI
pF3my9pwYDpPPhMUs9iMpH+MLMeji0BgY7WVsjgClpQjqfvQU7r9Yb3iDJOpe/zqLVlaOnSWXy2N
dGufjHI8tjNJTY3xbcg2cLA9NSZoabp1+Uv3ci3P3IoZOoChy7S5KaPooUtkpSuXgoGFPQimHLCb
0YqSU+fzUXNhOLiGbBmLiKu+6nReadKT/oiP0T1+YzfOrxDgqBJCQTXbzMucifrFac5BfFd2QG7F
X2QCMBj6IRLILc/mD4wGableORt0Je9jIkIUvGLNjcCpHUnF+cUfZVSct3Wyd/Ids7xLDfKQ5E99
XtYxb1kfWrrEPAHNTTiym7bbi/ICj4KdAqB6pHQSQoSFzg3Zmb3Z/L0O1rA/8lYwCf23IhNQ+WuF
bvnqNZBCmZmoLHxgXF5m3pbDh6ItYHlROIJW1C7pZjaStmoy73BS9dC0Z5sUQZ41ssq+iyfxGRsk
KXJ+TthhIYb6DrNzrZeGzv7nlrpS3cq7glv8YQ2miU55awZeP8Cucb0GjgwTz4i9Duesth2Yc5Ks
W2LYAm8+WvRzZyiyvQwc9s9/ad4uRLwdBRPt/cc+v6eJQoep0W0JkJQCpupR7JSl/6PBwBdGnMIr
SXXAEr3GCRouYnwJ7if9qXlyP2Uc9Y7XzJkwECAt/edNP5aMceeO6rFj9Dh2QD1SyekY/REcWDEK
oFoge6xNZ1WhElsO2wOUhpfZCwSdLh0T8AKaVp7UON4/9c4G47cRt07ihRjQwjY7bkIfgB3IgCMx
YSaKoRTO7VBF5aLOxND1tstvNDIwvpCwfcF6noXyim00eUVwVKT0nHPcwiSRgLaP/WtGa7e6xkBw
vX80LgJaHu2O0VQqRoBdVvOe9RpctGXQLe9d6kUvHUGKHWSNdahMhxHT7GFsFT3XLe0LSCp+gmss
2eyPDeXV/b7yMKXb1mhMzhKO71Ikxxnf8Az1P9/weGbgu9JRc15DO86PCc7Zw7xB5x6yZuawngKF
gzhwHUqjpRVOWahCVEqVKtN5gb5hpXNOS+MJt+WTjpJdj/6QB93ZH1xUfRutHmVxESGhUJX7KVwZ
/0/b99R36sHTKCUC1EFI1BjIVXx4I1+rkzctWycihEVuIP5gf7Ob1cuPR4X6LVCMIVD3JBcP8LUo
x5daBXQAlW44WWbTRJZSy3wbTH2QOHe/sjchROJ+4Wvgy9g5Le3d4gSMqx8gYPBWSWv22eB5jG+N
K0awm8RM8GrFyonX0mCU3bCIauBokIrmeoDxNuP+OCTahfW8kY26ZzG6qMOhEf0zvGEynX8z1pir
5kk1EUev1KsS+m526G854ijCQ66ZIb7zD3GsH04A+hxexMbMkpLpBrLCS0xkqWBfm21k/2QWUE/J
KJVmx9imQ41wGHfS1kyE85I5jsUr6m3GcfupBF64NYH71tdbE/mspqfmtX4p+fOtfDo39UdxZsEW
XZWdoV/RzcCJQUh8A/cnXOTZNjg1rZtLiSGE/OLyytDTpPA1xBZKLWiBQHyGM9D3q3Hc7fved7YI
/wdUZOca0NCj06WgY/V0Nhfq5gX62PjTr1hWauWhsGizm3OEFACMSgT23k5rMlr1JcHDyBt2yVO1
LblKeGJ+1TJi5jYWrLpRZKiR0oDYIP3AAWXVBBw3aHHRvwexfmX1Ya9Y5DAv0qhmcxHcrXofz6Bn
rHZNIpb6Tf3rKu5YfIC0NjYYw+cDT4ZMSVYXYpce7TAP+oyYaeuVnhI+5tMM6VgGHvcDz7TwHaHx
2+e/phODRPKznv0QepNDyDIIRHPb8GaZ5VsmPF99OoUITNyPNuYwKJReqbY6b+3RrxfGHPhcAzu+
VhKHOIh4rNQHQEsutBuB4RQV11i0o7gL6SRYPlXv1YRXJYLKXkZjEuubEHkIVz9Z7L9QEfb0T7vm
fVEloaGEkTlQqT/M7xPWVojZ7Pc6Jyh8vu40uqb5kCvpFC/T9Ud5ReyexX5bOj3OkS+WGBv7Zf1R
rnhHm5VUvUn4heXfrmZuNlAhag99Aq/6AyhBpWIsVVdFvr9gmNw/J+if6HQo9cOhsRL9MypW2MjR
g/KxbgQZCCoN20V1NzgSTioAHnUCfP8tHmA0g0XdGHaRqdQsjSEOzNDErdbMq5im500wCevVwsF6
r/CwSWmicIA3yvFT0GsJ5CmauQBCTRMSNdf4x7PSlmrGjFBVXj0SeDua4MJaVk2KPxrrzWJ+CgBw
J3CQOy1BUGWp4xFrroFy6rdE8C1G3ICBhRGmMd3N/0nKDeBdgOqas1WYpAkMWLJWuYdn2mTfibNQ
oCqnC/8L2INZnMJYFLxRyxtWDxgXXSwrpFfjeGaQ92IQ3bwlmvg5qbt9+M7KqN/UisRnmZ0xwvn0
H3HV21B17GrY16ySaHtOjMQWtu9CAJRoOvFqc0hXCn7ffpbq2Q/PTTGPz7T9t2rwYParA4g9hNgm
UswpGr/sefQc1173hs0udknZuI7BtkQ9f9he2p87fr9YapNVf6njZUI57qWcTRqrMEdk7gD8tWBU
a0+yXs9Rh7ohJ6U/Q5eOZKsrPh31NS/b7CXMJnc/YaJx+661eUhuOUwDwYd3vFyFEdNv8Dzg5n7j
2kPGLWGq+GUtBk7LigBJ6BcBaL2+2Hv+CXIfs6OhmyeHNz+t2MyOVmTkvDPyHYnR+Li+dcHe2eNA
eaa1+drBbk0mi4mDZyyZntMlkkLIzO9Wz6VrSRUTDVHDvcE+oCy2gazEOaAuR9tV1qRRM9tmrZhC
2aZxc6uBz3QLnNHwSA81g3TTtc3F+qRL5PnOeNz/tGplHoTBZ23GCNnUwryJlrKvdRvzobunrmEE
T+UEGmgEIiHx07k8L2Fp/sMocDp4WIWIWberwd8dBAds4DcBKMVthgw4nR3OLdCHKTel2ok16RuO
SbO7A2R3mv6y8Oug5+jmLbPN4GtRqAkIocZVEDpJp+OUw6I0yDGC6D5lOzmX/PsLbu5VNN41VztU
sveo2li4R0gL8+dnL0jgeNJidbtThY19t255U0ZufhnnOaodP4Ot9HDzfhnPABUIHPYuTB6TTnvi
WqMhO0agiK4GMyu69IhA5PxuGjPEyCJzndHXn/qayudMVx6KZeMAmgR2MpF/w7m00a6v3F5BcSXj
f7enkLzeRxCGOfgpe6MKX8U97dlFkd89bvJLl3pVsSelqz4xmDBLBvkPNFjy8Y0Y1W7VKhKmLnAo
Foiqka+Yc+VC76bsDnOaB/VUQQuNV+RCqueVrMGLbCQZSS38VdT51cGEqlaU0D4Ga8MboBtu7M3N
pFG1ol1aWQqOe1mYK6CmXzjDim1etDzk9WTdzFFO4WDSvKQ+B5JIrYmW2OWeqlVQWoOhfYq49pit
tBHltIvYq0YhxWgqM5i7+0WO2K+a9IchofUWhuxnsosU954bIJO1NQaol/yOEFpp/y1uviUBRn1p
DN35Jp6H58fNZ37CRFRCVOd/mZAY4ljuxM3gPBiqHHlvW0voDCB1LfqFHH7qsOFA+9nVkzaRf4Tz
BYFN0dFyIinsXWYH2Gyqc9W7CPiU+0yYX5J+KoRUxsoCVdTVpmBkjCqk17fx+iyS7KD7l1ReIm/4
+yPezSabwQuLIeYXbP3q/GwmeJ7LkdJcGD2uwhdE+Xh4Nvp6/Z/nqnjFRzCf6UXIAfJri/n5ZbdL
SfPT3B35Hk4Pow6L72dHgnSbtrp9WFQYBY8vi9CY2jYRoWf6dBxzHFYS4ePfv6XxmZZYPfTTHDER
4hYEp0RmtRFkfo/QAKoicVXHcfe9GA6U2vkkwsf2rpJWPwm3/jEL5Ib998CQw82Ugr5vIRIIqbD9
P+yCqfEVX4dMuvTwPXCSR19lFbaTGGXcs3VKjCMZmSnwCNwZF5jrjDSCtogOQexRR0+h0KVM/QjD
gk7U+P0zb2h8bWFCnjuGG3L8xyokNtNT74lxZSlnv4JP/Dp4zl6j9BvuRKdQuXHcpBua1E2nEEED
87ZFPkUJC/ximRvRcbJBf0/zMETYl4NfB+/GBjR5ooQNWt6qj1UnzrWIItbkLMGwa+zA/HU+rfuC
B45qJaj/BktIlnNnq6S2dBM61vCG88+FRa3bTcLtHtrn/2SdzjUWN9vRR5kwsxj5yhKjLP5nOiwg
HJib4S0kDNaGuHj5S9ew+FRna61YQwIvDVM2X5jlsdB7Ubhy5zQB6e83v9b9vBZY5FJ8tY6rpvxr
qou6MAaYjHgbpwpXmkdDBsN3DBzanFEQ0GTXbtBP+ysnGYwa8SKcnRCY9Wmu7SfpQSImqD2NP4/U
ZWfkS9c3k72cSkTJkQGT6sxHuvLB3IFGWIynIlpc4xNrI1qoeYwazpzw0CkUaYjttbRbIdIhfkQX
74nWPHK3+P8g2blpu1gnsXlw0ZrDbKNwva2zcEVRY6F8c5spbEnjVjykU3711OpFF7+lgmdordqs
W/kMoJAo5N4H0pnBlBjips7AvBNGwGfM3wmQ6FrB/FSaut/Pu5DhRhmzd4n+Iw/V4gGzhTyAP3tP
dcq/hFb7CiNgU+jpb+kYGWBPyYa3Gbef3trCiwt85ORLmClMNt2Qh538Mur+yHsAsBNxuKI+Z2Dl
1GmmkSFIh7tn3B1Zhox+cMBC224PUZ8QpBGA4k1TkAVgblazQtSXMjh1pNgNlD05bLwaYJyUVObl
pXE7dW39765JaYlD44MaZBBY3/r5dKli/IdCdVQa7dKiZF6YpEP6C88BcdSGuvt3KN1cmYT2PCxI
HrLO8BtdBQ5wfuo4uDD8pKktYEajVTlCo34Gu3cI2S/V6CIaagDglqPAzcKGwasLnkQH/UdxoDBL
nUvP31dZQhoD/iMZ3T1aqqYNst6Wku5s3N4Krfrd54lFfOYsz2HEgQXr1wEs1u1846FQiTVA8fOa
tjEgeDzURtyODhW3Oa8jmylMVF9+/4z4CKS+wrORNWYljYyxfJXAz6Rp8FMar2Jw1Uqd5T73QGUh
Y/eolFoqDn075qE5Tyld+4P4axkGyVukY+7WVvJSv2YqKuAww0Nr74+VGmRtrqrAe/VnOjOovQu5
oGZ0rB18oPoLEBEL6azVK79J6pGaQotToU82AvinkhdfT7plgVB+NCrXiwE00sSev30E74YbHA/g
4bmZxgu2tfo/nV4cYNkC+YpgKD2w+WF5tWdSA3YAQPNgP8Dz8L0cRdjPijqqsPsX6KjMWiQd4klZ
ewgDQtbD6n+4aL2sr1HFM1c6OOd0yV63eXmSFEO7sEVoykNTwgBydSgovNHEF6kYZ8p9xQz/1kp+
i/4N3BOvJnczgr91F73UBIzCR5IK6v60k4s8vYxeKOpprNH7xYNdRTnGjhMki6IJWPA3Kw4TDDP8
VSib292DG8GFKkZjkvpyi2rtqVfDqUng/VVzymse11okjfH21o+ORYTb+YZeSFxPc2XrawapFif/
0vmvJBHYU847F9WlHlwVM5/06Mxeayy3gvZFNNFC7rq4yikAFm3ynertaMV6fi1wpOdt0uYXcRp+
nU7GI0Zr9bEmv/HWiaIL/GiiA8swNC1SSnpXUgd4culWlKc+25/Ni8Ss5SpkXcOplaLWuFWuMcIL
tmmqsoTxNxPiHRP/sdyZr+8BwZfQGKu18zLslz0+gs8Czi+pBsCGf9NHxbIuuJghgusJmHRyBxbd
6yO3JoooszednSqycZeD0+rxJap6uVfcpmNtWnMB6ublcKeHHTtdj8kXDtXKPauGzwEj4slyxbcN
UxD+2UHvBXRZu1UCtNzOIB+7q/JXnZqk/EMX1Y9y2qWYg71cMtzTRfY10xF32qAIiE4nAbeT+BWq
srUdM1Oawgo8OcE68+/YSTrygkZZknIu8pi+cqd9wEhErlAqmAZ/OEcvOjOQdn+k5891kp72jAb+
gVaeKzERWOn/Nc6mIBEQn+6IrDs1+i6HSxeCNiNKnv7mV/yPXxc5/BTDvsGlJwg/ZGmA9dH3GVaz
b/ey2FGjFAZtiFUMFWONFkueBlIYEBDD7pQMuT5pSMyQzNGUbGkwWr1X5429Sdmw5OoDocuU/3Cb
l85ekKRIYCPyKGKIlLUq5CpA6E2F5UKccpo8apm7JvbbtmY+Sh5p9HiBZPfUS7GhqOW6jQGE4+dp
GW17W2aWa1ScO/sD05Ua+T9R7dtWt6eI0TjA3V5fo/lzkGR6A2NH8WDMHXS6P/AvJYl0JEnXF4vc
+uJobfeY1xok3Ef1PgdwikwS2uovRQKjnpiK70HdCmyIvkaN71J8lMlvVih6O7AhsmzG4pOblxLZ
vyKbvog3TYlfFvuCcE/kwDhC6tkojJGiCn4XqP/zzbrT/6yVYrCTkIw31fF6bjAql6Q+xz7otKg2
ZS/AqLjQm3KeOgCUi4sALAxwJ9eGsRK7bmF1V93rq/n7Uh6RQHnzB9xY3OUBnDiGY1T0QQsjqe5W
RFuuOFkJKRomxHjcePDr99UiiUnIURt7Xkzq4yGWiVIk/OQSBCAOqAt87JhTW4USEPdQzUwgMxC6
vqG7FFzG6GkdmkkgUOrLb0ScpnVZXK8LNUXsR/cX5EkdHgEWNWy3MZ4jpigkXdY4jlnhIdQYsP2E
3/9f9pQSAe+o1HOzqvwmRFdcTg2RjACHoVFo8kPcvQknnOT2FUtgWKP2lLk2dipClHzYFYtHV9BZ
IULcGpGQmYAJPubbr8Nrgl/SQpE4ZlV4Hsvw4KcXLgU4yUD28WMXajTENZ3ABmrrre/svYNz24kr
2sy9Rc2tTWwDJl4+NR/FgOsPj7UozOR52fKOO7akGnzDHvAF/R5rVaSoxhZJvuW4gSlpxjuLoEDD
hzlOF3Nd3HTUhdvpJyfN7MAnQR1kI3yu7eNSZZWvvS4PPbHMZOfgjZqz/J5SdHd4t51dvEhvy6hX
FuFV1Qjd4+MQAGgO7hQsOAygjC8/B1f3056ut/TKVPQ+4wI62MbF2sZwVJTNkDGr86Jn9HsfLGFg
WhRHr/TIP6BPe66ineiU1++Zrbp3GlEFdlVGhHha6h3ISQXX6q02X9vABAP4PhxjJDVN9D1qgpeu
JNyykfMaBqC6bZlOAgrJN936pQKMhKkTgkzAthoL6e68JIZo85qcPKfhEza4PHO+j7BaEloUKI10
eq40K6FFHK1UzNxejkuI7RkI+clcpaiElfG0v7UP7Ef+D+Dw4cIs+Rcu7NxGLuFtLuXudns4Rw5L
Ql9Zfw57ld34r7n5dwXJl7ek9glokRJ12cuyr9e+cO5P/ulP3V476ruS3R4eqgIfAn9B3zHg5EKJ
7RAIl0yHAzaCnr3rQULDeG/buPQrClbVEPLIyBRRg/Jpp1AGuWAyClkJ2IaMUi9tY4BjqQOSKGaE
9XfrwtgEvOOkKTdPxZxvUFzkJAPVsmi4v5DP73+OLk1mEatCSJVG4LRAMa7K5kVXn5umAT9Khs1a
IGsc4wedNgv+5zOS8VjYNDyEHOKEByTWL4NQZ7bOaPQXajpOyKmOL7raFYjvtb3jiCfLfOzCvAhl
yI9wumAii2804HATXhnsDjuCH9NzIruyBzX7c+8bgYFjMPr1TvuyvhehCg6ChhHNzCGSasMmVeX2
xzsICqKPj+86Dnsl7xxWdaklj+c/g8mlZMDutLFUMeTR3Y8d8fKJvPTI3QHTWEVXdRPAGVPYUZuK
bEVaSUZHKWEJGMwzvsn/kH/RtBCmczmdOHSLCiYkKaWzGXH8c59wvdmbjXUmwJ5DWVcE8oo8lv+s
agis8OY2cCs6UbYvFpFh6WGhUAKNY1cdey7wdKTiK8rlGiv04N+xhTk4VKCp2bfeyxtnruVbxH9Q
VTW/kCNa7frtakpAG5KhZ+EKfvmL0fkM0qizetUFvXqkjzIRrGwdStB1+AhDCdlEuV9Jxkfxnr8k
CzqfXN0T9FftsEjBLzbLFPYJSH49aK4dqGvpnsKK4fjQ6nM11sFMkgkyTAxKCw/v1cE5/VU+zK4c
fjgsMjxr6XSS5Mbkrz7i7SxrXUaRD1ohKaiWIiNdqx2jCZJP2w8+/T7UviZB5O/RXjTOnCV6gq7V
cl5kxN0hNxp+y1FMx0OxqLMZRlqQk61wPSlLtl/pHPI6MNeDx8SjVDGADjxompHXTFMxjfuAfOlx
I/usHg3S+ClJEH8/Dj+I/W+hI4ShwaYWAPXLRei45vUiS5aYPpDVpG6Uu/By31djb8OkdomqzVay
rRUY2mB7WhW1doDcUhUlOTZ8N7KwAS4Y2jMYICAcBRg+KKz5vfzqheu7QDORnsblIgzXo8H+5EGI
2IBOF9TmrO1EwLwY8D05igguMuRN8bRuKsbgSd8QTDaC+7Q8yTMgEMk9DtpHulnfjRBFhZ53qCmi
rYjABxZbfKP+BqDsw+L32zWQ6pJ74KZsAp+nMf2uDvDHna4efv9PLOkfoymwI+SRUeuAiaGAwZQa
5d5p4ZrE4DQSIDOTdN2KyDrJO/Cc7l2unl2DtqYsuJfOz3KnkZJnKdeCLN0YUJeO+aCcqjYnwlv2
TesdFlMCOIpEkR7vXyQ8ycgtbU05t2ajcNtnLIxDhIQR5IP07T5Ik0XsBjYd/ZEwHpNBHXBAlaOy
oIrA+aCdXi7QiLwf7dlyoYklLLCOGSqKMSJaQopvX1o5DaO+AMDqDTGbqOBua4YDB6nwDtrENHS5
A6G006jvCZN0w7CJ3ABfkK/oiwGwALIDRapMNYwQSzLStFbEte6rMW4t/QDxtHwGILRTG6D7aux1
voc6bOIh+WBofzQeoVoV7y9006wDmJ/D7B+iKf2PUquFHPRH41jbUYlU4ywXHEF9gQOxUbkvl1h5
EECV+w/4ViFqL1xr7Sedlguz7vIBqVihMrJoPW/ZFbWxA2M2wVzNCWbzk9gRyMdmPeLOiJmFDBJw
TDayePmKF2dfzG5Fyx6U2ixHLKzbqAOtiJ2IPddoiTyQlpMo/7uhhVg3IdsKq6jsJPBT043EhkMJ
WaWlepNyENWPxJot84lo50jJFdh3Bcqady2c40GqvbbOBzmCixOgC9hGKmer2hjb+I7NBnptzrMr
jzL4woZRBazYEQg2hh8y5CalDlbVFV7bGFYRpZNi/9lxe3yH9TyrEXy174YFhJaOcUfPGKfdmX8i
q7V3ovGSP6L1hKpuz2/4SSomlxTO2vme+Psh6/V3UCYoX/H/7JsFM3XCrytbJqZpCWRfr5GY+BdR
q1UUT6q62GJGQRErHebrJwM11/naQjzFMYzEzF9PwbvJTl9doLcxyjADzViWE76cKW2ZvkLlLywP
JFvNVUoh2L+5Y26DZ2ScZJP6Z9X+uEmSiriS3hX8k/DkUBwtf5d5fdS7pP7XD5kP6xZ15IIfWIH3
vWrmGHoVAsiKA70HCB7jl7hNhzt3CWP0lxco2Z/eMmQ4/3GxrrVbsF7zWhvrqaatUiIbgfBbNQyL
LtjFsHCoeu7VEoMvRLz+sZAQ70zH4lmcX4SkBnZHgOe1iJSHrU3OrZXXXa2QdbFKxfbEAr1b+QNj
UKd11NHbCYIzThYXq9ZYhHw5lkaP4Jp766zBxCBGOA94kD4HRLxs0KYqibAbXZF9yN9IbLMeYG39
LoNhYcSXERaZz4CUmg+bDC7+QTj66qCAzRuc9eBVR+1ElTF9DeQ0Cp9+Z6Xt5ni58bWKUrWRaWKm
fGIHmOnn7IRyvkhgSYZc7is+ce39pyJTdx4w2gYvYhYZXKwNMnob0A9lqZPhbgvFO7T6JeIf26I1
6/6z5501wh1y7NiNjH+lFUkk/T14raIuV0ZVs34MCqc0tnjw4F3Z6WjBvmaU8OMH7B2cmSmdLjab
gC0crEZ87ZUDmPElwb1Av8wFZ/BT1nHERtux1ktEDpDGtsTbDp8Womita6x5jCFJspkO2YNIisno
rdbKbc4kAf66coekCUml3/DfVBwZbZYdloDysj4CMKJjUISH4n7nFrSVWOSGr9mgDvn4eYFOZjYr
dLDtMCu2bnpaCKIvLYNMRlMXTseD/a08ZEQm26X1uZ218NFTBcfA5RkMKXXCYlrONLgD+s2n6f01
xVRBTDM8wJvUTcI4gTcCzdEc1f11oEk3c6fYpXxORKbz0gLVbUsa8gTgx8gBGccC12Z+a1aW6j1I
IwjwBSGcvA5V1jZAcfL2pAbn6nXuAyL0DCFZ2ssgA4+bLALsEoeLyY/9x+/+Q6GpAio3Vt4ThLF1
GdpCh8nLcCrLYPcmUzGdlMj04/Loi5SVfMPpvTmGItLt1k/Ynv18YKEMoaAf9ozRN+NJeS3v3Fnf
Hj9W6SojFmRJh3FzN/fpfyis6apsyTnRRWJ0eR2COXIanpkyIgpmyI3SeFVmmZpsFKbwLHIDTeoc
jzTyVJvu/FB9GYCt93MUNW3O31iGa9qUkg5diRGUx5U6Fgxo+4x0AplDyKMDtkbpnDATShYadOOt
psgeNS+LKZCEGUhtSJsAoVl0M28Ubue8koTb99h6r3tI+1Mj8pJTzyN8LzthG0NWobKIUZ+bpecP
fIUi/pKgmnEdtZvy7BpZ0+pKP90JXxPxWmAqwuqo9vZn3vMTMznVqbHVmfIJln916L9FIinKeG8h
MMO0IDL8udFdfFm/cksQYKR+1CZyzQGiKmuqQKobU3YCXKTyoxz4WQpyGaX5xbEpHdV/hEcCIwVf
AGxorBj6JR2gUjQJwT0uqcj7tCZIDQEjXfVs+03TjAdSklDwyo1QtMBJkyC9ZdSYyRzGR646Q2JX
r5LwCvAZg6UPWS4uNJ6G12qDWZ4jp/lR3xZZl3ZpahIV/oc9v/rt5CdgqP42IPiVTVAoMQGsJHCg
wKqdjvIuj6W1F3A6Ecx6jvRLduQjaDW47lbjRVAjChkkfxa6IDcXyFS+rHww5KF1klWf2DwycQGp
cvnTUTUnvXh6RNuW4u+UyFYNGKYxkWYZrektF1dTNrbhzpzJaMMbr+Efa+2GmtaUIPi+Z6cPo2gV
oGo18uKiHjMhSYQT1TrfxL8QzUqLjZ8iO9bhZ0eyyuYJtqN+eFvu/QE8m/8FrsmmIVE6j/rvD6/3
ksH/OymhuX6ZDgnKyHVXSPH8nAMFiT0n3kP62ikc/qmEEOPQXv8b31FRjUGAIfzXw/QGSWjK/CXD
6LbnIM+Ow14V0eJVWKnNnJw0w9EH+Cxp5YJt+7Hxg32txcEdLmdpXY17B63yLnFgdNRy2QaFzmIc
PLLul2YGrsPAkOW4uvopMGl/XTJAwcbfZlJSIJ+3MejjMYC3g2/irD/ry/VVSuiOX7S+vvc4w523
V13zurKn7g49lgg9FF36N9Jzw6Fa2k/yfQRSnGEq1Nj9mebLztRx0hvw6uG6DIXOM4FsdxRQEzYt
ifmusHmbWXjsfEhVM4QWN73cCTdKcYFkkBaO2uNpZfzIre7mN0sBQYNKqYThNYTmddAMZYwDoq3b
iJ0PfPTkrUmSvw0GBGLIBZ4xFkGJmXhobMQz9YiITXE0NooGAb6A2FWbsuASHpUtSukIruVzwRB0
KBA9owScKEn2x+WRqezRkXPGmscxhpZ1zQXkWGAHDOzVaSnXDU8np3NtS+nyYQM5ErJ2DG7tt+ID
KNShkUf20b+NPUgndXR0eNJTM5YrrpItAzcKCt01hQUEmVetsei2oQkfvnFzKBwi1k7X/k0unVqf
G5xyf3gp0W1q1yyyx9WXaOFw4cNqZRZQQozCiSLiJ6B133FSIt7BMHyvd1xlm3rkBaepxYfckfY9
Cl9td5J81xX1CXpERlblanu6wyUKA0jWY9Vv1aOm4n8h8cSNzn3SEN0EcNzknTm48+2K1Qg1drsS
jwS6/ezNsl0fRwNvhhHnr8wxj3jB3lhBIhuN7rIT8US5586ihbjeLvb7utpULeRmcMN/CThwCg2G
fJ+Zv6dTCgj1HuQDYbVB03yFrzluqZDDN8/PvPOl2cUYEeRrGtmnf7QmXvZsd34656CwopUfuLnn
QGnK+oge0hZZA9hUsDTiToK28um1kD/UJCeTwd01yUpQY6AzD7XRfmhMsVpO1jr5r/9OASfLWvoU
wMqCTaudBGvBvAHmA3770cZtEnZVmXNH5JzSCgCAgc3y1YPYnu+5FhQb7ynobDwO7z04KLUMmCG8
DvSnVmRWynlJSnnbK3i0htoqEEohCVtPQr+FmDxqqXvM6nAFiyqCGhxdgcStbS1WASSfnmbRf/lZ
gulY5qq1Urd/gTnsdPFir7uo2nROZ8b70OTim4WxFWxrE8jCnA5C3tXrPKgXJpFmzzV4vjKGYUKc
/7wm3yYXvUWijYo9o0kfMOk+4KCK63iGs71MKXZUjSc+2DRAqMgH+bfbSGap7LfolHmBi3t1NLzn
j7T6QRrmaXqM68fibmUVpmAywlQLnDCeWtwBcuCR3ucxTYuxG1tN5sLuCGDpfqgIhbVSh/t6lKoz
drXGATBej+/PauMJPxats0hYwoE4tdvMtJHru6ZW7JbbgFP3gP7TPPHLljB1MkpnnYFs7b+tF7z3
0PY2gak7vacx+zeTKQ+2Vr2QDTT5DYOsDzXbOYk1+4qpqZZEgKFBcMU1732+hdx71g5Hp3sL0RA0
70bP8SeiatYGlsDUJ5L7X8IddPIcWGi5hDvjyZT38JQKkD/OOo7Lg3ac9tRjmDQY2Vl+QS7514KN
ExK94ljxqdLx+1uxpDFzfKyov4G77SiRc+XKIfn+GMR55mSMV0A9C8ilif/YDs8bYh+EiLDEWjJW
rWA27cqrq9TPHnoITnK8eFvuNQfrkivuV1lAyjWpmRMA/8MrbTbZAr8oCKlIRXTcbzs3rfabsBCt
fmMjL8DdWQY0zp8rm6weYRyGPB4H4axPP1MAK/8w+QL0CFBDQnRNZp4pjDhcx6RqWNMIiMP2MgT9
iV5eJIkpvj63+rI9DsAvm2S2apEp4LvGJCOPgUExicKPmzJp8n5j0tQgM/ePzQxIgsXR/2ws5PmZ
y0o+8L/gqF9ItKSSJVKHGtMo1NIrKDCSXYPKQz2i33IpfSTynPcpgVIS0+S941zP7yj5wIiBZQGW
vjfeLPNrTDpYpaZmfpMiX/qvr54g9IYrYl9Y8U3TM3TLmQCjM3998JhUmU7Iiqq0+A9e6Ur+XgQU
uG/sXxCftf6BH3WZ0bMR6BBFxGj0RvLOOOxF+FP39BoQJ2EpICmdh6/qbwiYRkwBb+/rhI6JYBT+
UeAAzpKLGIJur2fmN3qtXryGKUyVcasm6zfmGAyIPH/p453Rk5VdUTREUpnR4eALfsRk6tFWNMVa
iz6SzxxgsUPaZAFL4q/8NfjjW+JYUwpzDDhYV1Q3CLcZUj+rxuMozXnXPyfhXre14ZRz/9U7BEFJ
NmP595ZEXB7tiNrPtm2a3XqTnNS3NEhaDWtLrQKjBcMgFkWP/TwF3VqW/7TGGXSSe/vU+2+mg6WQ
e+DM5qwhm2eIuVmH1xDJ6cDYXQl8zXPjqycwI0t25ctoI0DYMC6XAYELDD7tlC/illuo1CM8sHl9
EoMtMmKClONKh7hq+Q6HK8DiXwN9+PozukN1ybtVlulPsKdqDs9AYiK4oWLzOsCILExEw7wlnXhi
nDr/cR+b9osomPm05gkFikWW+iXfp8KS5ONMYBk6aUMFlipJA6lnp0VlOo/7hBX1OT/s8HeVvwFH
Ug/I5eW0b/odubH+F8gQUGlUVMev6RrQCpwff1TjSRLD/yrRaPBSQkT3wwkj8xUMjdDf+8OaN5b4
n8St+LfyyslJtSBIliZCRUUF+TL9zhOKZNsoP7OOK/ZabHQEMVFlKUHJo5g4gfgTTRDYmZztTQf1
spR5SPErdhb+BSK9q67wP75r2VrRSQVRSuf7K3p/up9aZEil2pgiqqOUSZGBII3YDOy1pFevAO6K
vduTmeZPrFi+wX29nYi/sUtz2NaOEgGJUa861BUOttW6FSecmpm0gGZCws+6dIazIQiOLICdVfn+
KRu8U28bCqu1BJxDTsCzJ7TAz9I+cOG6/VcKjiR92Iqe6KTcCA+02q1jjx8Ou3oWIAX1RXpV9cOO
iv5zx2EGlf55SqIAizosudoJV7DnmGvSbpg8OJk4uLAS93t9mg3ExtmzBkBO87CQNS+HRCY0ziyQ
MNRR5AFyRGu+fBcB1qFyn5DC4iyWpzwPngjJ/hkTocmoorP7DhiJB2ktJ/Gww+RSSCXHOAQ6ULXk
On3AUZfeEIvrx5Wgnp90FSFOezaEqQs6Gpt9LPfiyS+3wCuadLIOvtNpad5HWUmX84t/xByuOs48
AuXcCUylz8s1XJRqGXHoM48IoiG7CJYhblDw/rhM8FVlslx9rEeCVYK05ahdKdhx3q1jrN6PWaW4
JjpGSRvbN+YQc5qiupQZYlsIcTycj5HMlF9e1gkJsB29gFJ9PkiOBe0Vsd6zUsY3RSRmNsnLLQvX
f4qXY7ymHdf2w1f2pyY8y7/Q5UhK3E1RBccIrSqeOFFGcouU38g82oYN/eN+v34CbUFLXt+iJDaj
TVqq3yj3a+abU60MpuWafnrtesN+CIo6yDuAU+nw2WTkSgGZUaVkqGusnBkMwaw6koRJWKfGAfJC
LQwWD7sJs4ookVCkW+ojEGs480lcolyEYhNLMoOy7GUICJQVyrqDiTR0x+yaS5HiImrLoYwuBDXc
SJj2hWrY0X+L/zPxrqFR37s4a2urxiWWpFj9e4vlO9DEy0Fw4cSsfo345DCVuqEm2ewOwZIglfIh
EvDXJuZet69N2Y7YOc0ueCaeGrHQXxky+SwofOXBYkRGqKYbqNBocGK6rM/FpKQxxzhhJnIURlRO
YlaCm2O9ypITH8L+94A+8MJ+MrHVscLU6zDU0UDIjX9wIaEWcrzrk6IMQpinzOyvUnH0uG8Mh/FP
mKT8UH11U4RjXm7UtHS6iaOmHGXYicFL7K2k5C85Ak3haJp7nGoBaK/RgrjMMPZQDRUdJTtVCl1t
8JDW0zKc6SI1Nvyjv1R22H2mr7PM+uJHbtz5eUAWL8kFi+jF6Tm+ptfOnyZXrM5op0HFNzYTPozo
Vz7Q2txatseYtxIkWcu9ZdXSjbx/u5UlcJE6SBLq8/ZZUvBvPQiRmzNKqSSkVVD1laCB9M16Uj+W
onvOwQvq8g6lksQ7q9abvps6FO0e9skWGYmWA/ObtB4LK4I2ooU4FIa/9UYqA1RfNTg3M2E6CZ4s
X4l1NbhWL80cwRWvCgtxzE+LDRpVs+J1/zsMjZGK0RFdaif5vgA/aHsk1Zic6fQf5JvxslwGgS4l
gtiiYw/F0ddBOXxZI7oPhS9XaBdeRTCVC4PAxdkjKpSvRpcF6ntCQpiWkJkvu+cs4mP9K0jP7vwr
x4ZiIrppNdbVhT8E3xH6m3K2I/2FHvbucmbqIehcUs92xG0kYogWHYXRMxKCdqo2dmLdKWimkx5D
7FOVXkTn75kDOw7QCC/epwQliT/Nb3X+1hXJXRROqEs6CvU4mgGxyBAOWOusqMvrt1EZFdXXJssH
Z7c0ULTT3uE9oS+jDIcHON3lfDTB/IXeJCSI9AZcxKj95tjwTi/TRnLyVMTH81PPS8TE0ewUio6P
i/IgNEpH7dRcMipxPIXp9VIlFNq5u36Vl1aRql2O8xJKAm+nEEMP1M0aT71aST+fzRBPpClROeT6
sabKXyI3v2dME7kmHSpmE/b8iXhPsV7V13jJukulnkXEWAslPhNn6QHsSCk3oGmSyMHaA1kfDDjD
qiMtUsdu0g6UqTPmb0ellPEsEYkG66g1D+EkTHGNiySwrI1bBiHSbSP1g+7nJsL1d1iv9VNonNr1
9oQlVYok24ZWfJ1n1WeRlK8R/IeBShsfJhr5ie/ek0VGBpYBJ8QoI7R7NI2fMlvsukud+MJ0VZfy
vflLCQv25VXZBetbp8nwDHkPBuXUGKubHWbyEXFXbWNRXgS7pkzPgw9zqMqD5dVKhja+Njwx+mHK
DcF9LDw3YkEYoC6C8Cvjg14PoIT1OwRTi4K9HWVe+pajwkLjy+SS9YXabK/UlIVemVCTmQMPKEZm
9guckoXOiydpotNMThtnfGauO9MIoRJixdgAMzw9Xah6UfS6W3dvjcxgRu2xN08WyerSzSQOMXOp
T5MzQcf3oR7HLNUNgagsU45Vg6qQg+6sWLkOtmE+eRa39owTUn/lLZIyTamXhtC8uC618lioTIKM
sIojYoTD9ZpeOp1uW04b3V97DLYIcVQ16jY2ABGSctP2iW0Vyn00zB0ZzbkapIuY5eutBOLx8rCV
okHsD9+Fj0XdpJKJ/W9cl5tFk97phDjzl/o78ebB9/UaKuZCSDzMdg1rJSDH6JdNrbBTHGs5X2nT
mLmGtetPAdR9z7xsArcS0cDur1SN5IsWjRzoE8B1dh3qQMHSgX/g4C9BWmSFZcSzYu2ByF9H7RDM
OVxG8ZL0rLnq0vzIRO1tu2uOiU3jggSonHLJDLyJZXsN5MLFnamFTXJHHk+qdPluFeF9FTSUBFUr
hXugStzaTuN4Br58J4Xxmx/PUAL5qUsgCtaTb8mwhst80khb5RBB6AnzowyN5zr5elu++4f6rbrk
0K0e36sifoEhcPCpAlo8N7KyHtjdwSVy0lxzOpfAk+Z8+sY6yNFbi02e+4tFNo7Gm81Vn/v/DCdU
wlJYibPJ6Axpt22zfv6w9AQW18+RMhBRsZei6yHutI5pRLzSsmyv4rlj//oeNgppu9Dhr+mEPb9n
lurgu8KwEHpEacn0zBoQWB97gZCjyt+sGcUmMLNYzlvrOF0xHLbWDpFNhfLGyAr9o8rA20WCnFIO
3anQ1pgNVC9afZLypR1m+tsgxmIXeuiJHGt8N2sC9sMKosNu0Voq9w1o/2nznUynaFZe87GH3+zc
u39ywWPZI6cG7cVAYq4tIdj6oyiaAddgwyZMjCll+/n9SKh3emHt028EjLmNzzemyR4xkGXWa1Nu
3Ud9gA4B1oanAkV9NAKis8jbnoHoVKL07uyoEfmBI+ZrDqwN1s2KtxATj1AFmgcoovNUKtQyB06J
gd1Kblx8Hlb2lCziWLYRGcGo1WjHxsMdiNvAXTSXs2Wdeww89rrx5dw8WhbNPlMRLmADBau4gWOn
Uwdj9ksgA+l4zeRCkyJjrA9lsIXQrfoBWdjiANi45MhC6mMQjcGkiDAUzm5Rb2L7zWpXm6EvtXD6
dyhpIA9tty6Z+VfxvrRcP1x424bmHjdHovHH2CFbhMg9yZhvFcQq0q/xGywiSB3y6mYZWp5DqLZr
qSFJTxAOfdS31xZGHjm3YKKaYx23n+HSF+kn//1u8t+OxZhMcCiSJ2K1bq4XPMosYk3saRUO4V7e
WL6072rS7uH1ot5bD3KC+unAhnKvuSU1WM4zu/eIvtrRRHH4PGqFdwiEyRyCLj3jOefZoeRcFopF
lpIWIQp9OacFXTOuoGNEVbtAxI+oK5lgtm7tU6g9I/tLe8iegaoWnywL2YcCL7TkUd0tzM8NXHLn
6BBSAk83F0B4Dl2U6r3zE/PhROjZEMyrueAUtzF7RNh9/TRGTc5lIcmbbZmFuTYw1Ph9s3Cz2QCf
yZJ2kQziW/GtkQ8p5nYprxL+i0C8I6lYY26CLEHXKn6LHHJ5w5NSLf5cnJBkcq2rmHjGJGH+A5zU
gGWxDEfg7kQRVQaYtK+22/2qgI5KOGKp91QjQBL4mdg6ogr+5UCv9od+yCjTwfYo1FCk1WnqYI7R
8YZ9hMjf/GQQcotBw+etaVVUIsSJHArLbGRSnInyv75lelnue6sQTYAObHU1pUjo9h3kUS5xNHyL
Z275c9XjGwz1BVmvsA/8x/d5glAP6B8n4N+Lb8mMGWDJtgN0cYO0yxutWm2gtKrla3c859iZYrpp
BgEAP7lClY1d1P4D476Cf4wZCyQvvv/4WpxfTIVG9EBlGc4sN5cFE4v8O3OpDcquLI/ZIYbOK/Ec
FAiGjveDETnH0aKK8PT0/AuX8krb4uEByFCTu4cecxuHqGoHHXHBwWcYE1SxJD4Mhsvhny6Yta0w
QBREcZydkogBgpXsM7AUhJ7n39liVvWFfdbCsNzpF0oyCT569jsWYv+GCgp+aLuwOv7YBZ3vCCg5
ofodYY5e+YEHqwX4odRMAx+ZN0LBx76R/EIrACVD3+3D57kNUuyOjO0kG8beCz2qp46nVHjSe4pW
c53pV+pNnECnHu7NDT0qaG0zrpVirdP1SzXQQtrIXunDMX3BHvQQwIc3Vwr32G8odIffMHY0M3Ef
GRUTCzTyo1WYfepR7jiehjB9TlreLKbo6z4tGhn9L5yXB3t2bkuNq5srUE5+rOZQIdxEXC/P4Y+n
BwvqmVJaXYq9T2JLXF4ILS8dikecmmj6Z6wmwMriTi1aS7Z2HeMUWl/Op7fDf7R5nAI1a9QeD7YX
Lnb0SKunpZFYHx6Z+TxTCgxRRf2/KG6/yo/+F+ejx5CYaUY18vD7SaLHvXCYH68H1e6dxbM4T9is
jZtJufWXls115fdznAzxk9doFYpBb4nCrd/g8qD7rb2EV2MREHQSz7OKAN3/Bq8KvVq3mvE3PuS6
e3eb5udNMilhCthH8VmdLmbtPm1KXU8YBqcsayrYnCfBXIL0inB9s1gaF+7x57o2YcJL6VE8MCDr
DrkGlKlSIZfI9BoZgM/h79JttRz5R9sUvxCBK7m1bUj5rhgHfvvxcDcQ97waVDEw3ZiqvusM/jET
vti33ZYRumGadDnYX6D9lgUZvLM0BROc29RQqdD+tDZzvJipuIAK8p0CY3CQBRNrJavNWbOYSth+
eM4ea8OqAXm9FTaUUqzUhbdh4ghcqMqmV9FQ0UtCItJ+rWDJUsCvbNGgqYeCXiyUAD2pDfYu6HXw
carb9eHEUyXFGJ2xMDEHXWFsLp6IRZhKe2HVhugBXH75KGdCVWdHkX9CROxkisdVempVnjYGDS9Y
XBeinDBYf34uLh2wyO/VbVxRivq+1MACbfBt3j2ztSTM/XGcqfBtJn6us9b3r5yad+QTBjT8SOrB
aU3Wu2QB65OarMkM4PUAJvhrnuZQSV06FutipYlM6tYVxcMHw/Qp5xsxXIOw1h/7Xrp9mPeZW3nG
J4uu6d79eWe+FTdh7mycDJWaKqiS68QxNwWjD0MPjGHORgsfjDxNOEUXAM/a6BrehvUIYKJUYrWW
GY4q3VhzLEtnUBx64TDG/V69OCG3Tn4mdGyNoaxnUY/cQx7/7d4lYGMVV5Y/lgoUFMIhAK3p1R9D
wZyNHUru+nqGej12V/mNycGtWEzUllhspkVyCUlJDH77v0Dbb+WLzNB56EDrQkCJfUeBL0wdJl1e
htAO5FOtpObJO0ndgPifh+IUzAJr0O6S5wXk1i9aZ9fj4nUA+sxsQm8nj7SaT4Hc2vAM864v8U3+
/cQ5bKeSH1JAEjfiynDmbe3kQv1+GjDV5XN7Ta1Kl1JsxGgE0GvMRSC+IvFMvvp3uDdu2XpvGeo6
zLwPHzIhuxNjXeMfgMtFR0p3KQthDBR3+8jKez9ZURuOZWnOTzT9TPWyFHO2oPcRCBj0H5kuhHV2
n1v0N38eBpuHL/TMc+GNjRzIeh95IVb9Qo4OkyiTt6CZPSD19nas3egL3tq53fzZSt9D/uqfohxy
XHruc3gxq7T/n3hxbHhC+01s3C31G8X/bAuyrQqZzJVSSV0qNpPbZi6RjAgosz04w20MVnKCuryD
kFAAitnXuUdMznRvEyWGwN1xs9zZQpBG6wl4nFxXuckJtgrRipL1Zeh6LJ/N+ut3sN+xQlkMsjYY
5uRR5w0uYQm2wMpnTee5d91Dmm7QppPVMKarpjF/Ydo9svS3ae1NYvXs9cgKc2fYZeXqvJUc4DNn
+oYxLLA9vrOywSMYKNPqNTpijl8OzTJBfunWQ5u9z6bA1+d9gs5jCRaRlV9BnEKOJZH6N4cDlFd/
LkMdjVKprCADrei/eYQO5EhzxCfPmHkDX8muZlIUl2F/uIgSG5H5Hq7cCsYNV7lFqqd6kypomfp3
hsORpHNqcNjmbYEdhiddfVUeqOszFkQhWKO8MuMK+gn+v/1K73/rNmtD5MTvbepycIJWhU95EEbW
6D0ZwWQIuNs+rrFu1C8ch5qB1a/hzqtCABpKNR4ClXcFHUhZ5lWJTLWo10e9mkTCT+g7VDT8P222
xCdpowmCh+XwEkyi8fkzVKertb1RggKknpw4uRi4nka9Xr7mBuXZ/UETJUaILlYNn0GhTRiSVO+O
1XWmJx/iuCekJWEtREeLb9XSYEXSBZzw3Ojv+IJTT78OS/61qg2ur64Bl/REI949E/sW1qKy2+xV
zwhzw/ngdYbgKHLuW0oZXkpNdehnbiuMBosI+t6JnZBMfU4pc0u3twGW6MVzgkwacxlH56G0fOiI
cTUVOCgA9wARskRnBu8KI4xxjBjM7V7BPYW7Uqm3lFigXTmDs1Lvzzxpa8epraH5kEHm7x7vLP7b
r5ctt8y4A9zzrmY3+pwMuBweLFW2gIMjAvgtZp5qKCn0XXDn3nHzVUJPV1XhFFficNWlszHLin2h
ivW7RmIZspDJCwLwagjKoCnv9OABetUyNc++sAf9W+3FXUJfiWMyh3KdAFqTCsOqMrfQEwCbVIU+
CDirHxhSy2ngnxR6cuqAKBLL5gJiJN+WxbkxFAhj/uFibqBtljEmvnbivZL8YMLotOPFLTgrxsio
ItAn2D05ZM61hhaROhCWWqbVpDcNqjTjn36i/ZCTbz/8xbNpqHLhjrduP7nFt2fLpExmbvyRwLCL
dK3/t9eq7tD/ic0x2Qz+NEoXcVZP9++k7BLl1oEXrZh/VrZIN/I8GlDx2ZuunoUNE7irN99XR9sV
tSwxDH9MUINUcsAu/v2WUUQjC9tkl8KjllsLBR9+EWvN7Dp2FIXD0BwMN0KD5C4aL4U0pLKLOBvN
O7uXT8UTG4Sfg3n3WkBGCurqtH5fa79ORrDGmaYN6BgyQ9yf3lVaNrFnh1fEO8XrTWPzOx8jdZST
EWzGxENEl6/ZC/cMrNqz2kZLPzaH6KrRUqI9Xz546oVwY9VW7KsHoWZfKT+2eh4u8nQRyleF2KG2
dCC6rCrvBIMNX0W2gMEvIxTHXFPpZBifZyuiVP3uPDCXqdKPiN1v7kQ4N1wR0Csv5jYwOfzq5z2m
yfnFFFE7T/GweeOw0kCa6kzjnIEhfMM12WchBWegUFn61abIO0QfPHeHnCfgPoc2tRDArJGsNEc6
hDOVMxV0vCFElB53cxKZpDtj3xVPboDCaxwC3bilO4h0Y1W9GIy58u78Fh0uUWW70+n5l2EwdmTS
+gqjPxWfVsDH7v2B/5LnTc/cMh55D0qo//dphWeBYnszwQrtIQ4PJJHEFVn/Qq/pS7bwE40YeNHK
Ri0gEJSz1tyvKrpty7A4tntoIelWQABBlBWBb6oz2S08TbV+jrxTuUpYNfZal9jMXmjCZho1gra3
JMY1WS29k/0JFIIxAxJPw+zD541o63Uyu3VcAbxKcac5KbpH0ULKdbaZ1anA01SPpm4UNPI5qn1d
FlWrtr7jxAur/W6DxBFW8VsBr/FyznQGjaEb13dkKQVh7X53Gvv1e0D4ejQI+xya0Xx0jFPaFBGW
fdipohus/VeKYGHrM3MNNv+NubRCNLipw29PnF9h85A7Y3VDOulbNgHMqx9+SeRmbOCzaZDT7Ud+
pQej9JPYBsqOF+7w51zdgtjh5BmebWi1VpYSf61Osa4GxNi1yBP/XuEp1cSmF3EPSQc7aomEzsfM
w/fja0R9lTHZGTqH5QBeWCjFszi37bzbi09611mS6SAFrjJpcaf2GuBCnv47LRcndLET63c/TIil
NiOm8VQyhj73ozF8ltjPRfIeEPHr3EuitpoYn8pd0bLzqe9FssIQgebwQDDHxSiQo0KK7EqQgPY7
oaLVAiDpU/VVhCnQPd3xb45DJzgr+C3uuKHsOM9SonxTk37s/QtHqDCfzY4Ml8jwxblxu4VIqhMA
RTDiY1V7Ghx5ZOJlLIq0VHAPqmZvFYrrJNWowhcUyKK9w9we+PUFj8PZhz8fXqvU9NBJnd/UeCl7
qvsak5II7sWBAsTncCLWvU4BVA0SpNWcdfCjS5IzlnEv/eybOR/meixgiZQLJOmP6hQKe6ZbFWz7
jrek6z7n8pqSz+TB8MSUwOfds5VQQe9KrcHE5ribyRZpfgjcc4u66AtWv7VlvZj+o1EWoHyE2mTD
5BkeoZmulNVxZzUP5OkoJe76bXyJ3lYk9esZ4uli0zCUrnxc4ag19rS29GnJUv4sUzjE1pNzN/1x
QCbLwRZtFQ+HKqzZryk6u0x2lJyKyit57hlkn/s8Nc+UvgwOQe5ce2J3eIxpqm6dTBJYZVDdUzkL
8I+juXa5o78qe4MTckmRbRjeEfAQ/oilDdJKr23bbdVJdZkdS0OenLM0q/Hi1dXWXD4Y+4+RKH+n
MOGnzBEqBrKdiKkdob8AIbIqGkqIYUCBpUaiWBw/f4pErA0nSvbEgwz5ZWWVPi4QZYSY20LSUWty
qHPii3Mqwxb1cPu+cT/4xiqqwMoIg/Xg8sYb0Jj91hCvJJqvDxyrgvSSIjkkCDQcnE21/aVVZSxi
6Bita2OvGmnjfIlyiie5iOrDVshJ+PPmpUQvpexV2oVA2qZlVTqyDSj+E8qCyKcpoQed8wVNcWBM
68F0r9kVXP/oKVN28jA8zlmjAF/Pf9iPDTJM7QpMQ1yZWQ8V1jGWxk8zC0T1+BNalNml2Z6GSeL7
h4M5nC2Xmk7FZSol7vRNJazQ32DjERaYOxQWKlJNyriJ/U5XEG/yZsUUuQwAhSxDYazKlRM+vP/V
WFItMvh0qWha5IOWFbHWi6+IAUIBUsuY1puVDPz0H+umJbhPsotzhs9YurmQJN/rBHHoNv6TNMzP
IH/kHR7v81/0uPDPoSjcwnxXDlbD0GhEKn8+nUGrS+3Se57+cwyaMzUwI/HjX6V+VXiMg1m9k0Mi
sraJbzkSll2EfyKQIB19kK+oRiidHPfR1CYzxaNwEYaTX+qhU0pZml3UTtTYkLX70q4geaIDNrok
K1uRHd+VbDfpVxmbSjkPLwxC50GxdfaXCRhcS0iumBizU2izDslAKeaphrzCUcQI6s7BdKAKs2bx
EiVq8YqtMN/edT7H2XVEaWJwL7sBYfRHPXN4xL5Stfo8gKQMD1BZvPb/yIiJ1jwxMxwObGDBsLzE
uqhPmQ28T3/LJVdMWQu24ZZ97C/0EJaLQMaOdFjMPk5NUg8BQc3ed3Yxhg3nI+1bLKaRqDn1oVfs
JVAiqum7KusC165tcCD/eLVq23VXLdfpVkcIuCFNxAtlja7gxMXr+jmsw7ZHQnEP3P8BcBlm4pwK
litHdLWnmzd6HfUDsebkreu0FFzGbKxuSSVj7A163svKpRldBxnTWlLVGKMnIBbNKf7dFDi+hiyr
o3rx5jUFXvrPHOTS20qRfQxphRmOhcagDNRQ1qBcWtF51FnuP8GA3uETfChtUXbxKfJgnCiqAd1F
+QS3X+TK39mze5cWhx6aUVq1P7ppo829v3XkLB9o3yTFPDbFMJFSc3q/lnFqIJxG3T+wiXRnozri
AgqUPqHNOe97aIJFZFWxaYXIn/2AwIDjQrRrdFgeKSh85cWtLVKO1ty2N4eYe56KC71FUDK76hk+
3779yE8YYFIKBd0jBgH0YTgVXEQHVknOqqcF1VSb2e+AkxVE4z2+JS9MRl+r0O6P4ltDD5bUap19
4u1lmTFux3ThKz/rxJgIZzxXg6TwtNwF5en3lqosVMiVjWYBHzPExfWVAK7V6TqSjzqg8kbT6sqt
88EErflpaIzkDoeTtyRWtBV/CmoG5K+pTAzbAl8iDRBf8mAW38JfUIsuQUGj3Zog1+ifrK15s/5S
C/uuOxQigiNYeyw8YBS/3E7n4nilEMsUzZ8pL5BL/dYnzkQqs3WSn2rXBo2/eGKR+gK8lxA4j3cF
NjEUg0naP4UnfmKWSNEqqeChdaiIDkLe1Zwpyl8hMd4vtIQjnH15Kh+xJDaAFM1MkwzXfNb7vMIn
+/kmeUY/xmVtnd084Tgl6F91LQ8h1pxueyU+e62UpFihsWyKfczPqnXnew3iwxo8YshfYX33Tujw
2PBzGVqz5DfnUfY2Wf7D+Amfz+1KkA6NNzFJmzJSIsJMvx6pKCC0j3hUsMC2wFlGSdHNhiwtMVl9
8WQdrkLzOjJCYlWewaygqDh1V11u+xo7xDtvHv57HWFrcL9h3fMihwzz13kkH6NONWP0/T1pywm/
+UDl+rDuOX8P6bqeMIjfpTLv/6nEL8gbk3WLkSMEaFcFWtMXk3vwMWakFlfYTyu1qDqN0Oy35+Vo
vvHK9bCjaK6bLM9eIY/IJjZisBUbkJmmzpLct6vSmN7lun1CaCaWqk1c0i+jNTWsn8FOYRZ5Hact
ynLqK4J7/Cq97mFHLULkja2VyTmhTnIksDAYtcggb3GHf9Rouzv7LoGQi0dhZNsSS3FcgbW+tVj+
T1JS87WspuGmpo5ubttbHBtDjzmg/r6gRm3Lh5/sYwrNHByB0Yw5rbhP54XYpC14deY+CaZCqUln
gypICBUlbs4op0bHiPx6MpL0bRyT1GdTFPA8Nf+Lj5vqvyncc8OgyJr1Hnq9b73BgLYkf0bO7OX6
Z77+rz0CeH7RnmXJufNRYMewnGYiIE0SFSHqWYWUsV01RyLkf+eebNozuXZvfDXP1B58Y7ZlKrgF
nEn5LauwXDGPvXdgOPBo89sqZwIQyhK3nu/tClY6huKpZzYWUBQalnE9LsRUEEHNoUN3ds/F1SO8
FEctPovdvWWGWXloHFfngDgqS6DGKI1tN01dpVlR3wafjddAOIIBlav3PLtkRgqz8WFcClrUR9za
vdLGRuk0GvHI27d8ugTnSa2JjFBFNffHOFlTiHGnZ4IiReY/xdjdDKPI/l/9OQDadZXOdzer/9v8
JmizyX/Ru7udpDguTKCOdLq3UryOFNUKtsNJ1fBEg1DxW7N7WnXsXVli29pu6wjt1WSOwBjLarXD
JV9OIrWs5bz7gua0e0AVyH9oIlW4N+Ebu4AX5mHx2SJA6Wrg8ZeG5tjTvhiuUkBBm4djj90ZRmoH
D+cGTgS676nN0X/ds8trFWfv1MdOQIJ4T5EhUTpApl6LMyjoqWfWTVMsOc/3Jxfo7Nj4EL3dRIHV
ICPYkS1gsBOfnyRmZc01JgjcG88JI/pcNZK3WQr8XFQKFD6J6fQOHRwXvCeC6Zzdt09aKh4NEk5d
5WW6UrP8qv2Vh7hN5Q3SJFmr2E1MwDWru5wGmBucvDLqsLRDeaMMwJgxY6PMlN3wDJPbfwVdUeoT
Omij1tB8UeK6uSgvH+z7l+v5DwEpW1fjVPkKkTOVM4aYXNud0Nssg45PVfPuawcdLklUCWqPLIyS
Zs3+9JeMqy+kdEmqFjzYnarvVDCUv7dXzAm4oEuvJeRIX2yKMaAp7KU7UrRbBtPC/HFJuQVWWEIp
a9vLgTeiJI2kdNrgK60/+q3ErPs5qLPNHxcGdiTL474+zQZNWo4nxGW/zGXMBsKB1NU7yu/8IEzL
l8pHnrzzdZb5iPhkdSa7vTM6pylEgNunceMaEYt2BNuZoQ5alt3JPmb/RJ5GzCfKrwsqVZX8lNfU
vJ86Xio8+q8M+P85PTq47g35lz46q1oWjEdgYyrUFLyDaNfbGdORP0YshmChThwxR/w1YBRybwy1
v3KTUMLeXMro7r73jl4gg7QDlxJ0gXWmpRIeV0WdTW38TPxS7EZzTlOXKXRjHH6i6RLo+f6BXFn6
8fGfeJ2NUygB6NZrt4bzbU1T/YPvHuSOnh3VeDjlrT5Bmo+nmVx4Ty6T7lszNX4ibabVUf7LL8Z3
f0EyrseMnEIf/hieqMC9lrMcUHgbsjVah6sd4dZqePtctOvLqKkjO/7MF9ZxNJQlyYIzpg3l+I2c
LihI0WMGxrBOCw5EPxeqtVIxlyYReOHBiM8xnhEvr1fvFEvNM/CoWertbqkRC4L92GWZlU9m9LcA
EmJNsb4EOAd0UiKI3uFRhSb4Ep7y0RNSQ5+3Z8hVt8ILqejyMSjTaK5yQTC/3QnLTPCa3GpIGsnY
+nl2QwYqs9TnUEu4nZVr3Q12LUaM7xSFyeV+eW2tG8p0+52HAQtsVVg7f+J+tbUmprpLO4KxraQi
aes8fY+E7pvWaFK9VumTZwNqlRlQg1S545uhlNbwcCBlVsXXzjBQ+3Ndi32uU6rt8clpxvZnhclE
FWxbslfucC8M6h7hqnEn0kR7rNyUIVo/YHp1CN0swvV3J2AijnwPOxGKyzv6N4XU+otE5gIczw3O
cLEdcni21qNGmxS3Kg7PbWNJQ7kOlk0ftLZnrz07RpugO9l4gauxYHPU6cUje0QXLqFoaZwXo5pj
czKVHgOTZ6pWrLApdCgbHcOPWso3xaLWse8WhfhicUVKWN20eGJv96aPQKYcD36sEiXV1/dvQ4ca
zFb1sZQlOvfmtyR1Tz6eeJyVqf5ysDluFcG4agp1koK02gSHoWwLRxIGkt/TQz6gjboKSYVLFQbz
btdaQAJwVEw4PpNZQMmLNr1q7ba4ECcd0LhYjz/nLB2v3gJX1fxdch4h18xhxPjOAPUsGfM5h3W0
NHWf+EDHu03BNb7URakgLLciBelWgZ3PtpxgGRInR9tlzgspwAFuzN4SYIQAC9M3uEKiqdWMZT23
yLfQ8Vsfe1w8mBs8cdh1uiRPMkN6BRbB64XXw8u9aztgDzLt5EQZgUCBAMuIDXgtDlGVsRAg2Nsd
7BPSP8XjS6rQtDUO0eLMQwpSFMFejHdbIpJFEX/c5MW4gQZ+eFxN/P55MOlzJAM3qtZgoYcW1+6C
vAg9mQYiGkQ1jby66gN2Xzrys+u/iTjWTFVNnjJuI7DZMWExNOpZLRtxeLXi5WLdie7FAbriMu0M
zH0+8g7F17SElV5BzDnhk8ozfUkS7x3TY6CrdKXcD0PyceQCXD9mBubZRhC01KhxS7uxVhEn9mUF
kYGPId+J5MiuU6areBzHxlcfi8ouRZjou1okywrnw7V5aCwISqKrrM/I4pX+JqfyjPLq5chYOAMN
UKmGbeJv0yxqqBK99qEHa2vN5xSBOfGml81uH5a6vc3mgDrDxxMDZyW1rcI9ie9vuieHbgXKXa7d
uXYxdaaAH9CSYxhqBf4uA+OPP9+mxjnnliYvaVERxSnOCZaRO5zdQ6hL6HlgB1iP5e+Z6Y/ScuIR
Nxmxfztwgm/ZMj8pFTJewCFch8p0+tYRqDTxWNam90keQ138UF6uxxX7S2yAYvXRp5H1lYYjR2DY
+uors+wuOHHssVSQEIf5c5VOKrszMSraqKqZN08njfl0AMq9fYubBgMuhrtq5RSLbh8M/EDEjvAW
pEO6PU/fnirIZPEHKdwDnJvLng5LXJhXC/5u0P0fOK/CMFAuDmk1mapmGCYcRdHSlhy73eWroRgN
Ds8HMcTkg0uYoDjurjlCOEShNSe1/FfmW75WVe2VnBWxj7TOhEYSeg47bhBrRWOq+pRyqeckxYEh
8t9syNRHedndr8S/foNNWtH4/kKTVqWzv5glKtQ8ER7g3HfihKhHIIDxuEnLDdPtwpL8Pi+pL57p
0A1OMwbwTCOhiziz05wIvYD1OMqpUD0yP1IO1U+loy0KcxISQKRRnu3+chCxXzIo3DBB8a+550h3
4AMSfnGyl//eGr8bIS+4ZEETzgxderNxoKAx/GXb9CLNplXsoDTGESU35tOPr6882kadEsBjszkb
iiU0c45wnC+Adi/HzaataoHsumJbhmIPMLJ4qH7TJX7AcqRp3VRDaUQUp+e4ckQBzbI7TuWFJNjv
dQShSO2BH6pMWri8NFoWkUgId4adj6By9wvmrOpyUYwS2xWRCPOW7127FjiU1ojHA3HGTsXq06aJ
GtxkUt9qdHjOWuWqn3FdEDgH4tfFlHf9BrBqMPraTGWvFL2t3OMxWGIWnUGvM/LteD3eF/rONiSW
zAzhUHyISCLCil5rZHf9HMAkUBLTa/A4a1lbUrJ+zrLcKgMPlTkuVDEGf8vysgK3nw1rzOsq2T3h
5iFtFR4QCi6Pfuo+2RQTWOWHFI05kfRFWw/o3tQDaku5xtryYSicPRhMi/onP7oSQygJArs4dY3O
zDPK08AM7EeRJA1cfCYyB0qZi94wfdaNTjNizOlnkJ9HrORTVzQ+11wgnfZNsjRUhFKDSeDXmFHB
+Ma7CHJt8PWGAxModxEiRByu6KzhPMX9AUoJavhQtYY1nuiSAUxGNtcKAcG36w3wtd8Kb0mqkPJE
U0LvYPn18Kl6jPCYIeszNZB1hsMdFy8YeHlwrPgERewSOXRP0xzy5SHcqFbD4+ZhhuB3mY3hHq+f
Ua5o3XZbYToaq7LndXUR1vl+VONQZP7KSIq+WcFtVDHL0JZFFvCiwZg7Hq7fBFDT/Nye7v80M/qq
6e1OIEPpcvxTWYcmSuEtmG3g3CzkR/Bht97oeTvzl4PmauaDFAwULkFgIXYWh4yFWiLBZyjLKwAF
S9T5X/My6DfdJiZAg1Q4HyifMdR33FnuaYsLPtKYUwrCDUUWmClm/cP9wxZVDBhIcQqcmUDoZs4l
lfncTKVbhJJXa3OE0hKQ+Sn5Lti9z7yvfZACmAFjYM7XcZ5IGPpWbpKNxpMWeR5oEjeH+FdskTI1
WGQ2cdYb4BXOrLoj5xleyKeUpJetbvIwimNfmD0PhxZmq8GXdzTGGsZvADN+zHjhVVYqV1kokZSP
wL9UJ145iV3+46yEZcN+V5HVZ/SzQO1sdskWz2kliquH3onGWuVd+x2vI4fyTPIsacUP04RsaoMV
baXzYF0K9kvK2vDtbIB1Fdns4o9VGkhzHJ5kXKPxW+EwRbDSuH2F37OctLCLaANHxvpkHfQ9MtG8
ONrVkpHFZwNUroTL/OUdke+2DTDwgtmfNNipOlVoZAaRh+aiD603XifgO/cmZYDZ3K482PbamVty
LssIXbtZirj8iJP53UIagQ7TZIrQSdpDCnTO6yhaH72r5qUT7VHxQJAquqoOnKmriZ+Wof9bHdkO
JrALwHAuxFMBYlZTuSeBjDVc8D4rJYVVUT/d6Ed3dfQc4pZGNL87k+2DelU0+pzrAVElOKGzeeie
4NxbfylzPV34CKVivZBeVndEe+05xXf8auFDn2DUMUm5YgahWHPn4ggYWs/+CPv8Zw96UnSbrtWY
4L7JJ6E3PaLFNb1Ut8qUvA0zeB/O4QZbYju3fZTqlgPPn0MKX8v7oBB+EgpQbQukBtj0EeIgolNE
XZX3mQVKqM40xiu/uZophloYPursViakxGdctWK9qu0L1hpRLy33fB6oKWhO0PzUM0/63vO20SkD
+jqvSUnV5nqYRXfAo1JBivoEDzcU6KiHvbQCs6KtI+vhVQGGe9BliAp8Y3V58qvLMGmiM4hJMEl9
TYxZqqW6Vz2fcXoBPha3prMHSnQoHLby1ViwDIC5D5v+QnO8YeNKHxU+eXE3pHtgX1vwSrvjGinZ
5F8r+EosOcI9aCC8sdHqk2lZti6vXpPdH91tLKXpokZFSGGUtMSvPuY8Z6SELLS9WjTDnbfEzSCH
CCywdT+jYuKJ37e1y8a0yg2yLHkihwc9psINNFLm54bhGym5XaRhqH6DlCiqXaLgjrkoq8lpFB3C
xq6/wNCKDIZ9fnjAK9wc+v9VQx2UbTSS2wcg0OanRUJWizpKQJQPywxMg36pkdRKOy0DqSLaXhGv
KupqaNB9M2tyjyZEau9OJBbDlasf5IQ9QgnZt/erojPGXEj0RO/UFZQSTk7Sc+8pCk97veq1S04N
Dl9KBoCaJcZ9+AOqnWk9RQ2W+Mz7/l1hnk0zIluhLB0JCT4AtsjjJSAa92GiVtutlYKgNv+yJTR8
XrUlj4KH6UrsMg3sy6Ss13/pewSgtIvqi6vH8O6tfnB7/g8ZusAJzOQNPvHAy2e2tVawAMK21r1s
Y2b4tS6TJGCEV34ZiQtISrVOjSkEon/LCiH9PpEtmJ+ECyDMRstIPgbyHcKEtSrfp+P3sCd8lbDP
OiQpXXcpeDYWZWhsBQOVtW4116fDxMjU0+NPnmXkUpW89nORRMvMjopEoH8+3vwSCNTBvsYYW0fA
8kNaS+4+mDUwyET/Z2T1Nrk51eC+N7tDstc2yocNYavtOpxF6NCvRvv34/dsuRJd3gnu3FvgCReC
BiwQtX0zj7NWJFWA+d2xdlQrgfKf4//hapEnl8fk4hHha0QZ89/JdgRngES4JTbOwxj4Dnta4VJ+
BJIW5vplH9aJdx0GH8UmRMK7CmFg/As/jXpaAojCcfI0AYBCYfGRHex5gksnGKmGvCl3PN9jMLZN
tQZaHz6TmFn4oUUwyuJ1xGcaTL6I0X5qL32lRsCug200glqn/Jzb/77hO+RIWFtbMGOEaRTriJz9
nzquExqnSrolnfGtgZtWMxY5zmatTFvHGHWQfFboZ2hvm1x8QyUo3tR2w2k1aZU/qjdEMtvFBi4G
+K9rd8BLeVRUmTnGNmYV6bGZQZL1WK4Iz5v6gJUJgvZiMFMIeqAjxo/qguWzohOFbRS/wUdOm3Er
UrHyQtE7MmrFDK9wi/NsJ9lR5QSlKviKQTK0woinhrhfKxal7M06fkVUMZzudimFG69NmS7BwQds
+DD5PrUzkKa0M0IW/Ps2pbNix9aD6nENpHwzAjEhSXhU8pfR/27M8ZOSJUvxaY4eXt9YIB4lCKAQ
NCRBi00pdsqPaqvb+RgAdzD/Nayh0++Wh8wf8zNLpJjh9VPDGapLMn06kOOaQhNHLbd6h92xRhbB
hcLSKQJt8XSWOFTSidBLvZ5v4ecu1mKAeg165OXHvCRj3OhWiDoRMVf5NXZKaEeasAxj5r3KegEf
dGYJHgeI6AmbfqvFm34+lyWxj37LH3S8m/a14PfuxzrVpcjIY6bEJA12od0yTHX5pUX8ksa6l7f2
cSgAcyC4SyRp1LcO6whG63RQdGj+WHZ+rpWfJTjbmSrqhkJZjYD6GmeSaqOr2sJoKomyXRuTX4dB
0tezYXX3DkhKWnd6A6nTrqvEALzVlyugVkBgtIIa/Zimx0JAnUZR7eZYJ6yqn5U9FHJlku2c7WHy
w8wkWg3TaKuLTil9lkxF5kXdGW2eDlRfVG37onoTBSFROqW0UxapBP1ALmWKITmpM3qCV2uV0NvR
U2dyNFZFkxLB/2MbxoSHi2sb12gbFLKCNo1l2OxaZ7eTH3e5WYqLr3NhIbEXvkMggmjKL1P5sWwv
/Y1r05dMmCJrJ042uvL9vSjAv+wvJNKHF2/kX9CP302HVH2H3gvjunq5Va9xq92b+aKUki4HHu0X
j52+0yL5urKmp6ueJrOjaPxhwz6DZWhnbv93eefna4U7Xi9Bbp3H1F4RcruzQeUrUgPY0f292p9D
2J+FfNfi1Wg8H2wx7rqxQCx+RZyAE0WDOoV1YrJNy9pfq+dWPPkiZ0fU+0KUX3VTqwvGZzR7wlTt
X/yrSvpAaIrLiD53slBmAnxS4HgikLfcOgh7LJffxJDW2bGOgCD1NjN2lPM6lhEfYqG+e7mcEMV+
LI4yx2boqZIVfT4sYRWAIS0yRTpYYPBBZT/Ahj3gvObGauIVcnHmAv3ULH6le2P0Cjlf8iCO7/Ao
Ews8LaM5Bbt93CkBrhNSvoJQHsHS4FA0F+rRubboIFj7lzaAv2RoIncuj5YAaNdZub5z9JM4HFVP
XTsdjO9rr248TdX1OEixdtw3NiiwIXmNxr4JPHWXvzXXApeFPVx03uvUEw7o65RcIU31buxTaQT+
lisQAdPB4UNskgOcT1ttrJZy8DrxdYmqorLWhTbKPhf5RVS0/VI9Thj0nYnwDiscDzUFug+l0Dwu
nFQ5OhxQ41NkVs2ew5GsBCAZNqeNHrLg1DZ/uFPXR3ysDpahTthTMYa8tM6UM/D4N1iBXKP7TrrV
CRla2DvHHhGsKYJ5G29o1i0vfGhKnsnT9pJdQzlmEC8uqDQQksIP53M6VYiT+MSRIFysXP2vhNQN
dOfB/bn+kn8dzuUBx6drX3cc2USwFnUruRoHqcK4YuPgSQESG9m8EZu2owmSK3rg+P/TIxC7Gr2I
BVpjjBdVEZE2pf+XBAq8RNpCZZszgMxNd6n4tzqevXee73S0T30Ty4nlSwNaMmKgduCfQLRVBHv3
jMhO8FzFE5kRClidL6xtWBDg/E9ofxSNX6UyV414MeLrSEDkh1PWBmYyY0y3kxyustkv6PHXCUmr
ch9tWswTZJYqkkNLLco/ijoArzcEvpYDuhvrp4f+hsH8fGYozJLnstqtMtHl3GiNuj07ywM7XDTQ
FJ3SmUWPEEUB5UfwvAefPg+n5EsYerzHnPlo52UFiCcT8bR5hKlAdbsjmLRl/NqNmKWsmUAz1Utw
gtoMcd8cg2Tq4eHNc83vTEgmNkPCMCVWh7JDgb4KT+3b5xzjkT3PG9wDh2qiTZtarB57wEOo8/se
FYzgorFiATZWCEWpltTQ0ou1/DNyMdxSb1vfSjshez8vUjTZ4cFPtmgH+5RDrCnoM3m0Hm7UHAwi
1O8+xf5Z/TiuzH5amn29LeRhvuOX6hHrgQ165Wxw6JMhh0wxnD6zgOq58dBHf4bP6cpYXJi9i8BH
cbB7AKx7/c/Ru9m3vv8OdZBi3C+ReR2tU6y3P0eDvD6rUSCIusUqMuGVr3NhnAywBa1uiw9EEp2K
n6F+09x5Fv5UKS0PO4F1EGzX/C2n8P7sLX3vGZzGfY9t+oDABb/a/R5EW82PYQypz4DsUR75/gy8
9j5WG5g6JEOYuKx9rK4glfZXRBpqBOWVafqZon9nJ6gLZetDU6pJvQvGjFewElnA/JFt58sD8rYi
E/DBLXgfkUdAPg25Yov0SHuyxImcbJqKH6E62pQzW03lSzg/hahqNzasC2qarAkkXSaS79eBquMC
EYMR1Tzs30ppkjlBoWfeDhq/8irR2FtPqUjDcPQ/BlpB6tvgau4SwcurCEvz5g4OT3xsT+uZd3ho
4NZFnR3vvcyNQYJ0U72AiLK9W9Pq34Kk47Y5puRUEJRpc0YhMd+8V4U9qwTsUtust/jKd6LxyWzR
iPzeM52RJva3cLenY/x6G5gesl9B76JMR52X9Fv84W5fK1BzV/JlEHYmYkt6mmguHStcFEw/fa1o
TW8XCKebWHAmmIG7V8tH4pVnGN2E60YR+p7wtqD20bqjBd+NJwxXO+HkBhY7hRypEi+nKC15nCKg
5SJ9tDvsvbyScvlVoAjc4b0jb0m9T85BX+S03eb4SVXCbz9MJsyJg5zcleSZSID79sK7Xggtin3d
ieOPpVGUCmQXVU8MpLHiEWzxQA3ZCW1PYUBQAr4RM0vbDECjodHRk+fz3ZOiR7DvsKVFGZ6PQrTk
8fJOcTyoGCKWULz2HyzcbIacg31QNsgkBO8Z8aIdDPpD/2+WUtfu6mDHS+28//7KibKROvQfHTZ/
pUlOUqlFyh28DHsdZmDplZAlSLgtW13jhQDo8o1LBLyF6ZDQx5Qc/276GLqtg/48DlUoxxglZaTf
sCTgTyCgun+a1mfHm/h2158oUO0H2aKFm1DdbWgWfagylfXewUtFnXtf69hxMMzK0e8SPssXPrWr
tZtWuEEuaFvL9bCbsjOii917fpEX1Z7CsQHtenabJ1KbAH7+gGXZr9C0g9AD0hfUpxyWFgKgDclr
tRwH9juWJiLTw0dezOd+dlPq9OIPf2pWoGfhB+8b1d+HC+lSqDz7QTcfBqMbEbXnn48Tg1wC1re+
5WeuUGfT2kxlo2JihZGU5kpfzSdWqDIxuA6Feh0tSbJlrb6r3/duRBtxOMRreiCAqtm5bdkNb4Ri
U6iaFm31Xuxv/q78FGAwl3zDjuPCHrtmho6bJCyaL4URaKcilPLTM5EK79QY9X8oTqOtdASf0KzI
6t1fmpny+cQFtxcCe12VhFWGnAYDzyQHQntqq34b69PGJlu3KtMTW5bzcdL4xYtzYYiSRcYOYPfl
A0ZITxhrHTY/dzEUfrXNYpuqYf0LDA5s1x+C61M23cp5aYZBlPAlyQePuz3LX3A9rvVgH1fi8pb9
7SU6zl1GblbYwGc4joIyXawLGw+KYXLTCmmGODUArxKfPGIDb9V8qPGkE3NVpPAu1RhpKjhwySwH
r+ont41M7Pdl6GdaX005Bo/g6R7NzkmUh6gUMLe8i/KUjRuuL5A6VettsrCiY2jyPm3hc3m0BGF2
qWdMoIX/RRk47xtajUUehnNypF4/CQdL4FKqYkO9SfDXfNOxDjmM30xLVqVfFQ2w+XuLZ5DjEgT1
9PetX1xA4yPbAqvxglfmv8Wk/qOo5XurSgmFhFIpOFUcIsNCsKzjON49cgLVoQG7FFcWVzbn0N5L
0Qc/xfT+dANKFYwvZm29d+yu8+jmrUqfmsmnJ1KpIsOBHYiaXNP/fkEpRWDC3MscvBB/deNlfhYf
6uaznmRxuAMJW1DnClreiPEzLD5MeibL05TQdUxQ8BH6CPLm0vsaRwE/FUyi/rc/lRat1PIGsXV0
eNFwyM0E0GYVk6LUW3a6//yfUvhPXQhPSOU9Lu3C7MggaPgQwhAbvjCY6Z7rQ5y/kVGZxM2jCjfq
xkg15+zDwX+2KIOlU6pj7PXDiLl+gVYLNee7VRbbIlpEGzep6kbIFdVhNcsMN0YQ2139vU3LDNqv
jF5aWQuTHKxHIQh9DHcJBgLyOnY00ZnECYvxenZkezpn1LuCKbsfb9ZKX/+2KUt3hoaFr39TNa3X
rAa4wWn3qgUmaSgbHsa0STu6fxuM63og+yc5WQlG22qzH0MgpiHZStvjL4Nz1wGTdtm7/9Frb+dW
N2d4g20Y1nPAPan8IqxltGd/vFCgE75k8ztVszVl2nBwL+/t0B1MXOTnohj0M0HSSBsvxRo57/Y1
SvBcHwDcpjQk2wHeL3Jw6NwqH0d5HIIIynEG684JFtZc1TdDeOlQEXannZkUfb4ZAbWZnjntim15
Yk8wphtd6/sj0RfEDpuUpzsy2Gf/vJu917sYrZP5+xHkNDZkqbngsBXO/NxefUOjeSK3ap4wmdFm
9NJ44giZus7qwtYenOGg7GB2OKLPuhfHwYixKaYGLNg8yKUOLipVn7SX4Nfy9OuxpmekbXL/zJf9
dFLw7c5ChCmc43NAFTmcgYHLKGuleA0ZZrjlvMdO/i+S47TsXjWNTBgBAQ6TdWI0E9M0ruKhHVKQ
sqdVAqlR9HKgkAqLDbjqalNqJG4EAtRpNVWNVVkrMT6EF7LFOPIPBglFogYbYL/49dCnu+P6Ukxm
LHSmlENDJNSE0y/tdFGsS/hSPJKCEi5GKCP1KEda13rgpOJmP8VFLp0Gx1BQUcmD81D+a+GxWbpK
VuGsqsQXowrIvFrvpLvbLs+awhDUFnkXkVsidLjTJRau0bpmxPXDl8lwyG8ztAf6d4CkItG9X/vF
9ho5Ai7cNUjxzONwXs2PgTCcJT8VxAxOmSoFrYcS9jt/cB14YockLsPNlVbGzQ2yhY2UwVghvMx0
u8jtzbGN6VCjFisP60/L2Bj0rE5BdL+OALqleOnP6gV5x4Cho1qPZMjz4UjUybijArKNTPX5uoyj
eeBX3Bv9r5pzmoFHlqxVeU0AxucwJvPHzT9k9pz/hQKz2yON3YWnZGji5yBzCtiMhEFod+gKtl4e
Zhww85sd7EKsyIlTQ8OETdaCgkQu65f9vhlsCg2CZ2E38F1fA8rMWiSHX4D0M0EvEC0DqHCuoDPZ
PrtnIWiWfBHOSo48MGXSCm1BKp/zD3FI+57Imkna32ZMJ6Uf+kqj+GmwSJFitL718aC872L4CeEJ
+f6+MvQrJsYU0Fm2uPAynp9vN/0FLrGd6ZG0uMjeBrQU7ZV/lpCz8O3uvKo7rFzlkZ+eacOklhJ/
4a0IDxtBzXcVJoYMlUKdQEgNblRVP5cwu7zFe1PrQRWKHAXDZSCg/T6kOgzOzf6jTKaFjPNK7gfR
yJc2+ZSXy0MB7/NjO73RWsagM61UDcdhDOuDInGJm8cTSieVypI8nEJoPZ5/6HEtzBCU49ic9+f9
wT6yoI2+OmaQ94fGmon15gx/bKhj2+o08pAZonB3dEJa6PiI051KO6QoqeIRvMKukbY0ftH3JL9u
YNfUc3TdT+rdLH/7v8sO87bF1LW+1NW5ZOD10tUS/HISesOg/EyoYg8qdgJRtd6XSTo+xu6jpThd
DQJE4EsCZKr0yI17XOZigakvGr/JA1r+Xa/1sKPBozaJTimKgGLLFyRXgweqTFHrWQzvEgVz9/Ul
r399hLKheY9ElN5/BISGhVCpQQRyh10lJqGvJoWsyIgB9lCxW9CDxuQ/guuOmUqsmTWOCW9r41Iu
BYNxSG5jBGYnPCvrfAwD95/f+rtLOAGx7dLcFyE/vsWJHOMigySxq/wsgk+DI1Del8yCRjJcwpLQ
CEWEAE6KVjELJcgqAJ4CcHt8dKLnQBhpZnqvXX8PJHkpAdgF7EYdEYMtQnXJlb3qvsu2FjdlHP5d
KorjLY8b8d7Dmr3Ik4oIVeVN4z9YwGHIo+UXdI7Xiw6RxKgmqHi0ELjAbC2QE1rdafBNG7loS59/
KcrmkxacMNECqQexxejAoiRulKOZmuabR1BtIxeM4IuVMpks1YC4fBQfDZZpweWJ0yfNX9B6/HGk
KopsPLshGNVszPUig8I6gTrRmO9Z5yhjd5RUphNRA9Ab+K+5kMUqEPu5UmcXQPJtg8fjYcAqmpLT
eJ9Z2iShhFQ8WyxxYCUBTnmNLxRZN+piP3K8WzZs2y6pJsrx81rooVVrUJts/1OeiQpWzJondVUX
tImJbfl7aK4vN0vHpMj5N0NV3FgWIn6PFcetOmsGcHsSX0dKMifjey0bUJgBnc8obYzB+2dichS4
SJv5FqaVObx8cIEd0e3D5+qqYgfG4mHroBLfQG1mxbwr69aLDHBP0B5M/pU2RCIwquLdQTIepKXr
oU8AhHc+ya6otQEvXLlJYNCe6hN7gIX9sHAX1xPyQbeLWauWGXatWOqe+hWGZSMszwT+pMnQoCWQ
B6MfsWoV+foGWk6E6Z4mzNqpynnmjWk11dCnIWKfMWR8x60iBcS6EWXadhSr8cNRHbq+15/0FTDS
vgJUDLinIWsPaOUjI2NWgpV4FO+yC8mfe/70P1tdgBL9LmLd3c+QtaOKo4pShZUf46nR38GENTNO
zvRhurEU8L3AriaejRTgSwt0xkay1W7LPqkzDQhk7khgCruepp1lKSmM+VdjTw6IpZEi14zkUA+P
+BfcE4/bup7saDkb1+VRgf7tkYHKgIFwc+EExRRJmymjbm0VlXcKPIa3bQ98xNn1oKG6QtY1KDlU
Vr5Emid5D/fHF19AXs37bj3JbVCvvd0NlJjlSCFoO1dRWx671VrQJIZmk1PqyiFTrkRm5fWQ030t
6Y/QKRmVFtdBYJySvyvjVb/FiIyq/qM2vr56s7rdujlRId1VIybOsBZcF2z1fdhUxzXFD+3gau4C
jpEZwDlSNbwcHJO7GUQndM9CYH/lhI8bg7SwioUxyKaCAQ1C9TLAPdx/y+ZlQEke04/5zLpT/g3m
GJC1t3L1WmtDYh+pabi5bQTRQ9ouE8Tx1XWoScZhJAdHqA2GWboSDIupA0gMmKo0x2LIXucJ8s0N
S4KplB2rcNFQiIqi7OaudHNepRuy73GsWI+yBD2eY7gBSurLc9/MC0MqHrevFowQlELvNTUO4rYJ
UCa63XYCR4ETyi9zxoDyAtIMsFwanfUNl4pLNhFi+3vCfRjc+aLvVO9t2IHzN1BRryOxbBp0Bpss
jD6ETbjcVkYGn2fetkfRWDNX1xQgZrO6bvw+QVhmDpu6ZL9StwZ67SzNT0sGeuH4Fno8K+WCQ4UY
vrlbeedKRfqF8fiVdNBMuPzl7vYbExL7vT6SqmduLX2nQXBO6Po84Q5fWfsNjlLuGXBeAVf0Nqb0
fxcDg5bdJHe3zVzMeRUChV1K5Ovg7b7tiC/MNhvj+z53ubDiW/nT833isCOZe0KhxWOeP5bs2T9L
O5uD8k/C3LHlLZHsMsrqfU6J4YrY2DmbO2OeubDzPI/1/7ktZssVpXLJDrACk8XEwYIQpjSWzd7u
CYxfIBJns0E7FAAZ0yHrgFIj1Q0/Q+1BLqcCzZDnP0a7lZ/cQ177EFkAiWLJV2T69r6tR0gKE6v9
FypuNSFwz+8cQQFHdxrZe11MRf4xPZFkztdWwVrzGxXDn3xa+vgY8L/MBerBT1jKTSHPyXzhX7fu
H2fuDD/8uUPFhJIkuD8g5J0Zbti/sVgr2Y2P3Q9m1JANbOaBAdXuqfV/xoEKcVV1+fX4ccz1MMoI
sYN+TJnec6Jfw+hMNRZzlI3+MaAmn3Vn5IJ8Ad0YsSAlNdX0OnCX8djPbChbvdN7f0Jyzr7Xdpsd
f1FMkCrGt5N6JE3IoUn69NVLwVNlPg7uCm1gDKxLCx52e+Pf2GU1A99Hckn44XPWnbpngogWlCp4
4C+B8e/33O9Mn3qWaEDRhdb1i3SYdMFdf/5y3mXZKcsE9xyUvfOpPwfXhF9KOwNxlNxDCNrRhQd3
H3Zc2b0EBv9zHZNySaODYT/2sUjTMcK5RyPOEDVwY4inlu1fvNQsKq22l8yegA6fNNr8xoPGi12E
2GnIR8lx/LGrb2jrcax1bHQIGhluPkGVLgPx5Acpr3tliWTmpgv5dOQQ1p5JvIuWvru+t33dFMj8
X/1ruTe8SoR2V2Zu+sksDjynpKqGhEkt0KgpA4adbZMrj3BpFt6EtbvcIYwsdYFLEWaLAk5EWmyA
O3YC2FD5Qtn06sJogZTig/aINzpjX7TrUmVSrefHEk+h/ffKxtBmAj4/FnRa+n6fGhq9PeLYzheg
1b9wCHa/8TffFoRx2Ajz3ZBRGhI+pDf6XVOgmFrzb2MFvKWm0vTCdh6Jz5DG+o/ZjxlO6rZBL01B
80Vj2dgQBt2DacrmdbBQkQZlmvka9xqgrnz0yyHV/b1yTUhs4rXrYOGFg5D96mJgI+hL2VA0u6u7
JQBnWlyGJuEeUnNvUzAd9KE6pr69FvKzo1M2P58bZb24jK/WUOiWZ0ejlxp7gMe40cPSHM6XMyY6
uXZHhF4eMMx0NSJu4bSd0WzHuLw+C5twjgzwwzoeT95U4pukgwgqrUWYIBV9IdIXpNhVuf9+etEW
eKCUX2fgPnCTKiIOX+tBA+E8VSDbwfjhavwpHZGyAbzXNpZJLjhstHKfD3WxR+Cw6fVOJCCGHGUR
2y8/cfD5+/8OZ2rI62d3Xw+jz8hqBVP/PdLa6+9Pw1bJc1VzGD8wOoZHnHXO48pvWyfm9ZJdYDEX
UdxzVPzVK4Iaq+ZdCwpxHO5vXPc37UcqaLt3oTMcVr8NOKTAt6e3+ciGWz9u4dgeqKphN6xQLmHc
ABcGKZtxzMV7ZwCfMbQh6AdTM55h0LnHLeuyoO27Bn9LnoUVdgiAa0Al8iQu7f7xofEQfH4PPqyG
w6+JZ6zgvDvw2bu2UAGMXnySJ78YTnIolJqQxRazTjrOU7qklepfJ0IF2yW/NdM6Vcc6JizL+DBj
tFClXCpbv7BgkmxZN3qamUBDoMMyUSA8UNlx0+9vj9fpLZs+UeuK8IW2v5mwu4sBaCrgO0xv2B9d
sjMIVUfTDJ+96GTsDt8xkGUFn+hQKxPuq/7IL1AEJPKf8jhKb5EicGuW8Iyb+Mvz9s1iTowuIfUP
cqhUyXhp9yNkfJMcYPUuwRdJTpQ93PyA1MJu20MpIOsH/QSxZl8IVBuE6sdMBmmS9eUamRncuJKw
cXqDr3lHsHIXUg80PnBX2SPfeo8RbWf2fILz7xMJNhbD15UPRlTUhKn7Nu/pAr8ZDcj58XmYasQB
LNFuBvZze9JhK+HaA4+5002xsEQjfxJpdox7qaOXh2Xx7XxyDEO6sE7fx3Chxi44owl9y9hOpRv0
q/GALgZ2Og7AEEgzNK1U8Y4M8cJ61kxZKulhYiRaHNkwPOOTRNU20QbT+v+ur9DDIDOfdbv8tcqS
/3zfQckVUOs/hYgNX2Js+iyOuDFxSXQQShmW43ym2HZerpGxICm6tWDCpGk/cQPGk1yojdvj1ezG
V3XMGgLJhdYCjTyidZv69YpyvUyykJvCwxwhDtuPa28AirEXhFYQ0hUY6zXbtaNpYZwi6HeFoUi2
cb+6ePWu6JA35iYznmY8hVbPD8850GGYA+QDOc+UldN3vZdNUGVqRwLYJpwUOLkT3LwwKV9ZixRv
0IeSchyLnVUxWhRKvQEcKULTcyzpbsJMLQ+SbeLvO1j6euEB3+JaUarxJWdF0hhtDT3BvKJoTCzb
emcNrF61Y0r5iptDiPb9z1kOMw28z3DG/dmbvikbkerjfj2hZWpQRKfDF1yJe4/iZgYZIKRyL3RN
yfYgOuRSQVFZkCYu4M5iVA+NCYfRfKYQWido93gDzWMRxPYG3hCKryDvoNY6vpXiuDxoO+KB1Pn2
JRDxQYDjTx4HY1bp0KD6vegmrnmDQcgSmB6AiZPo1vS6Oq94sg8rFhzqkUeTGtqD2j0OLl3/1ddv
AS8uDuGBQKJezxMBjr5FiH+vEEED25L45S6YwrV9thyOzpBV0+APl1XF+26sCTKetwZmgbuIVWcl
PWsSHuTwe1+MtUua4QYvy5NVDaWJgxqIrwnXsS0wlQNxPyc3tHTwgE+CDC5TWAImxH81vYEOFKAF
9u7Sn/+rQdB01T0/2UsXkmATEPCFDyodw7JAWmfjPGK5O0IcC6Y9o/K36qUVyIWD1LrVrECChNPl
HoCkoWi42W5rkwRh6JJXZ3crYvu5oJQG7KvxI7B2M2Q+v4ySlU2ZTzkoCUOT8ZuJe6q2TN0u2u/G
WhVgrBHoIs9aIeor/TWytJesiUEUL8mPn0btxNkZ2xFQq4lpxKVJCgcAaqUaExVWmMJgB8ft1BLo
b0/ebkBNQ/tavQ684xOov4Gyp6dxpiuDV2YeRzWF/0o6B5JhWjLAZru2dtx3WHiwlcSsuno5RCnp
/tiH2OWI+snxKnNrQVZsqsPBkYhYJuHyu5Et0eUIYHA/0Xln0PyPUrafscfakgEONuCH5k8xOxz4
6SK6rtOqEZqkjCOTBaCqnnUVMeo7VpsUecwvV7fWXvqbttpE8Em8Mj6pHCJ/Ogezzk+N24KTOr3Z
5GupcQQLzr/hYTg8SHZI3gbbIeXevoADUOUoeYEsVgth6HgdrTJpC7Em44aG6bmYTi3YJ6k87cQp
hdyLPYiV8dXkNVSIXwAwrcEP8AIoyLaPGuTAaPiVaOCyHO0eKNBgIthk4QLJOHgev6lfz4Xh2who
5d3YB+xLywM3S3lNJTB/2lnSfdABaxX2dheRPHGeOX6MgW6zSwqHTpajYdKfdBHD9LBDUNYeeyp8
x1+78loy0ZBJFhPneiJ0GR3sGsErt6yBsg3Ck7X6AKb8lOEtyhqR3rY/5nSwTkKo/CO1obMbNy/k
DgXJvo9R+oomQoy6lGDaJKu4qGjvGMURDcPC+WMcT6BKDziSLCF+uG9SnagXBzfiF1cwemPa3niP
snhhU9C7tlXMFX2uZE/gHUQEqqrMdCCvYvscVYp3Oz0EBixrSHRF1Ya391g2E6gtU0ghrHZPELBW
ePoFYQkOi7qXnqTS3ZNyINYWbuVez7O/h4TL9eGQqcux0UmUBiYDPQb8Se8x60xeNAc0I2O8Smch
XwcoJnfgK/eGEWPApF+3JK/5vrZjqjkk5E7qkzVwacywtrt16C00bzJaR6MrVmDdAW8H7M1gVXPK
IkK3Sm+NcGFrBmpAJt2DXXOw81Od+omF7izOhTgwga6qTaeAJIEwFwS0wk+vP/fF7AUO14cQBdie
oF7OrIzaf2IrqM/YW1vz1lbPU11b6adA8VVo6RzSop+7zkA2LIBkm4J5I3vhwt4ce0+Dl4Rd477Z
nNL4VT5CRQLCFNwtzUvf5QnDIL6GNeXZty1E28JOTTXyiGAQ8y2Di4MiSoqk9lpKeXgc9KlUYMQ7
rsYQRqXnVii2NFD7/whiluXQeWb1kcFIYc1EAvUwig5g2blXVR6AHq2IYKEm1FH9AKeQBdQ67Y01
EB/hO4nStw3CSgJPYwekm3mGvEsUChJoyrzLVAvACkXu/qO33TeiGvOSjsGCftAQLDSXdljVm+tR
8sDxx5Byi9CmqwU0EkU2aHtM/+3E97/Che1mYsqbV7KUj5uXLM6nCrXGXlWOs8j4jpZRcwq80Rnq
6zSobxKQH0jEiFZGuNamcOerBSPdLVZ58eyTC7gHjEuc3BFklY4eh1V44rg6t7OD+QYPfayJnbdz
HmDhLJhfwCuexMJJ50JHmcg21ZX7h/PuQpITQh2gX/jxVX7OkGjjfyW30bBFzkipIoYKjpfAj3U3
eyaBOZOMPTfYqLB/usl2DucpBDKZm9EmenSSi2pDjSkF2ideiJRnKsu0ijRkC8b8CS1EPZLXldDf
yXvWJxUjgifOHwLY71Hefc2FwvopEg8XNY5+btV2sLcPHxTtXRBjz/V7cGowAuezDv/YDlYVOveZ
Xrh8XbeGWipsBnKOi4+FY5r8qz2htWkbMAWKa49jTL58VgwjWti6I9+IGb1/NkUdn5nIyo2H0jrV
7y8qgl1d7YlT9UviuJGs3sQcYJAKwu52djW4AXp/+JTsYodH+8fhZixMyaMBFMYfGots9aRU0SSc
V2JgTwnnVnvNSUuopJLIKJUGig473qaRhuGaXmZ+4Zz/gPaq9HGfAipUnle6FoxKP8cTU0D3i1Wy
Bgr1+JoI0pjBtS4PxUkXEL/3K10PH2+cOF7MG0l+ym+VIZx97kLkKEMa7iHrRTpEFZbGEX7mHtOv
N3dzvqYMOFoz/wu6Fx8nyuD7ZRpQP+8rTBdIKMLMj1Wo0xmSvmviP5JJQPoQeeFWz7Y00WWWXDgG
912juRZXFvy4u3g+xpi5Ajoa8Ew8KsDnp/Ov6kFlQw7pEUMpOdgQxe0RZKDwftnIJVaSs4NVrfeV
jQ/PZb0r67X35vOwLUacLhXTaf+lpBLqAPHJYZGC4eCSTN9zq6eeQM2mQNUyh/z5jetIKmBK6NHZ
HaFNBzNy0HFe4BObOhMFtuO/6lpI5DEbx6IljiVKnTCgPSMfZOcSZMoCUizTBmJruA5IvQIHc4EX
Kl7G6Z4ZQeTsrCJGnkMk3ReRbETFno6tbPs0+WWN4bfv7Y19x7iCiKh4dr4Y+k0aQQApLZYByUGz
0qXlI+ozlGWb9t3/UyIDhJedTl40hlBggEN4itqMZpTcE1hCGpkLtiPuoo+kbi6DFHkGjeJezQju
dC91kXy+2aKE/FsYAcItZThNcLORNmlz+z98cVs1CnBGkMMAAMDFmbIPDFscEWh2Zalw9TnZ3pbx
3RRNNKCSj9xD2sjTbcrpMhcUOk+YZlxRT93krG0ChK22QoHIRP+D3A+YFGYQ6yG4uDR50pAl84QZ
+d73b6LDa6eMSbq/rdtBlcPQLWTb5GVTcy0wGqftE6DKERS3MOXw+YiSSukt0g4aPsFHbVleNqYX
UJ3BiOpOtdAQi3AEo+XtP9M3Z2TIqUmL09K9EXnKU9/5JYze1JoaHpaoVwlz/b/ODvi+v7ywKghG
x0rInfbDl0+YLRZwP+wP44Mm+ba5RKdksPicvXmVS34O1Xr04imNkspoG2++IvASpsARkq1qH7wX
pOWokJNe6alO24qydLtt5gnn8xkkocrojiejNzUgh2wFHtWBl4AE+fk7YzRRc4VMn5DQnuKbHBDd
Burt4bruWciJStfAuAw2TKyL0Jc26U+Em8x3w9wKWXyYov7L2co1pAjlirufT3wLRq2/RW5MZovS
xwhRahZfsGGoj/vGfeMj+4VZh63Bw2MefQYLXYSwgDWq6LHrPqQhQKD0AZpyIoExgyWYq+7mZQos
TIn990QeZMgoVXiiFpm3wTNYkYL6mS7/BG8/kF2I1/QWqgOcj2WNFPcSVpdEG6XBWzFk3JOoHyJR
uS1uH2EClrhUvjk8oBtdpvsgt7YWmaYxEx4ow7QVxij4SBqp/DxWRVD+CoLprYJqwKj2UgRWHgGp
f0Hco1Cx1bh0fBJo5EwyCjltYSqaiMgjsZ3QbyaQ7k7dwXT8z83/1UsSIPhq5kt1vHojoV7zeXuS
VGEW1geXVYo3OfKfxIhdbQ6U5nPvjaqgfbfJZuf9+D+Qdl/Tbe+Ad+31tOPa7GqcTC4X75TabLqR
v3gRpAPm+QXnMdJqnnqx2l5sRMY6TKLGd6GviJfB2cXqmZDPbqRClE8isnpmb5HQhH433+xmho0x
ZHnA2gHGepYKBUyLYPqF/6861UMrBUnxJ4Ak4mtM0hGCWnYsukbGc1JJgp93kXGqpUdXsnT1KiAI
om1tkt8TpCCPPRX7oHY9H8SEgm/BFpFW0AJqzojqO1TL1KUlzDFdzRfzWBLZTCvo1nOic37jiE4t
4knTDW1E70zuPF9q1VXCT3Y6sFUigBW9P6qhC8AjPX6HJOUswIZowox/oeB11XhB46NXqlsFBacR
z8zNdJILrisaclSoGe614ifZKZ8Hu8b1rKSobDenoG9WCnBuqw4AG7INqvpk+l5fOdq7ASKKYYMh
tfh/ujjDFBv+Fw3WxHmCaiWo67SPo8wRJFvkJ7AJ6KBbjMiydLhhADR5SWV71IgbBgyfqJfSrbEe
8AuwiJsYBwkJY97ctGUdprj0OKwHXVSWZaVSS1Etuh6NVbYPgXficltWnb49pr+P4sFc0r37MMvH
q4/eMv8P195g9LUT3Lrf3u1MTLjDZ0davb8kATuGTg2UK395tGTKNPFAVOsnqYRUDY2foRgyL2ns
lXphbaGyhf12aYKye7UaZobgjhd6QIFr87zMct8LABbJGtHWNJ/ya2VLLOmThCJeYgXlash+mNSo
r1E8BKXz+w/LJGV64fTSkn1KHb7VUtqWpJENfg9fre4HhYmEMn1YyX2rFA7AIHm9fS73jxu3+9+a
hFQjqrnhPxXbaUIA38jpwJpfGmtdhbJCGAfdZ0szYXTDgBjYUY0gqn45nwlF0fZHH0eQYPd3DmTV
W+0D7ox1TtWorJCGgFKXkvOEob9cfHGN9Meo97QX6qsYqG554BlI+5H1xfYqHngf2jmtDZIJtj2n
VdE5JUQIMNPOS4XwRq+aIU5pYKREufP/BbBBu5rKtn6PalQGVX9Xzok4f89XzwngikMtDQSp65VE
FQJpnM3wDmotnhmnhaZkPz39qJlHkIKkJkPAaNRoaDWlU7vZL7tAmJLIR9biJG12BsTmkP1oPbrA
Q+7ljts0AarkFGHurQUEdlyeuMyHGlrZvnU0nbZTlA2JpsCrzy7XdsTVrhS38TipwcLw1lUg+ElC
noyKNovmcfPHuXM9FEkSyxW/RGUJ+/IPFfOG6klddmxBsVvdGmei8Fcfr/KbhfcYkwAOWnI0YwJR
eT5Vf91KtEqAUCbRkaf7NbosDQt2E9yYOgm1U+xVM/YKm+/Ie06QoIT7DG/t9TdS9W8lpSSChoKp
+/RBuHH5Ggs76vq0smV/Eat8tfZ+IT+giLibyX0ot5pg7G/ByxJ/OInxDMm2NSW3dReNQ3yUucKQ
EJEwfqf6RiDCtwD25PA5tz2yHI6SVrJMalwaQXnHOv98ZJfyPhzzkHTzsra0cGM4eTd157yeOxl1
UrzKQiZdu/UwOKMEUWYl6CT0v6a/bysQSW2r69txoG+AHzTQBqQ3RlzYg4YYG5MQPbOyuF4Ddtsk
kMZhrCSGJMzfEjB3YQe2KJALJXfZzmVaaiT0UEy+qJqUe9dTtqAgd4Tq4hkfle8GjK8lhbGsWaQB
mtRzoVmYJU/PwRkBlnlvXVS9fk+OjxnVDdn8Bl5w/yccbSSQl3zhD4W804qOEQS9rVf4zd6TtQYO
TKHgdWXikOVqbRzR+MG9xMHU+TtOK2wMRImcLdtXdVxRmqZfcyg1X6DyQiAH35/gILvDH6RUhJ09
aeiDjvgY1DVgHXUjezzj30tfTNudfh7ncESzQ/Udbszb/AVkmL2U1pcNwTK5FUYL0Z0RybYSSjz3
tqcWwlao+bxNgNpbzVAj87oG4C9tcVeelbtoc3YegqazkPGl+CFMf7sLbVkgFqi7B1x+RTLFeG4z
JDVDpFiemGwu3FuPu/OS153/bSzqn6kIgwWPhH3noLYx7Fbicl8Kt2bqiIwFbkz63HsQ2YJuxCqQ
MQ4wEIIG8DjtP2VHDCVwGZMDOGpqhaXYAdQMnvCwmxQsq2SXtk7AdfTxdhaax6NPuaOqybXYGx6q
J2ZNF2bYfcwsVURTAx0FVm1rSJpfHo9qOEZf5mA1pz0ZXBoPWc4c6b1Ce5TpYSiZGbKwC18Dm1GO
075IR2aiVmHsGrYXXtuD92v5svHUN5sUBgS96ljY3uSWAmflxi3pkwxsfnCUM7dXdmmYtLshMSQW
pGjQNm+arglfnGbNoztDv7n+og5vdOnFBkpLY1BMi+qViQdrez77TIUqXdz4KZ7+2younyTJthyp
C4Wit3oD4X+Sy/5GjqW4BXJAHE0tVNioFE7FnO9SIkiCZQROHo/p1b2MCYjnaF0ollWsBdDyEOrT
8rZ9ca9ZuL62VP6nALrdxIfMUQE6QTsj1FZNkkwrzcjDXHmFG/3EDUDoF+A3XmfNowakC8HLdhGE
aHk+uqJLW7QSO8NpNXKrqMfFyAoXnD5b6NiEPtzbAgRW42Il6wiOZH3JTNb81AnzaBhD0ilBNIIy
/qxGO3TNRNUYdCcx+Ki6uXu4Ys8IyjooltqUPKadVS/fA8DUIEA7hbey7N2RanMF2eBO9ckcR9Aa
wmT6nkpfsrvt6/cfm9CyZWQpdSPX8+VUTdG99PNNqRjZwo0eLhnYKfABXt5fFfec/0iC+G1G8RlS
6tdBI9DeCEZfag/Le0i9fWltA9OTA0hrPGGKOeBNsLXv8kpWoKKywDwlsMqNjC1uuhh3jHT5CkcW
qXcTrGjTw97G2hPymHezQfPu+apeha8S59OHVwFWG4pMMadTQc/WA/79oLMgI8oAxIKPDHgvhZzF
jRC44iz3So/DCb9TxzHgbjqHHXXfgmziHMV/dRJn8I1GBwHkEW19BnPJJLbf8ZKnWX2OodPSpQsd
0vg2mQjHfNvLGKAMvQrrMywq9o+250CAaz7npLg3pgeC0IycbbEkDJgj1RKlWvCldCovJlumApPK
PaGx2uzMFt9ssdhI9ClUbs3F71elC7QSgJ8vEwRxUTF21Y9WfDSCAtE+nxohVjXCd92L+va4JtGS
cgxnXRZBvuNYraBUZtPlwrggRzh5qjxmAKMoTkS3O8thDMA1FPk/XY3exLCeDtoElcVfUhlF1aIW
cX9+7TNWKn3FlaUDu5K9wkdo+g7KdN4wvnPAKhAN9C+ml9mvy9cHIVD8y9Ccon5UwJAbGmhHppjR
XFDlikcNgMFWqv3UH1EcDOqUTvWu12G2edT6WkVQhg7DYbCK0mtkh5++Crb8Fe0elvT22GgpLfdh
4yzAImYczZWJCll7gZ8kOS8ei5mC711AdoJ4xTF0SeIxxnO2emAlaZqfXJDcF14XDubjVHXot/YQ
/HsTDw7deXnhSm2r5jNcT7BJukLeVOVOfXgisCxXWx0YWQMrp05KNpreZ2zAkNb5BFlng5A1FlhN
kEmYGIHLFH+gcXzR4NuHDcdOpX2KY02rk71PSjYhoHX+Ky/JRE1udqc+D0fWFI0vbwYsl9kjksY4
jmYkv9nfa23VJ7BnGoYifcv5ezjLs3xPyyPqajKNojh+oqHVp4wS9BAlGE++dRFDE1sQivsgaKIe
S+gRa8idw/QgvtUZ0QI02IVrEATVlTk4Fl4p3d5he4BoShzENztzdxu/nId/hJYtp6nh14uu8OfP
s//IVcV+Hx5EDiBonhH5HuUlOEsTDOruXENl8RqebdwZcYvTdvPII5OvE3t5SJ0rBFyKIUyzX3sy
uGwuenLRntkjZw9TPuHWE4mLQNU2Xp6H3gyJ+12FvIVn8Xi9+MKmF6NUy1DmS2wSIcabZGRtO3VF
JxYtqNN/S2JPGE6SLsz5lvB6+EovQh8aJ0KJF2GDkX/1BOevvXU8ii8dRK0vduosvCU5y3k8kW1l
9TIEObysMHE9x4cCka9FuDH/umdK1q3ecH7qM/ILjFm2RFW51uxDupam96ciCDMr/f1waYpxjd80
ZJF93yYN/NDPh9wxWUnsRjPKbdkEerQuMBR0mq6UnNuIYDi6S9t3C7Wu2xOnvu4/Qy4oOLcI4+9B
KZcBZJCbMFQdBiGBhdDCZdqVujmR5GGDwTyQAg9n4u0gGeWdAW2gAut2LLl6y7kAJXq8f7WuZsou
G7rWXmSVGdNhWCzUQRWWeiwukRRfyiHE3ds5AN2uyOfKhg/i+J64sTAgXX4/t8J9LvXAJNZunsQt
GkEXkZ2A33/Aw9BbRS3UffphIZSX13wkK78r4gf4YzremAMLG7HdIY8/Y0LhJ5PNq3JceAaba3RS
VM2SRevDXKm1b3//5FYR5DOkiq7X2zO6HYJbG/+g9QneAJ+c6f6XSSAd8qs8DQI3EvqrbHHrikg9
Ef89K1P/dUAhdiO/wbdcRWPWrSEO+ql5bj3SksNEAh/prmjEclXn+iCqjMQSOb7HuptR4HQtBDYX
2OQ6D6KhGswSnHCTHUlZo3q4RUBM+SY6zlaTGoNzIjlji3kKZDhLUixfnvFvoV2F0nCuVCkYjNts
NjotT3HZBbXb+oXmmr0ULe2AowiFueaGijtiT1++uzac7OqAK7DzJ2+UT1c278wMntgM42ffUEjo
MfggveHDpEnkHBB5JIwJEwICxcCV+LJublAbxZcakkhiybdWJXaZs9bdNxmyBbdYGhm0syhw4yh+
+PzJ1kL4LJVAwhNT+WlrA7SYtpTWJma5esyTQ4wzH+y5iXz42t9pCRhh9csPTVaMth9HdXrMjbaE
5J3qV88Gz8ouctdnxu+S5xPzqhQR04aLvR+IAkkPF0WnJVcck7DWqpLxBJSJc2DedHO/n1ApRcI8
izXvyRQ3xFiYUnt3DXgIkOWSNYq2HBhafXQM5HqiSTmuM+O1WQTEPW9tHw9By6egi197kwVy29QG
//W2548XUvyQ++ZoTFUSQiRNr0KbVwMaWgFiob6fQjUm7pdIfQ/4uBC8TRQm2AZQx3bdjmLO93uR
Nyh7Grqsfv3j5yUAZ21rOzSSAZBpgjAzfqe2Po01TtOqg5E7Zdx6ialMM7I0b2llMndey+qnIm/q
aQeYsqGarQiHsG+Rv/91X6hRIgKWj6Xi0zWgoqIWRi7hFUPIeYk4UUvWvnsUOE/+cACoSoFE3fyY
sNanUDONfXTvWvooaNvQCZ+2WxpFM6qzqFWSkQH/M7IJBJXWljRwwLS9mrKx8PcMNMG1kefpEZDX
V5Kj1yiQl1N8qTV6ffelzwNBbzDn4F/jLlTY9XWj1J7cEvUIHgw4IJUg0X6b5a5vAGMYT194GDkv
0WvKV0vbfAPBZGH9VYq7kPUXSKHsH6Bh7fWt74lwXGM71fXJ+FPoaQsMi8yry/hkZZmxnep3PH1F
Y0sCV2agnQszZtP92MrXAb1QHtARKePOCgriQgfnpb8ZsaBeM1bV0wGtcsBV1VIq8ZbVwbP9onoY
ZT8okhVC20TImF5Igg6mlT8KEK8h871GRotGmUpLoTILOzNaHqV6rnkj7UywtjDz6DndupAN3Gqj
rCzMqN1nocxqBNsBD1Rpb21REo7ZJkkFVkO72CRBFWq0/tbh8ALV4lLu8lPaI4u5OsPz/AOJnky4
jD/4T5TAn7fL+mNLfH6mDsfzXcTsC4dukNrqhQ5zGlYbxxymJEdEDxVB/RVfO52sl+7MSa/34QUc
E+l4gXiO5FIaN/1vkfiWAl+FFG1+e+LPru8n19B4G9x2e9vOggeqBfC5nA2Nxo39N3Mia/TZOzqU
2VpXld3dUqGF465rk+5D9qcCh4zWHImPnE4ZFvbCFC6ivL+fzfHDw9sQmAcJ2EHH0u2i1T92FNY5
elx2U7xZToF1OJV0MCgKgWZO2vN3RPA6obgRrMrfOpJAzYYxllVe4JFueXSCu6GC5Q1DXi6cBu0M
oHFjbt629iRRYw0/4jgwBe1JygJMh1QYjJsUNYAXKlXc3ERs5tW3bTIapQgHFXFDMkid05E3DVKU
lm1mYzwt27qgnIkpi/UNr/TmvV6wZJxxGSbiUlv76/L4zp8flQHr4ey+AIWbPAOF17VOgj+vp15x
9OCj73T0fK6Lj3uuBe9Con7MIrU2AmA0W2CraglmIRVNqNjdrgAwDOCbyKHg9Vm/HO33/JEzhvCr
/58Cd242C1lYjQ1sFaCmV49iIn8bHAONmRvejJvK777oZa/7jRYbxYu934PT5MayBCXPHDenvoC3
CTSiftmsTy/97OeKmAY+6hUrNPNLGVqblhtWikwqESR6XxH0Vyiss8ZRIr5NwQZK1jquhGE8Mpy2
RL4nlonge37zFhhm9e+9Od/fFZH7J3V5KIirlU1KDWf4LVBfzJ0iFw79K9NgzzHTyMGq0yAQ428l
i3gVhlpjDovjpnS+eunsSpCI1tEYQ5XwSNJ1Z+MSfi23vr2HILMnGJT8KeGxEnUdeyrDrnY5bDfA
4tx1qZOCIwzNOm4XjkUwOmgogxdKuXJ/FwiL2jBahk2eJ5dez868ZhD7NkiexsK/sMdpNDW8BcJq
b9DJ0yovgP6Yz6NxT6qVZRzUOGz6LwYmK05ctFqpbOtG5hXgKfMh0DmWn7UfxZmwyAxTYuSZN6TN
b7tZ/+JSwUzpC69S8fc5Jqw/XtZ6edwelgs/oGcWBK9quYRi9Nl58a+jvHP0UZqT/uCpxL7m8ZIw
iufL9KKi9KPGLEhKWHIwMz3qbfdno2eaTAOSh/cznNoJG61JjmokspyhfKQsOsM2rggqMOVMQXO3
lMFPp8BlqOAGhSVb2y+sBMpw7QNZKegV9QFt/x5r9c1E+uUn1snf61QhSWYDc5wnrni6z+TQmC1G
pF8QGMC8moQ2H+cBy1leOONsk0lspkNRL2XzXXWVs9NhxzYx7xy3bH/Cmy2t9Zf3iP86kb+EYlaN
kq8j5Fq/qUIsV50lN3rKuspBx4a0o2IA1BhgSLvkFM++D0eylFkbXJGMuv9YYcY3ouYx8ScHAErw
JwHi+vkI0VGoCmO47l4QhvTI57p11AM/k9HpExTn/JaTaBorN4XncogX29KWUQSWYpXW83HA2CVr
s0IiDdmoMYn3FbILkVjDLP4L8x2yd/SX7YP+ulKlR/g5OI6Iy9bESuk9latuKwmYf15I36uMosk4
QDtsblRmGbcaXfievxLhwG/dXwzUpQxrr8u3/Qj4nHcUAQaehuI2WZ4N/NOJ+3VkjDzBqfUclUCW
lotnsewr+QgWHeMLN24r9yehGwnQqNyhmSIalhY+v6clZr2FgTsduqjw1iEG/5ZqALHNHh3o/iBx
SUQgXUcTFW4tMp87P4WaizFbwuI/uwwRG1QiDywimdK2tG2wuvZAyzxbTuWQUGzScmcrBSP9IuZh
sevEYBa7GN5u3w8deR2VvqC9gSm4X2/Tra3+PLIZXAMuUlW8tc4VVWRdRGQ2a/j05k/OwudbxxAW
kBMtlcGJwmroTYIwNZacgwFPo1pt4AFa5FBkd9H9UvvOQhlTW1ajdSiOPx+dO2mHxRkxCmk5LzxX
mMselpfnjQiobdGVzefBCuDhbn11/ezCLBYaUTF4/k0OEItoxTYVHmyyLMYlHXtADrLCMyPOIoWq
pEPYPF3X3zwpqRtoCUR0Mcu0LkpsT5HqY/Y7uIES1QD2CpOt/yHMxh1633r+kyXWj4GDgyouMpfK
WfVdbjHzoIzXiwgdwKUsJAMTxWA5GA7OkVZJQovk/dBIy0tzZII8mHk0RBEdYv2vz7bTeCry54ow
hjyO9r1RIp+KHz5P0pHlTUBf/9820gndhJuVv9uvLd7GMc2LJiVjkAA18bvxT2n86dhRfDfJu0aF
9Aj5/Y6KdmljBJz4Uy/Q2QYCAyL8i41MeJfzthEuNADzSjZ++LKSsKzkoZ7xWysadSXwPAiHhPqr
0HWufp/B9vJiUPANy9067Cc0THeYCpFj/gM/5nXq6DWgIt5xzH+0BaU6o02DRhRWTf1lyy2a8AAa
rj6TzxwoVrQnLZ/RM9MZRUgwSnh+uaGLXtyxYPbV1QM6aE6PKvQlc+XoHUEA3rPj6mLScgd4aAxS
kKBJHPHg47G1qxa2/n6MKejFw1bymRV2VOGEG7SDrPik7xZonwhSX/GFLk1V1l5/KaRXBSf0+sbw
T2/z/m3MyAIqBfm5KkUU61MNdlpB3UiRqrC0ZJWXusYmdXj1A6fm1OWQKeG0+YV1022HPLar8k5H
9dl4OuQujGfMGd8IBF0990I5muODH0hXgq9H6d6prNFjaW8qTFXvSKh0cGXuByPfJY2hYso2XynW
bMa5Xv7PMYSMIrt8BIfvtk7VoLihfwr9NjZT62Jx27qzYCjEVCV/gxd8IP13/eqUZl2/YEjIpof9
xLqQu3AN2CagGj2+6DOEy5qj0FTZyomx8jZDjyLCZ9xXBo+AwCZOkQJAa6XDZrQ8Jdl1/UOoMkk8
2Ab8E2Jx0WHC+DEITF1BQysJKUHg8k4fcOYN0QWVFYpTVJAjyAmWcRn4HLzCOHaMrACLSS+LH77p
NpZfhFNbIx6UbIutgHIC7+4pRcbl3DTOJQgjORJrzIFHkacyKKdZzb4p2P0ZG68iGtxLC8oVVCqQ
EFNlc8StePMTM4hPhWOUeNLZ7m62bxnDBqf3iFbRBWzYPppCzsPerqDYJkPeWkq+56a8jB2H3HKs
i8cHpSWi0gYOeqxPlEceNNMSIMcBsWoEAkygfgJt0ycI5hX0JS0Xpomxby0vDYruD6pEUcQ4Rkmv
8sXE9Mm4D995jOn4qVXRZX+iH75tKveNea1RfXo6GvRm29Jk3aJe8zF2kpxPDSaJCMrt5aXGTmNY
Cc8L9dosVVR6cZfjyYa9fw993Ccag3Zvuqcr/3cpH7+mkVytW8sBVxGwrcQ4olLyZy7u8cIk8Sc7
jc4QYuTBahPC0x3cqXg3DJY/rjuVnRRx86uK1Hm+41DPZiWbAnZqwfFKo1eg+M8C1rOIhKHDqSUM
9OJotS6gJ8TDcNwx4wpO7ajTa9xuYTpMNCejVHfdgCwL+FJ3X4YDrQgIC6h6BUukPZ0FMCF3H6Ue
Ot/On2jDeu4K6jzfGsS/3vy4fUPz1BnflPAJRf2bJC5wA0ovH4ZH53BIhd1KQ31D+OG58QuNXkhs
iJeq606YEY3t96S+oC27RjtaE6Sm1O4U6avEEZtvMXZkNUPgCClyLs+bEQAF9R62GDrFoM8HFhb1
aVn9BUQy5FvvbXG1k/nal9DrZzBww+94LbcXnVRtEy1YaLBIvfcwGH3YAik3x0jxHgZvAqKuctaw
JBmFzEYhy7XDxDFvL99ibcF+HujRVGBbKQ47+311S7NF8FBmoVmZFPbcRBlYQpSteBBx46YaLLLt
Q6ayNGRGBeZ77E/cvFWlWx7jCw4IAYZSUTywE8zpj9QFiv3K5P4X1HNdEzPpDad3Zj3ujQLICaA0
7sP7j2k2V+RQh1C6qGj0LBVwRoXjoYotpc0710vg1kgNWa3nvPkfAhj6vWwcj8z9tFc+NOe2QIvX
eGlraYB/IIqNvdoIUaSzKgfeZ5agXrWzDxgWzLdaKrh+fJISibtzcjaSiws7CVq89OLJHpR92z69
GTQsYX2JnZ+70bAD7xeSxGtuye4WT43wpg10vQyuarla+DAkDtRcq3KmCEXO/S0XvABSHZ5uzLFr
WA7vn/mGCR2vZrOy+8vpgmVFLdHNwgW9ikZergIUKgfCewRNlxH13/wUHvQcRyfBTSU97ZiQcP3J
Eol7dpGOoehK/0UU5LL+ROtzgEm08pC/58auEIR343sMF5oFFB0SvygHM1MNGbHgoPMPTHcuOisL
ssRCTNm1Bc1IJ4BphEe+0uAYTQCKlvU3tRH6Iw87Gcabe8JLP08cva83ZcrNnOsr2dAp830VJvMz
VxTXVN/Y5kkHruDeMRrZnJS7T5AUHjnSM6uMwMFgqccUksnY+K9FUFIWhab8BIN3aiLS7uQg3YQy
QDHSmr8RA5RifPd+DTn6M6g8kmTNPAV6GaAk/5XoP0fRzCr5Cp6M9VEBreDzEEjrL1jYQmQ1Ueg6
ViD+dnNYCHXXeNICQSN0TtAZ9sVtwESoZbuYiDz5Ip9wCl5A5rQYpcdiIUWvb/7bgnxI/6/YVHHT
XZyArk2d3oxJVo4JRrjYKlpUMCfsWp6MOIuyE3KHmK0JHtPgC+8G5t8/RoX88kGuN1XxGb+Dwnea
7HMxssCLJVQwT7rWGafuySkhTC0g93Svzx0wz/Dl5ZL91CK+TqMdxgJRzYSxYwWWPxrqMMbCpjMz
K3fSKGpAJzvC9QAMOlGBSTFan+zBYxxF4eSBdf6tm/87fSZyFbhDrjERI0ZCuHPJ2krcpEeGtDs5
Fje7/O23g43pHmkL3OO7oCMuEFRi3TbHvIhW8X6eOA9YHJGJNyy9ewAjb2NW91Nd1csvGejbRZi3
6AinwqjXaJiuvEuJKnlp/AhhuSLAZt9S2OniFo/ujctqEK5xFptEZUu8qCNd9kvw5OORaHgiitTO
hUeWpuQLhqq0U8EDWVrIudmROu/PS47iuPlTWLARWJ+FFmiob7YGNvHvT0y/XjNNh4T1HF7fhzWs
YaO4+GhtZLwGTlYqOPynmKaNnmlDJHDyQEnQmjgfiklVcI+/uGL257A1381F9N58NDAsuA/TILA2
M71wCrtYgenPmh0rFofRpHcXWzPhRHqOnkYVnAEDnraqw4jg2paj07O2C3KZzb2YSIR+ZGKLcpsv
QbcFhxUtcBA8ViLrgXgtpjbS5t3Kmx1q9L/u1XehmFrwkjor9gQM/034OTJOqDnl6nCDdCCCLCB+
GZt3VQCfm6cnnrdYv+S/bkAM5c9m2gRjJlM1d8SEchdjpbO46VnGf3bqTh3rBAY5ldnHkoeRFsvf
S1aFAmfAVlIwRFSDxEahuQa3/2t99+gm821aAeWyyNU3YAHackGYmeJNr8CUZeyHVfrJGsh1oTBn
Abnj7gv1B0JZP1gbhwri+gQRHKVs+9JAAbKjw52F1S/1SwUEpEFffgkgWk7h096iQP9GtImtHBS+
JjIpoeR9djaHbOpb5KBtYpCmchSbrbqXFs8oNvdpAfTr8lCrf8pLO0EjIuxtnf2JtvQ4g40O0KgO
lzX/oVYip/tA8hrOpb3lYjx4Pe2wyrVnSpZVpKir/XUcCQbn3hrAm8kEuhZHBUi9kWZ6Bkskr7UD
VYaM41v17HMaeAOZ6MyTsHoQqTX7xM5iQkAmlw1H3BJQOvB3hplIRE96zPtz6MV6IesRH1C/2zbN
tZ8Q1ViLrl4SjeIG2CQIrAPd9x4eV2BhpnuosOT2kHLzzWfikw5iwU7BN4bwh6slG/IRE73Xpy4n
4uAKQBtv3cilSUj7H02p+BDZ63qr9qBEq/i7HTx4OwbGNc3Cnvp9FA5ph0QFCMrqUnzQhGQowBWC
GOemUNh95rItToqILAFcvY56PatTLPKnkguDlnG0E8HkuOBOAXESjiARNJoak+q2cQrstCT0CkxI
VyEfNZ0iI5bOmeBq/Bh8bRinc8hRriACCielPLdf5m73dhCfCgiljt6msJObVbXd1zvTyKMmamVj
P8cWifYhA1Iw+oaRmXrifz4qn7X/ejcxoisWI6Z8CjCOX20hJMPJR8rQwCdKW5D7lldtQrmsm1Lq
O3NjXl9M5sCWcAOz+TYLCMp2WQus/Rkfot0CTsMpYboA7uR6F5mzJryv5CHJ2bHcq3TyWP4X9OCf
Gphvi6v9MW4T7uHzdXKM9pPwFRFkb/L7N3sc+aS8fJvxA0Gc6eQggCa8mjxJx9OuuzolYKkBQIRm
+aTiuUfHWkYdFAysU0QFP1pNw3x54csWYamJhoF189e/5owu7YBtvZz0Bk66HwpVPXfyje64Br+u
hHFawTz2tuqsI28sigo8Lz00YCWqUargj+Ds1yT+Vk8VnHhF99Bib+plxu9kEmx6/sxqPlMhvbne
7zhA+NOGYgZ+h7T2NeWxUzCtVtR8WjgTjuAcoahIEjXvJqdijheaToC3y/Psncmo8bboqJhQH9Y/
22jnoulK3gC1Z1mprBUZu18syCj5DMLDT0ZAUMAP/kcXWy12DtJfPOLdE2kQrjjo8iZwAknCIvk6
Z7hZ1w0Nj3VgObCbn8SWHjcPWyFx9X/DG3XRZzy/s3rh09fU01BjuxrxSYHoyLLTija4QfFEL9Jz
y22Ts+107x9iV8DHY+eYowSDpSqV5nhkPdrjIzadmpETH+vsiHLavzFkCs/5IdD7x0hQkaWPbCrt
7K6SSd6M+CmupyL0yxZlsssJoia8bN793nvFuZG9b0x3BxgHF/GksLX1OCe49ZNn0paHWDDhZOIf
5K+bly1FJPcf7BJV3N4aRNnFe8OeX1Cgd0SwuPjLJ+PsJfdI/vglAyLNdNpJTSXh5IgwA+gOy8Ge
NNEsnTtFTtbIIeIAUE88KhPGl/y2FyCa8fk57ET7djXLf2IyzAkz8DQNZsFYY3QFHrzY6RJNKR0K
NTdVuahj4dj0lkX1k7rkUqjyvGh9ROlyF/xkC8kC/LJHjmVLbMj8zRGeqf0+V48xJAj+uCSvYeLe
j/qM9AWQGtTxBH8AfGQLgMU0DfovCGZG5iqoECOP+lchcpjkuQFZ9qyzqZaxW6gAmKXpPgulOUWh
+/nXtqiGlWiL39XMBvpvMjbIVXIaG9ERsuW3j7QQKSrRq85arLTR5Jd1pC1gh2sZDYGttn6TEnWl
VVJIg0Cfnt8TGQ+TPuZPONp/03YZx+lzo80HxIKTZT+yok2a9yORAZ6UW/GKVVQypggW9UX7PIEC
3JxffV4sCpQ1WgblALAzLan/x6wqbe3aWV6wwuz0TnZ7Y/ACP/lvyjUdFnV4NLGaLsDqm9pTqr9W
90z3kjHmDauBz4N0k8RHC7gVRQGN0SIz7DmtIbNrAiBn+QAUoJpITmxSAI7+UZCD/6E5GbD7bIIv
MwRqL3tgqpPkVmLR6/HxGvz4nX76k7yFXqB8ZS37d2Wb1RoDbLZ1THMF/gwRMn2eaWJX4kv2ClCo
t9l1SkVEAF6THniDEchiwTqB8c4LToPNQtX1pEj1l2hpXETfvNwqv/MhS/wpNpkSHGQWvJsN8mJ6
CGFz7QdoAm0XiCbH+iOHhegdYIw5GMws+X0nIgQuQnE1PwNeDhXPX22B6ERqND0HJsj2DY6z7YY6
GEgcmNa/RF4lnjeyTZv/YyUSnAxLMO/QC/A8Ra57DFxrACg9135J3zPtSVJuCKfp1JrhrJzPm7sz
bfqC/nFHOx1cCtnh/unwBO5ypIuWriSusMjWisBZ6N5k2lQ+Hk93KT78dKGme1d1IrmzqmIS3O37
OsCz5JrzkRf6UnT6onq0YwdT4/A8t6FmBerBjkidQXhWDPnDy3X1p7G75YoLV09LzTdgEorokJ5b
u/TQ8Y95IxJ+16/qGFJZPszyxD72z8J4/Qscoq0mLk7xYSEQ16JibFLF/m8oAjsteIdQdmgtMvlX
2xIBvaAk1wW6erYaEqu9HLQhFfmBxUpqifw27arKt1FbNZlAZZMxPSNGEFgnqb+dB/hWE7ECrZKP
JRhJqsiayOfOkjUdp2aL65dL4nW6zPkbKFcWVy3QYAJGx6eRA8KpRu1dIwcB35G3Pis7X9gf/VOs
CzXPmAgr72LgYtgAkvRnuY+vCbv82KItocNFZz0Un5N2o5o61YJfW5Rlz5aL8yc2qPGQtAggec7H
OGOyspM5CQWdVh2wErPUAUSJQDzpHsqXud3krVwV0DUkhu+6yu+MXVCuCEmj0Fnn/9h7kAkYQFHs
qJE7LzFjWgifJk8lW0tiCVMXC96PebeulbPhhyfsmdmUz885y7TsmXhdAWXCbhCvZ3fnVYSlMMgb
1gdX0hwPLS1YTErloV1waPnN8irIJc8ueSxF4Zz5xqEcoAgzQdM9ZOrSiZkMeRTthY1Y7BToAFq5
fgy//RfAzcEDeoqfgVnxEwIlbTHdNC/QvgC14WMl76uFfNasa9/3MjuHFwlQLQ4jg0lv3lddB8Uu
uQmKy/mob07JHEA7aXqSf8vsGEfBGaY3YgGJg14NpRijNyfFlAVFQ0kJCUyN0+/u+JVw9GHHw80k
SwoCTnntTV8/4gF8zxsWx3pejcZYtHRGIq8TnnZw2+ArE54g/EhX4rNHgp850XzSCA/0WOr6AC9d
R92hg81GIxKpb3tWuoOIKyHJOXtYT6HgumCKRFPiu9TjrW/hQtntXtNJTKhXBheH/bjFqmyMGwUw
Xr6LpzHlCYtmgAD1ctLBVQXgTRPLeAsdNOjOi4nJ1S+T7JG+UTFEGRaqBEjMHMRrQxwxyG/RSJh1
nSY/J1W/wz8H4SCZXN13OOU7e/e7jd9umbTGBgpZv4IsrgTO4FXnziUg5SH7azeYU/oB+dWTOwg8
Es07SIhHbuk/BRpbYN8WfQsy8J9P/JOMaIlobAfY5h2mJ9uL0MTMbe97NYey5QB8HkY7v0UI8dVL
N8mtM3k7BfyJCiVZ/1Zi86JEZVMkMoJK2oeh9VGdb24BCbFSN3qX/8KtqeobyQ0Ep9DKnsiATMMv
1FHXQoF+iLzOlZjQHpB0lXeQHa4tcxHq7rdnywz9ZZdGNzFi/FIM85SG5FqMab9AF6V7155w85cI
9MhFAloEPTYUSF8HxA/hiBCZlKWnokudATGEcaPaaNHYaU3hdP+cOl+A3k8gaOMbhVxfvwAEx2cJ
QRfmm2tXCpIAvVAGZoDw562kbbZsOMnEdeKgrkztS643qqvLTPYrmWWUekWzevSywGnFyHgn5A7g
e60e1ViridRxJd7zCw7BqsqHdIxeOHQPTEMGI20qJ/FzM1IcZOxreTL+O1cFoeYVuwcYT5EaG729
RWnjz88wqDQMRmd7cIOWyN1j2mOzqxFmKCN5X5UKuHVYvo7vl/0N8vy6prqi2DczEq+W8QFuTY3w
Q9hNhuQdkL6PKTdt+fkl+iW7BaoBA1UdyY53+eMBMFeVUZ7y9f0rOVmzMCzOzxj2uE7chNZGtqUw
OjFVCWVdY7yokAkp8arCd4FjR/PyHlhG+ZsXKXzm8vyiGkQnbED9SPB/hNu7RcYCOSXPrY90XCIF
E3aKYwTt8/C/EoUQyxn/bCbaMDx+XRY8TdlClZIjMEdSUpvOHcHFVdFXZLMqYMKfqcqbrxaQcHtI
FaK2KyP0bLrJnGJ8w4WLR2vzFCirA/BJtcH81DRwemycjk24rvECEaVCpOcsa59wkXi0KK3OP+Yn
bftKFIcCm9Tja7hZ+2TX7uHvdCYiijWyXYqwH41zV7PueyuTeTuDzvIWsvSl2w4mAtccj9vEY44K
SQnNIQBCU3UsXIGzUZGZIQaetGXlPn2Gj+lpjFXFJT3wYv++kdcLPVAEi6ZLN5lnRM+rj+7sCgY3
Nr1ncssFslWpN4sCkFWrupuP8VyBbwHUHCv3XJA/60lD0lXChRSIaKY6TiMtnWPtSXqMn0zp6P0o
GCn1H30Mo3Wc96BydV8zZlcQ/L5cZbwwDOHHDn1reixXcJG2u284jSJPmH7jZDDdvKDUixcGhAy+
YHssFx0M2gQnmwPuj/K1w5e/1nqf5oxTZN31aKYKVa2H94TEY5zygQ+iahb5m8oFru8dz8rjAt+Y
z/qV/SpISctJ0TpqFkeieGRqPlrBpMqWFjbnF8V4By/EiaklZfB8cLT/FhPevO72jOJEAmcp8R37
c/Leo8U9/DBZrkT5Sb3TnZrsbtGireC+sdvQWsT2LMnVEgWj1JqMKeyo88mr272rx49CVhzumWPG
/pjWuwwBxPDs8797wsE51Qqa2jH85Dweyjllkr/V0uwPI8UOA3lct39JqAFX95+aX6A2rFogHXLV
6bK4NBNGzHMv14goraz/K4sPxodojcSWVbVn/UNrAqguAI+0tqiEH8X8VnSWKL48uYt+grCNDr6j
EU6EzTla5/dX5gB3S6RRSuues1+S5MZOA5QAG1XZxm9gD079+kykHCLBj3SZq0v8EtPs0qcsoKeo
GVm2lTPF+CA1ENMeqPBMY3ROLczvIIZEwnTaIQ5YMVOl+LFUuSfzpUsJSTKbU7JQpksOl6V4Ol9g
B0z9sYGrxMjTdfaxZyzEg6SQnxVdTVGZdPCStDK3jhk2efhCmYpKoxKf1jy8TO9+8/9wRoybTwWZ
yeT4Q2h1o3UzNEnizw5S9R8wiusxnwjEhViu8ayHkPsBtL6gAw4belxmJdneuGI1QPCHob8JyKad
MTNGQaxDn69I+IyLBFhXDbspFTnsB6/q2rXDwtq/uCVqiqeYKmC4U47ZifJH2w9BdVNlgSBC1rCc
ZQ2VmWdakiJCDEgxOegt1rFu1eIsb8ZUjpxoQi10pTUDSePgx2NH0BHxYmoR+O/zJhw//n7bl+Sx
h/3AWylZaj9vWz6NLYlsZMjYdSEGZyAJ4pke2G9vLlevytlNAQWd7KtLhCUNsA5JDS+gKWXrslOx
EQ62wnolbjEs1d4JgpNDL4S/u90poJONo3rYAb3S4jn1k+C506wPxPLQsnPSaS9zn9a2thpiK87c
m9KSCTmUOCtlZ+PGYNMyl+y0eQiOaCuQgpFuNEW6Ddno9GGqVcbKLY8lonqMezYnvtWRKP9Z285r
pP/hk8XTQKnMsRI+b3aqx5efJhaOX7pWuTveg331dmJLfFtwHDbb1jgQKSPs/z8W0vl8KUd/EipE
DY2+KMHkJK+03SekAez908OPlSe6ou5C41DZ97S80H/vSehTXZUEawYQNof0PmX3Jm9N/Ttr943w
tI+2A0QsaTTWgg2PREfdRShDO/ztD5Bp6CcdF8vPJG4NsScYnHCDII2W53PDRBJLwcLD2L2qhC1x
YusvG0/PgeGZKANnC+LyLgn+lHSUgrmemD8lXc/hfbmPzrWh5/9hWKAR4ee3hkunH6O/fNLi66Ru
47yWd1EdMZB9i5YuMWQDCPRhrf89nDc6bupmMOS8u9/gV2ebH7crzSdQ6LxPOCKmRh/XCasK5Qaz
AtgedOmrbCBkfJcXcMctVgtmHhjsiLFDqOgQmNk8rXjjlI5kjQvsW/bGRGSFqEAb+iAN8Cgz2TsI
EsrYYUmnUI02+rITIE4pOLdwOsGgiOEJRwG36mTqabwYfrHfj+L+v/hooh9350D5Ajfj/1+CfhCD
aaJqR5Dx27+vcA/bsL2XrGZvlOUpGV/fN2abB13+z5FvC5hXglasYa6aEvM5gQVFlKpxkSFIPLS5
CW9eqIeSe7q6lpl2zYjPMZulbceVup/2u30+MVf/T5uSkWTFZmoHx3EsyN42yljP901NCYEm0sCB
mDPpOLYkN4d6a/CiZMzwUyp+XbHUnqVrQcFd/eR318Mr2kVn+W0eCDuz2REpsGBT+fZRfTGnChMV
B8NrgrEY5EaSCcEwgnnokKoRQaOaKGJ5+W7Q4fHU73iSuzdQ7XGbmpgItn2WMtwzqkL0xGAAYegS
xrERavoVR+nXvBd7xpofx3BBt68lvxQ6IpIDZT6+iBfIC+P96rU8OPx2a5ZZ70KsuLixvxhQcZmw
0yqdZg4rB4XMf/ywd0nwwL2Didj9BlJ+4tcCzw7n5w6W1JE2hwuJEuvo8HBJrrAjPqE9BMUZDX8F
DeWZsXMJ/ZP2D9QfppzDLqWEcj5J+2A1KXnRtZ9uluE/hlc2gLtrcpiDzM7X3M5/PFk5SiL/6+Fl
fOO5INVgWc1L2Yhkke8k0nGl1xA6u0tRVScGn4iLyiPRjgLW8qLYxwzGmk+hGg2nbmEfA5ocMLjw
e/DXJ/inPm0O1CM43jBRW0IIw2u7M2ZcvUWOp3fV34qOSHD73HWQqGlS3wNQvzYfKJh7zHYGk2G5
b/kLCz0pK8S7USS2kE+Q67rxNiNpf2WNGEKfgqPuY7cVGM8GHz51HfRuc6fkThzXTZXqY+5JIHHQ
94hU0+piy1MW0xyD1Y10GE9mWDqn1cU/ijEpGTy2rgRvF3MBRnxkxGIuHF7vEWvHsHtkoellUfUD
ozlrMoWxb+i3nK8UOYdAEcNAT9tQq4TF+/9F71IZLh74KxhhhK6qlsqHLAVADSQhvkAA7WdCcpGD
Fq8Xc1BT1f6ANy3c26pboMf6Gb1ylBih9/43BAkxhB+UiaJs5F+1bzqtkeOyDSJY6LmJrJG9YOOL
jzwNzXFw2X4mENKrtR5vrwgsRULDvjdpMwfiTAI0VLtVQZ7Z5ToAeCarQnPmkDJhpnYB1vzFMF1z
a6zDxTwTJ4C7Rze9F2piJwhOiHxW8K4IGwGeONfwY4Vg65OoZjFNmwnv7qSoKOHM5qe5urXoTLJD
PQssNb1XZxlZ1e5Qw+7PRubEIwqT8Wvm89VdfeD0Ovh0OK3yIaHzPqb2qtMyDsstkT9eQYemAMix
uXMSXJ/IFxhD1hCNn1QnNYmIoJ+qW498pWP6Ji9gG/L+OJ2anNDqZhjEZA5+/L86BYOoJKZuVBPR
++hDhPgBSLyn6h690oi0h3cGAi511QWLKbE6EAagzE6uBTXekRTMDZ2GbIkMIuC7vOiV38xoVoud
vk5jJwZCptK5rt2mBT2K2FjPb3mqcensRrYwjtjd3pe1hnA+0ng0+l8sRgIox+SgYqJOxB51Z6Rc
pwx9t/OP74cTgk8ZyZXrVSIvWO3pYE2Y2oVUAP00DWdGieNXaolAVuiMH+I07QTklayAyK+hc5eG
C4cTjxoIFSonBkgsuwX61uGm+Xz0EhcsTPDJSoo69Xi+ncIyhPxfKwsqtdJLJ5Aih5X/GNwGLtIU
ZtMjA8oGDaiA4CmyvVsWN7Dy33gMFA1w8Tz3DoutPrVAejgP9LAYdFYnSv9Ih7iO7F1Ahs//d3L1
DT/H5aQ1BWhiCMG2KEnfWgpv9RcPYNu02NrKOdzb0Tuw7Ourvx8iQ5Eyp2vmfdkquHlh7cz94L4i
fWLSEOl9smD5p2AsNxZBcvj+iS+GPfYlT6/J5i7gZKsZ0scrTlM/DK9QTxpR2WGdNNMjmLr+BFCF
ktMN5YKl/kI9sZIt6/3olaGTpRy4okSBnwaNi7FjA8VSU37TpZ6+9cV7M39Umg47TWGy5fw+f/IB
05t6TdHUGJ5sInnQWXtjrWuBqthQfKNXhv0NLTSoxPVpcpNlAxxCTeUG7OOg66nyZKLUApOAsNAX
X+up0TcevHLgEDuyqXbhEX9TAiDt0oZoTLplNIktSXLNEBDKYTyc+40o/2TtNC6Bs6gpAoGmBW4+
Vt64acPsBOiv+41EWZezxVc8KECvuzNZcLkN4nJjXdzpSICpSn+mY3fzoPFtaKDDWL9nFtXMi4L4
jfF7VQRbHytyJAEDEUHR5t4bQ/1JORp8e7V8005JY/Huf8BqFvGAepzwatOJWkhgPTN/jRv+FZ9j
QTZZ8i3TffCnEAVnIv1ElyLXrkTySGPvAMWUi55VxAdwgK4qkIENUxmJRBeeo+sRVagbsp5hFoGb
BKqqhxivU9yB6MilwFzEupk79711ZyD/nx4L18vTZXegvb2n2c/v9/JQELGTEemV9eyWMhKMfZdU
IqRAPaNsDi6um7A4OTnbyPSdl5X7x7ML7ewwzQrsTol2rSxA2cV6TpUUt0PMdUBLZTglQ6Gluw+3
UY6N/JzdnASjZbkV/OtiIvkwTd/GgNYZ6/N8ZYA7USzGBfqJ9S25HmYrazMngXnD6sRuosxTTujd
CqrWy1cM/9X+48d8OG/LIMqh1WPgv/4vymIFRkzwIlkV0WuA83NgFHR7Ewbwsd6c3Nt5py9qRTQq
9yPsm/etNE8ZJyn8J8R04wKEWU4SHtqryU3HzVMDD3+ahdK6sf5yYh7ARfdDgqqIjVxa1oz9O7ii
ZnNI/QoTmxskqO1+J/ytsgUGV5PZtjS3wbl51SfQ644CboemKbnOsMvfRlTokUcbXsQkEISFKtKV
sGEgEqW+PvRMlzjsaeIJosypA5FrMeTn1LXoTHjAl4wUQcZ/tkUe2eb22wDrKjRXmtqfnwoACMh6
pJGVk2iHT96aYxVrTrUFRj7lQvhKa9Lp3xxx/tywak7hkZi7XbCk5Lg9xbnwobStAunziXh4EBmT
ePj8GFhtuX/MhtntYTIvOp1guVcfNXcV7p/4iaxLSb8t+6/85M2QYJ5dAtLqkfhNuA3Kg6CaDstJ
LIb1wunRvaR/HAmzLGu9xb5b+34bTZEa7lI8wsDLJqdS+EaPDRMNmTHKRwlGArMTcNcz/HCFMct8
oKMtm8ZIce7k8o5jySOzNfuJhfl42dqnPAQHHNwwloHFcIKUUkNBNCrypucSH3mcDOWCPWvvnLRx
o5aQ70LJ+LbJJxJQT5bT6vZNaQIvuVChvAoyHgbUwAligaa4yuAH7627M7bgT4IhW6QlLq0NKu7o
mE6WbukTBF1WoktAtGmwdBH3DzJyGssAulmnUXIn339N8Zih6RSbZ1sglbVX03+lBJAysPrOzCgb
+Hljujli0xOL1KsJkxgVJiRGvOIvzGsa4ipwqMOYVLosn+SxziWVFbQ2ALKmY0D8DDp+5y7IgpPi
9F7PPRQ+niQp2acCBVbrETy6gVHdEFtc8uh5sgE8IjydX7BRbIM60iaSY5p9gwFS5oLc+Bwc6ozD
AQlFu4DTpf1YkIEtS6SaNNC14dPN6VMXP1cprbN1v78kMmx/0qA5eOVXtJrcv2mqK9/K1gZbzZvo
F0YK2lvZY9qFKlj3PuTyRTLLk7H83LSKlz/7STDrwibp1+rW0SsOxJ21LB4NaR+sQcyKeauSb0Ik
uCR/AEbiMVNTBLXyIiGqQ8VOQDkBypFIpdIiG4e+PyV8D363Rp/tN0g4iLA71jflyE9iKG+ReO+Z
GgBQlbltZjikr4wYGCLcfwBbTQ36llpVsN5yf8QKgyePKRpVrhYCMPWH+Tbh7CChw1b5Utx0RsMw
J7mW1Dxd/UYAMwQpMtdsj1v9cx8w3YJt8VKm1mZiMk7X2TMHXCD+Xj5Ca2uOAfx+5WEPV/LVeT+n
4VkLO8QbNjdfhUKlMUXjzsVmYM5f2HFA9hOF3pylNgkyQjrHxpxRDhD8hMNoaCS6GgSwLmeFNRC1
X13mBSbfVXC6P+JZ6iF21gL4FJv7L9ZliHzf5gR/w5KB6D2CfarUtCKKMpPvq+krnyOAN1zSuabc
/fkDG6fzRti/5aRRiEbnxcvC2Vqm8NkOkpjNFBUJYTH+lxwadsA+smfPwahfhZE1VlEfTXfV+2gh
6A933pOWrgDRPdZf5dUiggYXAzPtOO4RwlCcDJllkwykj5gqJEGZmCrVEcUf4fBm+LhDwLgeIz59
2M8kDO+skvOibYSO7Sw2+FkIlyxk6hObVDPyuC9U5MMPuyBC5RZlG78eiPgOS/yiU+lAO5NSHMtI
2nqMwU7wsAl1663LckLBWt6M7OIXrjcpWDqo3aY2bd3Vhc3dsOYn5RpB/YE6Un4a0tX54ZKTcrRL
4H9tTGvGAXdKJ0wlF+z1die18MQx5mFLHFQXA0vEwUCFItlXg3A5+CaWXDrGHRIrUqyBS87II4xF
Evw/fdeoRJTYcO9Z6Tvaac1LEkInGW1RTC5ANe5NU0lvGZW7bMjB4WsfF5LRESJHFsSqmYBqPPIL
FPFEheeRXM7YrzhrcES0OmlngY9zAlyg+0PqKSNBmv0FCrF3M8UDW0qMZD+veAyrHnhhCtkT3ECv
+OOetP/crA32zbBcMCRL2sndSY8tTmslUhAJ2lr700IICQenbqP8ahuUCL1EiuPluvA1kauHhWTp
4Yqarw4BiuOj1npo+CJvqUo5Yz0HvSedX1t1mNQqToYTN1AgdclGPfUeD/GmkUZLO0nHveJ6EcIh
EhYTFdXfhDL7Vlo1OmDqgiKEu8SYpMJcZ94gtzAXhN1hp5dAKhHJhEuEIvYu9kPeAdKKlE55OZnF
4J59VWNgldqsuXnLdDNNvgOeRY9tVTYjnBwR+VR1/py8Mn9cVy3lU9OC6TRKpiZskTgmq1DTOMZg
fl4Nh4uUFpz9MLNVlms8CNNWPRRwFJo07Ogytg7P5RjjlRpGCPJeaprPnt1g1dpZW89xerBr9aoR
P+lSztKld6eZruZZEu5mjY6nsFozuoutXel4VoKCrjBLdi3KdEQaupoGR9n5Fje/+Xf3kXoPetUE
EP4yOvxDf+TEDhZylkvL4ZlOgG+d4ulQkvLsPZAxNb/GXejaVENgrVxIzwE7sjicm6jcLkY5/mxf
i3E8KuXRoJA9mAe4idsFQin4Y7B9NkNni+T106R6JA0HN3Cmuei4uwcS7hHBNn8m90TVinfOb0Rt
RFFAQA4324lmvvgPXPBYfUC99WOBVKgD3kBWhgdQdh2RetHfSf+toJL3nmO1X4b2YmEE2jw/SfE9
TSDrobE0O12lXDuYrNmImpHi1YaK2fHOdANz7gqSDD1EnMNp/etiM9L82sDR/lcOXBgZUwTHz6yn
NSG7XZ8UY4yklqi4zL6WT8gL91WxcUT8OTNdNID5TyGmk/X3SBHpQkCzilgn4dyx0NiU0lU8Tgbs
LqKvcOO82NqwTXFTUWwQUgkyzW/QYYJCDejd8H/ZD82BaeE6PBF8RKxawmok3XkNG0bJpx854dmn
n6zZqRe3NTJm3cU65Kz450C8j1nIsWrMVOADorJ7Wso/8EwP1KRdxxkzxyUD3YJfefzBckIVvw1z
hCn6dvcGw+zNSCfawZB3FpxcHfF5Oec8FL88oygE2Cjc+jGq67zzx0G3xKG4nkvP2F+tWqU/c4NQ
wRJgbvbfFtXGvVKWqF9fh1HfYkKPgIP4CmhRjppOhJYTMW+upcW9NkmC7jB1VjlLQcjBqh9tFZg1
4f/lvjRBrAzljQPr4PMNh96jzuomW7rzhDVcgGibIwhFCKhqbh6I9HKnhZNfSZW7UFK1nhwKneeQ
H25Db4UZwnTVDq8GE2DL6NR0tfI1Qf1Qx5ikkaDFM4/u2bTdufu5JI1PaHNgF0kyGK9Q3SawUmrh
KIVphV71jxephwS7ewJNyB7vECRFwjyovFUUEnN7s/jholzxsxtSKKAl+wsGYy0yyBmBbgkaBtrw
50vi74kMdnN5agqRxyBto5nVpHmowxUEU/AX7C2hRMgkHPplu49m5YKp9D5N6sJyKJqRTSlCB4VP
8yr0zmbx8O+GpvikePM6hgWFvClGdMYVTcbfL9CxemThK0ZAtuc3V+66J4koU1rzAaBy/8nIzVmp
Jv5/KCSBgXoIsOX1bqhiuFzNCj2YaFT31CSWKsHM3Ia1avQmX8vp95yoJQyUnXTvjyf0TlDo+KYT
DTEkFUoDzYKytvJx+FiZn6qFHI/kKmZbTWZ7wZuZF1XRmM5lb0smldn11Z9uk9e3R0kHRRb0i6UC
pzZdEzE+63bUSoJZc7I5rX3hwdsQ+DnUwRDFANczF0Q+GlvQ4nXr77My2gRe45Sf81hkwFkm3FYY
6q3ow9c441fqzQVZuCwtwk86g19EFnkl357RjQCdkcornIaVnsCdDouJW/85c8Q0Zx73F3CLVGVH
7cn/mp5XNy0qYVHzyi4fBf5/aulikAI2VkGALDPh9BGnwGYNsBG8oCKklDu1O7PmK8N43Uq/fJFL
LMDgrQOfJCsb2RJryZzyw8ybY9fB4jkbHYYRkHL0obiNtPJAcXmKOpWnY7BYeOCYufOCK02+M0Kh
Edn3Rb/TyfVrAs4xEztlXt7SNX7bO6zjIrEHwyUdE131hRLZnCrQHcaiJjaiokRE7q0wtipP6s0s
eJODP2qtm7SVF1A/5R0ltJEIVdeMABNNUTRGQm3DwoLMvJpnVRouLoURkVKkeyPjjXOxxs4FO7p/
iJz5SCHGyGTI9T608/pi+ZSUyd5RQjsGqk5TbRwvC1oSVcTqujuwDPuxIqjPShmEEjNtOeL/wekU
sU5Y/8a7SrbEfsa8o9IHELe7SQUnY88Az1Sag12vkV4m8n95dv+6+Y8bRX/5mIKwfBMrF8Cvpo4X
xQyW57A29j7gOI5+EA7kaRara0kSJs5B8xf+sPyg2JyYUZ8v/JVlOGBsc9taRbXHehaAcy0m/sCP
rsx48r0jzvJuuEdtDD8X1tfoaoKwfzyYYd534faisA3/UG9N14oIlpUmXLlXoykVMlaHR7sDj7db
YeTah1/9mqBH8B1LqEINWExXrl0E3m7civ7qQoB6Zv7uYJWbEyr/XeOxUKkjUiOPnPR4N2zYKTCV
OZ/YmW1Ao+1lrN2anfRUDPtQeUIizl26xNla0Yy50liBDa2eT9D+klxKLO35iU1yihCFT4iF3UI6
k57J9HS0k3P1cM+xIGXYzIKe6KV0UJP9l3So3fGnNKtKldFwLpryrfHJZkxSTbEY9vwPQN0AiIT8
/eWU96wmPbsJ5mZYKkF6u5acBlxqWBVu57N4+67Q8eyU8VFYy2cHSt7rE4kBZvOgwWY8G1tjUnU7
QK9MNL7Z8SYv4LUq6xfndTdyiUozpoPxkHdXa9WVr0zgPXXlEWN9q0mnPSsqDTr9pi3Z0PxaQhGT
+MLqf2NN5G+odrIKyROORIdC7nrvGgqu7jCDUI+dNb+Dwg9fvn35q4Ov8mt8j94nTjKTKZLZEdBO
rXckt5oBuY4TyKrTZkoYmWzhlWSY4gbUXNwGcmSbMqDyG+aVlyDZMsjd/XxqFg4qwAhmiCYAXTvp
IECR6AnkHuLmQl7NG2swTJA6TdZ2xnb7pSHxa4QlgTacHUtLeykGfZ52OIueE1sZWcUMucMyU5lB
p0KpTTyn9oLrbKrT/BUZEVZwcdM98nPlX+9NtHc+wlW+q6hlVxI9cfNENBm9uKWI+Ue/Lp69hF8s
2YHmoqpapNG4wd5AVWr4j1DbC01iWokJT8OfWB900DQJbdkJb00gOGLPaXv9k8yNCQqJUvLfga48
xX3Su/qdH/365wRQ37vi50kZJxNCT8TuYdewFkDmUO50sR2e0FixRfP8L/q330qm5dFQz3Lr/oU1
1Y7J+i1Gxq2jv15wupkKYWaHYrcd9nujDoThR6Zw1S1fim2S4Gwb5tfXHO3fulGcJveUe67ky0HI
xQfP+Yzo3EZpE6erQfExv7zc1WNSpyou53d8fuRpuhLUfgA6+WwTt4C33e8YHY0hVC+vDSXu3tbM
39R8UAFFXeplMqJl5FcSB5iSGMda3szfyjfp0mR8h0CzqVvUb2DfDnVMqaaWu+XmEugbY+E2wV1z
1oy6x/6L/AGL/idRJvRAIj9MG6jX3i91bGK1FzYWqwu21MVkAyT7qM13oTBXg/SNoDic9Y8XCr2K
7L0lHsPOxMm50jvuRuaVy09IcU0ghcCJPypfFeehU/7wyyNz1BRv22xrESPwFjg0ffh0BuPOLVIw
fzEOO+qrhUYKaQJU0SXF+4sRgtw1JDsA/0p+YUbr1OWWk4pZl0Xolr6sW9x026OzpIU/1Z2pAY99
DG36OHGg9vx4KSXwgr28enwkGMSoSc58bHaBDZ1iXNG4VH57fBB3dcFaAVpjtW9Pja/7EbIPGVJ/
UmxKbHTGPjXfFLoqE7jf3my36FgA7cggSSinSsL1RGCWjxI+5UD8D1VZyYE2ynM7N8emUYauAzzl
zF8aq8fhmjJucSLzInjuE/rLZMg5tSr1gkfwgSyJuPEkyQkpQv24DLk5ae9hsPfkfrocWN8C0ITi
Qt3LvKKcceL2xqaIEPmXOFa05yEPI8+QltvG7y2v6IsIaNVIMk4kvlf4xFzbmDvy01Yb1aMBvFkO
NWwrQ41kH2xSUUzxl20681bs4gfo2a7FOsL7H1q2lf9hcCVGmm2D8MlWYAyLfLvL6lDhv+hflmCg
+gFlOeh6tDBT3zsRKmiFGubUm7MBJGs0OPUp/sqVwgvqDwSWeTFZkgeq5dcxxCYlADoHD6eKwXck
86BcTLy5tvzhQe9+WPEUThf7Y2ECInDd+UmCLo6H/qLcSQvr+6DI26S5wd4LugilGWy1EhcJnDWx
PrFzl5VZ+sOrfveeZRYl0dj50UNCaDUUxwsQwBq9+n3REuCNnzxUF9KOgsqxG8GRKIbsx04w8Hjv
pmAK3jzV7VN5sU6+YiZf0t6Ln0Qis1F0V0iBSVt4Ea8dW2MMCqTtXPHzYA3cm5TMNLxMqz3h8oyQ
mq9+anA7mSqEFvl7earXPEtPRkAz4XSEE5WymxfVygPkck2FSSINMe/jg7axzzIqsyG6ad6eXptz
3gcDtNQaLNQpfZydF1gWVz+QNqwYW5y//LtQtogMjx1CKAxL1VYZTdQfUAfZeJaUovNaAzXZxTc4
dffXTJRwH1wBRG8fB9olUFWaMvLuRs2oN23u2hg2TE0aNin4qM6R4JMrluaSWfeH57LwxhQsOhyS
Norn+VcypSQuNWWu3CQx3Lig4HGS6ioTByFBlxjE+ITy1zY+lmcbTOUqUzW0utRhjpgqm7hkRhRq
cp8nJ9ohnXbrbGulZq2UrIS07Oz7Pz/ZNdbjtSLTsPs98oNhK/YiWfhUFW/ZXDWCOTQWgUq3Aa/o
3wluGi4zrMopiTz3D73/9BizxIYtAjohnc/qGzuk7V9ko7iTHg29E2wS96iBbrV2UUe7XHA5wvZU
eUghRMMYxsnTujVY6sgwTthOBwGahl7LtE6zchBhSrYyomPqUqHD7z56BHp/CtdQ0hTDeEoJbSgc
J5wqUZhTS7EAd5H8kKx+ZnCrC8X8IIaOKnq9jzN42z6ipdLJA8+TxTgZpcq3vDzgZMQZpSPsNW4W
qBsAzpnyhWv4OADM0DMakKi2/FWNMTQKbojpLIWUeHx4XRYIs4Pyoix+PVYdGod+pnSHqAxqhk5e
x+vgKXcia6Spb8IIceunN0Dcnf1AIwqydUnx0b+ZN9jfG5m0TPQge+12Y6dwrT+p5u3CO3NFRmRc
QYVfYWDUekc8pAYDTPi/mI4SuZbdM+dW1no1uqd4EJtUbBjbIdTi1Qv76UIjRyKxZNfLBj5GDoRo
M9gw9aZCVQimhDLSL+bF+3u6/XMJ+wwVCzOxlPPzHpNb3vnu0rRpp8bVRI3iJ1xXKGbVtm6RFps/
0zCSqkA1rG6uynliuceXKwBx5E69z7zr8n6/ojwMbHaldyxCHUijn6Hs6VSs6G1Lrbk+EwjKWRp0
QnRxaqRglgGHCLMMrgxjYD+Q530nfPPDdY4kvbntejz6Y3isLmoQ/4m72+SPxxlH2rTse+nmR8Pf
YGfTqXLTkvFSXZPa1QQE0eL4LXDKFcQbiE6rPXQkw8YfWxjckjKpelI4vtU1Q9wJSazm9wmxflrm
SORIMLFMeDnPwF8x9b1HkWYz9+NxDJd+AypBL/D4f1uOFxPG+x6ND0WjhyX+kh55NcSL5hFtL4Tr
KWtL4UmXq/DR3dpskpU236i9oRqarIL81uRhnLFTXheU39yiFcmBr7rOgXI9450AnBPt0d7EXzUB
kmSFTUu4Liv52maJxYPGC8ceayZC8AnhO0fdW/m2Tlj6XHB6ayWRtGjj0kCOVSGtEGmx7h8uRLU4
dUoi8nl7LABZ0cEv51fqR+WPPLeTecqhStNe2pYAN6ABe9VW5UcVU0m0TcETtAiNQI+W7cG6/Npt
4MNOqbb3F2pq9W3TxZ0j8KnbBCi/q718Im4kHVJS4hgxKHWTel2lJYH8DTh1gZkqQFpXj9VA2lZu
XAElWVDkw4w/XaZwi0Y8TYedFoMNhibHO1igRB/1fvmU5b2/YZaKB5YcOt1wGmt2cWN6MTvWEHGk
Wf0MfXqYHOM2Il6OxcPOHsWn4oebbK/brk21bWqVo4vlH4MmCIWU0Up+lSYE9ILUDTEwm6CNtJme
/KjQncbyb1G0+Y7HiRSz5YGeomFga2CxBJeKBuLDzYvrNMn55H+HLTRxw+rGfoptpk4eUxRlJ2tz
Jm1sM0rVAZAOrielPzhFoJ1V5R6ffmDQF30kUQD05CdS9XmvYS7xov1DLmMG3855fHZiFd6cclzx
ggBJJ9g99wn+hZ7tdveIGW+dsBkXynJ8s/ddcjyqJWnxK97pWkH2XSahRcMbjY4aNs9SY9iTEcZR
OCuei6DT0u5+rE37dxIuCJg5zBIAXABV+SZ54yvzlAgyw8Jimrswy0e1vLzNpilH9YnRmPD/IvX8
9NzVnF7PMAFxnu7W7Zkm2tTwRbWy6RrO1kfsJ3VCRGoVUnRse+e9fZY9zKTD+w5IwSjRgiFLelg3
UtR/0hXlzJyR1Dul+xzFyKVl4WgubLvXBpSsI1LxwjOLY6Q0n7EFIoE5pvDwdwupGXim4nV3/HXT
l3WX0Ebwe0V19gED71cmWPjoxGufVTMQECDEj7tviQ8Vg1/aemab6twdnV5v8Dyyg4IAnol3BUkg
F1dLhXIuWMC/uN2OWW9znQeO9DdZFj+pXijm5BISZikhvBDXxO+l0zMiOUdbCkyg0S6VrY9tgfoG
34fCECZ5GAvK4P8pkc4cGe/PhWe5ShIcOdl8K754dnv/nHDujN5xzIMkqYWYmQx7x7QVyLEQdnqw
VMV2Lc3Ora3Ysu79HTK3sNfVCyGi+DFyd3q/EZWCHQv1QEnw53nxYpFSM8Et6GrtX0Jmv9C7cV3u
/TrgbOHZm5yuo6YSGTLrwmH0weLZD82NVwjjVjZzlNV0KZ2ZmMYAY9zLv6xbDacfwfMH6+XDowsf
b5tw/tXVI4dh3yNrmAGa1DiVaYocVRN27eGrEWk7VXD8UxbTjSf7nAM8lpdV0LvZJPvcpqXikwMC
Uy564oBqeqQxzyEGcvMQjWgZpk0IcH0dIf70v3P/quwgMDs3FkVP1waq0O1CfcUcRAm1iv8DDGem
3fRPRJtF1nG3yWrsIcXf3UeMhTxBdHV5OeUNes4Orlwd9h/IyxDptCvr16BzcLU0Y5Wda+4QjyUo
KXAdMmFQUKGukqnlQ+vnHl797DD5OX9i6Xguw2K91EW+V1irlE68vq0w57fxvlkpkAQ7U7OuHBPe
ljtf38GY4TS6JEkLtWiM3QxWUs5C1HBxoqoaCZYF3RiAk2Co9g4u4aneJbF2Iix2Uscc48/W0xGS
c5yY7L9aV9xF8+Sb5uqdF2bn4ZdVz2orttyTDNC2xr378Ks4g+x5eOShPMValdI2CGYEEsx8C3SN
tSzCF5YYj5t48fKomwihlM1EXL5m+EKkLe1WtUKcTfFBDtzPVOvQ5I7GCwABETJdoE548AE5sXI9
YxgT7hjYtZJ3wlUy/qfVyP3H0jRGeVXL9llZcIYcv/locM2fCH7FHu0b7EcU9vKI8/AvhqveVCYS
2ct5Tlv8uteRUd2p0wbt6UUbx7acjqRcdr3VU4hT82/uXpwU8s7BF5fLPhzCJB4TTRJC8KXpx/ye
VXxdLHxGY2TcDf7JVHctjaOQcFdHmpgUbRry0jBfgdu/eJH0/mbypRGWPr7ZuXb0z3ypLtb38JT9
V6PUhYE5daAo1Fe3jHdeIoe22LH6JOT0J9LiuxuztI80i30cV5ErjCqYUXro29HpAwHx/2RG76hS
BpKO5S66hfMDYAk7lgJXjFfIpdk9SpLnrNWnJpjV0/ZeTFKoBUNftgbXZIfpRMSgFoJkzI8ROuv8
Nz8u0Pt+Lq5DJqJw+oqIboErGsLAAa3PapzcaIRpQecszp+zvt7FdyebMpF2f0HOUrFYzQ1//PQw
Q3lXa0Rj5NoeFJL1cToi4ZSMLdjZB0F/U9ELtao6RyCUiYYRzSgN1ug3FwB3O4MpGbq37LZ2i9Nl
aOQp+wquTu/FCkegbpxc4XVGtymLXjYOwAGZd48bgrIghEv3uMrNLAzosV1R87ecWCXGjv8QjAdj
J12EmHd5G3WwQ0e+JjwZFViAh7h5HszV/ZQUbsKPtiNzlGp1Hj25ciPaGN9jwxsI+WN58BoHsmuD
Jt2oABXMFyNDMpnJD+o4zr7twqv7vGULcBdZAOyWaGzhAmGHsi/C/Mibdmaxx6Tn7pi1/WaHucrr
P8L27YLbtqB2FesDNlO+noAbM78TIG6e368xCzqSvy3vaHnPIWFtOxSu8KGXiQyq9wvV05VNuncB
Ir6i6vfID9GYDqbG0isthmlLalrzMlpGqY56uS/T/qMELz7sjElT7QCYpDIkyY/UD0MEK6iVVFrs
zs9P36XrKj+IaKBibu8Me4C1hY6UKXxryBZKIaLuikAPrcJmP9shBhrrE2cx5El+bUfv0O6OGKpq
6ZJAAduMxGPD0aaWzVy0B8oZbbygf9zc1mjLPvafdMW4U6n+kSa9XphPAXV9pU0Ky5wOsvKfkoGu
nx3YeU57xb14o6mvau/yLQaQhOVFNZja3olbzoYjRassebE1SCORZ4kaPw2n0ba7hiWQnKEICc2X
BMpB8NmDZ0FhUE0rVZx4JU+m3RY4lD0EhwSfofR92lng1UC8Rmq5wZyOy2zKzEs7vrSh+G+s11Dk
cLVljKOx8fSDFHWsoTTz/LnZrQoj90xSxwz40tIw9SABEDQ8W5zyDSXNabBxFTL/IzkUvzmrZh83
euHWywKNc2K0uHaXtBhT2bqrFp2QKYiyisQp8/VUe4ztKpjd16aDlQkYog0v1uzJLQBRiJuYVPY7
RCB55ZOyjC3Fs8m+1OmpamraZrdCzjkF53Eme+Gux0DyyHYgNKfgqNkWd3hVmXymgl4AO6eWc7LW
+ynUeBwHKp+WNunvvCNGjmIx0WAAmQAI36UTBwnJJmYx9esF2PbgnMaj3nbAaev2LZIbLfWO4ZrD
+0L9HkxtL22o7pP49bey9JccI1k6ShFQ6K19ww0IQUsu96DC3dnF5qJWcKiTHTtcew48FmYm9tzO
xenc3+teaPUZ3UTp0zyt/RzjM+gtVyHOsAfJotbQDSq2Nayvvw7wFQGw/grVSWBfJQcC312UL5dW
1VXcAaIJIlr0bPgzbav5QkryRRo345N/e6wgqyx/eI5C4P+pqRBSquXTSA9hSh8Xtzr+/sneULTH
egPBhG7Nfdssj9wmo3+bB8Ll4gXjEReRjzr/kYr1cOxUAYlmFKH0qvu08fM2mV4g3n7bIv+BEzNo
Ovtql3A+rXucG9/fJxw+4zdm95vV6uk7l7w64x85uxQfFcCYFk/nsVNNFkH/7D04EPFuUaNDj2C8
qC4wR7zAVCdQRv5ifJRzoKBAV/W0PkUAlcqo1ogeqqyz/45Xmj1FQSegzEGHhRKDzjX54rdCUk//
7vKg/3AxtSADQ7Be45y15XlNGhIHDxixYRHYPgLteTdJyXB/JvEAgSX46fD4gDnVyloOqIHNRVfX
E+c9RTqop6CR5AhqmtNhhd3rIw9jNHGACNs8Bm8boPJw6N56y8q4H++/bae/WqMN4MIqod0TV1r2
kracjEhdfpQ3BoIDS/OJ5K3oL4M8FhxYGpxbtfyXQBT59NvO6GGszzRBecTsTCA2itI9qyB5mnTO
2O4pVeZYO1O+Udnc3WldwAY0mqkqlIKk/3Sjlukkz05eBfsL20ThJFTmJHCIPcEqo5WFtBPPFwKW
Z//mDhqUf7r36Osy4MlmTDihnf4D8+YZM4slpqf38QGzxAOPgHTpcn0TgbPnS9CAB4j/L6EL3Cm4
UUhsWg+/zDau2xHEwuqK3k4KiaFEwlZGSZNZbhqEiDJD3MAuvP5YtReqVb7JYMYgrgJdTEvj9XOX
Ostl0Bmyez1ghEQP91icPuc3xTq97ibaxQ73K9TQqjlA4tO9YidGenmPhA1dvj4I4zKflhxu+FTM
DKX06yvb/UTGNFOSFciEqfOxZ4VzPHw3f4BhJ7MIW0EPA+Bfej0XIA25mLIajoaWFuOdCAhwiN0s
JBz8fTPKYhefTQC1ONxGMN+hzcGHyR2Q6yVVNmZnDN9dSPLx8vPeqcIH0O/R7Tf0OComLmedl9kS
yf56AkUnXaOVCA2qI09qQZIxPof1oc7a5F88TRgEHOCHyX5yWFWguP/o8ZEFLKUfXPTm1GbWnDmr
UxsYGtjXGil2tYC1OIE/eQMM+vTmdcmAolmmZ57yDw5ku0Kzl4nMA922+cx9N0XisqjcHrc79pzG
7p0AafY6VHfyxP5q/g4y6vvwfuq0vejoEWvVavQzhwq5oVRAZis1Y8b1oHBjAEsYvNS4l+Vl7JAg
ajusxiJqnNElS6gcZIqNPZsp3imN09uhRzhD4i29Q90f+3g1AcwIY+s5ibEaVI4XTwLqT7oqMnl/
3XI6Lwo5qdfGqDgzUXxvk6IEi6B+0HAv0MF4bN2eG63+97Hw8AJmsXSYWotpCb667QkjcJaq0LIy
8nUYtRMxLan57h2LvnfKkr6tTyDFVLg5plxkLZCucyu1hBXVRmWcribpf37ElNJzomV/vrxxmkJz
DPYO29+iiWcwS9cSpkDmpSAeEGKV91fFsyfUcgn/blg7BAzK+nH60eLEjEUrvX+iguhht7iVpMPd
vCJFtkdu/z4dczSdoi5jRzfr/W/ianl5LpmI86PjWJHv1EJcUaLQ5IALx/SGSlecVpNmzScdIezx
QNCzZmDyZ9/wsO/BmfVbQ7NGVIolX69CKyzOC1zIYZNkGqhGxjiUT17GMrbLgJnlZx6Z+N6xmZ6B
p3hJzRpTDL06PnvgUUiDsHgGvsgYA1a9C+4U7+OCJtouHF0En4teFDQ9EhnYB+9DBnZ5nqOHDJk6
sWxrQJiQqitgMrvtp42YnjXTk8KGWfefp5Da46Pxz41a6j4+TGZ7fgLLIHDtp1IqIYkRksLulqyV
IW17jXw//WHfEKYF4BvJTA5ouOJjap3x5qauN5LFY9MiduAG5Ot54BHyvX9sNFBowy+1TBbHACan
OME5nv9XwIwkat8LYbKrRa3wQcuZTG3Fz/gJBxyZfxpgl3QJctdV5ta8tTMAYsSLZUEd5YlsU77f
nPFvF7hTyBkQu4Eezc5OthwA0fRq43Zcs0oUOCWuLLBppqAgjcDytwOICXrOvoQMwhNo5OqfaHG2
DjkOt+DL/y2TWtLWFBn2W11qs8LVqnSHhEfyzRjx6HBITUZuVVMJN74eg9MV99MEZmpQ4OLgVyBc
Zwc638HNNlY5WitSIOJvN/buAPzV9pgO1oTyZHFANBp30KyFxl0Dl5r0Xq+5fgMjYm07C/9ruPth
i0Wf2rl8WHPiAiclgVXi2dUFgRro0lLUwBHuSLO8sQ5FZ8WQp6XiirPEp7F6n4KircC3xgR5tjp2
3At1wy/dCk43c2rLP9ul7+5xqydT93fKDBLZdLe3t/xAqGWhN/8t6Q4LlFYSYzVVegvwqKJ1O+xv
9Q2nHcCxVg06D10wYwRkF55JrcEQXpi3ndcBt6LR4eDK5/KMWYc2YSkHFjv7osZfM0xHElIWaG21
TqoNqqsHBTqGIJx+L55BhmFgm0oL3cnY8+a3DFxHj/ECnlTTBNFYfqlEfL3NGxSx9JTMX3alMm3P
gLVwDgORIgRegp7zgWyrhw5aI5+TxybMSXDKy6SosZ0uQ6Frgt516LK3Y/OY3V15MHezWEBkUJ0U
VKu58XYajVIp2g25Fmat+1J9o6q1VIouA65ikoqjq7OTl8RsFFTbXAkxO9D5nfq8YIMcoF3nXMpX
XfT0B2oMdsO27A0MnEblmfAD6EgOEKAmifNaQiPPQrbkFZkbT5YUO1iRhhp7HAvFRJ0SaWU7qUNQ
lovkNngj1QTh3aYYd0yefxlaxfDUW0uB5lNaTNqhC3gEcgCRnNKyKPMI+dy9gme7gghQ7N7tbhAA
QyOSp5r2jCTb3vyyENxDYG+B5lviYk1oIEyDdAasVeLikBMI7e3cij7Kl+PW+UT3vcx/AehaELca
aTFrBY69a5Tz2YsHSzZhHcp4MzGasmymrmaHNCXtGsuZYNAplEp6ZAoNB1kBtGvbagyZigLUZ5ZU
57XGTkkl+/4i53M6UrJn64Kw2gh38auBGKYFAFB24KJvxfFkk6cGhiL0jB33S6BGuVe5GrbdcPsJ
hiP0bnijrqQu9gNeEHZyF+BagvMCdQuwlcyGrFOYevPmQIwwDHrWtgZ6eqUDSZ/J+78BtN+PwjvF
/KDd9i6VVj+7XYswMEwlJy3/mM2mKk5rLGWOfGgVJfzSnbkiDNpMMlAg3jwq3ff05OE3+of7MLki
0o3JrvpiD2MBEjy8XVp1mhumoaotyVDifUnrxD1lF5kJcp0vlIEKCDrKj39vazVGyLjbTCQeQkjI
rDoxTHkoFsJfnqxAvmbGVqQ3uUskHy5iyJ1kqacau7EIzYpFiEconZ/fxB+bpFQYIYIB8ygjm4Ng
YHb45MRL6Hn23G1svAoXVkkI4ZwtYHflJqUIzhRUZYxntI2+ygL1whDO1kgYgFs1pKVJSDlyI4rH
tE5gRreEJcIBaEUhKWx4ZUXgRRkzG9MzO7Tle3+qLSo/eWjHyzkU5ZGPgx1BA2VOnstyI8hJ9pv9
ivaYJbXFOr2dg4t3KWfnUQ91WqoKzCVeux/XMEJgVDMnZRtKMKWtbrMNfx2fSAyDo7VZsrDcfgU5
BdH2sDV5sVHfNtNqkTFebgptSllvUb0iWT6e/OhnXwBMdApexhIUgQiIOQrHQeyeXCXjJDYdGR0U
CtWD+Bc0CDuTFCl+XymMFKQCFOK7LMXHERulHd+ZqI+hyCRo76uhwiLAYNaVpWA2NFwSPMFspFea
ekdrs7mliya6Bx2GIOasAUHfgF/z1Z0b8o7Dr5v7W7hwejgFshpR5NWiJVy9yW+5CbusFR2KNuGD
uQpsY7bOIBPVD/yOyITa2h5P5x6MhQ7OXSYSxOGqOqkfurawz4NCF5N6HP0i0yH5i0BKmnYHaPwZ
6qLlxcRZ276rAdbIfj2aSj5PLs+A/1h4XXySDUfYQqhtq3cxgVxfy+9232Jarb7JpwYKT+/xhoQX
z6DK/X6z1uC/qgfTAbeBAy1PBmiIJbSQI+45LbXHB1fL7E5XvTz8YXjKe4M8fRpHYZTZQMXmPs8u
rD8rbsyQuKXmUmJc9NRjbqWyRn4xM/eTj6DhQkNNVDWkQ7P9yz9zbBJvp2rjgkMzOndPTtg9IEy8
VbGuasbOn4xtcrftdyXaKqsiIFbe6Kba0nJWfCGpApINjhAeuNcNmhpXpxe/Yx64SmfzlkvYcwER
+krsxk+BIwIyuDNLu1xftVcajCjFWCi9baURZFEZKgS26xMv9Om8aqe9D3+2tvRqOws2cNQKC7o7
EbPttcweqYIhC/VG4vqNIHsbZOYMVDAGSrPJZRm+LmAUKgZQv3FJMFi/XPbL3uU6Wb3rhg77S9wX
38dse2+Hakq0FMAVW0D1zdiA/b0M3wfESYDF/CT58rUN2ZExZTpgeDEyPY/5ChZTrzyFwVYdu/sW
I9bdTHqwmQ03kn0q9W6PFElWWIEvJW7DaMqAwAbE8GKi2sQgoJw2lmu2aB7ryOfxVtmVWuAZ29ZR
S/9l5mLyKi3ODhUKjcbvfvBakbRMr+WD3BG5gtOHwY30AvCA8WL3910nJpYEY7s1QNeIXdQs5OxR
ciXkTzYyZ+Pl6TlmSXDCV5U0op8Td09ldIpwzg/84A4W/esNoEP2h3f6AX20wWTtKeq4HpUAhWoW
E9pmvMkbF0vJ1YUBhYws5QGObnkMDZ72d/nVyan9g5dNb2vHWm7RPFdiisvjWmQN4LkTW+0vvHRn
HUhmga0AHNIdYMr+JLRw4HY2ZDtRLtVUSKxOF+opQGmJN6/I2LbK7pQYtdVw9uQ5lsrfHQyRDE1g
yl16btOZOelBGnGvZsZoU/SdWI/VnLrAuGLMliLzzujQOUj/N3KTEI9SA96vjKDbCDku5jKBL7M7
4zwkt2ft+xn61c+Tj9vQsKWK/48pI+lvweuBkon9eKtutwyFpi9zVgt5T0jWl2msNUX1a6wbf++k
dv+XuAPdxSdV7nohQQTZ/DNkzXKEgeJ6BF0QnKv4qWwOTGHVgzE0MEh2wvbGv7ZQzNrdwKrcIt/x
WeN9L8Pfw4dvcuxibD0py2jlPUwKEr8E+ZXMYEVgM7WVlzYW9nxPgXIb8e1eskP1a2WXTDRY3ss2
Pef5/QaflUAadgzbPcHGpDZkWSCEugnfTVWV3YShXEUkkeGcXTBOKG959lb1UrKC59NdD48KLSow
wXYbJyE1yQHV7eOMCvTjBvzjrZMXqDVQ2oYc1myDuHrBYqn4WKOXhgyvDxOfB4Wh+hEZx0pbPZBe
or7meB6LVomdt6kHeb8/YqbBs3dMFO6Gzr7lECRpwZI8Np3CA1uWV92Nt18kYe0tpeS7h60hMY++
f4BT453UZWh69fnEM0uaESRAETov4xQzPrfld6/XQIu3ncnViCht55IrmGyhmjO4LSryUx0Lb/b5
Pw/ElssyuyhFh1g+eETQ+ZNuauizwUl1XybihsWXgE7GOUe/ie0J5JiAOP2LqIk8JScA+jcQvB+o
d2Rg6BEXi9gB97lwqzV3mWnaPk9tCooEkVJ2ZQL6k2ziiI6jgILQPKAS11bUtUhqwB9I71irHS0h
eY2WIMSsLlBM7DD3PYZm/niZHphQ4DfcxpyTW82OGuKgDcP3ckbv3Y/bZO4XiaFzGvXdQN+Lv7QN
lN+km7/UXehkZWm1WxFiXD/tg472fLwMhqHktw1Jwba6MUHnuhTeLOPJDpZQ5WGlu61TCTNCxsKs
SSRNYPnjvfkANpI2wAo/IhzZ+5GyIEWalI2oA3rgDXcOfAeXFMUCMbvk1lRPxAuWK227/RXv4v3B
8yIOCYNsMd00gGlSgUwosPOOcYJeQBLTsZvECtvgFXAm1fLzuMBG80V5EB0VhDi36czE4lfv2Kdf
xpRDjsPCSS67IhW9hCGEX2g8jiDhz65i6r1moN+LIvMXezJYy6k7OffTjtTEilP814fa1kB4rWey
1FHXiSscVIbx0sUhace4WjnIdI1GSnr0qFHVJpvJYCYnu7+c26rRAphtCvl8AMPAobt9d1muKupY
lcpodaElInGcAznTL340AtMfWVzxD+FeCWJU/Bd+0APNnIsgQhXVt/Yu1KGZ41XU/YApgKpDXHD2
cKXZiGxfX99+IRg02DRnY30lba0U5QK/twTVljL54/D3y+PmY99cIl0Ll5y07fKo9RbaRZQBFNyu
MZ84oZuxYW1Yu7qfZhX0dcfDvGl0sEGPbTMs3oP79AyQbBfrt78ewlyo/1XgH5O8Yi3mOw44JHO1
uKCZXCnbCKgTdQYpcWRyabskKg3mGMIN/Jqoj1RRgZkh4m/DW+yThHh8sORpnhDm9PL6M542gJON
FojqFekQZ++8t5XQV2xJcy+ZQHTnBYtmhtEMp+8KVhvDdxsjWL5UfHFsFlhp2B9eTE6pex7HHlUp
FryvA96qrfali/ChKhVajWbySyEL00K1BOQ8t01P7uwAy4WbT0K5xH1LVIcuZKIraPKUhXq/MUon
SU0xIznUx7LPfjzNh7bm5u1mOOBULr0+gKl2yRr4CM4l/M+Yxte2KIppmB/L323ChgE7s66XJ9wR
pkZm7MGTA7Btf7DNBjwuS04CuF1eDEF7Iy6MPH7/2L/lFK5yn0dhXzGMJEm7/aq/78uz54xgMSiF
FPh6Pj6QoyuuKDW6Xxubo5YT2w9ZEeSVdzJa7PZaTl36LcKgvNnkB4fZPJ5h4Y/jDccPu9u2JLZr
tYFQHE6tdvPplbyj377nnkW5bs4l2qFraylo6Sl0sFNkitOZD19g4Qr8p8Q3N9W0r7IdpMDg913D
7wJwzrlrrcMjF8JHbp/6OdpOoCm2uPxcMmywXCggc7K4A+RI7hdlpf00u6btbgCU+hMmh6cwoG90
olU898IMvzAtm8BRXZBezb4PHdD7sNiF4ru1HGjL9oLHQpKW1Yc5Oz7mh1agTl0Tzg5XnO2y7lLo
Ka5TWI5wxoMLPAgOsN7KmRQxs+CpaAKRwMZDA2q87TZ802192s+H7zRVte07fkl3WAHr5RAFw/5n
7F9YICUjOR8J8dVP33R/Dc6mOreGrF2HdLY4UT9WbvO7yrRZxFLkMZgdUolFT7apZ+Xu4NqdpTc9
9/jrDsS2VvVwSUXlxmYvmNdDt0xKQcVdhVk/7dns0KPIrWiNe+pLUFUocIsM+bxg07FHFrB6DPsB
tgcMGCbqFu9kfWDNvNYnCqwKalexGFJaz4SG9gA+mw2mwZs3Z7gKfuvFxw2Frfw0/sN1pE+Lx7ph
vFdZFcQFvke3ZdVpOL36dC5yU2q2rM9z0laca+j2yRcqfh24OYesNQ3KKP/4ScdSDE9ACl2XBiYc
5KAj1WctJXfFt0QdENZ/GlaFuTcEoFv5L1OH5Lf1jjTgWzvO1GlgaLt9EkUmZgXo/X4LHS+wZmFl
+N0p6/k+loZUb/pgusz3GjSIUZgaR2Y7KVwVPnzxZ+eszIPS/kjotXE81nxIX4yd1TBNOVQT7euh
o7NwEHw0mHb2BiPIqyhFD0BtXp/18kOUbv2kqVUKt3Zjv3oYenWSTPwQt+DBvDZgO7r78o3hvguf
qLHwtkJxC3XSjeeLa7rjXSq//su4FwbmKHL+fVSrEZb9o2VXhPI57tB6252tyL51cm/RhQGHMl0+
yke7mGGG9c2Xp7lsP0OLiyez9FZpw41pNRcFSIbK7wj0yFsNMF5XIDrD7FcTiXTOtEqqv5dOVB+W
UdcsnBy2WDR3tSwR/7db6HS3tBCM7jH4FEm8LlCS/16PQVc0xAxGsBpnykX7pIH/mZNtowqnEDbE
g+CcSr/fTNQKQ7IH7qBvS7OqoInXvX6DCp8zD7WGTY4qRETH2WZyjJqAdnIfRORscEGkeqO4Dcaz
Q9zUgT1J+6Vc2fzwRS9kZ4It8YFAWZjch21/E6Ixs/isRQy8rsD7XY1caHItsG0rvCFtznmSs+o+
JUeu3VMmyft+IB5GEC5KPZIpv4rXtJIHD3Ijlg+o2n7J1Ul1iewunxitrB87o9bPsszV3xxT5j6u
WfiBusXuZVLrTGaqvkDYg0NAnuers2CbyaqEej6zo8t+COFdc4KOPXPRQcmzKXs9szdRIp0tZ05g
9kO+8ncr/OVktj1XupsUvosonH0gz6IMBBUzrCX80EFpDhVwqzK05BoieyzYeA0kDlSkZgNROUiS
Il7SjeHBjXWMNYVlI+U//QrVq6OFoPDP+ZKceI4vQc62g6IaadTRqldRS2l4PcLL9C7GVHLbrar7
Z/wVO1OsGDfCMhoGopB5LrKG/OMHmGKS2ESPhIgqoEkFK4+2+Wo1ZBR3Sz4FfG6c7V92Y1tdlcKI
052j3U5yrf60gu9ceAok+d7QbOPWqlksYXKOMtCDPIFSqj7ZFocji3gX7cDcEIxazzPH7P16WdR2
nIwnfmNdKTFklyo+cn7Fsj2dfQjThWLmHVfOB9lExw4kCeoJ5ONV6zFJesxtlbNkfiHl2jhHhq8D
dCH26gsp2p5PrconS8+9FQm51fwBSxsCzp6Yd5GI8FylbHxbr6adzRmSzlrOxpTNZlgtyXdahTwu
Fko/78reg9Img7MCWrKoUM4yWd7jadDXPYpMl53vvg++OG2iGb0/qewOir/BSRec+ZPDrZmiXenD
BwSAPO4g7fsf964OcI42mIXn+Nf0OoddWsPd2AOpjewcAHo6HAoJu31ziT0QUJ4HQV1zAyph4s5/
mDn+eztoJ54UYnLq31Ct80EjAprNs/TPxfz5VRa2SXoeEAQClDRHOYJ4vvQNNHFwLBSWgII7gnJI
S513sVcoH4cfu2055cdqdqGeh1bo3eRM52xvITEQMstq1NeyoXhYcM+Icd+S+bTriOZUdEhFS51V
HuRb0rJzG+alhv+j24kUNb793uDYmMXls4KtRr7lMBzvq32JeG3HpTzME5J8IlEJ9wAF7oFeFInc
kQqj28K/CEffjeA+0AIFtyRO6mpmys/kd40u3uJRk45TjbPxowxKRqUw8JHbqQjWowDS6iQFBmCX
DOkQGQzJQOoLtdNk/D2Ankvd7BRKfA4Vo1epzzVgAuYPqkc6ldLgRjJFXIwP1y8rWTQOYW7GJ0Fl
QL+ITOASP2rbz8M865jRhhzMb0RcuJeUxC0fT+LZsf0kRo0/drUVJnuL/4FFX0F8qHnJbdwM5JKB
J++8rfUGnYWygjWJ5BezNraN85kIKrWIzX2c4lkyvyUQR95SSsREX1i3ujBt6BZED55VeppVwMKP
q/aCQJwPN301yjSd8CeIX3bru/XIanchNSLasoWaLZXKop9rtlbE/uFqGoXjhk+ahbnnpigSG6fl
knhPslOQI38M/HrTzNMvkRLkqVMqPEdKeW6xgWDOMZ/guHhNf3DNMi9oTTPKP+lV/FrzfvQuVhNW
AOiwh81xCHLROQkTPXNMmnXK4c2gYa67MW27xifm37TOXXwC2wFy0mVjYIsV3cnQp64DQJo5hpwN
ozxNhoNXxvxO2/UucxqNspWw8AgpymzTnt6hMYDgwmBHofvTnOzYZAX5f/aVXsMp0P6qpZ9U0m9i
mabaZ6iPjbtkfITwjklXimRuPWuuvUdb0EfC9udaBPL4ZFe3LMLtYkvGe8tDfgiUChHMNgJev9ZY
9/RXxsfpvkSajmFIDKkoUKd6Xo8l6x4IltcIsiVB/HiPrbrt4y9swCXconwHuVSII7XABEQba9iW
BawA30MymEBMpBu88shYzRMtJZaDtVcjIv8zU1KfxWeYUjZ/eZrfesQ/rO4eiaIbZt9rMZ8Hiy3V
Qfd+C8SXpKj5T4qn/6r+BcSGNHunSeOmww9/3kQ/G1ZuTd77BUDiV6QOC70P/7szcHXI17YcriqQ
C+LJH34PDTKdB6uRqCWBy3+BMHeO3I6FYOyIvmbbqpe/XRUFBNrgFjroxkF1hPU8zJ4ETSNj+HrF
0weNTlpncKwf5suRmZrKrZT2dnYc2iqhR95EK5K/L7JLakUNO6ntJ8MykeUyNa0+mYXHezFOSz22
TVVUWeXAS2s2J0O+lHo/ad3pniAfbt+ZPKAi3L0IPDAXh59kgqC2R+R4SXRP1fvBOM9vwv1Bb0Hi
owuBju8Wy7hpEQ9Wq00Xnp85xHTmIQVLpydmjd5y8R/3VLbT3wuwXCoHaimzMeTUs0ntbzoP+A9W
IIvZ5ZdrD2udGuKxZ0KHr9Ro8hSj41HdjAtdPMpFfCvJOJz3BUe4HZgButlAwCRoMShExmTuwaYm
2vst8GwD0qsuaGg1wQnOMyl9+qH/0zjh5uUOQsZgfaGusgy2yS4SYbjP0IEkeGjJ60z1oveckULE
9J5yPaOFPxXB8WmHhdQfq93gXu41DKW1E37LAT4FNZn5P3nqmm0sJyMLUfklZAvhkaN2Zoer92yP
LTN8nIUk+wUlTaNGk/abrom4SVsO+5Kd4pFoCTTjK5qzSz6/IfCJmqlD49n91Aq13fNOEMnSqGbF
f2ROEMOBU8CT7l/qLD1GtHK1rQzTiJQCKvmaCVntuQri35flEYhSlYjUz3yZo3MdenrDURwvxR+G
EmD7ysqa59E31Mdcf7b6wZW3yFbneykxdlasJU6IlXvYf2QySs7zXdgu5WJgWKW0jCi+gpGEPxlA
19IeZxtHMFTqzbv5Z2NN8F3rFwcvS26jBTO4DoxJM3feQJL3gBbhDvdp5kwoLGfG9M0uKE7ZDzJL
M+6ZCFGOn78zxhVofTAkbNjlYqVjllgmcf9L9gdCiZAKzXJ59jWT2ZriV6JSCowqrDfmRWbthHwW
b14HS4A/PGFNeS0D2810xebzlBOy4VIcsbEf5qxL9VRfdhEQgo4GR2Oq+zZB9XaC60O4SVv7SVGd
U0/9k1Dm2mAC28iiwR2eHgl4HipxZlZzxvsyF4TlpsJ1s4k5G9r+S7LEpB2UZhOUiF1aF+V82NjZ
bHhUi88BxwrOgavPlKiZwUOq4AH0NLjki77CsuOknbyyZgjfzXvr52lbKJTk7cPb2/E1HAXVq+V5
dxKnPkZ3DO6F9BYJEz9789x2eTtDCVLNsYYqSYLVisM0Kz20fICnHoIK6ElN+tXShrrAA+RvDmBK
LZX8xhMU50RXKucsCrAtK2CM4ygY8FKJ+AylSS9wqai4cPaHWVqi5NF4nBxeitD6sMyDEvWRiE91
Ssp3DFgC8iGw62L3vUG4XawqIKnPgj0wBbiUrfXOtv0OW3RHkF1cL9Tjm1dMVg2UOZQ7RElxbu2f
m8McfkkKIgIahQGa5kt5lvcghZGVhFNKbC+eVUR7zQsaiyFNkD85mwX7gvUbCjQ4yzkuYFbFBp28
/Y4Cu+goMkWxW7nUf0urKIZ8LnWOmeLYPyvJsk2ia9OxGbiOQ+n32LrVl2noZypPMhGWKmRidFGU
3l5VpcooKqJX/bkH8Jsi079wM8IDygdgSWjdXDZkkVXNJwYAEpmKDFmrW3E9n02Fv8K2f2qwFDnk
8qanow5GeN7xojc4BdVVGUS1tFtB8yOWv7wLGSfvuJsCA4fX5ZV+URAbDTapwTomoqXPguuMr25s
0ijT48ENfeoEqAzM8MHNCxNKKKHesdZYlOscuzR7WcEBu33QnlAuc+Mve6cPVeBo/dUOytGnatk9
pwXibGI/8Oq48VGpGyk/tPbTwYcskcN+0etNMfAwc637Zp+H0Ges1Z/K+ryiz0DpR3ETdVWlsWKc
RzlYXmpRh/kDyD5EAVZMo/BNI/9sdMaOzhUko9wvqMRvWW9A4utWHKVEMEXvpMHEpe5iZ3dg/rEq
C924/hiK4zgSt5KpfbS1HqYd5+ggMOaF4/H/e8YOsEqnrpqWSNlqgWAGLsA6MS03whNMqBqV2UDM
X2RrhfLEB/oJDDbySV6h940/0N20HAqoVVON0+bSdr/1onHJ37bmlXnn7dIMqbYm35gEP6BfN7zU
e8BczVQJ+ttClx7U3Y/MSDmRu9n0+j9fN7QU9cC6zLtW/Q73WySfaGV+eY4vP/Fr1Zp1vZJ3noIj
sP+M7qFPn8sbmc5Do3JQngC95xEEPuWTiX//mCiTKmgR3nPhv8NjmXbYy5QLFphpaDLYhpjr3ILO
ZL7Hlu94xh+PFbsPoeLSf9opPBw7YYAQEAszURKgjUkXbYEDjdx/h9TnN+E9GeNmQ81DjHfvtHOy
FtdYkDTuXuoiscLc5oleBiUgN9b1j2p/N5mNLwVXNhyDi7lzw+WsqIT8/a2yDlH1+N+nwKjvDSXR
8/usom+NutJrTsg88nqTDNcg6kow0tciuhgrqNnvWXTNNTt6l3zTRIi1X9HFMyaYCl3BSHUihfFP
jFbYW4b85o/ALFJchUvg1Q3eKSS4LAGd847z6ga7P7Mv88dGNlBCz5SCBxfO3xpRfL7lCQ51ujjE
9xCjRI/XK8FpoWywVK8NlhkRGwaqNoSDGlc/8SN6O1CYbusEQWtBEVlCgg9SP3j5o9KiqJEPNQ+g
rs0FE5TkUOh1YPeA5bAmvsvsUzafFtuVQiZr+2aO+ptIY4f1MErkf6lrYdll9ZlR111HgQ4Fw/JJ
A/f9a4S1riTIGJnHUhZBR6HLm7WaBepxyklHp2QDS8tbTJMuEHt/dehH+NY07GJPKzuKO9D22q2Y
Ow29MJFGDyvpbojIJG0QcuyQJ8qhJX+GdtdWLcXtv+X8CjL3QXWefck1vQLCsL8aaj4/uOYvorn7
pl+I8G9xBdy7NFaa6BWqvTidvx87hulNvPM8oCLndTdmuYXou4vwXfcl5q6ZcrIxHD4wmAJxspF8
BE6qmU4w6DCsAvX6qGDfcbmrBlMbbjLNWXpCTcolCMsEuk0E6Uh+kbrSEuepKhHuJodGk2IQYDNl
yPqer843r8C5Ir/B6+CyzHruD2CGT4TQ7I2ldvQ7aVpsWimRocZuLaH/n+v/tWi1P4ywX2mqkf5C
eY/EXZ++/stdu3BaxLVKuqzkIHJqvhNeCr8gsLjINlPOeDlqsAGw+VFYgQz5656mZxONeNSnbfDx
WtocOtYqdw1soF/nbUgux/wA8ylnqFMDN5ard/JgaXtfG9kxm0A+5RkzK4nF1/fzH2tVYyk5nVbh
eFuLunvOn6WG+wZttc1MeW72McIRFRkOz8gMYFOPWOw7bX15xOsZrXS6A/K5RHBy2for+8I+LUzT
N52/5EO5pB4wTG0ZrpsToyH6arMZP/GYHbyzDFX/FOtRAlu5F1gqHHOatz7wSyYrVe3SOeYqw+Vd
og+nn/UIgSHsln8TUUfu/uNw/s0VehZdwbOirpckF9m9SeQqfjRHc1BGdOmEoghgvR4emwqci3QQ
8HTPJiHuuF7epGwsQ84dG2ouNB0AYO9d5gOg02EhG8yhO/Qbx2rdOggd+aW5Ujdht4f3yloGXx0Z
LEy8ty8oJR7sy0z4Eh0lFE6jl7CrCsOcgJUOPFtL6tV6A2NjKZJoyDSHW368TuZop0kHfp7FB3Tg
jj/lMyVPxvU5C6autPzgI8oWhNufGSsH9VwnBi9metUh53M0TKYpM2X6fOHaixTwIbgGOBPpt0DU
l0UuO9X6rfuQcQoBu9bn502St2sUCDjMT0/VFa0QYti3yjPahNyuV/UJu3smGLMYEgliHUtCckFD
8WS8DyQe/MY55KTQhJiGemrWs0t98uOIZfELlrbNMKqgdAE6biVbdj2Vgmrl5dvfRShHmengUHJn
DKAi6QxgWaEXngNMSyfxPtAmKNi8/5Wr2Ul64p3rQg0PGWXqSSPtMPZA5MRW2PCQ/aXKAvLrtzX7
oTRMVvynKBGpIkqOV3kfp690ctsmiCe35GQiyeEpKhlp/+FRAh5H+hFgrDL4GxfIrv6JEtGMScRP
zC+e2EE/Ygqlat99f0V5auj88qWeYu2vNPIsDDHuQCXswJcAZcYRZmD9t1oDav+V0wicg4LtAiuF
8d2Ed0an75TfrYtLZtYyPT5PjifqCei4Yx8QwUa58yOpl7n0o0hY+gFDnb90sn4Xls7nso5Ad5xF
yCf+xJwJ6YRFHE6EWnFaYio8xkP5bO2YEvU0oOx4zIsdfWERl4/ZW2uZUC4dPIYjhEiW9FQX5FK8
rw4FHtVdRwwHDWBIa9F6fzxvRu4smI4dOyf2HZohbjeqEs3R/tZeRJLkSyejFsRFLCReixFZdtI8
p3xWQbApJQOFrZtJMLQ5xmswPOTGnKNfIq8mkM3+jwOsxJru1P2Z5/7/0QZ5B7d6i1gZLOC+1izg
38o3HwDwreusyTCiWjYIowDo00VNC+DS3sCb7AwF6C84C3mPQCbna2AvQEmWDF/29ySxohvNHzu4
8ufCBsFOQ8SwdhhzaHF9W+jINpjYNc34j/vLrV6dEEcvQ8N/WlUx1wyBs0n6V9j6EkOzc4IO+QfX
o/Eq6JUS8yLZX2BK/Jk0bZbel2kocDZiy5xNzu9MTfWCK/SXUy8sbuHCcIgpSdXxJrK3CY8yPMjO
gspLmzFLtF81TeqBFz54mYt6KjD2gfJzBx97H2W/n9NOOSVwTQCd8LL3TGsjyh8Q5SuSBnP3Y2UH
Y1zQa1smZSnTs4hJIdlmSHY2p6xr1T4aWdLdDwhYXgnqb6H21rsj8rpaRWfyFFPy3uMYIJzyDVYd
htlwtyMjqlUlxg6820TEcN8dYwCG1GZ5Bk0TZNwLud5a5UUb5lN+RgPvnKf5zuS9zc0fopHoPOCZ
wOKmCH7K+IaCrfEobIDRGggUZaY8R8PaZYFTZlFu6/UsOc2EX46rsRoZUCvhgvuEjSqZTYUEhvSL
fjOxu+g+SvqKPa944nN7Gs77rdzJI4YAZHIejZ2I2NylnOSgK+V3u2Aru6kS3D3wkPVOujSx6bD/
A/FrVO4yo4j42biLow1SalW7/O/hr6looVp/r+Pl8hx6F5dYFyeACeV6hKLPrP4HUSbl/R0DtFqW
1TkxAyoYuy8NREKJEaCiS/7gEROBNxudzF62TDdTDonnq2sX+WiWmm/iGG2xsyqEjFgzNJsWNEBM
PKAvhrefGCAIPMXyr/2Oyf93uX2h4Tnl1n2/5RVkE5vKz4IlodVTXZXyl+5uXsJitl50mWO+g90N
DO2gjqjJxyRwD6AopG9hclhVDNTb9godJrlt/3I7T2biczGiYfOzjiQa9nQ0vrBaXe3CTeYs/h10
jEhkon8/8dMl3+huZXe6CDgPksoVzXAUDSpZxXKiyhOwjO/l2T5Afhhgay55nQJOnqWVp+sxyYd3
Hj2Os91OVTJp3tQ7QMiIpJ+7yYyMAR4Fc95hFUXLS1HqtD01PS7auO4ZMt+7p4MkhTo3Fl+Ub0nt
8BsvuAMvAK7JCopngp3fxEbEDdt7DmEQce7MXniY5CXeG2W/DW+66QHxVKhWKFzGDnJz9TUjAq5H
Y5L70CCrvGVogFHGM9ntwJqGlswJQLNcd3Mi2J6p8ErKXTKpS7wzshx2KpLAxYIdyZtI6yvAywB4
HPYN3bjSifDAzeLk8vAsXhmB4WIYRriSlasUGHvEP1mq/xcDd0dtqSR2mRvRTE2XkicnNMgMGwQU
MXWgv53SO8LdwEocAC+gh+daQkbRNG7aoydQonBEM9FTDsIW1FPkozhhDErj/uQOdfqgEUsRtKkM
XY0L0h+F3bNOxrNNwnCiCEcTgjTJUG8r2EK/yxw3Qe8yuv/pj/CZggu0d+WICe0xVSS1MyQAgPwG
lT3PoCJ/FzGGyUQihFupj1F56pNaFzqtsD11KI9vDkYf/dKKSBMkHNUbSELoC1JSAydtU74zj0Kh
O7TlVXXUf5LuxIJNXyZpfWm6K2VRnu9UTkzK75ZgC6wvT1NNfs9YHc38M5q30EFk9HaGz+Ac16vB
CJVbajD0wZbFG1IZIL6RTx5PoRz73CTk9lZFH4jRwAumxIYnEUkenar4FxLHECjZNmvijnMxCsRU
uqvT2x+Ek6em8SEdHuu8CFaJDoM8ujy6lhrkRGc7YPZ7a76lB6BaxsKGpVQGQYrE6kToYwROAI+P
YhNFJASN6vYOeNDHuuVgA5yBgNE2XsvO6CqXjqWvbMuroXv8vf3DgwTUHnzIUSskK+Y0lirIDs/A
8MkKrODpEnn95wvuJRIuIjWD59nastqh+FHt03GjuzsrT64vXd4vf7lob3vOfAPqN2/vrJlL69K8
o/uaIW4bBK5a0AtaxUQukcrqvEKjVJRK2RQ4rw49MobnBrPewXiVJNSkleqQ4XmSmIcg+zTqdkOJ
0cTdZiNlTudm+WrOkT0fRGZcKuCCZ9NXdWCmfTtZxWlB21D7+wvtQM65SRI+FqxASYyJxb517rFX
z+SS8haHWlpw4BohWPFZzDeAspO4KzBkSfJwZ8ZgqsHeDg+NysHeemBOPxsGYPZFlHiBcD5EcZA4
c+P49P12VBL09ORajraU2JqfNM8TKr+OiuL36ctFKLc75S3PMhVMKv6ozLdsanXdsF6L8zfSMI1x
mRMu22Oxui98RblRglSuGDti+CxiYTPBFVVWMxGUnV5112wNJaCWlvm7NB2fMLLMvYMdPdVkfkzF
CzOxx+GpR+hivBtCxhpJF5cESTCHE8WAF3VeA2EwmmO9lhBV9HKtl9mSMXRtgwGBzc8tseZojsgq
6OJ8oJ4wfW2PVZya1CbIoIR7+FLGlEmRepuX8Rqxb1sf5gY8gGONQ5Yk/P2997tfBZNTps/F4VRy
ZPg7Xm0yLz5CR6xfhXYSz/qhRMsCXmT7JawOxIK+aj+jHTTcR0ITD3sgVMO/VmKwvRmoJjU9cUhL
W4lVC1B43nNQEhcVP9VwIoh2Mji5wEtiWyef19VNAc7s8n4nDxaTuA147eDArKibb4VpfIAHiAs2
+n1WyHPw2OCOH+HDMIAPLRcR47bVZ38JOWKJoAih0yxX/yrfR7UIXCQzindoOrjbBwjuvD8tAEIl
90tGr+rJmlilYeauKKYCfDj/i7OAi4CpTkHokIE1Eb8Z4PjiWo6UuS3OBrG+Wy1QKBeRUG0wxUYu
cPO4+HejGHB67A0n5/kd0LkeE+LAoeYAEKwJp+Hf7gHDM72yZWRJAVsw41TeG0fV0VYeCy/QKXbJ
tWyvTVryti35wAWlj9DCl+lcwxgXkWL1zunliRuTb4b66GugpQEkoI7if69cjtc98ZpGDKdIF1h5
7LxmJkb5oTSjGv/XDTQMoMzwmNdj49X8P/NM6oTqz80kkTHSexejGgAyHtUO4vY7iEmYDcisQq/t
RHP9VTy9cTftK0Fpw/w4JUoaC50Q0UWAyqpjdmzoXKwmQmJ7P+ifEsNCbrlGgpQmArnT9OGeZ3dK
Ip1Y3j010ueniX+dK0+r1+ablADucxVANGWhTgjexUyFfxDmcVMx7eXRwDzDsQMVFlRf1QWUdvT0
eBt96kRVCDTL8tYvyCG0a59X8L2bT2p8vhUgX+1QdHWYK5M0CSXHZV/UR3peBIUeUCNGmaAaVvQl
MFTWlDEEA7tkMdSy7+zYZfoUGcyaR4+7can1g17YkYYgNkzJDHXnIKfljKMKgMT/ZYo5EoqzU7NM
ikYhuWu0BZdnQbNDdELFd0Es3lcrh0L5N21BOuNXgqIgp4BspNuXSBC/7RZzIicLK57IdAKpMJjt
1FOEBtzB7trr0X0Ae94Buc97jCa+tlZ6HUMgVXVHjz/5VeI+yV497XRjC6UZ2cWI2J5wNxi+4e5u
Y0U/g8NLpoDhl5VxIpssidebxdXzJaL/rtnhFB2TsDnVxjUXAdy9p8Cc3ViAOOZ0fkX9fk6CeJ9j
o1zepZ29DRmjU6yxsi28R4kt0laqp5C9ceZqnyM8q2jArH1QDHU6boqsT3g7dQdacYu7e63NAqoM
u0sk8tmuctKBY8W7L0YehmmdpMlUbMmdeIMLgwDWODMvob4+6wbUImf18mi4mqW+eqY31Unn14NK
4dbu9XPsztoXs8mayLBo2EHhHaeN3ExHqldxzx+2uH1h+ggbh8Rb+NilgOKiij0959hHevnFHiRx
wennmClAjYXdIFp+tz4KOsn/DXKWmEGqcP8OuGOOZidgncISgq0HdYXxAije70trJ8co52GirIfl
4+kGvJ+rSyJsBNfqOz+rD0PZwg7FnLbHeMvBQMlxnzLsHIpZ9HLWeLsEakDf2JRtYi8CJL7XqxJ8
uAD2TliBgiA0TFDk0SN8X2JKbXcS5H85RW5C/Yr8sYh0ct3Ktf73FhGukVcyiPb3SgLsHm1Kh0oD
6gVDxc33Ef8ZgGMU+vYLEOamG3HvTT2US4GyHMg0MdDxDdRIsEoIS8QoL03MV+VeT57HTIXQA1hE
05s5OjjZGlHvznTv3C3/ikqsNgv1dwo4GAO60AdJeLpoaBegrUv9Ze9RD4gg7Zr/KSeahGL/tx8p
4sYop6pC6npdgrBcO04ZGw8XelFrxeuzEKeV+Y9foBjtTH3FuZrl+fepC6s4qy9o/CujNIXtEAKW
ekvHhiCtAjA5nGPniS6tYBf5RJiHG2N5VSmNPQgmom2zYCB2tQ4nVzh5CfrfDOMo+61mrAI5gQKq
Iptua1WFOUT4E2dsyacFP7zUGod9hq0uixBzicFWEstBhzF0L4qUOAsE3RGN62/pUlv2FTN/1nfl
5mURn0PhCT9kiD2M0NvXj2U308Dtq27H1LjS2ouTERlZ5V5Hs4DA/SU3JHeT+GAF9yWvTyi3LylJ
CwNPK5GgNKFLbntEkWUkVHE01f+cr0Ukx2TsuPj5jaa6mI0f5GA8SpNHxZsTaIHfadltgeuc9KPK
jp6UL3Fp8Pk7j2j5K43uS+yATun2jao7KOIue+zx/7YrHDHFcV6gI658j6xQW58fRInQjTMo9Phd
aER7vZ/MUr1kLmgbnqsxMw23NFAK3LKqOV3trXON0hK9Qie4Xxtl2iHtlTz7sb+GYgjk5wC1cy19
E/rIhbJ0cmwRcXEa0+FrfWOy1PstSc1XiAg+7cMgioUHf+STsWzTekScZO/0D031lj1ilyW14QFx
OYOniYw4dDMPVThx4GkjZdmGRXjM0L5yvmI7Ek19RIwui0uYFdoIBYvJ/0LSTwwqz59aWnxy366b
qZgSZ5vSEY2Fnz0/qewj12mR9IYBqt5zG3VnBXeC9SaxXM3/qsmlVBU2Aa3kHdshiMBIuOdcSBT7
OP8ps5bFwzykr/m/a3qjd9q73f5NgTUPJfnaFeQ5Ary0X2SjgP1Hv2NEHe38dxFk3jKv5gkrcnGT
J/Tu4Q8N4ClgpbLPvaf7sA9e8xBcLK+qMJK4EZlXUgLcSVKeezHM2CGUxwH2kiFeHLCEYpYowpg0
6ZmOcTgUTbwrHv44GDUrtQHT/iEZbZ0d3/Zn7O6sugSGlkXdxir+lUjNaFDQUQr/2TLNvV2414MR
LcUZPse1uc4HemYP0ipGbSawPhBNn5+vSyML4iKDThXNreZzkjmH9C9peO7Njp9l/wmO6JELo2f5
UbnBwOjqLNvN0YvuC7cnpMfEGe/Rf8uYSf9R7PJodhT08Hd1dQPWzp+iNu5bFOkfz9K9k7b2Adv2
uP00YZhHOVSu+0KCjjo2c0FixnRYZFDGU/rYuXAa1ufSwE4v8eSM1t+Iv5wdUCJPgbfo6dZtcR8i
HVhjg3oK7g2pph3lBSLHeLBss2Ep9KeBeIGdHlrOB3R9Byn4GQvCJAwegaHhhTkd+R30k0/Zk1ir
TdzKbMvy3fq9OL0JQYS7fP76ZAujmV/rpQl+PfUTxL7EX2e04BxR9ycly828ns8UPeiOrkt44/Vp
VQ+3MEM9AaITv3lvTP1coWkmTwVbFQbhLCvVheoR0dcQ7DXQxQ0y7/UcRZ+n732fetCh+5zv7NQi
IFQ9sIPi4Ian+KSEwap2+R69DfpJpjjTcura74OWvJXi47fKQD5mra2digF79bQX7xARY7C5wF4R
wDy6ycKqBeXw9TUQcbiMQKLNw8PC3LjxO5kAx4tKANq0n58qWP0rLnedCBP97ly3z6V1tRl/hvwU
TNKALrlq1vJrVHjk5ryaMp6yEBJaV+MLzDwRTIGnjRozXLY7lrw32Rn705aTB2tCHcGNTfN6hZmM
aghg6LB9YbcwH66MCHQ57YiweJjBS/wOTW8DWSBqDyfeGaeyal+Mr1p444ymPu3txASzW6SI3F3b
9Ttg5YDCew07J1znV4QWuurIUQQ3L0fGcyDd+0WSf2HqVRShM8PJC4O3fFtZsVpJBr8lrJPfqRIl
MjTa17GQOBB9MXaGBUOWEJVzchX4x2huFfMd6En2nP3MYroS3r7oE2jQe0OO2JAsKndSqVvq6prr
z/J7wqCuRftAhoLjGSTQ0fT6ulWOfhHG9snUhvbYeD4guqPRlbB+S8DFYCGJfdLGEsAmwlY4l0Hl
KraBYfrfTt4Bfy/+d8TFEXM9X6vkwchCfiv/TyLDUgpz1HTYYUJHGDQCrc/iO7/kgzIBLy0vOTW5
HD/VIXvKhDXWVX1F42teO5+miVKOXIi0rbc3zQjYX5zoLIue4ftjs8NpnnKcpRSf7BC29eseXZRg
YpGUZiSibdUTddO+fEFGChKAkMoUx0KT1yi63s5dS0vUYVGFCI/NpBF9xU9KCMMl76rs5/o48ocP
XQBxzvphb4Ccim+jSbviS51RANZ4qpS49O4XFA75YbF3zOw6NPaO1EtNWkGb9HE+Dlf9LUUUH4M/
cgtwEfSnJeRJwXuNNATuIhwECoQ2Ra0kluy9ELX/LzD+nBDbajq01so+U0VxcHfM1I6/31V+5mPb
ZTVzg8mNJ+Y1gtUTW9G+MG18s1Fu43ITXH6r9gvNInB7R0fXfooxD1a3Yxe7IgtXgKPb12EJDLFQ
s40Xc6B93b47bC3S7CkV1/VMSUB//PbgmnByl8k66soVRkLpMNKvHq4GXwSrBtNBhwa4eqFqcmdq
IvJpGvIXtHkmtbeWhH2cMaa++FhAH7AzTGHnbAKaBbHrJFS3X/bKVSiZVJtgvpqr7NPjOV0odjgB
MTgrWekXBksT0AFeSGn06rmhJl9pCQHBZnY8mKFtha1i7G0lz7lMpYiRP/vNL0R4CJOhULesSZOh
36pZk+QxzIGug27OdOHvcPTH3yxV/Bh9NNvI1r5nrbRG5T8UH11qTdRDzOXTiTKAxBfdoHSsDFTX
+KE2mg9sAz5ADjkydHaOJmCPoKVGCnU6RkpS7wqz6sSXiBhywxENnezeBzWYZPVgnCRchHz0P6rL
tFdcLIx6UlbRoXY/WqMuua8stFxBZDjyFAI1g4VJaNYXwx6c++bssz+8XQr3vzNZDiLZSahjHPoK
lwxHctIICUuMg/iFCQFEKk7dYZqS4LBBIekYNJiFbH5CzKhjvIo8yXnV6otz4HQZ8izGj8mNR0qK
KeQEoyggs479BNzwGScxLMDAN7HUJHSRE1Fe5nBmovZoKkFy8mwlSg7Yc+51e8lQ+6Yj/EKs6upS
SejgDllTP54Kv0u62fVKb/PL9x5dbyo8GVFGmxqZNQruJuLlpE4srzWLkgV/YUZHAQ6PaAlxu5tH
Yohr/rkMaIe/0wIMqG5jjkyI61ioIgQG9nYOnzTJDamvoi9M6gPkXqeg3nI5cHuFXPhxsI563WNL
xLuqaPei4crbWmVwqWXHBw+GAUDhgH+rJmxAD9OTXrnIu49aZUWl0qdfQM2BBZ5mRb8Ztt3SwQwn
gX1+q4Ur0nC8YVdbDy/CkB8bNHIXus857SzOCjnirMR9cf6TqW0+0uTMD5aFeGP/rADtQ/LZamIH
SItCUNK1gKXQqlWNAg215hmv9yXzaS5ebXRlscHZMSHId8qKRw5kdwLsPvhJf3XgEtqkDTVt9IX1
xXJ3ovLcCx5SBl42OJFXzQj3AIlAjbUmyQQASQmFKs2ymULfPoQhefUdU9cufvQKa+TQBMWlyQaR
Jw+q6WbrA+yXApBcN8Q/+J+GTPcEPlNxDAhtNZq61FCImqFMe/dXvTgD7jHmnb0gR7OWODIpAvV3
W1OwtsamBaKyw2GQqxf4fSrXYlMkUdVheEK7Fch0HxiF7NN5wU/OWIGG1d7uw1fWz4FUVM1bV8ts
9vas63fXoE0o3z0GT2zJK0rupZV5D02+4jUe0YyUVdnK1RpFznLwp83ioklJw+oVPhzwqr3o5+/Z
QHjXP/uRhBaOgywwSuJFro/XpBUGO9LhWy5sTN1vliG2EGKKRcbA0wYczEpk90RWa8CIT2TxWXO+
sN72IsVcqkeAN0xOdTDMcFa7MGtpS1l7pMmQnr3y0Wf4MTnFYr0VMzwztn7xyjzZ028421DaGOAN
AenHetkFDAk5Y9BuIcrqBblP9zNVZGVwst0RNImMXrA069znVddRPdVLzRmvE99qd7nqlj2bMucb
BKFpJCLTk9XbUAgmfZmguBrwjwDDgJp/XD+xWOeD6KutIECCaMSv9c7rHrkp7b9FOR52vSYzRL8p
bSJkAIqiHTd7I/N+XFnfZNCMwkJ0/7EfYRdhCuilUIA1DOUxNpvPX/ceJaT65RUfw3OEly7of+cu
byUPUnGyM6QM8FZvqsLkZ7MoUsL69ehabJDzyaziBWbgtkl53FEUrFczaj3/V8SNZg+o9Anc7AWy
yEZfgctLIeG8hb/N88CEPp03maaW9TvM37+s3CqKGS0KtntebfZsm+G4x6LHQ4TIBDaOkz53ExMm
sEPlTFC7CPsbm+Uo2r5skk9P9oWFnVlrBwdF3U+XTxF6MgRUhuOX2AoQ2HV8IPtAmsnHWjc+vkQK
rqzxgzAEZQG3lyWGyqEg7DRlbuc1YUNHA6/D/KycGBtw86OlaSy2DmApsvzQiHaLG6R1WdAWVPrW
Wc/vduxsSqOoIHUXJr+JZcCotVwVbNWNqOCHyrSKNErBylirU+G3hcqgODNdTkH661aiJplPIZ/d
iiD9onxamUsFd8De/lgzcOdJ2vVSyQ25z5rbeYc6jQwqAk0mxTHfDBRi3f3wfZB3mTdSXB84xlci
xQNUe9MC9mbWxiYWAbaDevrLRxK+fKqBaoUPvhD8W9OoQ3hxijpvMA6eWODQJ7fhp0mcGFogheVY
NRR1DGBkZLE4gVl6tV5gPeAs1nZWqc5St7Wa2YLB1uz75cB+ovM0LB9uh+sRPwo6stpi/6OKGF1k
M1l/1zXL6fucLjdrrGusz6zerTpljC8w4+4lR+4qpDwDQXtdRNXbiygLoYytZl/b+/EBhlEuEFjd
NCqlU/jpwUgfeKMpr+I/ZZc3qyZ3MzK32kkF5udC5irrz+fHy2M6BXQ4z3bz3K6dRA4xlgYVRNIk
iWJMHXuEkc8CIrWK27MVARnM8CbTU/xO5pV1HP/pNHIg8CHAK9payYX3HQ9mthNNEur8axh66fza
USRnhYAlQ7iqEl05RvgFB4F83WXolZUejd7Zq0UGd8c5fuGPJZ/5f0HP+ulqEHQ2Q0B08AO+wAYQ
VqnHg6aoKd4lHdeGe5ZPdvtptuAYnqF2cslV3cRg5XrTwsDquhBJJcGM8ya76HkveMZatA91oVuf
UNu1mx0r/TeCXnNpwZVfMz1D08D3UuGPNfw49fVBDFYLcTH5MyTkoNxJKaaB8oQwHUfx0jV1zkNI
uG5xuMD5EMdesc114NBibzwYlh4VzyyxNNpzDc2V3WlWxCakswfNI9SLeDDD/mfP4jym6Qlitm6P
Ih+3ikD2l/F5qJVjCkhu2R0YuWUmPriMOI7ohOTXqbYI3lND+YkNo8QEdPRi1tkKymjdpHC4sFFG
zIy0DHpAwoIaxM/iuhUclYuo5xCKI1PEF8cXu+73yDZWT41tGgrJkKCnV9ywh2CPb7FlAE0QMQ8o
j/PnVO9JBiRy5XCbTy2JSUN6VhUl2wcdpv++Kr0lP1pdWyhPnYAMO4urErzGyhjC5Uj8ZvQUHMAS
arV67D+1mQtE4ZBFqLxUKx735PsCM4RSk4hw7ypMAhNMuVYQCEVs2leqYPUgzGcKQVBVaFA/Irp2
yN41eOaRz3xe5ngdEsfdLZ/HzPTvDfnsmweskL5Fs3on2SR0Bl3qGqqNWgTTLwujpxCUpXBIY4TW
oQ6JeJoVG8vaEiv6RmQEzdTP+SKNMqtrxvDPgc6Nq9isr6E6F/BhSNjtaHAXvTxRRBS9LynoVuFn
wtUyPZi0SvsJnffSIK04euGdliYeHBoQJttrieDxltmIlwv6DhTCLE5fsHu7UaIoff9sO2A2XXG0
EFWNl96jPyzSFLWzfJn4UYjidBRkPgBhJsUjJqXtR6a2dQZSn/Ckx9VtvtVoiKt16Z6jx8UCo3M/
l1Sw7QibpkMA83fYmwz15TqzIyNmx4IbatmBStYISuvBkKZBohY5agDuAlI13VJJyhiEQK88NsDt
HIX0nLqRHJ5NBbK2obOHnBmcBR4Dh6BA61EAAyiaswTNZFOQB6NsPDYDyzxAY0jPx2kUv8JLmn/l
28BDzNwj91wIEGfXRXCJ5YnENywmR8mwzfgHZc1fp4LJXR5WX3QAkJ7N9aZZ5rCWj4RW5ZyGQV/6
hy0e6PZLUuS1KwhqbX5mxk+Iz9RuzKHcS2BwYk7zqGKGxCQ4yvGlQaCws1QshqkOeEuOR0os5j3o
peAjbUYjSvs65yVo93ezydW2ICO3eSqKlltKzu8FUJKa0XY1LwMnY10exi+qhbITWnfyPi0yfryj
d/5AaiD3u9qCfXLssWSVXIKjnlUQ/KusdxY7NvWgfgIwiLesaYGjLngJD6lf5yz0SngjVbhCarYj
vLL8Q+7s11rY2MW8cIp1dqvGPoo6C16UmYC11IJv+2M+NuGc6R8d14Dmdln6LTESZ3mB7iCmLcS8
Nkv/YdWqsb8K2bmnp7OaTKUzYX+NOYMF8i57FGk3/U6AGnt1DXA6pgYRW4bM9IGLa03Zyf4+yArp
pTSUZvenMQs/KIokENHJvg92akgiBxaQ21RxtfyK1IMoD0gxNBsNNxx6GIuqC0QzSZeUFxz7Hc71
e58OZENr7muMgxPHlziaPiiaAK1zBCGFGX8Scl9vVPDRrn6sCtTTP5IoL6xu/kuU2UNfAPovVzmd
svrSOmYGbRRr73CdQNTESNMnH6A3/mriu1CDyAj6xKY1UfuMpEjyp5MCJUl3bqagbcV8zR2xLeJR
E4JwNUmUwTf5t2aSv13PEwKnWOkF1FN+ehyI0svBNQ6oVRbb7VVYXd1crB1CiFg60rofuK5GVccX
4PAaNKMjk5rGm/IWNV0USBuYjBWleE1l48hhafQ9KiN+ORcqbH9aoe/Cv50Q24G52Xivd2HiVOdF
odrrqJBZj79VMjbExhoKnD6JIivATFwHCaWEvL6MebipQht4swLG7AFfn0H/cAY5ECb5HJSi8NDl
BhBRw6qasmOiA4YONbOzEs0DTpPAdJslIMEY1bJwRbuvPDSTuxzPtjt5NsyY6XIcK7NDpoLnjjE1
cHyHgqHOk1yVVexO67kLJsnryVkzREOb8XPj1QnbI4WzYIeS8ThKvhFXoM2GTC+xhrAd2BnaJ1zB
7vc0VrSVRoGxKmdZ5gaX/PznDHwIEhrIRoHH4OaET0srVRkuiqoRmlQdT9x66chxSSL4Fsb2/YFQ
RthKLHunaRlRWITwSpIR4xRN7GOIhlgJalc+vll6Jzn3/q8jThx0ruDmXBnhRuCJ+3K9dRf79Ajk
yoELJDWZRyUGcrhG7ZYwvFn8dkN/r2KViWRfpKjZgmoViS2XDlB7MqEDhI9PV6VyYwrQA3e4BnvV
BFCkGkzSTVOEjZSZ28I1jYk/WBR6c21EM7yg+XPQPf8J0W4p7HkpeCcIfDSRtYXrJSSXwROsR85g
SdHF0ZOjv3VYsnVgl3bZPRuxDF50V6OG0UfGqRU4hKHfI0DPrwgvF3lFTHz9BJJq0G/3OFdfEOuv
QKNCDc8YI1GoivZFhaO4TI4buk37Z2k6bFjIsXKU+UBgFd7nkc0C4diQmgORjsv0Guo6r7bvk25R
VKK8NCnoTL+w8UxDkTcwvKdXrPIqrZuxsucFEYNCeiwYsueM6A1b/vtyMuEV0RWjuuJH+IjlBYeG
KSPzJK8oorpe9JtXsYzHLifZmVgHTnt41B7OLQevTFsWf0F+F6T+X7gOBHxRybh17eLZW8iFj0rY
Rz4rjY/GFQ0BtnZ1C4KRtB0K+yVnsraFJavN5L0MTHYNBwK+j8FcxlubbSQIaI6DmeB6vMWhUxvJ
SyayOrIoKLGY58sfv4YkO+gQlScO11zqZ8U4okoPwXlhKc3+RBbfFF15wFd/2zu2zZLxStLSsPxy
zSCRdZcwzJSbJTTJe1OR5yyTfyC2Jndqfd2dJRSmB/TEgQpOmse4yaIuo0qOGQwIGZsSuEg8ZrgQ
lXfxDnOYFXfpBB8wtUTpleBdEV5e6LjkMXzq75pzHHxQVjK6IDrE3APBDh4d7LeAW5KB/rAFaiIb
GFCEuJ4SDAmfCOFCjUJjTPB0uGBk16CGka1XKs0Ev0DL7K8L9msOvLylfo4GQbML292fWCtUPN7w
6u9bG8gpLkqFXlKtUfK7SAqlRUEViO9AJ/W6sKYoCiuWI32SFfnNcwM397UtXk62HWPjOENsiMRI
Dr7XZzR3cRT3rzXAyHDvKu5QfId3/bnnPRLpMo35NFOHXdc5GhUv+QCeQzhx8eeUANyNepRUKbn+
AOxiw93CBdsmBW65fyrpcNkpkXLO9Djs2B1PvWxi35iWAY/KQ1KSJ206zua7mFtJAi8UNuRTKsVK
MYL8nPJtxwjpLioRCzEkMZtzqevoZ53TR7Fz+5VWOXgCq96rAvKQDBIuu7H+zhqvgAvt5fEBbAd1
Jy9QBcDzDC4Fy5HaWGPBqA+dtoWqi8r8sS0WvuIWrKDPjlJbMM4t7MyknNM6fNgRLu7aqJvo8dZv
GkNyksDj/3OMSbvzvUX6m8oaJA68Arw02uIjSDh0Y9kWVOrbdmEXVKLK7p43l16SGh2Ae4AlWDO9
nv/NXVJq41WJAiXSFCU25G78pbmDCXU5wKprK3s7W0ZkJo8fDgkBtSQwOlip7uWGhda37jyR41bx
rs7fD2ceMw1+mIbE9N/4WcSQrrZKzV3DO9Y1EVsz8JMlb7tQsU2LLjI4lbR781aheNhgnpposzkv
5ZMc2MYH/FfvC7pYcoDdAMmYlxG8DuNTisrmMNR8y+yIDt1P5G6St1kxVnzz6HTXQESiyUEMi3LE
bASq2MRvAMJr9ndz683+cNX71OgMe7NHhq3gEd0t3q0+yzEt8U1Rg6w7HRsCP48aI7CFlqo5lnMB
B5/7QRAaJV0nx2L0xMb0UOagn+Qwj0U3g9cUDllWUFZxiwqmTLmq3mfXoIzpQl+oqAFdaBNcxKJr
Vrp8nalnC6jSJe7ChvaUSdaFg5ZXTMb4Cu1H/5bZuriDBcPChXNTOF+B7kkKDmvaoXyFl7+EEOPl
C+K2A91j8IXUHt87hnxT0U/hkcwSruo4uReIE+JQF0FcIqRWjkfTteYvaZWSJNKRioAyWyS2DB9W
fOEdz0e4od218ZpWwlvYk4RlLbr5TKZ4ZblTyFydotFa0ARMXmVLoYbB/owsb9WuISQgbW1ANIx4
WQLOotoDxmZy5llD5i0O/4l6VhPMWEhVuVFm5eHJgiJb1I9Tdcu22hk+vuX2g2gpm0YIDGOVZ9VA
mvGA/psCYXmHtNwzfp5IBLWu0b8OUJ+gS/LHa+NrMkRdPkd9G0yRnkOvrlm7SL38vPJXBxDR4qjV
nHDtnQpGzwkANX/wTX/cxFTj3o+LACYfmyBADxhWONsRtMt6cjBdG1qV/aokiZE1KOSHjLwtHVHn
xCEMgoy7CU0NVyP3si7/S+MjbpHB6Q2ovVwew3sit342T6HnOfuPRzKtGw3vDYBnKKr7GD4p9pH/
F5T2NgZ+jEWphr4yxIkXXeoP6B32et8otoukUW7cQEs8MxQLPWrWE3CTLYODw8G5265IPPz0fNHk
o9t1VDZvGRDXxXw44D1HKMSrvItYAysSUXDcXCK3QgSN7XQ5HDXqn6pNZUtDspGW+XfnHnmNv879
JJlc4WKnQj6KVYS0P1f2YdiRJm+RCCMQ1Hxw1ZaHbPI8doarGPG/BTBY6FiOQh/qIVQ+7RhvWIxp
Bdt0lI9uROxAg1hObpTqSIT0zvOLpdVofnen0gMEvNoxcvw1YXINqVwMe6r3I9R64Zhcgdl+06Ye
F4KZdb0oxkNTU42cOsGjgi+jBKRGx0Prgo5iKOKC2VS4MkKjLpc6IV3qtbSac8mLVMND1Nv26g+r
tY6RLfjpadqD1/BErD4Fe2FtYhFoN6w3jyfq8FUp/oH/nhHvtx91Ko9PoN++Zc0fpOkjd3M3tyET
VtFagW2T6lYZo+EdIi71G3DP9wX5x1+EzHanykl94C36p1Mmov0YVYppwUbKtMXWFq/rcYWZjqNi
uqeIiwNiz5AyZzHC+FO8AQSPSmiLPvjDS999eujru1PUNhZpc6fwhTNf1lqS5DEn/xcS87lJctOA
sJlvwfK0I63gSrWjOt0fdLUzYVlppHKuokKwySuGRkQnkwLqxei6CHPWR+mHIy5R4wNtQah9NXIK
T8MlM2AOt6YvpSjIWGniTfc68/QwKzJ0m/pzsljHVOyNolXKT0t0q7U2qEl2VNPVUtEpCRhTVQRu
+/gszf8qfujZhHYpALIBcbpBAAiIN6aVwyo1Ok2HrpzATwJ8chLGRFNR6NnDIWzaX2/d9mcnPGLH
yUipMcZ/X3KjT8eAl6d6SNnk4SCFFE/tqVHi4xG+IkgfcXYbwKicMYOm7aqEjYT5285k+jv+z+Zd
AADeADadaWz2ul9l/0XPFHZxEjrm9brXQS/AU1Az0B8vbPXPreR8XQQGNfrNdy4ytn0wth+ohfH7
X8viicadfOgMtaOtf4GQlpMLu+Qs9eW8R4mDjt8RFTiJPHQY2Ga0QBH+OaCZfYIVlsJgF7Ruu87i
RRnQ3YwnFybGyvR3jJNqRPYyqtPliht3Jym2GH361aU+vyYftCy5W4cgSdzOr1z/WOa21F+YNxg2
i/t7h3urJ2viQmnNYAaJrcuXHiUseklFM4g7PGytG7r05bQ4i6cBCDT1jgtXGu0n7P/qj9Ydc5Iw
UX1DmGVmGesWXcAWeVUC0iRYK+lkvgCoRMjl96hHaGgCQb3faRFfZFrrzQwwVSFBZmm7DoRPgaRw
cgR1Rgu7Cnau0DzgbnlbMiiLY9O7DyBevHMWk0IeDF0fiURf8JQk8utWLBKItCWGLa9MTTuNVATC
oXGp3Ufmhcg/ePYyELCd47fJ+GmJFke9VplNbWLXEdnV6cNY59MHoCHGcVIFO8okik264tgQC4pX
7ZRRUqdZzedAx+PhAIHwGlYI5/ie/jJ/RhwhirFXQ0c6YEOmwP7gr0Qd4It201/m+hy9jlbZgfnG
qM3HzVoVFFHqKUso8TmAYfFk1XsWOPnMEDFjee1gbxIR7eB+uDYmz+WpX8IUblNH6DIDVtFfnsng
wlle6vA70CrZKLMQ/MvHnvEIunEdTSB9ZeeJ4R7JVy/5UxanoLn3m491HMXX/EzyUVr207lmHfxP
yK6530h7Lqr7HzrbYkmdT7FyIJOHbbkfMQASuCkW5n7LLapQ97UdiVkCyFWs/aOPmbkP6yObRjVv
famCOrjR0DGX6dB1CHuv4uuXQ3hRR2tesE0wBAvFEtgthQGAOcZRQ3yDA66u6RWl/H514HlwLsV1
sPYSLeo8hjXOy5xRXkwn2qk0DavKI4k6OltxyHf6jk9B++MPLBUSMhqCeciaG/YbYsF3xPL5+Gfv
mZG6y23oZd9WR0Jgk7iP7zZeWhK4LFRbkUplDVp+9Vk4zwRWgGzaZ/MnOrmdkM8rfw4ptlKwxgxN
BL7jrC48IT+1sh7KTkSAqj/UmpAD45rrb8e6UPj5S1liIOOgT3UuYVfrQJvBbxQ6S3Ss2t47+Hzv
peTjQVa6quk5k713ocSvmXEYWEecZ1WgZ2KxFENSCa4Tww1EeogfzKQtKYyGwiY5d1ncvMkXMa/d
g+TnlgFstyR+UFGzxSkkNig7tBAbL9ne0dir/PdwuUfb8MNhrabfdca+L4xcgof8H9xzhcvtTuCn
ayGsAkgGu5Oq6Mmvaw3s1x39d7Gql6xMqyKcGEqrbhIle0ObaJ9Y2tmHWp3pnZx/Iuab3SrOvw5p
r4hdVJmtCrILIooAEFYirtKrgQhYts8jikvwMUB9wsgB8siBKzYgBpvqT97ryhdSUUZOGBWL/Q1Q
UzyVn9mOfhzbc4UMmhbukw0LU82wlBjUr1xnMAkhmEl04+eh0krViRZndf8t5+1yPVMHuc5/DVvj
mcxppU/bbfiZC8p2NmJ0uM5qlA+96w2ByYcUiNRSJUCCcHKgkut7SbJobmeiee/NFhTX8PKZ7E3r
Ue51pbhZW97QA3n6mNrqNpYeGA6cvqPlWdlIxrmFQNZYBrhIBd5ZmC4vGMliZU2pifK1kfP7Njqs
BZ2Mxe5rzFA0Kv1zXXFM1DpGZEZYmXnQs2DfoqGO/QqF5fs5mkORfSYyebxLkjZh3vSAHQPPVkrH
N84JH35tbdmFMf3I8eFQNsVqZW3OvEVW1fzdpNrrKvOdD9ofCFXNiNpwtyAuwapgds11GYFt1iFV
Fn3/chBNgMm1FUbfUj/j2aIk/sU2v7F+GjE2lTZqMoX2hnetBiPGpFp+B8jksQXiUMCh6prBlhYs
O18NIlBsjBXIJLs74h0Cw+IVXQbh5/wN1PhSxIZm4jurszccbfixzdtcxqtgUHgdf8KiDoo7Nwqi
ONLFw47ZPFCaIgtc0E7Ooc/zZQFM5SxabaEHnLZDIsNJZ/msbk0YzD3A4kA0AoUBGoWFkplraWEZ
grvPa5NLsYthVQnvWfYsSJJ/zuWHqjvwBQCEqdr50cA46yxEevLpaLPP2/JUeIWKrcybCwQf8Gq7
bpbDZ0nLOCKWLz2XbdkePIVwvntXhoEZpGLb/imX23S+JRB3GKyuvdRXVSC0I86CN4YvxDvr6FRI
yzxxL4JpJVdx9nEyyjlRDqS6DuDPRA9kPCkc/+7f50MMe/lPSMhsn+Ik4hmaYSC7nBr2M/lLW8q9
4mbXbgxoLuhssNCpe3bbla3Qw+vb6FEuB7Zloam06A3TJiCR79PBjWe05vPaMrXOLYplXSfQBtfk
tzTmLhZbZpNE7z3KuSdYKRci24/V+x6lxqsLjj5DDonCENz5vx4ponFqxBLDrQ7cIQbQ2QoA87Ks
MYWpExuJxfnklWD1TJPeSLSQ++XU2N8DVJpOv3Z8Ftp7Myfd8+j3JOd1VHf5QQkLnkALJDiZUIwF
2KqOPJAXZQgZa3pt0IQdlhxMgEQa0+dO7PLgAPE4q+KXEIaxBVL1fPa4/UXBTplus643xbF6N6Wz
Z6jnq1fom4PZNq8wcoDaVZB91ix4tH4JFGwaU1HvaC7rusdOb6hpbZhRD9Aj4j/XZMkNZRooBsgN
IjN17FgRMeMF5vyARZzhOAjCtv/Jt4G9TFzNizKNJEunnkZGHxImrHfszhQf9muXZYPqyiPIoAH9
fCIV69mNEEWcGe2jpsinJFy1fDui5YnWVMshYo+nRK6+QiKGsUJ6mnwJkZ5K7y8tzm1vIbfaP5Yh
yHKhzbeGn13dECGai97FB4zjs5c/uapK5uat15Ak4ESLUO1PhCZzZHlXqYxr1qbM4xi0EC0gNqb+
jem5kkU2PBmIxU7dS0710RNQbYBr6DBDrSs6LeqN9J/zIxkms3MRAnwCJ7IFgZNM6fz254wH7Pyr
4ZicOjG3vZj7rCtsyBtlkE/pb54csNWeQfZucQOmbr9mlJPlgcMmblUoFo1sQ5tBIuUOpy1QMt/J
7R6LTSvRQq+5j1hJXfSCyMe2aB/vQ1ohEBprV2QX5vYuLdhmJ7KGW2XrKFVomhFknr0Mv4DQDDhK
J88G+QB4fXASDOjbv8FwP8DIc0yEFClHycF3lOYp5U2bLQQx9ZlnvBPd3nvdShw9V5pUmMwEVoza
XHR03pb6OGaGpsAPewHqvQCJ2Joo0XQuPIwdoUMMaNRrkibINzz6vVPcIm6/HcTJqKMROiYqCyGV
4t/9U13+u5vLG2TD0Wwt++qXaZmP/qfsPVTl0B+eP4blWBkhXy/o7xbpoG8uZVI7ApvhCCxVuFCX
7PnUankmsgjvci2fpfKs674dUsCbrVkdGjJXQxgMwkENlKEWLpGrTnwNpY0Usb7SYuRU6RpbvRgY
2sOxi757qfkbCrrQJMa/twtHIWhScZzk2UemyQHdQ4ziNoP6ilVppafgmUT3XpAf+FWj+2kTXVEY
NrPkyjKV4TxIbBUM4P9MjAIx2UiyFJfOkeDe8lQCZwpRt1cwYPqZDgSWQKYWJgn9TyH5rM0SEcpL
H+h22GEPDBu8hf2LlBNo5g0F7ZW2goIprGjatOjpqKY44mXYmi2Yb3Y4RMU6hrRI0kDK4KYi1qdY
Ky/0va3vQPsXHShE5x0K2l8Tb0WPE+33bOzqF81ZVYIIdsrTjPl6DpfC0yyTHQahHJv/mwafqDgn
9BikB0rq3A5CkaQKuqR30XTixohafN43UVLZvogXtRevE718KC+aqL9l/1034g2KlYXd+NKB5gL9
cVDJe56Zf1Hb1inmKja5OxxZ5MQNsu1BG7JwvMlyEEjup4Re4mUieDHV18+t1x3brNfQ+jZm5Zpk
yaP68K29+Rz/7bTQdkH4QsyyLuDu1d4J3Wup4lb2GdTtDNcKk/vYGGRNl9VtTP842hkXd4//tt7S
NVyDczT1jVfqY2wXRlazF69AmRZjFbpNwm1KFMHi5VAtcPtWiuImFL+2teRUHCjHcAy9DIBIvHrC
FlkgYvZkMx28NL9cuNvr+WAP/RQRrJWG1y4bN+w46zKPn5mL2womJSJoKxmsUgRUBL1oeK0MUgiR
yq5PORay9+8JRWjnDn76SJf9ZXMGEs1hXMWwX4LiJPNb5hS4p3ODEuDitMRFUQML0864gMXQDBi+
Dyc1Bnl8l/hTQfpWbeOXKhMdj5Ha99bnUdZrwQseNRuNliKgSClseSOFd0+Q/KOljUXBeqZkbZa0
dWvdM2e2upxADDkmwqyft9R+vpp554Yp/LTsPRYTWliKcsB3/A4V5mrNBZIz7dMuWWnpA75T4QEe
+UThhZSodtJ/gAkwy96Qyc+jWWhXnWVlHwz95QpYpr0wNie4RVg5lSjeCUsmQQpmb4pxY+UbZl/d
aUtBC985qLqg55wje9sfYHNJvPZcvgNDOIsLQ+l2HFI1Wy6DjuqjpyNZxD42YMwNDD3tx2YP8Zqb
mm/InoqxIONgkEvLzixc25dTEHfZ4h54JYCazc2X6qTnwVL//JfkkcuGHokiI+PnV2yjm6jJMqEz
o1erFwVUFww6UYUR1fYS7sNhGca1kjLHonKClmZgUqn+KTXHjnUXp/0cpNtZhc1SWdjZf3ncFDUA
GzxgdEjANnhb708JhMN+81Ho3eAN78xfLaJqkSvzLLuWxo1dFTwLA6QOmL8eHTG/7aSgbvcB7k/H
IMzyXYhXnYUV9xULr+Rv1K91XQ4ej6aI8rE1vk4iV4URNVuwx/W1TBtzXAidIO9Hgj/sYEI+pN1f
mZvfWiHVWil7A1r5hvSfniz5UGA83YYzkZ/6aSznnIdRt/wVA96a6JEyqqC8uDaPN+GsuOuAcZ/z
f6vDJKSrJQMIzcqjA8SP3lFAagUK4Ur0XKaKBEpHaNAxoNPvGUzth54U6No5u8jKCbYWbia7L1tr
8f67hmtdcaALMUW0qv982RaAnqcmm/cVaZSv8DCZDBmiAO7bK6VTnOOEeGXZ0bQuWnpf3TaFRjQY
w9coPS/wxmtx7Y8DgDbuATNU2HiiE1CDQDOkY8GbIU68yBDG3FmKfOTND/KiBVl9v0q9Gl+JUmvi
cVfMHJzUEzM1gl3+xhM8OGdbmuQnzdNFPl9Fh6UxsnPqqiqtdf4JqxHDMmYz3WZ7toVDXp/+LjA9
4Yg5sBcSHgVGvbky1Xz1FAK3k603nHfky1yeuVh4pbBj2NM6oXSk3rcA+kdSrab9s9p2kFtjETh0
LDnninC3nXpFFrnbzh/5Syv8mShEWSQsPWKd1l2zWH6oSsRCYayeDwA82WN0C16sQLah3PRwNkEZ
4lgV2kXh+wqEsSyWrlWibYwNKZlz2ca0Q44UiiFXYcu0qJ4D8WS2X8L6OVdOUfNIEMPIZABtkvTz
shDsAvC7nDO6ryGPUkHmiZzEWAouFtrdQnGcUnH+2ZTctYcfnXmBB/LufYcvKX3Pq2L0Ci4l4OFl
R8OY3wHcFUv81/gfaAK9bppBqxMp+UJWNMBaHLsmKlYOaSDiu5q9fzS6s000lULWalC2OxS6ygCr
FF7iqTfhnFPim7wGQ45y9WNjL4jWDXj9XSwndG4eL4isO1RyoRZrlArDTHFm5TbWyojCB3hGRT9U
187r7SuUYMg6qw9GYetKjQ9z1/fDzvuNhuzn41b3ucwIJ6o9ixdj2GWXpK62PQCLNknyTCxFLtqK
BQFIhUVUuFVbXEYmS1Ri0vdLRCD+PZHhbyy0m1GgndH5Y3RS3DRjWLyRA6nx6SLUG4hfqe7Rd6Qy
2xpLzCx6yhveOwmPO34XqaQfoTbX99t6PRS+GY75ipFtanAcYCCvzNuhG6i4W+3LVJlbfO9D/ph6
my30+hr5VKMQOJV53Gb+jFvxBG3vH3zep99eKA7Y/2P9aUkde5M2/696hcBDWjfvtZN6PL61Lnme
hrKW2R17FhbjadcidDqEEmHyGVNN62+FuIbQYAmnmD0VnCamvEj9LO4XqLf45MS1n7lfx/MERCNw
JRM15tblkkcW6l39dIjmgWNkWyc/Wn2PbBR7oNzSSPTv3juYNyihlXXRCjmcllhpregbkfMCjc98
TWSPZiYxsukEfvTfVOB9gGKtvuUfUdXvApvrJuBTysMlqOLFOPITs2PcpqGADGfW0HvAutWNupme
ds+ASw0RQ1NNBPM0iAQr7llO/o8zxs17Md6h+GM19eQPEq6Z0Bod/gV/RS2LlJMX0qzbLfqH5dLr
/8rKVz68c13LRuNi0i6NIgJW83lrcn50p9Gkzn/ccB/u8Sm0Vdv6hbbNu4I4RXEtUDsbl5xNVESl
kk40pSH33+sG+R8AsPXCptyJvr9VNgHqbRWi8z6t6xgMRCMyE3vjzWGEo79acQjXrcMy0MyYE0Tj
Vy0r3FYbR3eUq4S9q2QdCvMHjaA/8nkLCsMth1ibH+R4cNJY/Jh8fNRggFvS2J15xjTQnelJynK0
1mvxjdiQ/2Q8qtT+YJ3h+Gvd8wQM67ueIrDwhISucYDwuBgEnf/a+2SlDCZazbD7n4RCeF4KHGWD
iYckw54Ns9QFGiNNCHkHpJuxynpEzOSkD0u93kB1KdzJCBEnhR47MImvmaN3WU8iNXqDM+zVGmWl
hCN1MwPSSN1GrFTDphqpxIE2AVFTDOU2KWurMZO7KaGy+iDWTfZnp2zMyAJWi9D33To4fat6CA0M
5wSCrIGXLI+21Yiz7VPrOv+LEnSmhlfEkGU/6X1sM19+eG21gikoquKxtJ2z94gS7xTD9Ub6Xr7W
Pf4DoO7U0tAUpyJYSVi/9KsJDNwekB0eV3Ao7u2AzU8Sr+NEybmH1CNizBeChgGqucbamN27C/D7
ZLi03PZjwiWajW6i3n+uH3ZCuebYcyDtQww8+/iZEolWbRsksDLOHUq14r9w2lAw4lebkTpyN1V6
dRzaJpvprGfPZinXimJH1uxLqHsAu9ruW8yl8Cy960echPZkZCBxbFdSBeZHO/m6jK+KD+9gcrpR
0MM11dj4usIsi/c2DvgYiD/UpGSf1e0Y3IztnGoXqgH8WBmhWuZYfwCJob0KR35vGBnmfdfGchA5
OqTIGa50xUY9ULgR7nSU2pqhZ4dI92kNQCPwfsXUUssrigBsXlcXO7Bja5MblysoAIPZemZJceLy
6ixa1nt55BfFxQYyJ0S8wp9SsbbxWlCwtCDsC4qfD7F658UtqAuuAffZjIUlHF5NYlEseuGMqwfX
o/4lHp6CbJUmRrvG6goUZ7oScollitzqHQcnq3n7/EHMfHwQLnc4c8HO81RPNs6LGfeqFpjffX2E
GnSiD36tWENSKLZDYQjEtGTSj5/B/rLaPcyT63raNXImr64fdZy6T1yQrKqfp4dAl6BX9INPxgnF
YTC3jQKKiBc2WptQeKjdM9oTZSMvxl1cv0RiP17BpWc8AdWtm3Ii9kmf5ilgj/RJ44o/jvDYtRtx
4TE6VhN4scOC3AjtYQMXSWK8V6IfNXqbw456N8toXF/1v1Pa7v5moJrzomJ4Plainjr/+YARYbBB
gabtnH4uI9boaFl5peizxvfHu0HvOuBWiVn2YdZ8OZzs/J45E50V3XjqS8228yt8euxLKuLk7m/r
LROJQma2Ht/uEqQ41TRann4t8VHBVJdDmlC7v9JYgHzbohlKzV31Z3f/oJF4W06k8UZXbs7x8zlw
SrUi3EebB5nf9J9QnpcO6LL4PC0cff0OOhaisISSyctnzhBLM4EayLbtKhf0SZb6tTllfGK561m2
6mPCEoonb58Xwjsb/b8EyDCQecQY+Cj20WF7dZUKTuLAe29JjM6ME/6N65pifPSil25xB9yNYcRv
g3FjgB+TDBNnSyT3vbZDqwHC5L2200Um85Xr34hTu3fp9ZmEOfD+BbJ8+0gShHU+lfmbZG8Rhtm8
BxJvta4B1f1XKeNtPrYoCwFsYdvHsorTjyG9NEj5sVjaI7b22p6J7vEnc6fe5q0kIJwCM91X3VWk
jWAHjVC2d3kn8QayefeH0Xqu6sQyLH58SMYadyR8tZ2hSO4AtQjdUiW+NovdR4XiOVAWK/Czxl+v
ic7L/uQv/vv/++MtHsxPoCKbqr3p1pk4N9/JKFZyvDnT4TOTKdD1UiS7oniHLnv5SkKoDBWwy/RR
DmOR63y34lfmETXbsnPetlnqmz9bo3Kcew2lKj2aSdo/tE+zzjEyKOUzNDl37eVL5SK4RznGWPVb
t+juvJI9ghcXFl7CV2n/6LKVG9csvJ6S07y2MFWYnOtI0Vdx9oc9nwK/itexAEj187VQCoeJNi46
z1TVTQTqyMiLwKVzj6P2Y7PS3OJ5cRN7oIakGIhvkJi0PdiPq0PCRV/Ok7gMBJigMYk7xUgeftPq
PSlYAX3C3A3DpTWGi56TWtI5EUaL0qX4m8fqTgWhb+EG/hUzg4mYbMiKrQ4IiZIj3BYDOZDdmiRG
UcbhTYVA96UFBM3q1xmla/5EqSi9RNfld+WXcx4493CHqx5iLL1VG10Jo5GLTAbX7XaoGwX6gL0X
NM7nb72vy/PQL+v5BQoA+1OMHQ/pZRyvMVGVWwgxKA0mbqaBUH2DdDOJrnj31BWJOcIgY/opgdfa
51nLNwrVBf6gzy9Tx9Xrb+dsXNzm0FFvzb9yqk+t/WbZnCDlITHk67FOWgM3leQ8xiF3CX/cgKVe
ORqKt4EwPvKnHP/FtmhcFR3gVhCQYb+Eat0pfCzVJ0qu3k07UK4J0Odvwzp5zJt/3dZaKZJc1V5r
pW7Hus3Gt+RHb+xCU+yAEiQSTmjdXrRu0z0VqeQseesaZJC4I3nYXyo97+PI18MVZPM6UmDFPcfB
PQ6uHxbr1XDSJGtpcsVplk3c8XoO1slkb6s4qjcA+GJmVGuTNSooQZqyUa9IEgz1ONC7q/XNQa4F
RR+p/qy4ZWZVuQIpE2ptluWa25LnofvO2ub+IwDcWp+o0ect/YDINNc3orKR+5oiFX0uj+6SmTvP
kxuCz2KOxtw/rKioq3nTM1iw4k/0QP5sT4BlzeCIYFNHFMcKASSpP88zFsAPt6NGutx1Ozn00qjL
eP1SYrJrqPGghaUZ9CVu119+uRVZu6eO4n4hNBGjtFeF8hMYJ4O2H2XSk3k80unNQFpZSMrCn0p2
nwRUEl4EHaN/vGhgnTJkf4aDMUW6gUaKbhAbITYchf1kdYvndK0qdQjlMDqu7As1ZTpFPxZAm1+r
e/JyTbmSvoQw7bGUZLxfKTEXtVvBtn54Fwt+EK9p6xfE2G/Jb46qM79as2yQOBxGn/j7Z+QCS9ba
5ya0VvtSKiwgemnQK+BkejDZqpQnIMYUaeKNMiUTDuN2acn58cDVqzWDCh7s8zHLQcQXMQgGgUJw
01nPVar6BJQOhXZ3bLZzu8YpEbhkCXjB6poHYAYw5idLylz+TkE2dZR7+/VXhLSIzQVOJx0a8Ut8
PF15iwO4CZ72hh5fpX49T9z4/LJoWlXFx8CqMVxzqfCCtY/Y3x9p3X30UuXVR2V2x/DPQ0gvtNu/
cL4WnUfAxIVzexYuEe2L7Ghl8F1B5hLCfUZbfVlWf45Ts2Cft+N5sggipScZO/UdA/vHm3Cf/DZO
1kg3JJuva0feLcj/msM8EgC6gIBE5jEz6btoXi4olQo3V8J2n190VWZv9I9QsLEQB+CUQHFDmXyN
VMQHKoJ8t861lkuZ2kq8TY8z92GroqRwJPZzuKzi25N6WbcBMABW27U+g/FKm6/JcSKeB3+ESy+n
rSlnrpk2Lbvguna0qJNwek9skNhh8hXJzMSoa8DA1DhsF271T2RKpeYjGF/md6mO/PLWZyzz4yKt
gC/zlaE1jKpChBblp/DE8cJFpNdE1NvbCvtK4gGqnP5XoyBQYB3aocXzIxpztACfxDWxVPw3IDlD
/0m0TqwNNv95/z34NM1elSjrc63GoBxRt5ALY3dTMkl86YAordKQBgBJYtN7gBNM4aRU17HWf3Dd
9mPdwua2KMpWfRcPKc4bp3P0CqwJohBeThLhhw+4iQvJYDh6CWIzFGaeMKFxAhzWJL9AHAdpxvW1
uZr4mfCgU2bbphbEaMuvcOqWy1OjTmdQoeb0e5AirKn3yuspKVSLGzG6T4Nfns4MdR9SqJyMWl9W
Hc95n41nBwvSHrOuXmPTTgMJz2KACA98XG5wg4leZpttpdQehBSZG4Qst8PJLWs4y15OjM1TACrr
+MSOZf+DZllhOSLMehIeFF7GoXFxb7pbbKdcwXOyaBmScTQYptIpcA1wnGZD2YvGQCaG73fRvhyF
r53zpznz/1imaUUcl8XdBiD4fPrI7CCit0AjDGvHcqfd6gmOy50PSqcT7y8+aTYinmb9Xf9vQ2Qu
TX0oXEihtYL7BL2SNRIJl4/MDPtekCY/5mg7yFnV36nUTY2qP41+U6jPQHK+5vX37eDwroaZGIfi
2gsVY7TAXsgoYpiWPtfqO7QpSF6+kbmDVOMpAIidyApo53w8in/q4ftNaU+MGvGZzBDxiFkfAiWi
z/axUB7Xp1MTlBbWXSFHNzIjFQIoBKZgiyeaHifdAtDxvzzvFC63BeyW8OSr7dsQZNlnik8lJaIm
9yT7GDkIaPjST+lIk0qgOC7OGSUf9DwADeQFC8zDHArDm6HER0Ev+Zc5Imydb0Gsw1/UmhK6edti
KvOMrIqQuFnP75HmlFtXWF0Y90RytIrAwG4LPl5i74GffOqrOY5BHoQtOxT6NKTzGJem85/gJ8Bz
/2KWybzcmyVbRKNMJxg57X3SE6Cen1dK2yUWKLppKx2mKd6CMkqzd7A9HzPKlS7QG+beO/L244YW
9J9tC4NeADR4xmoVAVwk+kUu/095MljIkHvaWzL/4EmKV/lkvpv9Q9c97HjQ7S7uLaR3UYroccCI
pf4kM1ybe4jsofKCwEmCSSCSnEj19+ef1QKiCHMS62e/JuvoKWHpK9+PudOeVunvIhmmoKWLKiOC
9++Kc+olP8UlUIkMELfaMo8mK0bG+h6nJas1qYK92jPdnFVRnt9m2xp110IDZknycOyeoEZaFlsy
iFQXN6pKwMdj4fZHC9S4ZzZ7YtW337TzMydJmhyYpjOneNz3blGYOVZk0m0OMkZXuHVeBg/iAswE
IkyB4Q5GpYjRokbpFqKEkhRmQbou92lDaU+bHn+LrWzwqd2Cbg/+c9UX0ureslMt54K7dc+G7Ywc
7ib2DXEp7jlhqe1k9ADgplqsTcukPmAAL5jXTTskXVNCoz2uQNlaeu4rnOtx4t0ZZAWFMT2N9sOO
XD+Ux6Q26DlX48HfM1CwxNPwG4+aSAJxJEcJNQeAujEJ0BGp4wx2wLbvyLHeCvWTUWySzzmpJpSw
lsLLnqVSw6bcJJvxx1dXnwwQqu1vvnepHfnFIsWopDn7jx64LNCZm6H7pS7C+bPZtLXvNqFN96DB
RKiRvyR4VG6VB2++Z+5oJ2MFTkNDA9YiB7dHxkK0lXqJCKwP4ckX6HAKVWS1o0fqvmiy/SEsjOhM
5EXE+GTKGtCYK/4HLMCjFiL1osihSokKrcFTd6Z3T330MeErr7mS3MLCk9Q6eXqds7ciqdDn2Jlr
BOp76KwA9EfD0ALH636Qx5GeVSaTnhV55AJ0L4CDeRDnTTAshuKRmMiCe+AdRbKf35IRvNDuwhIK
MWEfxvll4v3o/YOHYvMAl5YeP41Fq5ZDl6obntM10jxCYVEs4bXqV+2LeokRP3QSVfIzQXOlz+pk
ku8DNFhsUY+iqDM2pfKTCMg+BpGJVXOqc9C7DoTCNvKPB//NaDfs75ZvMPH+KXetGPQUab7QjkFF
+g3wqx+cjVI6nFXftPY67Ge2U0Rlwqh1gAT1TvLLS4cYAADTgTZpJ8w5HP/IYQ7JYMm3BUj94OoY
lwGH16Ht7OwmjOEyxRXQG3PwgHd3EBd4sgpWPaor9WqT11fl5RCsteCtNr9NEi+iQ3wwhoc72lwJ
6n2LSjmDWRauRd/UV8xIv/dfihRowWiNgy/f8XFjXzYx9pQNs4b0cLGU7SxnWPA87iqJdlwGGzP7
aMchfhBbBO0QiH5FlrC65ML5V+vMsB0ZWaGm3fIF++CQyBp93sGWvnuYV6hFsJnjhhXdc1bpYS1z
sB0u29ZryotuE1eauKkUGWDyxMU5ELMCW8kJf4Sq26Pvq3MpaxdIiXOQBzCr9O60AVw9xeiORQl9
Dha78TOBN8euJxoEKaUpLTQSufHzHkt+9vYRoAa98BOscCyoaXqGCNfvYxVWbFx5yg01m01y98O0
3JrEJjnhE6AqAMnT+fTG96GcK8SsIB0ws/lhAKRknWMySOC+I3ez2PAzGNlIYVgJ3gLayyAog0cw
oaRlAYtYO+ki9JIs6HEKbVNhGaYCBdRoZVtSQcPzfCAaffLC30vW3JHDjnoOIDrA5ZnBWFKQ3KPy
ZJ3jrQ8vJ3HifQXk6fLZgKjydvxd4own3aNQ6RCzgA4PiHmi0ailHrxq52i4WfWeTwUxfJkF9225
ELWclUscKnvjD+1Vc1MBnS8ebNNNVwPBlCu9wsJ67UkbnQ8ZtSaDwA0pDnt0rGa9czN3z6ktCUiC
UxMgm1I60LXNdbpU+57dimdFw3w+eS4hOwJ7EJUER0vfHRaH/DHewZEERKwIGAOwTH44HwHJGJeC
Q5s8yoNa7yxCsuf8eT09mp5nkhJVnaXkn8WvigaqOdtODIw6+z2TC5ZO7Sqq/Liob78XNRfkvQac
sr8wSATOKCHLkJzdeCeMpN6wg6u7MfM9TQ/Rh8JBBjsxSnZnhcYRJa5N82yfWvsNX6Qu6VAn9aGm
CncBgSXZ1Z+Dyz3geY3ArFe1mSHUsaarptgSdG0WPE9G8Q6HH6pU2xaQTOLCQi1dbCH4Z1gJaWvW
7El2Q7gPvsqUjUlhC2Uu7aycrvE1WBM7+44w5WtMUDkURsyCHPnSVToDecJWdkzrdenp9rZ7WSWL
Sp7B/K3ACc8P/6MtsTADDJWbINMrtQs6OzVG0gDfzHS4rtazCziRdijY4MLKRWmZ1ajViMLzo5pa
562PGjzyCEDr5377D66GaHV98QvaK3/Wo+87LJUAoN1jbuk/KTjee5HTfUUgwUZYCrmRsCGypejU
6a0Y/0j7p5vuCL2zZuJBNx50gyI35981IQo3c3cAWHFZNDr47Eo84WLpqvPXpDiuFrRC1LXK11UD
0e/0fM2lN4s6/bYyDuPEpRT7dMFZ5IhvFazNC0YJ1XlVbvSAQqPxExM7ufHLc+g5DBGEuS5w/zep
PgtNHdizPLLNkJqIjh7GmzUP/BC5q974K8F7mS0Q+68YqIFq549VLNaOYxtKSasF8G8CQawR39cw
fjVd9xuvcWEjyt09psEQOW5FUjIAqncah8nsI1EGylVOO6erxIY7JLoUXcIdbOMkdFPX4x7tBrd9
do8T1qS63q2PQ7h5ViDgEb4sTGyaRk2t27/FNp3hYafCTWf2fSz5FAu46Lhhqh4NsE5FxFzMZAiZ
zywOf4yO3N/K9adr5zBn9eqO4K0YnXU7TpXFxT8rsgOYruBeIezjp1XBexduOhOyMZRniY0leoqr
yHFykV5cZq0RfSz7fdO72Vf/ckEMdRuZFhToR/n7BsOGDMDt5ccHLrMfms/NNWSyTE2XhEq2luXe
Ts9yyP08jBqe5rXu7utW/oMX/VJVDY6RP3c5fw6BSAO4V38+JAm/rz6U+SWfPCM8Kk6FSPmtrkPh
6vMpm+u5J6pcovoK8Rs+AKU/ze/U2/Jzk5fBI7DrI5LxdzvMk31vQC5At5gbPY+/ZkD2SbgENLpX
GSgs1vFD1Orei0QYdP+ZOWFhM7PCYLnfWKdE2tSLKiXsxEg2yFJMKdRZl6zpROHCbNAbmGdQYnQN
5MJJrW1gSCjc5qNidLt6StHrCCmOpuszvG93WGMeOzsjSp5OJgzT3L/LIcpKw7HI6W/LdGnBIVJG
7EEMFthZAzQZUzhYzBHKODyMieOG8xPJ+gCR7AXP79Vib0Y7ifpKH1eh5MpEtcdp8XVy3z3iJpzQ
EKyNuvnlxAfbZmsrPVc1TWXu/R7Z9MmkWrLKdrW0AQK+lWTJb0xAMn7jMuPGnWss5kuh69RpXTpa
rrsaQfQoMl1MWQem7x0aDNLK/tqUNRzIyx6xuftMEIPNPM01JMieQ17ABtR15Vb1o+0hrnMtoRi0
by/ELWKBVX5yHqPPQmYpEUaf8XaVR60LHZhcc+I5z+SHuM5YxvkQv5AvUwGxglMWvzy7/X2yIBUl
8s9DtI5+fNQflCrdIg4n4T7ggz5Rfa5Q9oMS1lvSawM7N3mee/Gjje86rn3GCsbfPcPuJlSWAdTa
9qY0NGqJpCSi9eH3aPNWKyCRsuJNarmotrBUC3s6DYPIXyFPOGz84utoZR6F6te8ratMtr5Wv/Ag
LSit3DrCTP3gK7J5e5kH0m3tz4R7JXJ1U5ydA/ED6Ru8JMLoJxz2l5jF77a2XNrwznrnaA2/ekTH
re2fhc5JCUdfsGm8r0OJy2Dbh7v5NlqAxylCHYCoJvFVR3DOwVdVr74VuA+bp1ItDSVIqHAlYFD7
rVBKA3kERDr5CLlEJqxG6XyP3IYJG7vUwLnfPhcg9jl3Ks33JrLaGQ5Pe7bnyKQIJ3qQRUYjrgil
OSqXH2GY7+QuKzbT0BzmvcpM/jMRNRTfuDDDwcUx3vlwBa9Fv5AwF+/Sf6WI1uaFz9Ctca09PAUI
cc+VsZ//XmgnseWnjdDFcSjZ9+qFzawosiQdG5OjTDIYTKM9m2tRe0fyqQ47/5Ck0fzn2EhxREMV
MUEWJRq+Yey3nMv9dceJYyKjxDMOspT6nlVRbnEt8exFUXCUfqsC3n4tOy7VlCXIGhqQ7twuvw1i
GdvPJMKDvVkuRmWcCFDyb2RsDhPxJxGi+536v8Uh/FFy4i2degvY41rFjaQTbVON0JgNznEJITtM
azrPuTwaRhmPMQm0ddviqUEXXDFVumk6sYlo/J8vqpCKDHyRQyKGKjIWBXQb/t0p65ZVYEFpM3a+
UjIAfeKu9LkjaSoTxvmhwCRNVM1H0sOdxRsLbVmRb0g1uXyKRXuD3c4ovAup4lay1i8531LiDG8Q
EnG+oCbZoE++UJ7A1O4EpgpSawtjBaHPJnu9ircB6AgYIj6lYtdx/ZR8gwSA1MJkM/iyJS0sGKCk
RERHa1ZAuHbxtiXVrNoOvV5ud0sJ76H5BKLpK0/CiwCARCMVbcE9T3h83HWKWbsh9Tuf0eYITeVi
oedF9+sQbdUghF+AUrXO99wB8IA30C+BB4l2meG76p0oJ85a2KTXOKnNU9XU4V+7B3qwy/uRDD6b
h6LlgEucOooL2hhWpcW6hRfZQPpbn+NhQN24/KCdFcu7CwylT5lZrHo02ev5woBQ9eCw/KN1buX9
kcNgfNwtp+7cPXtyqi39BPFqeaavbz7Ax21YIisFgTvQTY79PXvgSSF+741FcixPUW4P4TZNAgb1
l0u6ZFzFo+jKeJW7EumD/Tk54OKu0dZiqSQOm2TLmDrkHfDGY/vdzqD4eHGG3Sux2wIRcSLpinZk
1eW5sl4QZHX6D187aCIettO26Wjgv9nDh6ROG4r4nSGyKGJ1zJEfqKhu1AntQvVptgeS4VPWtYCd
E5KqVSPKthxRv9b0a3u59kThf/jwShyIrPpm1DLAppnsJJRpL+OefS9i8NtJH7aVHau5F7HCU4Vw
Aok2jQISqNIzxXH1Mh42gTjU/lC1AZrSYqpYEoL8YEat8Ai1Yv7F/IpI8lIk5kPu0X/Ktys+LCUj
MA2WodSuW8QbqjnBXHhxL3LAtEdeeARe6rtQounzQuEpkRpuT+A7OZoEOEWEFxNrK/z42Vf3zemK
j20GvDu3ujL7DOIbetbHxjoTneZcbYnMqdp0evXZjYI1mHdfzXGAXf5Fr0ePzkdTiRgUXHXu2qVk
yCe+9mcwijRx/s2e+6MRZ76MR+cLlOW0a4Pvda6jC4OkJGpWaHsU1p0FVaJfymmiyD/HSiH82ClU
gIqRsUHeF3Anhn9g8YwhpQPDRwctLbet9UuAuyRSr0V2yGHP7l+YXRwO36TVCsCrhhYO9EUKIJ9V
lbBLyxTRigcAtK4aO1mAsLV+bIRCvJOa+7TBeS9I+v78u8jOP2ctOI4x3L36TW4uWKj3oFn6/1MP
hLasp/BOEQQAkLkAQvPxuzwz4r1lc/rCCzJFbQOykPiZt52h+d1LZO0nc9DEYY4tSRqjINO75gOH
bqTDm2zVF7/qDoOFfZorbZIAy86tWj5lOq+Bl71d8CSTwIM71SBQTV6mb7oyzZ7w8olCQOK4bIfe
4jaL0aRo8Jw5Vk8HfF4s/NeAjlgcD7YRN8LeHOWGTsmI9zDEpgw44CKPerSVZxqaeX/NMWfh7/YH
VRjbkz6vPKtpO+2b37T0LCLDrWHKhtB6lxRH18TfjZ49gS84PpEHJ4NeRfYgtN/ozFO9CAQASiLB
sIc0d5uTcrtF369WdqcD8zk9crc8bRP7lWRZzIg2qgIJPzRSEriSXXNl/+aBudk9y7cSw6TfeQLa
Q+JgyuxPSGj5ghc2rpmcZagiM0OpDOVpGsMtet3vtHLs2H9QG2y7YlCOqilgSOxWw+MMc4WivaEi
6bvuL/QT5Z5RZa9qfrpSV2StKg+0OGp+9MkFKq46whZsVNN6s0+9ra19VdKxS+FpSpojRjme82I0
tI9+kFZRoUj3ErP78XBvi2VgXonMabUkkHEuz6xOPcq1SvonVS1vXuwRSFTzmouVNVGP5qhFjMXr
MGem5z3G7OkI4AMrgUkqrhkci9yiUvzJB69PjMzl6YuNV0Ni/mrGgd/x9pvce5k8RkX2c8l7VU1z
x23xyDXi6yyfasDltgfvGN1JgVNOW6kZYHgUHzANkmnH3kCdGNlFoscAcODEaZ3hvrmc//0+yM9p
8qOaHuAPKpwdNLyeetEonA1oihTZd9CxnEQenS9g3sYQI5jErEFzsU7nTHUr+sjjtUEbMQLn8RGI
THAAG8nC0sS7yohnyti9M/QEZNJww3AvbAtq4jD1Jij3PNMxihSBWrZawf5R121ch7XhBBHDnlXL
f8GfGO2aJ/yz8cDdY3oM7dE2fohGea9GdGEUjJ08VM0bbBrHI5PGrlaSPnM3BOcjWwkpAfMhgoVD
uOzknk4QPiUSSGFlmXwJ5TwWl+d30+K+aCmHvbZfREXUCg9+sZRav2p25eU5GBQdAHLfgu0vede9
WdS76Ix7lKpHZBp/opMMc2TybBdhnBJ/HV2WDEkhfx4hggZxLcWK4fdfvBXmCP9dDZTD7yJd53Il
XbQJbvDOY7vuTXy4aZSEwvPxs2Y62VjOUDFR6MjYGwM8qn0kGgvz5x3NoCceBpBjLWkqaftL1P1b
AXj05EjSxlP96P0wUts5KuLMfakW/bA4XfOdKt5IROoQMnlS38yLuOUWK0Q1PuC7MHldfLKRRcNE
yCJ+nFvJtyZRPsKLk4RzuMWw3QdtjI18wH3oR3brKyDmYDHeqN8/vCi/1N8rj83LGQpaaPbKCJWZ
8tue12ELA61VSKNkVh8hdLDYFWji8dU1lV0GcXP/BlpCDHYZar3JSZJDt8h08lKYWMeRhhB201Me
V+wbZTInazxdRqod35ASHSgQE7HSdijbWi/ukVmVDdSSjOJdiSrNHRPJ39AzksoYcNP3Gx25vfsJ
4d+WYcSxeSPO8roZEP7lOR5WbtfwYaWp47rCn3GV2DXSXC3GVqye9pLXS0wgqRKUlCTxg34aJwRC
ONiplAM3IFjjg7tlazyldBfPrny3bh98a5rN450e6s0//NUD6wEtOiQxDehJ7rPt/tU5tE/sOcjJ
xpSl6ofp1SRUN9lRnzo3f7VF2Jaexv7mpRM/Th6GCIRL2OeQ00cStLrBVXbsbaliJ7/7PXDLVa0J
6N8eiGI/SZo6EFv43UprrgThKQjQyxlSBgCa5RiNwNgNNjSQjiiYdu/7fmBbCDxNU+6zwmTLXIR2
jc7J1Ie3Zehxoe5cGe4GjeLEw6KymTNuEaZhv+wqWsA335bAa5A2QXnz0FUFQYULHIj7P1KTpr3u
jSIpDdpKXjp/WH+VlR3tHPBzjSZ15cOhnk9msTGEUU/hcdistVYP0YEl7WuqOLg8hxOhEyGbxs43
gIOZW1dFN3XE5ypH5/uUb68sDm8GuoM24JQPR1nDTRW2BeD/nmVSQII6qB4Mo7A28Vr1JdOyrBSh
3xRMOUNyQdjeibLG0eSIwHWes2i3PuxNzHfIPnGG4tFIXBjd9c499xeZVn5o9L455uA7v+MxrX3Q
z+nEKnIPgk6tfayGFXEqEW5AYEOIbrM8lRR8sFDPDpp0E0N+HdLzXp/fstrphFe790tCNbUOLrbh
oSQrNyefcr99iaHuPc1RlfdWYmo+KKdPZbSN1FNXMv4lwa/Ie7hoBA9EAa+KnW9l19plI9W1eF52
uASotnFz/SFyeblAC+yxP3qZ/gT7+qxtAAzFK7gewx4IwCzzfDbpNn4HWs3gWSVjxg/L7E6GDO+Z
OAAdU4lL+uDCbr4rsG6Yz8PBD23xm4oK+r9nDbu9mFOU1wWhQ5txFliAkG+/02sC5VppYI6Oe6GP
NsiNlnKS0Tzwg3BUjzMgAV1cxL/cFXEF79PPSAV54y8+CBfhb188coosZ1X6MheShljBG3KywM0T
TRGcmVRqss5fYgEEgBwE4tdEzDjTbC+sJdmkgUXsXuz5LYTLlpXYnMuGZBCmghTGcEi3rjngYQwq
uCuMT47lQ5N+5vAvU9WlLB91TKZVOOtVx7BKCOb5LglYmxLgG6C+WNwcZXw0hXNCS3YpEXPb0qyP
t72OCXW4SwJPS/uTeWCNB8glGd/l49JbITAVc2uk6o8C088bRJiLsxAGgyPaBbYlJnKxCjWcghsg
DKlpT1LmNOTrqv4iKHCu+dloSeLBxXzVvGprlwfWtEQF8YbkkuKFTWItBEl2k2GIP/B+kJ4n2mlA
wqYYGDeZghoP9tVxMvfjAAwy04Rmqn4IKI/daQGUl0FNZtZm9s43no3qwSQmcL3JulWIAHi+mfnO
bNZdtA/DVw2viAtakp2BauvWOFVGPiWTFMgkbiqnyXMUSoJOW1FvoNFbTOzY4qcg5OQLN2jTlMRH
twa59S50oEMVdrO+lEITOxduk5LVIAY+nvrQYdeyKsCDWj/jXwVSXoIgDHduH4yZ3tt8aFCh8t/i
p9kcptGtlMDOzxVN9EnXim9BN2vsQm9Pq57PmEe/VCmtl0osqoMudnONY1o/WtO7izuX+q3HDWUE
purRe8LE319qo48gAPEqtbMXTh3s4JnnjZWprQfS5TdsLKvSJ7DPH2qnhHH4DBm2lZrnAmnfPHKD
QyBTwqVDttGd1TTSZtdyGAYnoclKtl64HeyMMeYPFtIo3STJQriG41knGPMCFTRMNDSB3jj5oJkd
w7S7eJ3Iul+InROV17RKpJJ2OI/pPmQgoa/wR72g+8RbIIEtraGlm8M+Z8droKG6WX6jNVeqDVL6
z247ggPPMlSdlqyX+BisIZ7oJWc9bNBZ73RaQ9bvHOn7SnRTMkpLkT7cgOFYtS1UG5eZneCzh1vt
qf7JgxmyANFTJ3ay1bcU+Xkcp4vNUi8HFPL4rLhWzXiEEMQ4E2zbpb0yYePd115Hsw6WcbNO8grb
zIt0pb+knFYCGs5FOqT8MGte+HNhrjH80qq9B/R33/V6yzl0CY4zohF9u5BKr1cEJ0O9bbQorZvN
MMufF4HeCqREGrCwRLPJYAupim7E7XLBCz1VGtDzrtpYVADgSvmnBLpL1Zbr7F5JFnCDh8lqbzbM
vcL7SHRDp4aPBqm6yxyYEs7DvIfKIRWG266Y56yLY+35TdIaCNLxgEGCaSSVnOWtXHGSXzigEkAJ
aZ5KIK8kUH1qcrOko0Haw0AtR3fWkUVuuDaKTynKKHtm/tDt5rY7HaJqN6aFmvBEVolE9wFuLiJe
tFq6Z6rKjlkjR6NBdjUKZv//ks6s1D8JQ9z+01n7m05t2EZsnA+vWeRbWdyDKn/8d4J5QQOOX5Kk
e8dhzX5C9cm5VT7BeTqCFXTs/nK1qhZeN+JwVG9JFGz7WZt+AJvOMgkPM4uZOohAt5IW6NEvIFc1
/VcD9uGV8gItpn/IbfH48NCAtSBcYvGc43TbdpQH9hPuZFoQhGLSrZXNqBKMqLq1WpZ6gxAuz+vf
F1OvoU9xQULQskCbAFWuVZEVAt4sNFHRdn4XA0Xb+j+CHDmzfs9HhhvW/nuq//rq73B0JR9TfGK5
8IDMtjo9vhDzuzzXCeSqt7FGLXIENH+FU/8UhedKGxdiLc8BCrXkKZQIjQbPVBPE5IrLq4rriAx6
QKqntTo4cUFnKUJhgjE4c+/6fB3UA1socNK7StThiVzDN3m5BVDV6i9ef1XaDgjl8SHZx3uongDC
sDxsnxoCMKY0TLs/qtWSkBdT5/AKwcr5aug9xrpc+BjGlfiamJnb1Plc90awbDGo2FAV9s7yFmXs
vbxhIfckXWSjcg1YpdBgTSPSJx1VsC5QSgt7/aTe8bKTokVwtlJFkLQ/Ld/2zI0qnoM20yIJNr0m
O0M7HcXM96D4zMBYoEmTm0XT9oOsCg5OZ/1UGCb3ZS0l9Yw84ODAQBZ0ehW5uj/RJ366CmGKwGLP
4GoDZIIinE68EVHHn45LmEbFKvdgT2KSLIGgJS6+19UzG1lVlT4sA5e2SaX5N25iQb/sDtCFg83Z
xhrny7WWJSf7/ZpO3qbViE4nUXVyljfftV7RmrDvcrxfGsaJHBxhsXtxT2rlsTnZ4oRsLj3WFvzx
XLNfR0merFoSQZw0eQnjFBP4JMxMzK+K/Yc4hyDxXuM/aU8QBqh310VWT3jJB/munpbyT6xWCGY0
O0PKyRNlff+Gan3hUJXG+seC2z0y+OPvD/gfGdq69yE8mDXA0GZsldJd0ijdgM4vsYxLpsSlJOPi
4bRbpiqpameqqw2rIdQ7uHC4Z7b+rDqmVSzWVcrkSegnk6G3Tw/Rg/h39gvwXQenOzw8rDSNgUtO
za502wQTa/fmKdTZtztZ515Fh6GIpvxIQjzoJpclIXp5q14PKmsu85m6rsQTNqyuuV5j/nVeSAqn
jDcqnnLufyaKJJAdDYE8x7bheL3VUqdgIOzDGNtCytOgbu3fucUVQ0pwHtCbayzmUEiWZ+6k5CFN
EpiMz0QHJk6j6A+wyXj+83wKd6fDWlxRbqB+T1LAtut0JZpE6FwFtnZyT67IXX3kEznNRkMM7Pz9
oC6hel5xghU1YVOo9AA0wAWhzuYWe8pEvjwrXPhv7CMGyhCUE7GXXxn7xVYXaW/MWXgMfzR9xBu0
MRtq7ZzNGp8YvhkGii1KRjcSRwssmLbZo1phxXCFOgfDV2WrlfB3SnrOGS4u4PWhdQVLniywvVfx
R0XoVIFrtJeiQrHDZYgPa7biGt6sXhCBX7Cc2vOaR7meoVPylhekgwi3gyj+mq0eQ2arrCeQfhWD
NJHlTyC929Fqj81Eh6/Fllc01Z2E/+WuHnumgJDiS2U8le7+AA6iPzQYDO30d9gl4Hiqu7kNcMtb
zjH62wuxKaB5rUbxiTTPTBLz5J8Y7/8lO0iBKCpkfCLruznBbd4Y+dZDricEmOSLPGIAfEl9xX0n
4dzdeFAlSRK9Ik1xt9O8S31um0gIU2cJTKENWC90C8H2wCK5BnBpgwPibvhrbFLEGBdlBomTZ4Lw
0aCUB7o3M0vEY5qHuLJHaHWOKghzeoDlUChNuuNpG4b2fubgLxgHoXH4ncIxqeJd12OVIeiR1uKg
CeAmwuEHmFMZaRIqQRlOq5jeVz8wdBs12l8RfwVjm9sqEEC+DUxohBWH1NHcu/ji0d1fA1bsQNfw
eoiskVDzzXEabSJY9CcHKbEUyOqXiUCSbfB9ZPUEzvJHuvzRldZQ7imWI4pws4gEqm6kZE57ZKwj
DFXSm9ticNkSPQq4YZHoff3ugshx4Fcx+imccRA2EG7uXNXfGIFes//GKWNsy6Ap4o/rPYq6rR3Z
05rQZhKwKuXR6bpNCjZP+r76K9W3oOKOUnD2vqA3irb4xcEvNIzuhwXUWU0OkHnfdQ/jYpAYsCZ/
xju621N354OFXvqj2KnAOW/sPu6eppcOdKLnX9w3btG/346M1YPPxpez//BFs3GRb4w986GvPmoK
hg7IxSKNX5ErMk7ALaHXrGZMGiS2WAUaka6+lqtg12ywugZNmhjU2GNXFMoLjgMOmzVLod7jw++8
wZuu67Tnk2wqWKsDnDpnwQyEfCuBAsQz30nlJNBhE/01ptuA0j08DNPfb8uHDLDRFGKbXV8O2Lx4
boAfYZXF6E2WBoojY+us7ddLmSBnqTSFK9tke7qHSqUnqGxdD/Co75WVnBakg2ZPBDX+7mMRvZfE
I80A5AY8C2ccrPDKbTEEdJDNFVIOM6p2BBSCGzF7MD3+n+Ph+tLcASSDdVi4eaTtRDinVskqpKo4
iHD2OI3Oz6QUujHJViGtXIabOpagicUvg7SVr9USY3erY+5gh+NoowO0I0ETHbrhzgXRkKyBPEnH
FI7s9i4k9Ug/rr4pU/oxLUbq23oullDotjY4Z8OUlGhRxhKwrzOScFZg7yOn9Xu626AneWtwGNDS
+WopFe6XMPFz3nNGggyNmSwT9sKhAyDOz59S4RiclZnfbkpStY4ZdHlKup4Do/cOGMt5rrQaNVAE
mnufszFUxwreE7K2okG/pvzXUeVazN24SF1j8Uicx7fNT/JLQVTBZ4AjGjymq3VS92PoApWA2wYa
fy/hS81a+HyqSZpMkaoyqmR9VVWy5oqNcI+0sx7RPTp+Ozh12L7gd7kbkI+1aPM53kIouJdaKgX+
Kua4QG5Aq9U30Hpn72YmXQFeTYRW2YAZCOpSG7pCHR9qsJ4LTN4zZm/2AUPcdBJhu94UmzrGqDKP
Fc0rD3BkaQzm4Q9Igj2UVesP3rTdsBcM6s3Btk4ps5LvM9wTcmHQJMUwDRoLKyl0MgDZJihME0RK
nwjnY8PTpjyNR35b4wc+q/erMaXq7IfW3TaedNaEPeO5i27zQ2NUHf/Cz7GCWouZInrROxUvZefd
Y052ZRNya3Cl3evSZUQQi6WZLLeAbZKnIPtQeELDmwYEz+8CTAdJXjjG1pbmqHj92l7UoxbiuQdo
1JpdQRXZ9cbYeuEoTsaMht2Yvj5+RIqN+ETWwqUn6i7arueOOmtfiTacI+gU746RQKB4G+W8RuAq
Ce3vYJFGEsJZsgyNPgCVXUwY5BlXG39IBFYCkTd6o0MGmoWa0FBbL3LtQey8Y0+/OESjmDoXnYmu
45Z8QMlcjkI4JDI+VhBmxLRSGLNiQotX9sZSuzxNnIGGTcI7CQm6oVuoO4ivIPm/kwC8J9sBwMdL
rphHRCdzvdb6gB/jOE4I8B8A0Zgpk2HOupAU/E8YynieDG0c7D1Atfq8axhTYySb913hlK6knkxi
sZN1F45BUa5FPRd4EBo0m2CREzCf1D3RJii9wloXj+ytUnSxBiV784mKgmGYUvpqso9ZuvQLi1Hz
3TgcVc2KnMiJr56RzmX7TkrWy+V6Rdxw5zucWPxAeg+749gUns0TvRgGI85ivASsHrwU8UiMLAuV
BO8r4o8V1Zt4QrduZU1R8Qd8bM1wvwsctdJhuqRoUhpKg9756s5r1PGJGdiOeJqu3I1LjbwqLwvn
9ZV3EtADXwzOIRCo4ME64Q8drseSsbEQyBJmEf9vdCM7qymFOf1toCtZgtb9ODXXmrg2dHP+u1OF
wUrbYLYbK7EIx6yUJBrEybMs4kpamc8fxEo0mTD8HJTesqY6IkMWo/Y4s69CM0jJegVbGWpvrV+4
5wZYD91jbKbAau78osO14vHk6nnIaKGqBXpcH/8Kv+06Pp0hdVW4uGSHmrTmaNvZzrLgHrC0QtuN
eIXv3gKXHWan5A/myz+CohARVEtHg4oMz8YXKS2MjXHTpJ8Oc8pBTKkWFItMG0Pt6xLJpYmNC0ul
DMp0+yJUeJX69x5BmLprQnlndt4QzP2eu2KIVF4RnjJTeTR2+Uz9T1fvCIqPadocKFd+Q877nLrO
qN4MT+ap9zCBeA+cgbldHe0hP57ct2v2VsXKvJnCzjvTPYlL+O9J8cSl1j852dmupidtITSZKb9i
1J9FHE4thYy6heX67kL8eyT2zG1RshcMTkS1qeUB2OjDQLSH6Trz30QJzBPf3NUAOJl/CLtV0D3U
CzRaGveIX4Seg8N2L4DMUVxjw4EkZryYPojhtfs0cFj8PFDeQQc6SaohKfou2LESkOyFzSdUuSdh
tEOo0hjFAjT1s9+AjbE+3CwgvicSDbgeISrgerrseaaIrevTFs3tktOeoKgMPyrVfmVZW5hALBtA
h+MR7U3qENf+RHcUo1ezq6sxc76IuBTACeGnIKqpokMW39yLEZSwDV8rYy5wlo3zBxO79OK15Ufb
W0kBJyzNWgZLViRWRIcAKzF1OudnbKAn9lhu7s7TUZuQoGMVIa3wrHotaSueGhXOsJGYE3GHQLyg
0vePFuFxYzUB+SpkOPqwNtGEfOvz2ZGJXpAf71CdMR5eIsQAxKmTewasi5O/iwcJmSK5OKSazQ+F
iHXT0+m6qC+njD/T4zZSmNIlX4ZrYLgiSbBnO4lrT8AacqsJOyPk0mimJfhwCjpqGfLn5GC3bjOU
es2FSxUQ5VR4zvbo+SGBeCBmjaZ8Xe56EJkBSk2U0s0MWtHFntS4kQzjO1RYRvlvq2LhA+ZDUOOC
oKnXmh/DAZyygtREBVM3cPVglNA2S0gDTLeAMldLiBMzz2ehtBft1MP2AXvHVSnJqrY6vK2OWwjk
BhCCrAjvrm1oS2sQSXV8ip5WxnpeyihKqOxMe2S4bBOelkczWRvO8ByXvRQsHKmTltEVh7KNe+y7
I9vdCzHXa1GbyL3rw6/TLK/K3JYnfxaboywT5eBT++MDhjodrt/Sq1HyFrz16xCuIP/5tsQUUav4
jMZCSHFYWQBLAAWDLG4hGsU2mbaCF34fArYQvTw24OKT4xja18wGkp9HFo+gNFuItR/uWmwjECee
i2iAiIzc5Uk2choc9b4/04dlWsvScjlIIFPzdyUbMWLo48/Exx+OR6JbWeVli9b/JLZH3kPJJHoZ
rM3+KdxP8556uTomHErHNOO9AqoWi9IWuzi3B9JHnlY7Le34A1prKumsQs7OIERDI7Ifaas5vqUb
LdA6/f1LWiZeCy/l9BUlYwugjKN2s1Q4uV8DO5QuOv5FRsJmJkM4UYBFbLTeIfn6qZbFDpxwFVrs
KNP2J6SbuUmxuYrDALkE7dnEy8bkCRwlgU5dFoVs63r/yua90pPkSj2aOfAtFMEJhmhQW9p7PcTn
kn3FG5SoMJ6Bavzo7CVyatWz3IvT0p13lNr2jbuoi4TUB2kqZ47zyJmnY3fJtYAdEqqYXdwrhdbR
0OkgvoSt0k8/htX1DDmxsPQYn8ZBg0OJ8UA+RMvHN3VLNnzZN7BUg9FXeED2V/q+WIklabA1Scxm
KDlU/FS2uXvG2cMBTZANRf76QFp46b35FpzcnnFlndokR8ZHFM5fxXy8RPgTstszcOWNFNK449gS
eOXiDnUJPtSG0ZWqZ587fPbtpfXTrooLZH+1XIQBCaAOm1AA+6OWup5Ff5fOJ5PECs5By27xV5N7
6o9BdvrB0B9CTV/kgOXDTK8saYM2rUJWozp7tQt+7pmQnyO37hzCtruBeQIFx7kCq3bJhGSxJzVn
GCaSQDheBEXtoUopU1x/l0Cfq5Z3k3QssK8hEXa6NSp2l/h2GmJiZaCn7u6Hr+qmsylg8MqdJX7h
Uo6LhKeHgqbk2hKU2Q20Nr2/2kERHDVF0ia6fOwP3umWFf18P+ZzbdLTvKwAvDdRFmOKU0WPU/+K
aqfoeKaVjF6FX6xXW5jqFPnXRayc/GS73uw3HdS8xVaRCJxbc1YL+TWARlMDsPi6rN/JDGkbQLIU
HboeGkacTVT+zhIOI6iFwtYRm6l1F7HZuLvtNILR4s4Y5J8JqDZeHEiReCMJtmmxb1Nar4IQNvGp
C4DC1RilEP82MYG5ld10rTvo8m7d4ZVL7lk154S1NV6uQPUYJqUGq6ZttENRmP9l+T/PnkZQqlMq
eYyE8VVzrfeE3nHEAojTx51PkmrH3W8294aIHYq9G4APARuHpnJuPeToV0HKz44R/HvXtH4CJ5+4
vIF4U0YOTjAYGTJrYpBKE+o41BVybi7+lfGolFL5FsoHVx+oy1PuUzHDkU2GTa+jmvVUkbHq2O9v
vvGrcihqMn/QURjOaPcMTMrjO97epJIGgndT9X0IHPuqXJfs6Miyux/od3MEvwwIiBHBjNSi9DPT
T/1D+lOX+JBl6YRGXHBBiCxQgOWmhbcOd9+ydpkwA9x8PpZ3jXqtVSSaszG3B1M5VjOgGHOHvtvX
jFy19B+rbQ20ZOsofPU6vC/IZhN+RLYcDcvib/iADEX1va9ZgJxScXO1jmN8F2ytLAn7JxFenjGk
aJsMeGgEtnPyPznFKxTKKYU6cedX3PrxTFxZ5jcWzyOglyeHBnKEDjK97KRKEqmQX9SUNP6hS9Cd
eg7IHJPgb/3VJz/4igSQRMblkE0DK/MUJQvvwWkXaUbOEmOC1XnNP8zS5vbZDmz2n73PaFo2F6Mz
dhcKdgnxvpRZ2DU1SijtbExJUzvi5uWvegZgBbc7q7KKIl5Wc+jctTkhJ79NXKbx5lA6KXM3nwS7
WXaeUyJVxSwPgJb9W8c5qzRmttff8wclqaCPWnEbcbdseA/25tUdf3Ln5LkyV60ohJhyeR4lNFaH
8RYLiSSz+Cy6Osc+G66ayj3FjGWgDo5GT5HVPj2Jz+QPau8vYg9yLzgKqOG26tHFbajWDFPyyn3W
kD+QrZL8GEqhDfN4qq7qN9AcoL/1NtjFt1i2RJOOPJpaSaxF/wODNRwJcnUrmA9BoRWK95BsUfOf
O7V7Pee2o2ujy99gx9I0zDhxpyGmlUsO3iRLpOYfFQiF4eBquYA/8+2MQgDopnJZzvijVIEeYev0
maCrcHyNw1tXISPA3yrRUCJqzluM8xYBY1cqYa35cS3azHGDsOSzW5eXEFZv3M3kobIhX3Zyn4od
Jey1Swd0yAC4gOzvBOSXFOKEa+5iUkaf/7wO+72vZe1yKc56GRO3irxPCFeUEsR5ENmr0UPWBx/3
d9WF5DvBkefIwAF+2kpm1uqHTjAKcGIVMSsawBHOpI/X/sXrtV5wfkY34k8ksgnO7IhC9kQxrWfP
2CQY6mH3rwajnJd4iUdf1MUJM0UH48AM/g03uD2iT5NCxNa3R4RPTztoqPqhwpuU/wnqvE2R5b5J
WWydhMD5IqKAud92zCV/VfnqurUc1s8hRauZKvXIWPWe2vE345DOZ/QwWHVjgLrWpzyORyH5WLLz
tCjl0G0TPEbz65iw9INy3M0QPijaT4MziClwluaYvpA/O13fXAwNbY6K6eRNnFBjBfpGRGmR7in4
W1XHPKn12AccztuyQc/4IcL8neiB1dUGXp8ih+WWpt4qcN1jttfPe1ThtQ0G/xpbPh4dIRT1SfD+
gIjp8zXUh8LdwLMjhQD71ZtHP+BbSQWSr64C0MJeydnAjBwzehXH4emRtBG6TFG5gb0cWzZa1ITw
ORQCCEyBVDkcScsH1yLdxCE6CYCJic+mKK+MjIwRxMuKCGOs5uqPdWCxJ0l2ZX0JwcPqw3dqNYRK
nMvdDIHf3SSpNy+zD3IcGduZOH7PimzPgFAkIMHNNLzuqI3+H2iLTfM3DJxrlAIPILf5OaKSpsik
GKYzJE8XMtnWs54ZNOg1xlGsD06/Cqdj9ebpMJEuNrhGBGH6X7kGgspGySta0rOBSoGKnsxlLK+I
8r5WqDUbX0gh0Qryz69CrwHZ0fdUGV6MhsAzdgs2dkOGBk9YzYY0BJLOHNR831k7F94iI7LRSv+n
PVDkKpu/mJkzNGv0myVqlPyxi8J5X3HGv04kvuhcbZH3nuHSbP42C01lh8r9aBGPuv3TaODezg6H
v0pnDOKBxWp+WUeR9Dw0SVmmx/hfVKT1hkGj30eEVY5mkZTxsnPDGWImwTRXyGLpYB2EYJfVvZfK
7c6N3VOztsRK8ypQkwHxnBeEwCT04pOIh3ypstuII7Uk+AebMMfOCnc87SgSkWlg5ggvWS0A6Ywg
tbIzYp9uPLlu34Z4RsPlwzjwFjD0ftrJtpY4EEFK/45gywQCqEcXxq7vDGMDOhJoAeltFpLxy6//
OFi2W8iaDIUg2oa4P2LhCLwQxyJcEfW4ldfQN97SAOja/ZYtvAQ9mCGyUBAn7N1+M9bis9ONiBYF
3v+3Hx+4s8n7qEE/KHempwITvTqnERerbmOA+8C2WoXZxQwVgsreZd6vs+1Le9DSpU0ugSRewlZ+
1+IzAeO0YvG8SVgP5OEUhTdSav2oOa0BBOSUJIo/mxvln2wc6dqVbEiuKOoFtPyaPYxDLhkBKtQO
D8ACSVfMhRJLC2KHpBsfrOiBTewGquNxudVV/SbVJnO3wQIiEGH+MSBn7x9Xyp/zTEozcdGOTNz4
irRCoGK+6tEBF9Jm0Fa5Cll3NohbCNuD6fTnuthw/bj2GfIFtG6s8rrF3FnLfiToYj7Ray0xaeW1
LIr2TRSilnDd3KmcUldAeXDRLArhFzdCfJNnybqacDAj/HXEW55PZNTqh3OB4D3k9Pv2k0LOxHI/
6PucqgPplPAkB8dV50O4nTs226L2nwfQFquoNWKBE53AInmQCcwcCSKtHVoUTdfQnbzzM9cWOtF3
cpBWSWLDtluHC96fdTzdSN3bd8OU6YLkEtiWEejsRdGWFvSlzNij2w+MwJvsBDxE0u4zUhruua3T
FGmbincxv5/GgB227Ii3JKS8x5+tgiRde2Z5mjwt7JRcZQgjbocdsodq7PFXdxnqdHbpobOATCam
tQFzT7yQG4sCFjcYkQ8n5G6cLkfTVORvZa6Cc4lYVUZcQCLQTjSzjWfpxCvfTC4P81WqEyecT/mR
FHomISLJdOo1B9D/YQZTHnp9RCgUXJ1sHMA1uVw+XPnWfDvQKi5KCO7NbXrlVX0PNLDbDScWJ9kW
TsMeeBIkJfM5+dp0jaSCrXO1Q1FsuEBlWok/MoAMIp0OaUkihGPT5tr7Gc9/w4KsCrcacDL3V5oS
KNeB1f6Xgwy6qPYwqmw3/Fwj2z9bocXT6dqEM1fuD6rRl79VAkdXrAPPbJsgf5By2nPvyuekaIML
bO8uptxrNfZ55ULoCm8O28TMVT0RZBHGcSyBZQdG09eqIbQU89UJN33/UJ434227TbXlLBU5JgFW
/AnYEbIZOtPWGvKjYshEGmzHyzLyqENIW/I+QDUJti8qbOkfaz3zVQZcqDHifxtJTkD+YXKK6zWQ
zELPISSa+OqrmI/C1J1sCIWawiP8bclYYVgtoVb49PMc6gDqft0QR7MsvC1pdfdNNWThXf314bz1
VvwBCenH+f+PFnnwky8qwHEfOeZFzbgUvSuaGMzhorGq81tqsoXlNLB797CNFOIZQ/cdf5fhyV1v
C2gJVo8mqMSDn5w+rdhkRJVhGGp7HXSKJM4haZEViSCSn/o7iHGu3BUpYinPz1rC2ZxkNUb466U7
9gidmqVCASWZ1+n1kMi4amwwNNTSTpNLQSfNHzCs7zq7UrrScXF3Mna/7qWLai6R5kqqnzmuZHwq
D5aNLn4eTbjM/Lm+SI539LIomPw9eT7V58X1ddwA6LEsVVbwwI/Rix/UVOCOfvlGoQ9w/mlo5atK
BFGZ29UYdIp6DwDY59OGt2Hm6cojpwI/GwFAYkT3UdQiyndkpDlYnsfuk3bcXvrV+RVQIseTaX6L
3JKJ8YaawxpjPWYG3sEFQOsNt8+GAC8V7Dj/cGCUE6A03VDV4K6heCZfbK+pblfl2JR4qN/Z1UqJ
flpFtKBgrc4gGV8VW2WQFeJu2WIwad0n/FP/G9t9JVkam5lMZC9//RHd+kDeSH1bsyl4L8kRihgS
2b8CPOc5WGqdZCxzWymBt7xntiPTR5dYEH976ieM9W2wBL+sEQywa0XW83B7NgcQljVa8TyL9YqA
16DOQATRwv4pVFCPTvCLJQZ7aYeNn/+lDejGSdp/84KoIZY39jMonCTbGpgRnPNeJka6yy/LTrUi
hEt9NNCFVdL70wlLZC4Ch3NYln5mkc23YWoO2TC/ThCLbb/SoZwUxlwkQeLYPB9RIZ75FabnZzIe
Sc9oS2l2dE9a6PfEa3rf644RitMsb/vXy4mJl5NlhNIBxKo/ujf/XOxnkIIThQX0NN3JBoQAnyzW
Hb+0KmeNUrXDVi2r1h7C36XuqWOHUDAbTrykxJ+ol+YJz2GrXf+W3wI/HCqe8hhJZETtRRwlibrC
VcTL1Rx0aLlxpIT9WHtkP73AHZu5ta+U5LvH00sUE95EwYKzCZ36o0kXwsSJm80m1RsVogKxOUFZ
3r9rgsdFLdlV0f0/qW0trSshvofNl6QD6se+CW5Zkk+7EJqBw1/Apy6pAN4pQlbEPiX0qtaOKEpO
IgzAujTUYKcl3xE+8uFZaF8YhwDd0xXpQVC5YexhfVPcOSeSWAssMQHYE9QnC612rkErEukQT5lb
PpYTq2jmA0bItSPj26SIIQvKW9qYnY30+0mSO/zuAMHL8f8fMODVJ4RLR8zM6htTLLG04s4ToOc/
umUMLD5xO+ASJoWz7qPsK9nfXi7ALbe+4N8qfGYJ0CzAKZ7Ct5wI/10opqPsDuuTUcpfndjPyKVV
VHoODhUtG9/CRHtY/GL3sjBSiI0/xCVJ1ToNKrXaOOd9loNGAZkgD/MHb1A1jGJvBwOiesMuVjeR
eicbSO4t1C6q/4juKpPA7cz/JIUAgKDCa6sXClDHaUQWidc+23vfO3vdN7GHFNo+78bpQ8lAIPSg
uhWHJlawBzdRQ5SGfRAeJ1ascYVz60J0wlUegTYZQxrg32yNxqFkciJp2VeBtvefJyATkIhsL+aP
IZgf4E0QeqOjZNvco7JwUNlhZ/w54oGR5E6XHalk8ZdPaDV8j/RZ8taapwQyjsITxI/FCk91Q1SC
Ey6Z/aGjoxEmDc7V6dA/VqdsRkPypA2rY2V0023NPd7E/9Ldodrma8vz0Wi57f8l/vOFc8D+gsl0
BFQmA+8AaBS5nuDSaIqpbIZSiE3mgDj+P/4oY/j/yhinxaU7Z5xzcwmzN2hSHjEy00yowpsTBiPY
iZiFWUrSs4kRIg1Pg+SBZbflfXBPnWctW5ci7rWj8AzfEiieYJ+SdmlFXlJajjDy5mrqtxZVZmNW
qeCwKnRbqAlk4E8RFvMLvh9m0Mfx+MORgoK0hb2Ye2Emzbyy54NfEGNp3I0EbBpN2oaHhqDMRKHh
R6crsWbwebXlyIANNWVENJYnewI5g6QAuQF71JGSfb47pidW0WdjYZuMevE1dVjzQ+LxBP9I/4hY
J0+PRdM66K35nbxhUwmg0qe3k8Xy4v00V8G1rpvgGdRhz3UWlGlYNtFjxDAWVrmFHJ0nR57mjEXR
v9/GfOGBBNC1xY1km8qDoaRBR5a6Q1vnC2t20p5Q9Aj11Osky6kPUTckG/qp/NKi7oQe0ofu4N56
r7z0UzfC8H1gnucWGdT0BNt3aS9Kvc+bfx0RBTzkCW0Du0hCn5ehF/r39LgfeNKWj8K+fjKPFKo8
uKfITikDgYqf4R6lQGoPGEXzAVejJz3kvaoeurpE7MVErSyncrWNQoXL6VNL57zkaYw0lGZEOo+w
uOnhtt3XBlzSQRtifGo0VyOAzJnPrM/WhcJ2oJlYL4jmtS1XlxsZIstG37ifAuF24ZqjAEHOQmcI
Fw3ag0JJYlpOiFqxsMtNCzDsokhJcmx1WvWQPHS2EdYaNO+bdh3j/Pqyaw0KHXJLrSzKtKEzi/Z2
DCcpgzQWWYtu/ACEjaMwVdLDAXX48vt0t7sI5Kc5/wDBs5Z9ETQ4z3K2l96MuUnG/94+9X8u1bvL
Pld4luk+6H5U0QZt6BWS+xnUXYitAVM5JR+a3PuuuUUAqp8BhuU68718HxUEpG1YBgh+/CjxCP45
YmetgeJjs0KL7o6K4GdB8J1cSd2taJonyhnmIyaWfUWFGq9/zJ27SDhUfDQRF/G73YtFZSaJUoj/
plrqE5uLn3ObYCSVnTFTDqdv+LJCgiVpbI89dPbSYDlszXHudhtnGCQJwvC23Nyodjc95TiqZQFE
epxTcicEqh17P/f+OAHFE59ZCnYf46Lpu2Z3iJvxwf5xtspdbKpu5MSVfRhHK+V0Df4typV9XNFT
ACFR2WEW0g7IyJr3EG0+0TD/QX5RVaSoZmd4aG8FDqlH0E8tejIr+Wz7Thc2Mg6Uymu1QVJFpUJv
dozNgMpZvgGX/yHZCo68C3Otq8ZhTbDt4ODPZy1qeN/rv/j2md6mjbsu7P4OK+veuakYSOXss7PJ
NQEPprFrS6hKgBQ7b8HEui9f4ALu8o64huM2s4qywHx/LNjKnosE7uA7IZCTuAFPbjkpkyqHeHE/
lV4njtYRY+doZsRF9swEfv3Hz6Om6YNeqWDtQD8q0kHp0Pg1ELu2tIurX7m43MvQs2mv2+Cce0rg
VOfnjicOsIyr7VRULxMIZbqFdNgxqntnxmXCTPP2/Bk0SGWUnxFFAbfICaZNqkcCv7Vclr/SybFb
tVBmoQxFvv543w8wIGZkXQ9bYOrfMZTGYTF+YJpY737uBKjY/d36Cqt2quN/jPAVWkIKo8hMYiyd
QAXPFFslwQjuAK9il/3W+fdaQUVPWZ8BgRUBn2y2KXOb7rSBISulVkBUYK/Dq3nas1HCg6ptUKA+
tvaLzKe7oqhfhbA21AF8d+OnmAdL7HLnbxYI0lqm7vycmeBo0KknyblhBTnW6RKGZgjxyt0evOnU
6n/kviaf67ITOY70nZGM1ERVAN1SNBw/yshZh58SaFDcWoe0P9K0qigC+zAaCz/N/po/S6CAqmMK
g3OYkr+K6bAwTIcTrJRQPdDPJIJSlkpb8F2g6CzWRYahpQ6I/JzG6cyH4l4sCWlhDgww6Vu3ggGn
P13M61bGUf7IjaJiowG4867iT3keN0ZbHFFrxPOMvOCwWuN4d8JqeDsHtkM5D5FZnXUHjSeeR6SG
D1JkbwMotl/MFpmdldjWNNyOHBNNWy2S6L0IxTmFCLs2kkJPdPe9i9Mro6nJb+DY/C1jy2DSoIQe
FiEEqBiiwhsylI+iLGC0N6VfhGSyPGvxM0d2Le1JETIeGHqiZTo/CrDktw+exPiY7LKL4O81+Qe8
vh67MdfE8qrTS9W/ie+v1Eq+L7A3S3ZgSA/5xRDAzOJY1kf1CJFwq3BbsE5jxK76EjIV28hnKQzK
n6m5wivtpxX+Mhgouo9hDyNErd+rTAP1tfRIm9uWToyWAEcocgZmft9zP0QZcny/t/0KZUwZWgV+
EFouBPiexlsqFCGbHwM4Kn6kgoX7SBqeRAup9lurJK8CaZUb6n6aFw4T2eOXdpYDfYc7dYMropSg
zAeJ7pnbzYCdA9G/oawTW85ZmHDl/qXUImuar0oTkOMMBlWXmqMIHuuwyk1IFWLloJKe9eZ8dF4/
3sM3YyDVa8nKZkbcyO6oIGJeWd0lvi0d3ZnMxMq8xwvcCqJp/A+StA5aQWM13yv1WDfSlY8Zk/ev
rHIjR1tfjyYtfBvO7t43FaM+xmGZjmSkesdT+aOWgdozCrBK+konv/XhdkUfSlHczw2N3kfESW7I
3ls2ydpWRFmb0Amqiwya/abos20I5nVdLllm7jSn0CTZbvRYIpjSY0fVju+Cr2Ibn6N5Jm0JIFQo
jxlRgsev4W+HDePGz3u5kzSigqhXJtGzHWHhqOU4njfGKVzk9JRliDjZyVcu+KhzFh/1hxcNKwqI
I3siZ+bT6ZecG/KZkb7+dNX2FiMxgj8Nm2nHECBAHilerpLWJuXdLL/KKqXwPM7Hg2E+VWzgNrz5
fvuqH2AmPyzLCQ38Jx1gTpnpgisIAJ6idxbnmX7YWceaHdD2zze0PqBUs2WBHbBOgdIpKAZBRuff
2AyO48SnKPVT6Avf313sefFbYIyc07JghepzqdEPVAmtvesnsEHXd6gUFLn9vEVajYS9nXSSGeIY
ESP4HbtlPImM5eybIrs7Hdb3EIEHundjS8wgpDPj1PzPLp/nX/qpOnXbXKvwaNF8UgJWqLn+yVbu
iav0DlDICgVcXgy+SM6k0J0bx1UkwFupY0B05Wm9uEj5JbcgFVbf19DeI1QF0U6OIBqx2Q2F68Mh
AmztXU3xym0L8VycfmT4zTLNnZM0dBvPoXoL3okn1d33bkMq9IDdL8E/v3YemRnAqmT/CQgu1uEG
h0mdqtBpPaMnd1LVpC3+Col7JdYdB+0Y72dOItg5gapYot/BBFh3rJlVvXsegQYWrpEVSthKcv7V
SdtxOM7U18YRJwbT23YvP7BZD9cKlhWigRINnd8XnjecPlpvE7WIQ7q02oyCE7PIRCD8aAlXMvze
8A/SLLdAIGpRsSDzklWxb78T0oo3UkuNDAz9ucifdxiiidM2anuAF7Q/McageWBkqsFlHOB5v0jN
n/UIeDTWnb7hJ56vvyyhehsrhn8cLOvr5tTuLOJx2R29qMEJfxRzZUN/H7WfSbC2PHaYxyTVkM1F
c2jekoKDqoCZedalLjdi4DmDr/xTRksFF2v6D2X4VC5Fenq9NRl4prN1xG7r9bxZdWISJkOtq4vd
wWQnXveZKM5KvVN12KSnfAE4ajx/QN9OBATTRPoD04emlMu1LRYUgBw0X5E81XM65xaXDftjNfMT
zBUxEudHFFWVG7vN+KhzX9oA8kW9i8eQTgH/j4FqaKOJ1QnikY5oYOOouYr+fmH/1BhuTtd6kEC3
DfNuzln6mf8xp4SlFMWOAhYCIRzbKY/ZXhWvJFCA9orYU+51TAtnzklXXSGMrcYsHs1zAuC4UYkw
jPiAVVIBwbT4ol6H2eEbBzxeDv0dQBT9YjPErsFRyJCgl4XnMwNzXPGnYZEhE35kV4unXO5OHQ7Y
f2FEwoEmE+bxnlk65WV1xxsYc9zHtI6vGlSZpjxd552CxK+wWtXthMo++E+Ko2E3+5VlffLzSV7+
DKeuI1fl4pydsMfuHAYVJbLIBcMqqKPbT+B6v3X+bSwOLojJCS3d8p+x2mNpMi+uougEv5Fjg9h6
vjFU6FA0ZM43mXYV0MgDzL9kZM61kAXlUfCRna75HCsuRW9OR8GRbP1E1Vk41BtE+0tZmy/0M2ai
DlqlWcSHBuHi/AhdN8cEx05zBUPNHCYf8HpM5tUNL0hJAIfKIViri5hSb5Qtnd/z8H2FZDrMxh2k
JMOEFBPm2JrDNx0DH1vBVScI5aVugChsTrnYUrARvoZh9pCvESVpB5OfdtDfdZX06W5wdWo8s7KS
ON3iQdX5d7+dZSwqtjIewBr/t07vPJjVU1GoamE0P0UCT9on7UlNwLTtL+cNNaWX95sfmYDsQCK+
jHJav5RTn85VuCxUhdcpj5uXGQbKCnYWS930MnY0RnW5W1nrv4Vm1OosuSi9CHPColMQ3I/LGuMv
K0BanA6Go+01oob4cTjSO/o8KPkt0/oqQ7BA2HOQcaeZpNx2xgwwj0rI4IlVpljsg4Y7mfbe/dLl
tlD/j47p8PCzd3oSqvfgF77C13zBsIVPaF0FibdDC4amA7K4JE+m578j156qhEa2yW2XW1/z28Wo
15YqWeNUxpe97+tLsuSOfUouVdasSXAeLXo6fMRMn4nFTxoFC8hhp772WRr27Jm5Wy95LO7IyjpW
OjdTLclv7vk3818CPK2k82f78ArITjlOQHptyXgVk5aPppntnUeqTQRk5L4g/g2NvYZ70qNsfhHD
O9GnDE8e99nwLrmGJ3K3ZLgxGAYXKBGUNjYYOkNtpdId6/kpgxWzM9zh9ygfKZF+WomJC/mxFNOP
I7nix+UirWkZRCi4W6Yp3rtLuqRONcwc3NXDKjOo1GM3ZNTXSGljmfCQFJl440+WOaV7by+6rtRe
HLwGoslL1tq1A2XJV6PU4FBPKuZnRvFpJYzgFJaKa4LTEgUaqlbbtWmx1+I00hRAfl00OXIspJv0
RxSi6wnsOT7tpbG2Vf1OGveP3vykyWERpl/WBgO6DPEjC/KmD2eOTPqWmCp0fFUj/m6TUifDona8
402aqAZ6PG/9SOcOo/KcGXSK2Kpj/RT7wFY3jP53nny46WFIDO8jFC81ax3gFgZ9759EhLTm94Ic
xo7Mynod1imYVHpxQPdRJwMRsA0LGOnvNcuaYY1nxBfLfpczYYBYZwr8JmBjkpoiL9h6HAxOdcxK
VTrOnHqWzBLW5DCPm7BRew3mTfFayGcM01Tw3aKf/Aaxxca8zXRJE1hRrbBsN45sb+X9NCs0kUYE
dCzTp9gka9sZ5k8KSO0pYPj+z5XyMpKTmjcb6tmz3DeHmwYWQhO78BDliauiCP7UjhVk/qmXbF1x
im+Ta4Q0dUvrtq7cp80gewXzJlYTTdqNc1Low6+/Bt1h6XkLla0wT9/kItVCLHvlD4zCTYdk8wiK
AROvdoiIQWnNSg5Jvey4e4E2MOJXQPWNRU8itcoCgtCTzz011corI7+A/0DbLQx3pE6qlbR43qM8
YzMhCAfgQtLML0DrQEJg2QZfBekXtT33fbjsIBzAW/Hzi06Dfz4Pn6G1Dl8CRkiJipSGgk/nKQbx
wn/cHcCHwm1J4Ro4DVZ2JqcvjA0sUGqvxruIV9yhi72q0z1mn6EAOPC86ciG1SI2D3wO6uCfqFyP
/D0rkSnpamKhQ7R2B8SeHPFkkTTPLGSZuuSKAu3oaJYcbtYEc5+1vaK5t91rYy5RT3YMrPEUKb+U
TQvJTH19sOPXkBZudQZzn960tIGOrG64Tjz9kjW0+m1SCg072lPJdGQ2dJGtvxb+U2mO4qbqDv5K
qbwM5Wp7fIUxVKo3VET2jdOuFJDWs0ljn5SopcjiITedPwv4ePMCXRnJ9foOv33zWtOTZB8vRAK3
uo6TnH21vk26v/nohstA4y/B3wlPmFd1r/F15dPOnl7VLbAHVcMlbH31hWX/mQbMGW07Akdc+rnX
2XOsO138FTH2w5se97OJW17eaLLuVcoiS4aLa/dWdyCxvAQUGrt1zzlz5w6BewoEXK3Ss3T8QhmH
P+J2JY/k4uyExduuQ5PNEkC7PTDTmjdsh5u4DpB+zrTbfM9Jt8jBJjgMfe2mrkEIeUS42G93XYXA
4ZTbenzSYuNsEuwoyJ3UUKsMsSeuqXFn/OJJO8YAAdWMnfc54jIpeL2UWhWfro7/CsS5dM3ggJ7k
pMw+jElorPat04z+KVOnA8ZMHE9ubyb1GAjie+QbUxUmfUH0hLDQWRPJ2qmu3XiOCpxFszMso0qM
IElRtsWqEjWv/O/jxfFFGWIIQn42b0KHlDSB79ybGu3yK3CpumvfOjY4UmeVVXHpBFEGDlLmQnmW
QUVaA54l/GG1/+WS/AkaWZyMXCdyqmgRztQDNTA/J1AT10IWkAWV+fNrXKCZ9DXSRSCkPlwwhzOf
oQwgjlSvhQqzy7fdxE1mREhuNgNqlqLRylO1vAN6P983Y8bfxP2lFoVEwfZtZRX+385mEMtLaU4w
UTIXI4WVgN+0wLcmXKi2wX6w4I0aqVStP7M4oEKHTtqCGfgwWKGIAjmkZUOV4LfZ8z8axzIHZDti
bvQ40BhZO7QybUf630ZEf69oMnKyhCCnSWWTTk/0IeZ1THV3Ehe3MKQlKHc2STRpspcY2vHW3u1I
dl8AEf/aug9XG6D0yvBzp7Ua4+KJ53R9CIyeVuwImg/FBqSunSNLo7muvtUafEa+qOUl2mqCjqgz
Tfn3pVLIC8HAT/NyFxzHP6xQmQbHZ2hcbNtVKCSRBZzecSbZY+LINpvyL11idaw/gScXJItG6MPe
nrla32VQDAC9sBM1UqhETl1sFXOWIcnUmBA+GFKZypu28+oqrxXgZtkpEga13O5jiA1NrZQ5+HUB
bszwe8UYXM90xtPAoiLciMv8lx9U4JGjLg4B3WKMKhtxdyYwi50Lwy4XyFArjE8IEX4yOzFtrPDW
RP6tPncOdHqolkk1WPS55YLPe3ooCB9LkU8C3uoZvVH7A2XiiLhbKoJAhS4AoV5tEyXTGWjLM0LH
1Cl8mLnijF4Xx+z2YDUsIHbm5/IMi/OUrTS/Swwu47zK7DEULtraXk3I0st+/Xh/X6G3TYOJj7KL
3AW4fkwAPMP8LA1ZP5jPRNFQ83T3lNvwACcCWNYnUzXqCphW/cyhzlJGltgDoXKM3m63nnZzT63p
aH+SjMphxRhGkSz1O7fBKkTNV8HjXafTUs9XX6t9X4WmyOl8blzLtEl3SqfNRcU049vLdfIA78zl
t2Lnsf5E6zmdgnc6qcT28AGjvwRxICvUDojwWZTyGFwV4lKreWTJ0E1SYwQHvttkfBxQLbD6rcar
hcU9DLQ1S9iTJhV9oXe9kXanqPoewJhrKsA0+jOlKBDRC3pFTccM8e6PfdP1hJrQUEu+cpoa4ElP
x9/AdS9jNK9kpOiRwZvP9SX4UsVq/crXg4PV2RQSKiIB8434oZS2FBSu0hvY56UrV6mkpy5f26bW
PAQm6khPvmFrKzYw8P7AuC7LR5Qf3cZ+/VrPoYQ3de+t1nDXQo+KDJK/76ncPWYCm6RL+9dH8s5j
0CIG96cze1f204WCC80/AyZaGWiM/3/q18/2XZfs6FR+yNBl/+KIsdSVqCOyT6xKGc61JiyKmBom
v0c5QSXLYqRJGxdYu9z86irhqpzPxPlyMGnQZmTcMMudy9Wm+sMRsBJLNKcLjaZCo3sX0YQOpp01
ovW1s9nldCcjz30jZTzmbFz/z4tzayZzTbodz+8n1GMtltzh/KPUjDFXa7/kOTxBU/3eIUvY7T6j
UmrupfQ2iV1lOlZFpJW2I14SPQnwObgLGL3DNmNRi6MVDGTp0VO+Z7WtHNmp+KpD46AJSrb8RHwi
RYCVB1bvCFrye4dMJ7AyF2bF1cGMTvsz9jZVE+KlzAfH0rZ7TOuEzAUNeuTFJFmpdvVVL9zCjjAM
Q8owYMcoPp/fW4c6ki7DvwZp/ANcscjouJ82DqoDoi3KBQjk3WyOlzEnpBdWn7RUc1BYlUWNqyUb
SbQyqCLNtXRWJfJQQG0njlOBjKpYVnlgNHUoQshMWF3u56K44nvaUIKaEOGvBs/pK/oqtTG3DGzU
jE4k4Cf965gLCqC9VPau2rz4d6j5im9rBrYhXyjiWTM31OC7cBmx0A5fC7ZW8E2tLWDKa47P1bhB
B9r8215eup7b2SYQE0P4ynjtW2XVwdHCJdsoLjahEHJHpyMBol91AzOilNufc/64oZbbdOErAXF+
TU8jpEtk7uqD6lV0YIDoyoXk40VPst5CNBp7aMC6QwM+Lu4BthhehZr65IVeAWYkDu6VpBnvS1H5
1UdgITUO4pn5yOXjV68e14tVoVMgwLkufWW+zoBGdEROL6LlFPJeWZALKUk0Hez7ck8Ckxk0D2ng
qlctyS3uMaLJQNp2uCO5OhRoAjtsvxc6uCaA8pU4sDoqOn1qxeRm+BrgfMx+FSjfZSxnSA4chn3D
Uzn+IhBm97CkbykgzMhMo3XDshjwjC35AkrAOPMf16Q9dLd697xfQRqx+Qd20c9bKPiTaT9mzZeh
o3Jwc/HJeuq21UTwppJ60UiYVlYqrtA2CkXoZLF6C8UNCnQjpeJd4mVt/Qz9f+FW9Do50zVe03QT
AzD4i+5DoWLts4031EVnelO9/yJOEKgJ/bV6kaBuSb1aOYjTagESJDBOpXliii2uu/ptuAFKPyPN
f7ohOJRNqHRcU5+Gjseq2WErLf3LPc95F7hSKjAykjsSy+V3Eaf7ImyWAmqQJGSERSwjMLHSNwiz
aov2qV3PVEnrYXLT8nnropxgxPbWcIrimiO3F/DkKQWvr8P5q+NQz3d4Nf1ejgconrafJgwNTH5o
fkX91E5c5JRL7AZixdlKIGWpV/qEABiiPjlN4lpAj6p9c2lqrf/f+amSa45IXE5SgZ/k9LHoLfKO
x/pA7YgF6Pmm6TPbVQaR6NCzOoiMgFKnTWOwzcDRwoCdS7uHnq1RehWZQjISS3sPRHedt4y/kiG5
x1sshvD5aOojLFKKPZHOfX6cgWeAEHcMTHjd4hzj1p4rSRxtUCxuKmb93GFK5lp+EfpyDSkJ1bLb
zzb8YGHOyS3v5s4uuGDLb8j5UQJgHpfV4vvQqYc/BG4X/9lqtSK7XZkZ+K47HxLLx2iwGUSt6blG
4NHI3BiaWwDC+moKRmrROzz53Dyk+l4UiGD3pfvR+YXyGCwBHbGVrFwlO0vMYmxiqAw1RScfoWPQ
C2kxIEymHoundvu/2ttMNjsZ99Icz0ZM5PzFE0Tkc9+ZWMACHC38YnGwGfiSV5ASFQntmW3fbHsc
S6nU1GbZ4XlgrHlYoSVkkvuN9Kz/cRm4Ubk/HLE1rVC/xuVILq9NAoaLxPvauUm2bG+IYMkOgSXu
+vWR/eF1WSRwJyhbv0dZRaFsMFuro8fSbSF3myByJgZ3/Y/M3mx33dYBpwr4brGR6E0Wngi1j7GX
NqRAbug2bKvHWuRfbDy0Wi1p0WGOLCDpp/Js+sTGzLIhZvGFqDlZT7cLmm3LKy7G+BUaoYuyZwKN
nmOOQioiqvKMmTA5Yrh0PYkwcMauMNUlRDdr+zCiHo8SbnIsuzU9MM9VxOtEYYl/x2d7IjnvzKSz
VKsVYAYpkT7NyYJ71gr2b34j0sKVWlGMrZpHQtbCmEkDQOUOlnBBeIxHeRnoZeR40WSyNPjULt3l
ckTH6c4DCFGL0WP6iZtg0V9XVbs68gSv4Q+eRUThRWKLNbAnKTY5uUAvTVhuiqPZrXUbKJtV72/r
jjo2pbT3m04s+n/re8hPubBIn50UeTsRK9lMg5yX9rR1F/hUi4d38q72Whd62zF6m4wP125j9O+1
TCS1Q5ZsgeR3aALLYZtDPYKNSFjXu3Zmjin5TzLskcTogC4oRS75r8h4eTq67verNnxJs31lXpeP
9zIcqlmK7V+jI5BwLzgdQH6HZZObMs6DysUohvXcBGcFZ2ToyGMfvLfKzWOSoOjjfk6y7cmv4sJz
wnwNr7zFoFLJvsKYnv5b5MbpMxVAwMyzrG6+g/V/cFjo9NK9fv02VZ9hdewP6CAp55JTSIyACuT/
VtIstKQZs8uoSLy/DrTVwDF3LCYaj60nZrzw0/5vhQ6oMC3sm9YHzyTyNZ8q3qMl9+ajfUM7ihVf
7rR/L2atisqf79aQZQcxlGWgRCS9z0TqAEm3whozbSeA219eCYtM63zEhfPjhj+3PuEuuvQTwm+p
E4/cMh918pZ+rDbvdej6gYAWbok10winkiDV93w0fA67fbCqGARro9959SXhfX6gARyVeSX3EbDV
ZnzCsjHGcAGepJ/P0mn56YDxSeWrGEIOR904PeoLDt+Ri8pdmdP01RU6gp6ss8L/o+hZMRMRNa3L
drWtdf2UqbGm9MIL0sam2x+mVq3rRxEtub0Qd/YBfubEE3Ut4WzoZ9t2aATwAuKn8B4eeTJ9HVYU
pIzHp4LN6imKkqAHXj6ligsP0QMa8QtN5AOPdr/CZNdaFsLj3tomwSxhQKYQBfhSifDa1m4TUwqk
hb50waTf1Y0ufqWRaNWYbpxlcGnM5sKxRl32aOApbsV8tQeaxUorP5xpPjEbnv/Ip2BsbCEDj9nR
Mm+TKwhmagRKylWEma23KnPnW4G/jCqnu0cDmVNb8SOK9o6dcd0hxr4s76bv40++2CgtgkFbH3aX
AcA33tWLiatzW0UmQbpvZTQzDrvJVdHmkDmPrrQTNfPiMxwVRai1ZFSgWiddjfJqi4lARZ8b6w09
emT+qAP7AJpLk52kfq5DSEa1G8I0ZrIUc0T5EiSD5I5aJ1/ELeyQ3pXTwx8IPNEun+OrUepmMUHc
CZ/N3oVIm3q86uey0cIjSJTxiUQOt1Ht8KW2zXB6PglDZwIOJqWuj+ZccK03iCkGYzwG/b02l+Kk
+6hcP9FlI9tkh7rMSzX6fx56eJnWefbcwTrsXBgdvakwvudMhFzX2t5g/YaJYPWujJlNtmklCEie
yQn6uxGc+QTwfEija4fPj7gROTqmvNvGa6PlScnhbLXQknCoUq4Yw5mJnE7aZJTkxiXjjXHzQkdB
u206h2eYKrYzyXe4GrKJnbZutYBMfkRliK+RVwjrBimLD+TLLfnIIITmt7agT9Wcg5VfZgNZM0s1
GAmheKXJlgiw6Ai6y+0ov+rbqLHVMP3r5/XIMWpC4scix5BH1aJpn7XZffjzJtmJjvlHTAuxzDLl
gAC+YHDc9SrBWspB1lmQkaqkB75x+onpDO0Z2Owgeqm1KKBQhrHnj2xkpdJBOLEWAmCsk3+1ZvnB
d5/p4eAsd1zu/G0xcqvssedywgzyA+viliBxICbhNeOFwoKIDki6Ll8SpXLl/Rf0YzRryuQzHOr3
sKwYK5hE3QFqwSrH8VHj/9hbgH7Aks9QeL1CMuCHdaWl8E7Cmw8vuTnUQk9AQ/wMxc4IyGG1d9OJ
m5SfDXfNfq/oPS/Mkc8jSybTt61ejeKa3GmvoKNw/G/zPdni9H8vIAQN9Lvnvu4HqWLSyvOJwCCF
sSMflP1NWdqS605l6HvdUnD+Eocb3h7rhdMn7F6IahsXNkJXigaqIdlpzg2nzR27O26230TCEEza
SMJfx6SZuSpYsnxUuVejUdIxY4UplMBMIXnXBTlu8VZBJBM1/li8vojP/LhjLDdNxCnN+qv9CEYw
pRfNtPr0b2IMp2m+50Qnu3t+PXvrvtsBv4vlnjRuAHw8PJmDjkM6bJMjrGNQfHp3lV8Q46cfRTym
8E6SxtFCo2NcAKVeYq9NMbtqK913hr+1q19TBpHpMmkCuyHKC92CiX5fXhG9cA3WDepR9I/b8iHA
ugROLZzZy2XY2d+s+/pWMGB+CpoyBTAFZznkOj3O4gAGu2iq4Z8L3pAjrkPEUuWUNSFUzLeXqBIQ
AsCZAAgwLkE3m+TPjcblcpwHOCw8bR+2vbygIN/J3gxDYykZyqW7G57H/3jOkfmzCXKYxbuKOH3g
S9G+lxBCfE/ea0oaY5ZSYuVkL3+1E0c+lRwIzChwMIR02DDGSWuZpzlFEg64GvwWu0OQebE0r9gS
FPO6GOY2ztGgRBpdMi4vmBxDZEv4uWFgRu4hw5O1/XEtzayGxBAhqEfeRPALsEfEO16BbImX+m1O
UxlhNmPQxwQ+9o80+tgTGwds1Oja60H3IkDDtqHywjeqfKb17e4YOJH16cgVp9MKXZHCVNUk5l2X
wmnZgXyNGhBpHgrxV44apoiT9dmlzpG81ZK/dAhgOl5HJQN/SGoV9l3eBZzYaiFigVpE2VH4WteT
i5xwd/gCsrQpB+Y8Y23PDGoLzkQ2Cv8mVhfg/xH+zFBATHxTgRCFnDd8NrW/z2JGv8/thv1Skc2Z
BwY2i5AEjKZl0IDz5BSN+R3pHmHphaoZcbO6HdETDl8z9nHt0JS7m0Qccg4L0saaidmDIw0/1lw+
e6BQ6jRjtvC/muQY2jGuR5FmAVStZB7au2HWZskfdd4NW7z6UCnXdD6jiES+Uk1S1NTNPu3b9goY
ZC94GpDmV0NH8vqgB+aPnPSfIsSGZES7pO84KSTk1yCdm7EhmNxHKcTcBdUiCGZqd+gFyRFVEXUf
od52TE9O8DRHHi/+qcuRoNVU7VQUvjqkIJpWE8LmhuAWRlqu+2sqveE3zkQNst9lyihFUoXq7QxI
iGCY6M4E0N4NJVWiXvpkdqTi0GF5rjeeCjbGJSxKGE7nM98ZpFT+cbV7BoChhjbuSJczosVtUWwm
WTJFipLRu8LWwapjJMtH3tk5CG7KTfuMMY/U6eHU1NFGU1ddhA8POSCjFfJa9b1LkE0jJNcUY/ZX
uwNqPukhhhfCkNmn28WO3PG1Tsn3S8tgGhSWm460Ph6lS5iqJqhDqjSX17JdaqlMCUkvhnI863EV
UALKUutWE3R7oBKPktLV+AuumOsT7jSGKSS0E6OVoN5xlvVZCtg1P38IRuYXvMMzobPen7+FEqP7
TkMCK8RiUnLaqT3SNWIrD1oGduQQBgWwfEXMz6EjeGud1vew7ftuYsONiaae64kTY7vzphnNUaVz
zEJAmO6OwBaEUCPfafAsEZpcLs1XFPImjXZWLbPAUJz1+vtRhCFbdHlUpdHtrR4a2p9cUVyc7WpH
02OWojdLs3efTlLRuu9Q3/VKSkjxN0YnP9ynC3lIN9Kbah4LV6CeqFdxMLBJqfg1z4rDsS8PfpyS
ozQeOgqvgDohQ72VAy9/oZDBu/HpkN5p0ZvmqgVJflxNpXzt13UcUw3r/iltJ+5uMbVCjZ0L+Tg9
Fwuxtw0raoWfdZKiyhsrsKBwQ4umX4us+lrWxTNmD2GTNUplSq/pbelYlvJzXPR6crFxj9UU+b5l
WJTyS0lbCy0QXvs25IKHLfgQ1Af+DmthR+PHqRQ/+/lLJzfNw+hTAZ0AvhwMCDK0GeNK5lqYr2z7
GqLCkUYFQPl12ZMjoeOS+zs+SlWo+30fk71VN8+3fNO+VQGHeaM3GEc2N8QJmsbR6hM1k/p8NU5t
ZbYCH/MKi+ynIM8msfEFO3G5PLcp64I2MkVnlvRjQsrNBtEI/fYywAeJLOmjSDSZlHLroKXb3qiq
vOzoKwZhYagsZnqcB6BoNQTX1NCTCohre7pD3rXZYmH8GgA7hTWeFBsjIrTLwa4jzqv5eshxa3e1
n8gBktF9hFt0M/WhscQR1+UQpPHTfaLndT4nfGsFV+d4yEGZrHLTkHiBgcI9xhkSrlBDX5UJ35JI
e6a8VpML6ErqvmR5X07+or4L1qHquRIzGId4BE1IlZdGmbjokAhjBKRAk4fezW4MvaXXonFeEPRF
bxQXH6D0Rdpx8XccCbvrSD7+zUJA+yE7P3bAclZAyvMxzC5HJYcBqzRWkaMtiSntQmf5VLwmq00b
sJdpF2l5c6j2u6+C8SUILIioiyeaoqRevk7Qg1GLnjhkihsZHQCQBvJKd5CKNdhYb8SzC3AmV/ld
GjuBqFde0FC0zqnSDzOKlzatnEpBAoJ3vARR2mCTS+s4mhyyQPbNc9FU6tkoiSoQGpW0PIj8LC7W
YNUL71aEslDcJeJRSoYt2T+a0BGDJ8z9LlxahPdHGc5+vx5pjxRUdenfZid6GJHSr+gPN47vfzfE
ch0mgdTLIe6nP09YGpdj1HYCQK1meASSCIwAlH7tzLBvWbMtzZcpy3rg8q7DMw/jwVMw6vtkQeGJ
i1vkd3HDbEEQsE9Qyd/q9Z2guOYgRf99lHIlRab+VV11Rw3ut0VWWtPMltYXXkTKgXKbx7wxl8IT
AuAFJZVM7u/MeqQGuYduc36KPUNKCPaPxjm5K31FkstItwEUGRu0plrDX0/YUzpk/j+Jx8Al0u8c
pwnxCXGJ8L9RZROdAyBT2iR8uCUOhvd6kdymXxI9QWkILvn7CAoGqNjKudDUTdfF5HzGI+y7rdqY
ChkobJmokFyCg+NjBg+F+LSTY4+oGlg79UccfPAfHdUooi9cRpQqD3hzYjfOMtzV1JgBnIIuSfa+
jh9IzXSWhP37BZBOAJMkKYjs6WyWz+uM8ILNxOCU8jW8CDvxcc5TbnbySLcKQ6iBT2yqishFxWPQ
ACQyS/GI7ttlsScZgtPirYalCKqcJtU/qsnrzxD96YyTY6PwZesvogS0sn/YECucAN2h5SnH0X0O
ouZFWJ1npNwRX6/vKFHHS2u5J4erolKvjrSx0ifFCBkUUUaQfGFtEUCl/4xVyXmvsDcA2LB/GLmJ
lP/prbRTeK7WMq//xl49BurM9/3sHEihvO9xw8l01xrw1F78AygY8+aPDjFhulKW+azmklNA/z4z
CU3BiLTVMLuyos/vi+Y2KobMQerfMxmRwVGKBGp8Cu8d0IUrrDmmh1lO4O48XSVb1F6stWBnry2K
daVq0IWKXmfGECwAmaIUTKngTml697wlSrLKiKMDyjnJ0D0P7KBKrWvW6Q5a+eow8+h3mebUTZ1B
GGax8QfViqXJ40ZN8VM+VCcAj11l9YTuqpxMKTmTP/hjy4PJtGUW8G4k9mh2T41qxHHBlYwgRdOV
V72mMbqCX/Bvb/Nd3WBAj/Jspx4R5DwOh10sKVXOpI8CaiC5A654S6HULE3wzIa7sTXwuPeZiS82
JXInTYNHrN9QaAL7YNG9zA7I9C0o8gHLqIUE9Yko+jPwpDaihQrKENeUcKmWss8cMLBhEma4YqUV
vyxmG1DBEipRyPEEYy311kts+2r0GjQIjuOa6K4YzrFJaWLUxTB40SqYktwQ9MVV+vTrW7Y7BUOg
pBhVJF5KxG/ml9QpDndQ/36xcQd655DpyJB/ux2Eb8TIu8g288MnRnc38GcBljQEbJxKPOLtGPQg
290STn5+sqbIQF0k7boJwOxsb7IRQAWQsZLgplquOTztbatt61Gfv0GuQ/mdL8P9Hcu9HfxaXqr6
ZKV/7U4netueSAtVNusjJAR3/1LzaVSyvUQWjk9R/NchniB+WKuseUF0zs/NYxWOpLmWiP6Dj5/B
VT9Lboh0yDd49Tp+LLWfVy048P6F7ZemG47QrqGjmkXtO+9SUX5LxvOLbVj85dNg0jfjMJ3PmHGY
Djj6JbasqRhjHVx5nt0tvlpWR6hFuxjwJ005XTIz40ewiONpAOPExqpqv0etOrBTOol+dvAsihSY
cMtVnMRuBo5eKkareDvxILTZUkFtVweui8i/XgQdymb0aAFDXN+fNtqiTB/8J+O/YHzbNoQsUCK9
KB1ftkAaNKKr8OdPcirKHVa+kTU6UVsNhZUrEoDGqORVCnQhN2dnEku3EQet0d02qkgBAcrY7Zjm
eXeW7eZGjpOWt3vPgUN7/wrydzaq2mk8o9oW3E85DQZ7cnnAnKLbZxT4UYu2M5tuiNu/bAGeicHe
vB4bl+fpF5svpUTuFhqDf8UVi2X9XE1xqsbFbDd9taeJq0S3NFaUBl+RkKsCidtcGqcmzw7bj3JA
kdxvLE4xAiI+oEnga7ccSFEb9zfO5GnUhcO0TxfP4B7N482SOwwxvjqigRYC4H3dDJvIL6mRjn+Z
YMBJnu64l96TcR+fyxQ9nJVAEe1UbmiGy+QmhZzRf9J4UfSjnLb5LRM8YWxmzV7gWC/H2fqEKjcE
klw0oZsHYB0V/Yz946JrOhlz/WyLNY+9d+QSFd+RJ0NgB9rHFSbOos3KBQXs37ZQVoI8WL/dXaFp
I77vygPGCG0aQ4DJXr6ZHILAlom47Jl7BAjPutMRVJPkOKhu8STCVkZ69ITGpsTxoQ+szgCQbvF3
5KyXkX33Q4QOyjsTTRnf2wF4fj2JwMmupfF47YtY4I625APYr922Zew9NnLz94RqxGEkJyltdDhH
rNHB9f39oLu9bM/fZGRAvRcH0ssQntS/eMtrHGuHSVcnMa85wBrIEFYdh4NrcTku9moFLFfRqEuh
NWGtAs3zNrInAyCnQF6eb/sSZt24u4LnBka1FRYQtknDV3hxVa4+Lpc7Ufhz7lFOcA6Rr4JyJstE
LC+B/z5G0F2z7zjZiqouOwPQfRhyit3h8AK2PGM5iBAVA9CHQkJuSddq+6AySTeYOXv8IGeHRh14
K0+nlV2aNQJ9xLSDvBxc1wjr98Xif5Qjjt3umiKQvEIdkTMCIrr3J4JJ/EjraLlSlEwT3rHpDfui
wmi+3+e2J7uoQ0Vm4wyMV3+Hn9gqs3zNxwEb8LEiN41P7zx/Oia1oiPGkEUDJOL6rbvWFX6SJz3Z
DiNII2zsmcpiwequ3F6oQw1+Z/iclBxVDMrCbl3lNx2c2sWSGgRxNaB+LjJ+Ap5nAQBvmr+MVdAZ
raeU08XbADTQCZjLUNm53QV8sPEdqlDbtgnGRe71Jp8dclyM1/26qC0rVU+k6Jnbhc/YDgPs5gHH
6KtWSZyjc2Aizo5hFmwvE07AzcMAE4FbTDxqGrP88Z+U4pXiaoUoG8DrPKBbfZmkBAV2BouXHLF0
GwjyQH7Qv0kGwwjrUsV8achYzslQhX/8EP1KIOsbpWaQL7glxSDH6Hq2NHr1VjYtKljQKtObazFe
7HypiVK9uHe2EZqVlaaMzcYckg+D6V5/F2pRmIOHhzKMyBuL9mgSgEuSEu+XgXon1RGk2LJlf6sI
KFStwT4SL0AcZCo8QvC2iZQsxC/7wrbbG90lgHRJMDzC5/rT+nCMHBegYKiF/qyLTb6fHzJZTiTN
9BYOyIkdTRDzheDxOPA2jyekotbIoN6TmAxYQS4XE/GatZ0jcKRukWkooJwR1XHlj5/wsfe5kL/K
c4vX2cHsO2Bo4d0quh9W4sIzSyV8Y7o9lqCFGze4W0Tm/9jO3oDhC66KjCRg1/VErqG2ts3G6WcV
d2g5b6EwQ4U+fD29snyROhgRZclFIz+7KpC4Vk7PqHkqDFPOHRBFOvnVdR0WFaN7LDgsBnYTiOlD
uudc30N/oQLfR/v5xLCtDsyV9h2A2yb53lTQI2WzTaCtAlfK7U7+gj4z2+gRL3fwxrogHVa92CNi
q4IYRscq1HDrAt8kSqab6KZ1wJARbpYsk5/vSgIcvFtZz4UNBEaGcG+gjoUEPbjmEVnE4YDtUF82
4k7+5+FCcs5QCrNIXr8SR1IQIGArr48Rn9VSIcCZqdY+YP+YZ46yrPg8PSmUuA0HPQkvV/W7jPJd
FWrSuIz7AZ8NhTb+JkcDwi2OaPvVLI3Y/eNpWcCXqUYnrMLw+E/jiDTT/d2W5Q+5clohykZ+EkuX
/iOfJruX4X8Voh/sf887G9+70lij22fM4gBGV52BBPj03j/bBZLMaDTQ1RpRK/AmKH/ZlZXzzlWt
zBPRHp7+/zM4LS1HZe/2ZpNrMaR0K4s4L/Q9S7AuZFaOqnYOtNJRnr69ZjdOO4UOK0PLzIlmyvT4
z0ltxfULTlXtJl/fgZO/yNY67L8UtIhkYytFry9GL5Zi8NkpH6cCQNrRPorTvPEtZagtNNpY9WaF
72b/qi2pn9KGsC+7+jFWwwDyLWnhM7JXiN+Jj9LcdWiYcOIvtfLxUsuwxr9qxV6f/+U8LZvJEKPR
Gw+Sfqan+ccw9ZpAVjT8I0XgnKkpeqxczlCl75KC1n4Pml49Aqix/fxF7DmCtpoZgzXOhrheWAKN
IsFgXMvmeeT1CmV0xofRyW6YeJTH4ONbqg0UeL1TuXP7mOavdl6JfvOI4m6qimaxTMyrqEaiBCG4
C5ZdQ2kDX4trTRmboYV4sNyten1KRwRkVIw1H2AJPEhjv8GgE73FVSjcz4iENSrsYKd8jU/9Fyyi
PZ6ZuFRjgrgDm1VSwGdoA2mEZDYVaHJtnl89frJMzbi2OKSC12uuJImXrg+RowGm1vrpylXezbLt
dj7JMQWwVAzCNOvVUTOBunYqrTnfVPEdaisy4q7KAQOPnAhTnYeWzSZ6vuOaTQal7Yc1SsUa5Vz8
09vp+vN437WQNO8Srb2AHKDbxP+m02wfGQkq/gnJQlKEUobqlyegLvL3bjysVmvva62ZFlDrkcDp
1nx42+Fs0jafLYylYDH9FXPYBMgbfRbjqQFE8Nntm9qGfad9ufOABDD9fHqWUMYZerPdr8rz1eNu
5i0AhN6HbDKJTmiHKaMh6ahW3ZJv9NTuDjONsWXCBFq0E3v/D3ISRlhzH2p4cq/YxiX8yT6WZq5E
Y6Xt90PoH3RtVa6TwEQW1D4uRCt492tPw2wsOVV6LpNES9UxxFc8NAne9z5EngcGA/xBT9+AiOTJ
q0cBqTZOYXYxlPNa7FYjGd2AHFk2o+5Zwpn3HfZ3fy/k90Jk5RAF5uf8aFuJi+U23dfyZHqVeSHd
E4o1DaS1kzYj+9i6bWM3wfDjvXD/1C0DpDn2cEjd3KX+ONvptuEMtWA9AgHq2pzHQMfc72Plyhm+
5j7Z7iYI1hYYviZ6kfTQmxH6hLygfyY/k6Bn3rJzK2y9HmhxcG6tvIPSxoJ9UiFoOOwl+dCC5dOU
8po7huQm0yx4NDEGWdFRIljghF61q3h9p9rzdtmrZkc9Jfq1Mx388flKA9svsDsPznXXlyzu1915
BtdrA09aYIGCgRwRbHfhsyljUyRHAo8rXpuGVr/QJ1MomX7lqsEAkxwOojUht/UWJjfwmJNxAK0e
zcPdHVzzcjjOz1fW81k/c7Gz0HWD20FvIjTMVrs8vwHMpd1G0v9n6UKfSqXRgM5S1kyNxalDuZqw
OxwV947d22gAUHXRcYCscWhGxjfsp6rpcaW5YlJ+r3evSKLhLEbQ7Z6BhaO2YPhkHt88PapmGLrx
LFqd8yW3ntDxL56dIpp005+b4TCelsTaGBwkkh3UGf9JDvEc7srXXWBoidKB7B3dsJc6ADS9SMOa
h1jB1+12qi2A3nFNETx7dlkWOjZdy7hCeTNgyhy3WeFvshUHFm1mOSA8W2M15SVr+if43NpGRQ79
/Gt9OCkflbZvOxvlsmycukgV4EvEMqDbNVZkD8WoJ++IXkf54pCXuRaS23ViFFJs8n/9cz3VAfcB
3WWBGhMElm5RjfhZxo3nbC41NHCv9Jb8mWUf1hml4uHzKH7BuGKXQU2kD/mnUPIdnkV7TQ5+WDRC
UeiGZGaaXMcrc/ol8AjUZfl7vjs0AqjmCBkUrM4cjqJ/wU8/wv2CQqciAqTdch30kdHBJYvBIVlP
IjYywsF0QMP+hgdnceC5iyjJspZSr2Rg/QTjMl6df9bYl5z6/mYV0j3KSRqsquEgc9qkdnDBt2um
kPgr1io/d4evSHcquk/awcFTJw3CofDCLDWM/4OIFzM+6i+ycVx6py/6R5k9kokSVMzUDHq2L0Dt
yESbg3gFYr+qBoX7gmet3a+PaMYYk0s7fjUzE+qk6uV0BjiitS7+KOPIcFOt1ZadIyrNRGt/6XCj
quXf9P2ozOOKWR4IYKE7pNdJgb/bvxM8oYhpxwFhE959TxGHU5cb9J7IbhzZPUHjYlPOfeqJmwTy
VMPAGdTmzQSIGjRcGxmBBWelwI+AZGQrysTfuNM2r7uqU8gFcOQoKnRKfAuGr0bn4ztHHJu3TKg0
CBdw3FuxWWE5Vj1t87PUSKRgUJ5pGmVKPlIXrmJAKeKVCbhR3vEgCevD/S/54yrabuVSIqvLucdh
+rFqEvPuqsxBIivItDFFEwq369ismKtc1suTEwjUb2NSciHihi50HNp4zbML+KLMX24z7kkPaPCe
O0XLgepmhDBEHy6/roQL0kqzdM7dvy7uwC/TpKILlNczydX/Rl214QofZccxYYSBj/LORI+he67b
gxpV2VKR0QvyslxVP1WA37ayMYSbNpP/MLhSLL1pclwA1cGNIyq1ftjdRBwh9IPjkSoQxNaqLQtz
1Sa7bWel5ZimyGNRV4+w1gnmsFupTm79jaS02Ss1cRvLobQtDoQVyorpXrQgkJHMjxZzjkwfpf/Z
jeNepAApDMVPC9eami6+Cg6yBt5JP3+4ZHeO/eES/qvqMoYgwnMEk3x1OtvzZ0CDuhS9RSs0I5YZ
3IrudCf0YADB2xmE+nnagM2Wnb3//m2YmkN0alN1fF/DHm4cizlRn+MFWSh2hwcMW71KihpbyPZU
rzYIPEBizmY6e34kQ9lSF2QUkbxKnXO+lGzHk0GYdDUV0E//b+EFkzJ204x3cqYAnQf3Wl4NChaW
7o3A04oR28VvxevNw5hKQhL47KnQk55C0S/0MOLNOvXFhymbx6h8dEPnp5aAXWxFEPCDBmMRSysE
LS0CbOz7ETybl2XOs95HjN/ffynqBC89TOhhg2IQPoiht4qB6OgZqRIyLcSzzOo/LM8kGxoQ8dAk
6HMbEW7sOe3kcfItMVO9EulRZUpqjwLUSfSeNRsPx4gzgPcK9XFQzOxv4lS8ZsbwP6h4dJPdc/Ck
Wm0RBxyamZJveVS8DKKuYqCAXV6enRgJJ5LEesBilkW+N3b6hmnWTWL0LutEqQxMBfxLqLc3gk1O
LjzrzFE797Deg8FWvjEMflYd1PbgfwWiJ3aWMVJEPWXKT86lfYKTkGh9MHhkFq5WismDb2m5fkF2
KeMzquANBT6rOrk2BNsvmBh667piARtuFSNWEVz+Ip01METiqdfIXXi9X0x0wL9+9aG/gWDlfLoC
SzuybWPitWrlLZ8y96RKRuZRgbd8kqoc73feo57v1FJPBy52Urf/YXvo03iybdfDMCKuGDuBdU4o
5zoNT/K8g/UYGsfR/ZAenqCHLy4TvqsrpkA/FB7D/WT4/V1r0MzZ4vviAcvAZoXtYV5yvuvfFCuC
bqyogEN9M0aUUXVLAljChCH6HiPfTBlPZq+llRvQ2StZj/D49qkiExEa3vVc3e5fUbivAVkpIFL7
TByxQml/4V3a5EuqaJk0CBopN8ttI4oNfZH+MKWrTNhd5pZQEpw/Kz6lJ7ct3mb+QDmtHET0PwFJ
bmQZ00YPUbri0GsJzpen5MXNg+1ro224yHuhOR1KBd2koMdryAARPwBLvR54lZJ8WJrADLEeP3Xq
yj9szQm317ikp1xgZHGB7abXhxYhhaAFX8+lZgpA+0m3OOzbsDCnFNwae5tAfteMjQGZn1lxQ3kp
+eQoMwsCR1Q2VIOL70VM9Vu3SkwUIxGHO/AXd5WBrE4xgPrqF28v+xasRboYQmRLfcmRz2T3Apfk
X5exQAiLnj84wVo+3aEb7YIODO5+H9EtSul3VP9wNA5NH4CbjfQDaLxpBrsNrUdZvG8zfh7FNGaa
qV32wN/9H3JiLDyZURyRzGvoMnaELKiQMHIEi+LRvRRxsBVbqjmNKAGN2+CXKtFhwaqyJ+O74PeV
TR6VfpCMIgio8Pw0HWQ4cdSynN8L+DaQKmDBqVAPADWoaM3nCi+oY59kCPOKhoDmDUVwsPIk7PGV
IQnoz36B7dHLXwMJqlSp9YQHHPGzWtgC0DpB1Hpb0SqJ5rnVMeUuxAZtVK3bJETz9474m1qZQgl/
VQvrk9frKFiIBwqPKJYmPzV0fL6IGrLMi2yeJt+rUUAbjVA3F5zc9vdTq4gQCgUv2rF9HDWH0mM/
FjZDsqKhsx2LslXNdwyiBesHtHL08W/qlHlmOzxLymteNqwAwPz8vK/fD+MTk6J/C67RJN02C8+B
v2GAsffrL4UTcqXB9DkCSkeOZ8VJ62bDshqFsZYMnSj48BcaE55QmBZ88fOHz0xgAm/UZgvXcnLi
KbDQbkUy/i5tDsGCE6Cabe5WUrm1rVI74kVfcz4STHvj+RhoFxk7GFz5Oat9i2r7D19XCrDDJNG1
j0ScXRvHDTvinA59iYoK6zGvWDoR6Dfhwvwtr99rOLC3Mkl9Ggj0xZDT0f6SXbWR1XccmnfjHX2R
JsoIDK+Anf2p4jkVMfMxnzJVe+5CXy28EbeM8YMVm4bgyiziJdoR0eLfzsukGETYqieb9pccICc6
4/JMq8p+6xfAZerGJToWc5533wIXTKj3U39uzYAm0x69WfjzUwhAunlk8r8s9u4SM74n5C1WOvUu
CQrMD37iLDan3dtHdJKbqygwKgrUSxbjXnrxnVk9VMSAhIHjc737Nu125nJjTSgKLE0pIVBTj3ka
qRq796h8Wf1WnlAZeuK5qKgsPLB1ZlFFH5jKYO3MYFxR1beo9wYDf+G/BnHE0BOIYrjlCyPAaaBv
nAoFxsOWe9ULtmfBl+4jN4o4VeRsg5A6Uz2NZWsN3nqlV/XaMdjE6l2yEeS2F2tfDkEY3WKjSSIO
SiDnHj3uz74bQAUlD3Pc33DnqGcCygdSfwf2XeOYbsvbSCdauxEvsz7MWqf4efzFoA9e7tZ+8wOU
hKjRpWgDfPe3ljWBAxd+jRZGSWOec4bqjeFdnZoL3Iwsk7kFvaKyjRZewQpqTkd8q3lJl4kJPb3D
nHRTCTU7ewMh5Z3jQypOTI6ekv7uVVWtdnoRCK9sQR9U4eBDj6EklQxCNjZtYebJtalulcJlgkB8
Tp88hrXxjz6GW/OFcFtIgZleT5zp37viwmOOkU5gimLeYzOmcP68lNt+PxvpdK7bz5Rtx1T1HDnS
mDKgY2MI87SXziT11ldjttP9MrPmx4chkFpXSIv3Unif6kqUiqdPh9S4k+ciMcVLTjJm/2A3TjQ8
OzG3/AlPZ3GQLOliKV/5RQp7DhHcPdI9VspA9PWnebPXVBCKrUl4ozr1bAKh1eVnG5iE60ODW1va
smxWLDWNoq1WPAgKPzb+zltXj34YNtBQzKPI8YVIE4j98cJcDkvlfCBoAMLuOrTZyJDxaxtUuFUb
YQCSwbTaz3ovsXlZ42Zvm4Wg3CW4J0jn7Nzcb0E1j7gSMJtb4WF8ahs68I1VotY+Jd/NsEEQ0uWz
HbOdRi6fTCl8y2iuTFP0a3ofBsoUocuxy/KXPx3zzuHNMfJFuxkas/5RInB2LouOlyfqK7YMqRLF
qaLhtDa/kFSkUeaLSsKqjgscLhQZmTmuGks1uPg0dpgLLbbiPTCFqw9YDVRuMi/7KLkg4zwQBguH
1TMr4EnHR5DI81nYqI5lXDbiM+gOhXBNr2l4a++0wyfQZP1G20eCiR2D0ZmYinY9IU8dopMtgroc
0vMB6+uoCAXbcJVGP6iqVpg512kZR+fizcy/NaQLR8xBZEy289S+34QYjZBA8ngPEX9QD+Rbu5eC
77F5aGb872Ru0PxjomwDvJagvE9JVrevBevZq+qRIasv1+3NoJ291mLb8ptOC2VP7A6ffLU+pIQk
eFt/gwZC2qImsN/uvdV74iUSIx8JBdjwcEKVNQ51AdfqyUYHV/wDzvi6II7hmOXVUVaIwJ3VDOKO
7EmJXCxG6bHuR5PAtwnTd2yjhRXpGipcC5HdVZFU3Z1sF7FcreO2f5V3gmiQMZUjDS+pvk/Gq6Cj
oViuEi7y9Fs47lnlBj/BFchvw2QqB1xaF43M9F3OCiCiSBg3zBENf4qaTKia5D9TqISRe1JUq+g5
BNT5sKm678kMtMhTuLlmfsV5FJj/jhoCWSO9Hju4Nm5VRc1MWCB9UP6FEQWdK/Y/bI2xoZkP6kVU
6jEWv0j4aj+1xYOUENsL5LH0FOV931aoctATTUtyB7g6JKKXKBvFqPeErVZnauHaYzU3Hf4hBI27
jVqs0lT5ezYgL1V03hVjO5vVv54vbUOMMj979zEDkJsi8BEF2D96s765kOcK9V/c0xcK6IfobIwx
mxl0zMc2PgpYf2R1701UEAV6d/8HNbuCdtpsrd/3Shwxnj7+MvfY/5oI1WY61Fjsk0VD9ozvPP8M
vq+PdK7Daa4yervfSEXAb7VJWYJxa9KeAubAVgZno8+X+tW4P2PTZ8X0StTxFUTnd3c/W712J4xx
OewDjHlsA3gvzWTPKvUdK3MZmRQwiTOkCxozN/xBHWbxS1iwS/KoXPX2HzTqUGVwIJJmePqqg+zM
+rAUeKI4tQO9rPjpK0FYTdjhHOo0isGyqpY2Dto5p8dqYRE0vJh19GvB4vFLlkMY8OLF+LNtr1y9
Ckg0C8QhzjSlBGRIZVedXWmbGKywmh2GlUJPWgtRY64+QL8EbA1mKMfCM2DrZJIaIypX8pTmyz3T
/GV2TbhLmfrZd9gIZd2Wn7UVrk+rBzZANIe1AK6SVP2phvfHJ8zHTB/B7e4wzonBRPTzVmMnBpvP
U0BxZxS6N2nFp8IwNemwLskpRr9fLd3sflaQ7xCgzv5bXRci2bd7vU5rImsdSsWHqMwOQe+Kh4Wj
TtWhm6kD+zGtevgR1Mc+OKqfZIi2MHb1TNlA0aWNh3uWZFYs+/4/BNDTQ78t1vU2nnv1JhjIOUyQ
ZNRbO1BhStSuBLawOSr3Jc+mqGYdf7SlZHwMukC6mzmJUAuX1kIaqMEug2hMbS6rMbWW0oa6npTv
Y3pHvoKToJtJ7kV6XUdWCVTkzqwV4lnpyZ23fAY6X15afiM0xU3HU45QUCi9pd7T8wKsPi22Vnil
jvzOSGwRK7orJRNVO2KgsXbU+KdrveJFg1XTZ8RVCpnpIIPkN0Ar8e7spWo2cAWkJkw5P9JNJzgp
FAq/Ft2/1KWqdbU08p4LCRmn6f2ms7WPmQ3pXy4mgi30AEijdmkp0mt+NLNPm3jUoe7ZNvGMGSVG
d9Q46nlXnVuQlk2KKmboAHVUStnkUFXJQ4ZNRXMotlKal35k3WUCfMocyBW3lbJsUz/YKIetIQyQ
PkVn8eA62ijTOv74xQV7vKMxjnWkJQzHJJfBYjKKzet2dziJrAV8FuYQRjhiFIhUu1yxapx/PhGI
B736kXe5GQ7OXg2IYkFZUPnuwJBCBfrts+vXcGr5T6xfkHuhKeam8honWClPTzOhDPj2sMRmK8Z/
NUAnDh14OaA3QwTuLcxf/c65HX6QjAQllGcqEuQIGZRx9iw+Kzmagw5KqX7Fc05ir2caSBU5hf7x
PNgeCP+EP0eNqarZvI3j3di1ZhI2jCkDa+ZLy/WgDaACYIXjEn3VFpWi790FjixJ+kLSEMSoSDWz
q8cnP2aqSxJYKjs4KZveS9HhV0fo6HttZTLFxKcXaYhSsRPUZ8xcLfsjy0oO/c8V4Gudzil2YQ18
a1WqL7InkMPhRAeeXkLyqccF1XbR06jgiSg+OXG4xyCFwz8vlyBTtt8ZQ1DD6xzEvk3v3ihqUY6K
O9UC6zgzOAXZwXgPvJwvsGb1RssyTT9xl+qAp5DgxSBsjr4uDvNAiJ9QIGktuR7+EsJFVp/SgOdL
8ymdADQRiEPa+olUQICmsVGyobZA7oM0pbgvygi7VdyPdRV7BfXXohOVsvQ3v82MMsFNNgWZQOuT
t2DX+bBO6HIGg+Xjw4H3yhjTnRinO4hQgGUtoNdJWyVfGhIGcsAk2Rkj/nJITFaqlxTYdh/8bg2f
qmOW9Ui35/EFK37Z+BbjS1grWSc2olHNVYmGP924aORPom2C64hPiuIXltSTMCMyC3eUXQAjYBRX
3SHmYmVvuBFsZnRAr54T/fgr0frjRYsYV9SstfIX18litoSorUUqpaboDRcAx3XxhB0s3e6At7qY
scFelYZwDXIJVLx9PKYVH1ICRorpo2o4QvY3mlrSeVaC+H6vD6saYrIlCcaqc9T4oQO9cKomT+VP
5ialZQcUaN3GHfMZZE5fkkgjXLt70twvzvt199s/nMsB6DUmWQm5A5Gth48QkqDBv83N2ViFcBgE
RVsDIlbgcjF1c4krXbq75xJrTJVbsT+BfBp+8ItzO/HMpCR6R1ddGLD/3kio9eszlRng7118Iv2F
uNv4GzFDqG4Eb3fAI9lWEYfFarwp7eLnXkRSr+TA+u+4zRA2ouIlEjz7oMNs/32prvmWvs8ydNIZ
5oZST0MkXp5WVK0W3qFb/cHXVVLnKApmCYtObOc3b4Ew2U3KfFc5qgYVauPC/cGCZvj+tdIHWItr
Sd+ArmNkSudh0sp4nGBYmnDCk0YTP8npkHl+tVvZBo9BiCbmXxi4bRUm+CbPQ01VdwM/g42bb0iY
77FZiO1UIi9K+lQ9HDwBLef1Bmh5gxrizbsCSL3O/nX0xm6Prl6+CbBdbGPC7k95iQn0UI3R9cY9
zs+GWXHHCD0CQ2EluFJCv0u6Tw820Q7j+mZOeGGVG77mk4YwFpj4ta+XLd77EOLrgw5s/NFA6L+c
PN7mDkYpxSPLbLdD+BZIJmNk9a6lUebmd5hfeYd3XldI/1eCXDVs6zfNcbpoWfI0KKDO7EK26VHO
R6NrCg3fqZQaA6k57Qn3GDTyLQW+QKuLOBo3dwOnnf6yY7kyhPD7YoYsn6sUcmV/M3Xj8+B6akKr
RabvpZ34jIEt2A0/PHRqolECI9JNkNL6p0Fjow3MmbGpd1+vUbToSGukSDH3JHxyDWa/skfFGhMr
6zyRD9U5TTbwwZVqkFBccEj0pVHNNoJU4q3BVNUKy/DoyLHi7PqL8kMFCnGwKgKH245HHm4Culzp
qCTaLUuOg6k8FrdiHVUmqA+4d9SEMKVgfcnNWWNqY4YFC77mhrXmABj7OsjSaMVgcNxWeONq+GiY
Lm1ei4xmLk4vOrv6py1PNgjGH3CAuzAWUg9l7MkUKXmEGx5FfXbWQcuC/gmQDSObUTcU26ZnrgHE
n1aXeL07geKwthTODXvV7455vTwd4AuUSabviP3Et+IOOtUwL8BBRbiVPCTBcuOilb7qAKvOt6h6
7bX1SMipWllfbnUXmp0Ja30sAn0YfwUdbcWn3J7T/PHqw3OvJ/QXqwWhNjBsaVDEetz0Mv00n9ly
YQ8G3NweXAGLvawkNZMN9K0ZwNLTtXwQIJpkNn6PFUjKhuLxDq4uV4UJ5/pUcBy5gBkVi9FOD4Qh
LpFAMg4QciC8f3Tv2qTP+k9WArTvGG3ngqTzfRLGZomol27SdVhBbBXCVURde2FQ7JYv9/5cmoi8
/em48NHa5i1oH7dkbU4YFnWwYYQsoVnxLtkuygd9OuzAUGBiTrKFBIm33xjxOy6qKuLGFCQYeyoZ
ncALuHFJN7hxuZLI/TOEplk3gAFUQ543DLdIjg/rSzsp9WW7Qz6v77QNXykzmCnjZU6gSayWmpRB
v1oQVrwiN85iP61ekdBs4Ji2bvhJRCPr7KDnJBbv1s440eKha38RxQxt2qggqoDqbLVhBJybxAow
/qmKOiH65UDKLhjyKsGAEIsOfsZgQJC7n6uFUb7YtoU0wePxoKMIv+zBmcT4vpOJIV39V7DGQTfy
W0DHka4Qw1F3SpR74dezoojQSZIQ1svO32w1welEuBm3RTMDOz+ldqOQZ+kFLz0Wm6JQx+hFbPvA
/lO0Pd5fLbOkwpYlkV8XPJ5Eq2PPf+gMxEz5MbMkVQn0XPiqfirXrKXkYHr1GNikNFecUBktnjMz
pCo499QHhqRqQdisB/N5In7vIhr6sTNe9r8H9Ys5bddnTk5jS+X3VVogyuOwkeZ96A7eGbHuphms
hQ31SJlAxWPVWb3XrGf+li340UCMIxot/pgpfQRZ2693UHLLtPbEnhnuDNXCjzfw2JPm85gyvvA0
878ufCbRYup1bcmMmGNx/bBxEIDnbxLEYNgqQrb9FeWZsmYK/BjAb64dbjrPidJks9NnQbPmXQo8
a2GrjS/tdjEry+/5Yg96Z/FPAa/PikIuWhVmmneMPhVfbwVS70ogFVdPjqTqznqebtstwKF2aiXp
x+ogFAaqT+lgYo5pB21oIRpAn/ADoRobfyygCvseGr1tgou/ahBzt682sFASQs3nC01Eq9oda47Z
bScAjemWoBiIXF0+TVyCfQDd7hz4Uo3kKQYtgIoUhb2jkylVf/d8HzHGkpP8RpkpEM6vV3Ku/eJE
ssgtW+Fw0O50KOpfvSglkNWtUC5YR60SJ4kRrduEqKtyihIy48EcDS4RJbgwoEoUT1/+2vEHTgwH
HxeS58Oy4X84H8s0BV/P6sAwO8en/3CFb6Ijq/o9IEYO5ncbT1D7DRXECzhEGpbWZg/EGvxyxDP5
nMr5U1SbqCa1Rl35dcZyKEVXzuryyBQwEq1X91Tzalh2dWczkAaxvqg5eP5mnR39GgoxxYgDhMk9
TAfowfnFCvwdy+h8uf5mCnOZFzsuPVxpIPNY3+MYxxcDWi3++q8xjRn4YRtFL2c1ftO90dzL8bAd
i1yvwdHTjY8oau7cF0x4IxinPJZgwyqwjAglNWWpdRFxUeewfgwY3THgsyy2p2iH+XZCC4aU2v1N
3yWYbeEqJ6prZyDIflq1nEUd8kuWTV5FVpyGBHKVVNXIPVtCSeI0dwW8slHOekYdVFG3xaNJHaVJ
RafDgpH/n1/eVoAHnLgfDErNBnaYN2kIDHrgGexOkygOueTOr2F/baD/2VIR3Z7iQcYDWQahBP4J
+v3aGsFxG0VTbBBokuWjgWpxDZ+fMOiIZSkyAXFMzF0ov+6aCnN9vo1AjuNi2udXgrhJLsQVTulS
dINJ706+yNJfHSaSWB3KnUsMXIkRCIGSk3NxMK00YMJ3XHEle35YjGTilt+GOdZHwntnLKFqdIMN
D+06bueaGJEgzvlbB0E/SrYHIvt1UTdWV79DMd41z2XwkuHxTRtq4n1Ks/x9QpN9xztKNzKiaFsH
/qGm2Np9a/u0pnXm3sgCN7Wy4qvmXsoOdOFee3kFX6RwL+/3zaNhdg70dOUcY4nWzYyFEj+H00yg
iAQMnE5MUBUKvoeGsk0PzGxAc59Rc3XcTTgcsk6qoo6kYa8pL8gF4Prt3DwDzu/O/HWqzYU/G42x
cyeVsnxM/JxqdoagANWSCzYmKfJFO7X6dzzoPFhu2RGQOZpcb8MGEMbLBachNsJKoeliztDUEu/A
dmb2ri5ms9HhLlSfcBherox2EUMS6s1eNAEDbwyFQieIo+si2aXzTqDxTtmf+qeOYD3xpu5F6Q+M
6fUdUm45J/AhwIWRoitvgHf1pVepSuIGawZj0m9pdXGW9j6bz0XcnPp1ElnsnmU14JktD4vmurQv
YthGqBB9PK53l+wwgw2BjTBxM7Tai/x6d7L8VrMlH7V3AUYvtfCNEgbn1+XKcsYEZF+83/vPrrOx
g0qfSujEDLWn0PC9D6w+F2psB4Nw0k/ldPncrrlP2zu/5kQlzECNYVjVh2No1Oec7CQWiCPGp70v
imtoaXymJOF4XXpjtFQt0ppc1121ghQvWkGczJjZ62Bc27oklIaN2HWMk96H8f2F2nxNjXpEZ6qn
fj8ENo6hFZG4C+uCdEYlfDsToRiyn6ObdiorHJdmJl80LPARchrijKrU93jDv4fcaReQWS9KEv9D
ZnHuPAftQiMFX1MviRNLwMw8pd3QlZFfTf8VPLvirYijByyLlqBKk278XCXZArCDVQAS48mmIwlt
VXokJAjHDqJw4iGx37F3Dozp+D0mAzB53F6JAdFD4l39C0YKtJ5KGCBd+4kt3XytzDakTOS0ipxF
K41SVESy4kQGkUK7zBPSDoB9x+DhLdf8jpZcYnzdrrotwcUgzWFueBZDXA3B0gCd1cXB+WYmkVBB
dLtoepO6ErqijeEDmsy3dPT86FAV2kX3mlGP1VycBLIgTKkwwRLJbyPxsPtCsdXCX6eeTB4nCULW
tLB3FeF/bp7AIRty4iq4hPzQk3lsW4U8PCVfgNhfSvs5PpmWZPvg+8ki2rxxJGAGEgQNGlIknKGv
WyujfUA2r2eCi3fSXuWO5aDxpvbwXB2bNkPS09bwToIOqOgtV89rP0dUhSOVMGfuozr3hY6rNKiE
onyYFMYk7EEJ6eR+KSMbYn61acH61TpR1WcOZ9wXOAMj+530MzCuFjgwSBlHXR6T6V1XsEmIQLhJ
BwJMxVVc3AjEX0P9Oe6HS2gSJfqVmlrUJX3ZB/FV1gX4RzkUw7RgpB62S9kOhYgUvDQ1F5520H5F
9PzgRAdcincQi0H6r8IHNS87K+MXvcGDhvQMUp/65lJ0XT/uY23H1rY/PSOXOXyL0qil0LDU5znE
UBNVri+W/vAysDnttGW2oza00EkvifSZkSWv/otClE7RORKSAT5bu9vgeuLmpuW+smdILaIHl7wc
kgE/lCACQpY3ioVxs6H5uS2G5VFs1+WmiirO3k/VpPcXMUP2l/IWv893bFOf2mt8Lb8CKYfdTK8D
KdZJvXk9vpfaot+dUVoqxUtD+j3GRKGyf4OIdtF1iNcZoQpIjKKFtH7FWxoJmK08A33P2QAJQWzc
desLB+9D0C/Un4lFjV1kcg/TxaR9IwNlw5JndKQ7CzHTl/qEHER0DT75bpD13RBFsAgCBg5o/P/s
EBZv7qGsq1G6WQHqgxfuY1s0JcvTdwom5dQ8GWUEjepyTjvVb3Gowv/MiqxT8Wc2RYOX49vo7VZk
ooTXzkBNk2EzdA8T+qyl5ybbhigSPFl6EK4PZvSsoVH1Zixn9fxvZh7hzK6UiNOety3Dmdyn9m0E
Lc8p3Npa2z554Z9/nzCIbklIweIeHRgrTdmpijy78IV5RnECxcJvXugzNGC0KrN27x2TR4p2qT8u
Pz19F7jbN8JqsZ1RHrghxvFAT1MvqjN88O0k37rSD65GYES+P73H5XHsu7Nyv4pBtA2Y4l++TzsB
MsgnM4N0ZRAbdltMrRzGV8/UZktvUoKTjx0CzGoYBQTUG7IeaAmMwEmkkwTGHgS2Je1AJXpsKGX8
C3T3CslEW1Wp+Zh9jkmUko+lOmfuWL19zXcSU1Nr7OyvbswSRkk0GDpHrCd7meGV4pSnG5b3v/cP
rMQWRTus2P/jqitenlbKhCzGBoEKjmBtY0j1VIFz3EewLAt+NtPwXPA/ykc82GR7uEoGPnQz+Np9
sKuLpJ3CVsL0fWLjUEFOAtA3UdJximToc9Fhs8mstFocYN99ZTMjKxH9Mjp2716bNQPxa5tzuzNF
ryum2pQWV0RbSJk4yqJ5Ve6ZmkIs6EQQ3IGvD1bHb6JbAkN1M61l+EWikYPy+ogLpVXwKEKH8Psi
XLJ6ohcJwifi9q4dMOWzmaHo9iGhkK4x7f5lVGuzSltxnSrtvAi7I+h41Ek4AUCUzfV7ymnEZ60H
pQ7iqiP1jk75KKB9MvQ622g+vqHwH1uh+yDiXGdnYKob87CyzQoB6cMgf7bug8BLKhDCOLqHWa1I
ZEEO0xuU48BbzboPaUlf1g9ig7m3k8up2a/G4WG5fR7y1OUl4qIbU69gzTEBc+U+zThhtghL9iu6
dSAc8N6a1XBWOLlJnBW8agrU25UJQlCOYsyPI07bi9RGpzYa/YLc3NURIZ+iIGNc3HVEZLwW85S4
yiu8ugoxLldQ8Xeat2MlziLa0fEUI4LC24XyJ/CAWatLlcmytBjNbTqu+A2TARjsbKsqtknxdPYt
EdEJXYI13kwn2DY17/9xt67AzzfMeGikmkumMjD4/jB3EMSfLm65P3UfrgDihpJi53VHVWq212KR
ma2/37rqjBAFIlBmKYwLPv+hRIsWFlsfvCaOsJe5ciIG+9J5kAEoYM88pSKhfDgLIk6mbWD2CFz6
deWBhAJxkr4FdSQm551o5uC2jyfWd7aTuAZpSLADm+thAML85CGDgU94ZZe30NGAThJVi8DGHNVa
OS5F1iCJY4ExLPLutxSN3UzK3lKJFvAlAHca09WSnGRe4XP7xmaXdNxMtpw+NyQVvon/cFnyOsjr
5KufMg1mE3JCbcaxRSuR7HlHcs/pTKuTuP+xBEosY8XNlvbtIBrH3Y7bn0WzdLbAoF+y11IYTX6j
0czWI7gESzB7qLjLg5DpCTBQbSozytXoBR9P072iL+tS+o6lTtLzDb5zS4dNxfmsNixMDFrbaneB
+w2aPt/zKdkBDadj5R8E6W8tg5bsoZxLNZ428spNIZJTJXnCepXVAj2KJETvA1q/8KljfsIxPTwW
soPkMjJd/Ltjh8wuUH8/+WPHDofxEK3j+4m9owqhxDEEnD60RqSmbBJ/+3OS5DsrYOhWlRZkFjxg
VFnrQYaXE/W7MrB1kVJacGQNg+CJpJT+s/Qwg+/I3a1NQTqm+fo+q9erNnf8MUZjgOWplAm0G1T/
nD23STSdN30ZqFKWOT6ZiHurXCFf7KNlCQ4t7uHKC94yGWzXc2P6BwgsMYi6RLdRM4sBLeRO7egA
xP99lIgZhOg+5FeO4qH1y2VmgKbJwgkq1Uc9isDsxOrR/5j02E1s8cgEAIBqlVyAJKfef1wLvOt6
aTrB/Gn3DpOWhQxcy83ZqaNATRLsG2YGyZyxrB5syB8OnxTzWPC38k7I1JR7LFGfSzNPnDXxc2/+
MFEHucCq29bpJuYKCUYCYB+UKCqH4aRipHXnXl637szVvKCf1dTVem7taYyNP/vi7d9DKmeQfASR
dGL78ZoukRGVIbLW6OjNQTWUsfMaqni5UZbp44CCmUON5MEs8o+AfVyoubVQIIY1eXjT6XkZFZ5K
NSsb3O78PSz6i6cKyjfUfjDbf6zosMdYRcBuXHohf3c06SfofAeDdcvcgnHnc0/d8yniUemJuWxT
c/LY03W9ShCvVD9RCKspaLkDejN0tW0sxBVSNE+5E9UStmXogejpnq8wbLgDH2kM8t4WfBlSbflk
r/TgIoqUHiZHcvBgNpAPBbgVnWuNs9V/AR7OXdWphOIJ9AzhOx2wxW7dCLd4Hp01KbyCfB3zX39t
vTirVnSPYXcyMChrrpxkNenjhnvGDwtOW2paSPne/NGW/ieYdR0CI0jdpie2MGk69P0ChgOiZjiG
fWpqnFd3WQ0T8opeD/Ko13nyO9/fDp0RrtKldseFgQQmsFYLJ+z6tesuZLRrsQp7SVudPsKVlKo2
d1Xk97l9pkTZB3+OMAZ/qlxC8TFYsAT0dllGOgQL6sTK9ZG+kqGDL6WtBKD/EJpHqNsI1yeOaOY9
IY7dEbiAB2LIbxEkRGvv6+BcNWFszAC9/m0/D4n8hZ2/E1grwivV5Hw5izLQClDL9GEuKo9fQYBy
vCf/btyENHavd/7/FCAdH3C18wdJ1azWN0M3eWPdksJxb7ZkDkxSmvHhhlJvdXrOlwEmTIdmN0sW
nIzdvmYPkP8mzzNUoZ0e+gQHgRs/8OYWxwyf3dGpxQ5WFqY/N8Ns/If7eIgziW9b3RC2r6uBfa6P
lzq+zs46+M/km7NsIEc4t/tAqlngFnYr4z05lJv4W+95l7IrogY7tFqJBc2CeIY8fBD1BFrTnJCE
ZF/UW/7D6L3QOhgQlSeAf67Foa1ATBdVkRApAiNbeT74wmOnxGBQx5PKdKlgQgdjUhcl/7uo/JGh
chNlI1AZUnU3OmsNMofAswgv1C+c1YZcv3VU2zWzcW1Hjsjskj/XT/dsfhRBo7OQIRtcElLanjv7
3KnQOR0AhhBY2c6TuoGi3XbAe3SrUgIih8OYyzkYqJm9dJtgVEegWjqKCAFZa3Lbd187QlenHbHJ
17OVcf/ttb281H/rDJzejfFYl5/ckex0HRTRq1Ish0IoAy2w7/ZicevovydNbXC4Tnw0ANtb+x9u
+EmHjgiJPULqODEXtoqAnAWF6d+S5+109hvPp+QrNzwM/jApBc8LF0wGOanED/qy+hXZAbZ57DUL
YXHnkyF61A3UiJwJhhmOeTQagfu4oHJBSBPegvcvbnzIO5Gf9UKszQugk/2vdVcxJqIO5TXlZmqr
wqdAX7f5yipXCbn6K6Iw+VMp6s6WIsq5qDamO+MG+1SJXv9tdJXMddusWmoeNk7CTbVG1fZoia9z
M02rLHnxXa4z4HB5cpbycmRjIPHCfBS6LCs7YDlAHHb7VoRvgnKQr1Fn++l7k6vpvef87J0W13Wg
ePoKaDU06QBLt8x0EGFFZnVfvmZwoOIa5K7JmLbON4J57eHBlLuGs7aAn5huu5ydDOVqCcVBYvIM
Jmw8FiO8+mh3i8Dg7lOqKE0XBslNC9JGxLPRuUNAjP22rp4sQMd2jmmmOHFdlitPJSGIs79XqjHo
Tc1ETpZ/t6zPJ7wFWxLUM3KhsHlHtZ5lYx8yl97NLnCQG++YkEhtAe/KPkIOtCIbPSrtwni1CapO
GJBqjCUhTelw4xfGpgefeuot0kXOc6d5sf65fn8ZWTaXnhAG7N629w2doWU9ykXNO6Ft6r6HxeFd
99D7KgfLrB3tRb3InX5/kGCNUn5/RR3ewJNJ+oyLKiFHPdnjC9VXi4ylIFB8GKO7iteD/z8stjjQ
yJHuXBj+SN5zQ1x8k6fE7wAU3lTMep75wrlHy+7ttjxDcbhbFsgz/SzlURtfFbC9+s36YHSL5MA6
OKzzY3D7gKavGwrSxpDx8fu0nBUr1as90hT4iiSeP04aKysqorUBZP40WBy9yTXhR0f1EPpPYJD6
KsmsgepJDuX6/ujz+EV/dr49oWLS/wG663JJPvfq/6NYgFH48ByYyE6OBDASYGndb8m85OgIrA2U
Mb4bokXsvTkYs/avwiX3euDCJJyajpele9xqi43K+jfAjzPNrlp8Mww6RfYQLf9Yiz452zRrVMbP
X6/YboE84hND++TzXhiy50WMOBoKmPsuHfjDVtJSwwlpeyzlr3rzaWIwnc18Y6bHEK+2ExjA3GqA
ZGd7eKF/MasqPoSlCNVD3fenHDff0g8KcQ0k7CAmQhqbvAg2fJMDsT6sqrn0w+/VEiu6VufsfkoE
TgDnNTKArRATJlO0H+pMAuPlCyghSTYPFH7C1f4o3gQMB+FRkb9uLLOXVtBtKRR+IPXwqDreKdmJ
PymWdNKmBczU837bJdGAT8LEiKx7Qd+GH3QKJTQH+GXf6VyTqYBHHGs4lnTOJhKimwpTF4YebQwg
PymhARxi7NzGhLnUdrO8zfPaTIR29YfQktmNGV3NyhVsA2YzTppPYBYXfkZjl4E+N26kKVFqrEkK
ho+F9/KBb0SxETzAdRe3SY1ouMV8VyLh5gYyh6LCSvvlGImaD9kbQ6zgm6tK4h2kc+oFv1EjFG63
LrbPbhjjoRxxwgbUP5cR0ZzCuvivtIPH3ddhCD8AW4VZ6FsJkTjJvV0ZP5mVYbAa3XXhwqy2QmtD
OL0kVGZYldII66gYU5z0W/bOmyd3zx+AeQnAnsYk7ledrxyBBqvCCz+Nno7m8qhW+95JqCTS+ga1
dZUQuWr0EjgHHnl1LPajn/QMday1y+9+1esg/jSCvuxqpOeXRegSVqxE2TxpvRN40Sl3PfyPyI0y
/CNsZZ3U5mZ0UoJzXHypsDHTmR8TNU4dZmx/cszdhwPzdNfEstGH4VDOCC1WfEVTcUCFvgu3IopY
8qG3/7QpCOxMWNxGtaXMLvxZOERBrkDhy4wEQohidc9TR51IMjWlQbgD5HuJXFL47MxyZ3dbugj4
MdBJT6moGDCD32lCUv3yzvFeaNnvDknJU2ljouwiMh+7sDUNZv/6bagj1igkHkSLeIX+/QoZQb2c
RIMLY2jWYeoKIzxsjgoNgIJfc/Lw2duG4BUZQKFZToeOfpCxXTOqbV4xXbha1spB9AE+wltPJrmn
kKMGB64ueeLix/vrCI4xwgio9+/JXVuTjJUMpwcch9l5yCNPRBgAUBXb9CzC6SLVukalbvVy49xB
gIg4/qZPJcjR+lzCi+2hDDtomDRh4uIYfA5f4F9dIpiFUfT3Fp8r7wwZ45T6Hs4/Q3HGAJBfk+mN
Qcfp3dsvw7Y5ipdvr7c/nKT5QnRvqaSKEAbUNaNj1AS+bdu8U4Hi7CJmwdnUH38WRmjrJXaI0W8e
GwttIH2kkaA9KmtACfCg15zl1lt42oQ1ERZz56ZW/Apm6XPVw9tCS5nRyR/Lhh3QWE2zplbu1AgT
L7XrfdbmgcQJg7JpV+QGdr4OZg+agT1UoQWQNGpdD9jCTaMo3dC8lCcQ/xylahS5g8wyWA8TvOyi
rt8TRhwGCFY0QihNy/tRO3558Pd0z0TvVj6KSIPZrhUrQkIApRuW9o3B+w6TF0iSlw7g5ttk9jSa
IFo3tpjm6m5MOStxYnsto58zpgmkEpBgsoh33tLGs94inACmxEzfW3Ue6mM3kCcBunINi7aePxFW
G0Nn+Ou7tto7PfChgOc55prasPMJaqALmfuqOQDmtuvsO6BrIZRjZH1G6fK3bASY4RnHqmEhcm1a
sdMnPlx25wsHe/yitp3Xui1C0W11Wsb0ExMExxYH/nUqDX7DqlbObqe/zhHoo0tyDZniecG9VgDi
AiTNjfMZu/Rwwnuuboym5ByvtN8N4CMVIR4ke1iIAEAjCieYkpg2p5se6VzD4jltdCPS6zWkRPsY
eLf82J4VCCRKLd1o7f3NRQzLku09srF1IS5XGRji9vYuH68VUUuyp6ImjUolApoKO4Ns0c8Kb3sp
Sjryilfj42qmTBohlq1OLZFIFrRQO55Q/v5iaLZCBccIha2wDtEemj5tnjH8NFUoVkSKEBi8puQi
x+fE9eVzGQVgMEzXEgPDVNyeXYn/YnDj7wjqd2OTsHGubvUknQeeCiUONezGbVFBQHhNiwwmXpi/
I6jC1wMilLdq5mnPywnpkbTScsjCoYrbYRJSMi/woQrJyDN8P42VRF9jshwPjxV2+9Ous0UFoVed
08oLhzWzeYu9Ac8mtXboFdaE8FpA5tuaM7jTPvbTfA3KIal2+Hb02IJjwMiBmrFkxvj5I2VWbgp6
t4XNsfNWJHKjPNH1PooP4ANTwfAJ8sgdS5VHR+Qx0ewDLb3RF4FCrQVI+87G11yUpwKXcmxWnkbc
i+/ss3OV1FdBbhHvUKnlwmK0hvBfXjsHaqRf8rpRwsEqGoQZQTNL0xEz6NsDhJYviN2OLyWeuDil
pvI4nTi6esX90UTYphLIxlkb6Az55bj4DUxtilMa9cF5BKnqO83mC4dm6EsjORhMG+dE9hViE8HL
Y3vfj41Ox0M1oT60rTVlYa5aZCublQgkUstC0BN1R5x9WcwDfKqGCJo1dFi9vxaFHMOUY2Kd7rPv
a/gjAXAg04cxV8PI7Y8rtGo3I4lGWOa8FGq4RtFiyDFXWWWXeFnO1gcJp6mdHDnEtZ9vpuad3Fad
4s5YTLBggbaH+xQuv+8d2mNDWs0+w0DLBon/qhIA6F+2D7IT4Ed9tJCaXVOVFUKu/qTSrc+atv/T
aCI2x75/E3PzXgIYDlpOTEZtofqAP+rgDi4yLVgIxUY0/9RtCrlFSebx7OFVy7w1w1cm2JtEvtmM
Fq01K2rZPhYlpS+uBk0uC/K0JRH+IFvm/EOH0c0F0BULYj01NKCH3aXkAMFwgNLg7193YaP9gosD
aIazHOjCuZj8PeEXhF/75G/yu7brrq1g/2PQ7/CRNJH75VO5hvMKT9xCiMOnAwhzLzql2LkCLZmP
p9kkl/yYD8u2lGA2+nbJjHE2wf2BL8rTQM0RnZ0KW/SFkz+gGqgG1cK292/FxcyYFNigZKDh2dxW
8tHCRIUfpk6+cs0+Ed0foWah3LT3oTucHKnzuboJ9GOBVFv2vJhZkgSDTNlDulLKjmWRhlv0jnPr
JJIxE+0BTHlK8uAfUneDe+cH9oZdD4bsDogJTjfuG/2yjhb/H4dvN536f+lgK5UWg9Dc7JjjUTkT
quDbmD0jLMst23OpDg2lBrhaBJCJ0AeT9xBFYgfuWD34ZuJxtLkhy+ZuTis1ltq/KOc7WXZ7xKzt
Ba8ThiUubeIIw7QB40NpWSR1N6II8nTCBCTDsSlis6Q+rfcg/kUREuw2hzJ/q9tDhnKKacvWL/wb
CARGV6sJ27w7unaL4Ugs+BESLdW/D6Mr53Y1+lu5nXkY5zHEBe9AE1IKKlIHvl4RvqIud450GNzI
xTJiEA35prD5WsuA9ImZ/TYroiuSSfLXRwv4a4TxPMIkWI7IX3xc0cE2u6F3uJnuS1TWRY5jVL5S
OUSdG0DuttxKpbD9akO48i1VEy+aaqxoGl54RGt/Ox7UWmYgJ4r/qvIS7khPBPVGjp+9thOUKfuP
WzTFmwvVqtjPqoyRkbojp4HEO55Bla6eW9a4/fwWbDzfw+eqfgW7xuSd9KSyq9VqZy0Vo1V+/yof
s0tazL2pwWyeb81tHtrKTpUnNJYZvAYgAfESewk/zZphvHz6gM732t6skM3rvxZG79xM8MtWi5XH
3MT1dDhwYlnc62/UpQiI6NVL9TEXFOb96dGhNZW+Fxpdh6MVTUFWbdJwfiukq3nJfdJgebybfTOC
zLkS99lSfmQEl4IiX5FmQo462Bb9puCqrbP+3zG0rKCEEj150GXicROgNHvLVxFbRUBN5rv2YpyE
rZ8YXhZeYIXesRLNcik/BRWzfR2w8YMldd70IC4cCC3CWGJCDs0L9LwBvkZ6g4mx/3x2CuB396l+
dk6tNp+KKRTtIluJGvlkqPo0vZVIbmk2t2TcSoAHo/QnlIgS2GeUwiA9PWAuK4P+ujVqlZ72+sdD
FQn1rnpXSMcnApxH+cQJX/VgZORvM3w9lW+8J4lRzP7FtgopnXE4lNZcXrMVTY1NVQU4nlyWtbgm
gzJfYJSPNSbwU1eRnDCBHDjb22+UiwQgSNV1W+1sLPAiaDbgu+tesNWH8DNmSorMmm1H8nG5aCax
vUOzjugTChVuH3RPMG0VmLe/ZvAn6NZxp97Q03PGnkERhqw5U8b29U5yFsazQv9CRw/UrhDh2xnR
wlq7utZBbYt28NwBmpVrrKn+E0HNAIPL6YCCEK1QJvcLjXGB/S65wSnuTe0+e4zFIbZWerOnOpMV
hbZNfDpqkT0/TIBzGk7I3G892TL3bCIWipRrq84EVAr1qannKlTd8tePz0g4HSo0ui/Vye97TQvH
JkxUXE0HpbDGhS7AJWZGXxR56VmYI4BVprBKdrXwkVTKExK2fVKWMKnnTb3PaclxSd58P0fvHyHC
NQ7+MgZtZ8PZhhXZLAxcaY4LWW21qq6gTB2AXnqnhG31eGq9XZV5QmHZ3jDrYKzEzwZzXCLSREIc
kbCaGBDRuRr9FRHMehfQYmVUKApx7p3RB8WgSlUVFzpH5B/1XdBzSQAg4oCVbeZ2brVIKoDJWprt
4GAnP1JrtHGmdKKK92BPQ4qz7kLzSBnnRWJhYSCcq3+bVhMHRElkyp338LXUmHAHdhhm5x4XSBGR
ZJSL0KGDb06PxgDeMQq9oF/kDLVsNEKIbyRTH16DA2PYcqp/ngTESA+OQjQeErjRYad+ZOfTBi1H
q12Lvv8cMteOISzDnTw4RVPexxNRZTM0seOHu9A7yVPi1tDSlMpEzi/jwCJKunS9nIOmncEBv7O2
Y4kHsRh4nSDt5ja8VeYlyKeiLPkdcFu58uvh2j8MGCMwm/vNJZfu4tH+ncmEMZg8CDBIBqpcn6sT
Kw7Sww9Y4Ts2msAFF+pitHjhz4j/gOdO4o6i6NkgB0EX496l4uJ2CAkoHXYqzyRhigCjHypW42z1
A1I6JS1J4cBGpsZzNBib7Cke5Min51ia+SNYQa2rOHBwSHm1NwH3etDUdOsXN2i4koFsvNCLD/t1
o8loto7+nbsiz/hc6zi18tqeQSb9qR3kPYwL8tFH48OsQdzXhK3YwLt1nLUFAsdPF0F2tpZaXfA0
l0tTqY+L40oEOt4rO1kANhjGllf1VCnrWUc5cg/DNJOznHSnqr0rcSHJ7I4KlbYe8KLdvZa/OmGW
GfNuZMmep1oW9VGusIG07+gHqCd8y4MFZW0PtBSViABaH2OyS1KeXg2J435x5tfixAKaA8hWg8/1
URxDonGLmRS0fnVzE937IvXvBHWjc9ZPb5IKPVds9dhaYTj4nW+zMpRCwFp7iR1YZDcDL34dfMEQ
VGMTG5y2puGCGBDpHX13jrOUabK/VMo0X14Abl9cWnqwD9JnDlzHZR4fsuEh9ZVGkwe85uJ5DFQi
dbVY0YlsPTke3gaedJYviiZrFZRQFaJ4b+MRpENR3p9JXdIm7+qrIkibz4in+jurd5ingJOgWSdJ
93ib9faiaWyRry65xH3lUjVJYDS0Q9rzFPLgvsHRCiBZiV4hsWAiMynuCnOjJTry3RE769ixc2ho
QzMRg798feJiSjSwS5+Mad+WyRFxS5DTX1VdVWwhNNHF7X2GRjDfoumQiwfz0SxmL3BIuIzTZ4G3
HZjQooJWvpPzjSur1fwlsTMhT4rsv8LUZE178+umyiI1ULbJOn9NO9YqKaPrDZXX4fint0U+Dke/
LJvXtdrVSDOXkS4PYICu1dZj61Rt8gneEX4dZD+aj4q8BD4u3bZtZtSY9aKWbere1C000v7qasVk
8r2VDPhOmRRffUyB0nf+3ecN47sSu/ItLYbRp40S+WEkUOh12r7mWhjs8dlX91VOOPBQjTtBuMlo
L/fP9qB96tPW2nnbOw0bUCej5sV5INVNSIS+12Ax6N6BsYleySj2tT3CnupANxgZ97Bp8WekC/X4
yrJKIX+9C7S7/9Q6cD5WPspkpn9bnO2EqjyctYwe9xWnESIX87k9wWT6FJIqLfuWaj1itcaJLRFl
d2P8S6Nfri7Y1YLQkQ/TUTc8yFxHIJE8KrY4fAcSvFibQyo55qAph68G5JFP/ratbJ0zdQC32u27
Bf4ErBLFUdR4AOv1r0JBuh52vWb7MLj55orD34KbXDqAOr3QXn06UQLOVQgl9Yo/GIcW/ROkesLx
F8gnT5WhDdEZ2CZJIbUxlNwYIvmdS3n55shk5copwnA+FjhFBHvb5BR7CwgZtfvOoV6bA472S8gk
CC6iRYq/Y20hwwLHHSI8lIUVtWnen+1rPeS0rkj8jrkAwE1HLgfqMohxViYEYqZWmKQpOccKXX8f
zcEDNtA0YqwONUr+a8/XyNR4bwgfow8OirCgvmk7KX34qmdsA9bYqkkUV5vaLQhNBzNw6qxzQKuF
ydr84rvlMChU/PHL/X6RzXq0UtAqBkkalSSO7aJms+iPuy3lIqlKTlSnx5hKxRbPEZp2IhghvY+a
Hpf3P04o7u3fMMwozUoAdOxIZttd6wuIcgogaiPDNQwePu7aDxKDdquKBvkeTi8JoTgNAHSqmyhL
II7FlzYfr1xzP2+JDFP7W6gDnu4ijzdjnQyK8eKZng8Q58atjpegH4/4dJrTJrs40JQFLL2/g0hb
yt+sCthTIZphPct4So8KBBW8rsexGKjgS/JWFcb2Ji/6fsoJIuxA2HmHhsGiCTqLMcoxHW8BPTh0
7skkzF1/GKFCUobsLwn2EZrKBvpIBB948mB4OkjBUZJeXFM5fXNx8tYWdKbZVQMJrEh4sDmYkD23
0b+a+uybJe1ok6CPOYZHQn3PMQgJV9OSl9qMfLkIwIQBmBdjDFdA3m0HProIWeWYOPv98Z2SvR/P
G+ltkIalhE2cDNfYjXZqSMBh+7qsCkx5JRVmUpKnnSNgVPI56YCuxK7WmMRB+WsnyP81r765Jac7
9P2CVq1AlbhrHp++2ObvrT4May4Q4ewT56nM8MaeJLiMtTcfKPYSavajwsnR5MU1+9HlFTI7rqsR
o0vhnW95qmfQDHWXNy7h1jjAhBBSS4YbxMDkSZgOJZ8swTVluZmagwRO9IYEO/9da1KxQEU1Bvdc
CrHng5KAkzomQfO9vjze+Y4plJK53O2QNAwBdbavg1Rkg1qUl3G7wm011jOihcLW0eu9U6EnYxcc
IHUt05jMcElzVIirS8cSG1148FUi9cq6MEcmDtQyzyLq/IV/0w2pF0q1LY2pSYsAqV6hlrcpGfXN
LGI2lvEAIf5YEY86VG4ZQ6bMe84R27YZNG3dT8mWID+sIaKszvzN5JJqQYdQTr7/1enmo8Z4qkP9
OB3dx5kxbv4Yue2oqIKz1fMTLdq34rO14Og46T8PLAqW/da3LeuZx2LvdKTsQlWnxile3uYMcYhF
NKj3p9V5cxzUlJsBbSU1KrAS7vLHA6dTyPNllS9yhVCyvuVVAXNlIsZN9vIbGEcomC/4rg0vXaQA
cND9hAIbl/Bp9LFxxDfZCxtoHQMnkoAEKvuDVN5GxXXVJP40m2ztFHBpXUZJL2gYxAEuVw1Vua3g
aiAhfnRDFbN554qcJPE1QWunlqzhSleYAo6mE91fMrQgfO022U0l0xsCc/CbEqUzdyGm7Zgqbuf1
kTOUYZMskCgRHA215sP2s2UyyUY2dYmpYLJ0MJbIjConhI+9QehET/701YWlpwomiTEE5k7e81eR
tnJTJ2WmymijH5t698kyjph/q4kYqyxJfv24CbrA3tkawbQVaH6EpAEG+DlnYN7IFwxFfbYNQsHR
12tIc6rLuE29be3G+NQhTE4PRDzl/uYK3wnBupHqIy98aFrUm825Qj06V6eopuA6gRzIjpocf9Zu
bz8yJeBcjZ6fU3Rs8Y6oqSkN7wihYUvh4mA00T5mut/4EePOM9WmIfj2fs5Cdwbqjm+iRMjAAYqK
T4U6abNSnIMSGV61gI8vdfDjUpYphlP8/MsfYtlgxHqm2d686Fmbv4ggt+7rz1k3aODBthIvRojT
Eh4CyFDkrPHA++HHKpkHOICMXr3DqpDmMYFdTvDDeEG49opXVGRMYzGvo5DA0tVj68JGI/oh0QlY
EZkvLAq98AxZ0QMn5ObTABl+l4bJXx1us/y5RpjDKNBcU8cbApXL46RN451F1ORCezDAm+6HA/Sh
IsFMqgQo27Et6gEFi3ffEPuNMTx6CLsT+GH2HZGOUZaSmlP//efij0VwRGh0G3Z/unn3Z1VMfOJ3
vjrGOhz/PU/GFMpdvDrs5H7czWYBeJuUWwJyc92YIYWOJg3UBt83g7hvnRJ2YBc8Bb9Ncr8ID+OG
ueQy+DMj8ymLZdqCTTwJip6L3a1dGTXIdr/H9ZCf7uozUSmlCPH1/tYhMiVg1wO1QkGVeh62wXli
1CVQ6+oBvBDK5dVWFH9rnPW59VolbKr/f4UdJD1S4fq9rLMPfyD+EF6zGYCMzkB2wu8Fzzd1pvjS
xm/+8Qq2R220rbyDzSEN8QkBFdSslPK5YEY1K6q2+cfiksVfEsqy4rR9wz4R7B6ez2y8Lj+3B0pg
xozUOJ/EkzTFuc342qFFyJJ/IXwfXFT+DUAzKnuJVFNvUelLJ4T82NP1s1vxfl0g/ChmoFxve5D0
Cuw7Q65U+lESuhFrSDDkbMhbjCu0wnu2gj3/0pTotn2kZ3hQkMf2Ib+yNdjeDIncMGOC7CTax7Kk
aypnFP41T5iQHy9BcJi+hX+f5ZSFgGcvO1Y8Xhas/sZTcVUrL34fHzx1XMMobPyo4EQYWNpR6jub
VJqh9Fzkc4im42v4zB8JFLDCcC+tCHN3idzbDS7nLU5xBgLgyiOnifcQD4yZJt/RsRE71147TQGk
Jdl0q3rbhHPuu/ntwMekS2mSyg0v2it66WPaLGNVmyLeuIjhzgiT4co5e6Q0HsXQuTfX2XCiqNuR
chSK19TYjWEt4Ti22N/ZiCU84I4WPDQpgf4+Bybr8XVZiECltqQGl3TVBykk/OxvC7mRXLHCC2n1
M9gox3G/mFAikMQ8oLrvaJSy1c5B5zns4NueZ+OrZsHRaYJoMUprhyJIQT35603tA6ALaUosoZcV
LHulkFnQ7n+Oxu7z0YaA2q2dO76PobSV4YDqvz/TZo1TPLjgZgDFpQ3TWlMmpS00tAugA3RoBqsV
KCzumQ/jdvKac05N1Sn+QR9WsAWrilN5988I10CizPGPJVaCfMSExMZNDdBsjFBrJxrjaUub/ru7
NAU2UY7yH51xrh+ZuMH/tOj2d66hKnNlJcKvrpP7qagjWtzqnOs2OrXKZY12DT5hRNqYtOA1MqYK
pRBn7BcVdw6SjKJZvoA6Tx3bC4k3FxQPTXTolMSjBgSlAYD3Bbf0caxzhPQH1oll81+dYCLfOTXF
FxeGUTSXGFkumgHFFsOWhS6QdWFTYhZOvT28bF2VJW2PNa7BhU+DIhJMejcsVkeE3kC9/MnJCwR5
7Gzh51vgDp3q00Q/gElrjLPRVp/4vR2wsA+WKO/XFUNw9KGZUxQ1FwKK5caA+CI6TtayX4yLqdRC
eB02+GRel8H1Nf6i4hSjUajh3abaRjhjd7QRCy7bHPXdb6pXnxyjnbPnKbB450p4E+vrWJLQzl+K
3i2qKc7EMBGJ0VKz+HBTvPDMexAaZvetvH1FL02WT61zemvMu/JOVt9ii+dPQNcwUxOVbKX3Dk1S
ylhb7JwbOFXhPrKNW/4CtfwApGG6lwpxik2dLMIxsoaz+t2/065s1Y7aZL3GZkM4EVgkjwh18k63
Y30jL3QHjZTysFRCaenlymJ/B61MprWkpsy3cf8C2oixN3hDbdX/dZQ1iGV76mbKm2Bd/HogPxsK
Nkp20BQ2JB3UvSjYcdaQAhhHjBqonqhNg+WQG739KiCaZD4N9QZYtDgGlh9/L3tVAJOeEB6i/CZ6
6wTj0hfnueHhmTOhlGm8bS2WJNqNWc7GsegvYrwItjRynSZVk6l/4AncfnqtPb3uXIqx7Z1kBubw
kaGzh6JI6ok8iTFnU0K5O9OCx5gBcpz2G2NcJgLWSxNDdZjEUy0ZgoSZO2Kznl+L2BJFhI/GURfh
c/Ya2trMCnmrRE3a2ZjUSOc9xLDSWkyrHZC771NOXi/COaSVwyLDSdoOYNjcs1N5947uRVjEX/HQ
T8HEsSKrztpgCBByFp5ymmxPGcV6+2rikQCEJtTWbAAWJPxZwVKSdXQ4Zz+55AxZU91K+GPMBazD
XR1I21hDS7iXIPljETdZDGD3ePua0JR518pY3bMYTAxejKBqjs4R7k++RwGmX/LX+kFwCFGNY6MI
4rrPl8WDBhXcG+9EpBn5GIa3C5APcyBOkVFB7YG2Nk0h2SIBEJCXueU5L01F+YpfS5MVVRglm5CR
jxBSRiK1+O8fdA6IjPDe+gEmoVHPRSmc5nrSjZ7W9qj4Tb93uF/Hq2tlYK3XvdKwYmumqxRmUxgZ
lqFdCAtOY/i1zDt9GPoXqdZAEXWBeYdKlzzPf9yhJaIwL3m3uqIclXNLQocUYcw2JCI4rvSyPqnH
ZhqCZYcupYEW7a7S8f01sQbmjm+egm+mDE78m8WLZ1dsAsmS4LGZohwLL3rYegAtnlIYqGk+BPvw
HWBxQtghL8aV5HgHfBZHK7E1jbkgEbtdKy0/RM+CCswcbcPIUb+sQKtsicctn9g1Xn6h2WmRfJ6Y
AVOfItouZvz/P3rQDJmoOjRZX9fXm65yVw0WiD4fuu6GxHyjHoC2DEi2cyKDo2rUBs5uEEEneXdG
2iPl3zLZlMgaigIe1nFhjIoa8T07MYSTmPfKLySBAk+I0ajoT+orngbLl/pGHd7NnXiAUbooOmJm
aDc5V4c1qWNVvpcDJDCISjGSfoIRyIcFcivs3B9EincqXiLNhLMvLPP+IYg5/f9KqYWTknWoop+Q
FBtxctTe5eG0fVz7jaOKTXIIcoBfXtBIXik/v6elp3i4GBmB06+5UvYNyU9VIf4L04wgvZ3vrmvr
KTQjX1MoV/nKESbdlv/PQ8TiOjJi0D04nYNEPOoThXcYKG9+4p3Mxn+b3JcGmkvkuZ+r+4hbjKnf
VwG8FbwTAI5mpngD7qWHvG0gevXaLNTx/shCKXm2AmXy8TqXiTw3l/Ib64G6F2Js9n82yB45qDPW
d7gqIHdhSNuR4XvNR5MxOdikLS6onfxpB/Q8stpWSks7mX1YKZgmZJ7MESp7q9ODOB550Fb5GP2T
lvaBf+FW29T6k3M6MrOpP5F1q22NZFIF1s6BTE9SUXcpTw/0iQmptdoZL151HJOJd2NiewDbyNNS
145rjmzb2E01lvpn0FJsVEiNRRe3YskFmwlM1KH1riS2dw2fAljolN3RS2GgQj4GLNzloykUMQ4G
2VZqG3vN5I0CVbaQDX42Wl9PQviUDPYQBz9vB3O/wKsTlY+3Jctnqgidg0kcjri1RbMMMMiH9jxw
Kk5gvsUfxeQEQb+UfmtKERWm9AR7OsIEvT+61hIMWRC5zvnlGiifVuD/KNfJtsjh+TXVPyO/Q6Rd
QSi93N0+o1mPRHtqpDbu096ReG1JPCUN0qp4yPOsTTPPuQuPHfUthIqlCNVKrYY9ZeaUFCH//Nky
bd3pG4HYYbHteeJXVdXvViURN59FXVu23XwE+jjaHIQcUWxjbYg5UU+GVELPhxBAhrhNP2DKkO14
ipaj1ul54TUFGM5f76rUWmqyJW2spnBihagdheQKCJ8DIXdls2x0fishRDFfgeM2iuQU6SIBgEsu
LSG6wbSSd/AQlS1eErFiO5PWYGDhRHno64h6gF+uBjP8yqprsBCnorFRyii2FEetMvPIxXBzTVIE
nRVZHrM7VIZHsP6hgPzVOtZa4vYs81Z97NLjTrVJGnCENp5eoCE0E41WW8XVbO4LD+/6DDs89jRr
iv4sf4s13sO+us1r5+Ceq76sh2MoAj6wCYJTyJhP7WIsmefI8TvywusJGEj1AT4iJDiB6MlXYC2d
q7M3hYEWBu3qGM5aTVEOTKXcM/VL1V9yDh93jbSk6VgquzKhiffXHZ7iGs8LqMJhNbPS2pWHPfdM
CJVqRVzMV4/F52T0VgbJRg157+wPNAinfciHiQEBvJ53vPuAxDC/zvkZ5J3Mb0p/0ncjUnIzDTE6
wBm+g6VMLMQG+HYMlGm3RYWUid2POdArN3ZumkGtPDqy7arOFvq2Jxf2/HfIjbxzs2U+UEtSd8Ov
ddesDhBSB4enjyN/C1UE5uDH52fR9DyCBZUFSMUH553eH9nqpgro3CXPlkwd14h/z23b/yficjXg
UztX8nYg95TyoCmLeNKGV4hXX90/naQCEjZY5SqLM+0ab5OFGaIFhFTbz4tKpYP2M+YzAJFTOQND
MDgkB9i+YDOesJxrWlnmG7/dga2eGG3y4d2AkQ+zUSgJIvadbKLTmscaPbb3MJGbvs6vCSjRdygG
M+YQ4mw7NwdwmPrOGnREBie8K+QAJuYRTuWuwbT1HPhiZ/9s5ZAsToFImOKOWIe39Q1gF6fmNUQ0
f0bVNhJLIMngFBa1uC/POjeredhkO3tf17n4+Qqz5r20hfP2qBd/4OdjDiLIFdjZjzKtEOTOTZqU
6LqFutuA0ytTGYVNOlU92Nsm+mQiYz7n5XvNEbrY0XSDopoZsu44z5Rc90mSf2McHSwA2eMVi9Ht
38Ni7wNms4Fw/wNJPJDuGn9V49PpB2iCkDrRV6T8Djp2aewd6t9Vsjdu50WQ5F4vV2/iqf7Tgo2g
qIstnH2io/qZLh+pB/vDsxnE6LTYJ4gd22pg/19sfPG3baqWYWPIgIASGJ0IIEGFCHj+1mhoJ2Wi
xXd+5pBkIzEI62c6epGfYx7PFVzeAeEQrWrqRZWfbTcPdbqbhipmx/cmiYKJP7yaH914hBzXsAPB
/LYfohmz66zfzyOYHmLBa8emIrYLYmk8HWxWjPnIvmBiBgjcqJpLB7N5dXH5Xovd6lEZ3iacCakR
o9MPdho2qSeXofvEXUnSE85ABIheOteX7bJlBmrKqfn5S0ZqFvJg9AjucCsQZwt/zzezy2qBopRM
8UBqkbmjP6Ad4/guZGFZxI+1P4x4TAJXIiVXBFK9x69jXr7kriF/EhMj/cNCy/FVr99TbFF9BXA7
if2nvFU5iSoL9Y/sQEHvofecNLMQa6S5sprGOYP5yo4ALvJTJgLUTIVJb/BKOSSCTFWNybXh0Kvr
3ytgFujmBNV5WbIGKf9YoEMcLyVWnquA7WzDZ/xxiUBBe/PIhFynDSOTF87koDa8yzJ5lFidA+JN
zqjXRfj2UVODM7YpMMPkJn/l4hy4zKKd9uL/zRk4d1OQvaKIULoyE7NcBaKEjz0EbjPo1pibqvFk
DC0xXSLLDIL2BP6666pdxBmaYcUOj9zKY9bpehTUFCAbkR0x66VvtH/DB7aFGQLyZY+WFMCzhcAi
8nczyR6RyLWsempu0NqIDA+hK5yvLkdrRzhy5tkzwKA58onmLmXcYc9Hn4pn3CwgdpDH+fqJEkGV
gNg1e2Q0KOZcyZg6piouev0Cm4l3dFZkvNBYzK99/Z0hFP0hWaxKGy+ezRgRKSDcCyjImrBhCwQk
h/OvS4HzpWU34zh+tSSJp9Xz66FxT2NxiwBW38LOYvBkCOGmuLVStE16j+5OoZTbvkM01fxtavsB
QdWgBXWIzdnx0YZpI4HNXkTOuU1al4CYxfEHl75Hdap07pUFkEQdN8bhYrw877ryskZ+kl9cN6l/
9nn9MaqqeOKAQXRz7GQBGgFXuiHFJ3+fERJMbVtSV4tSnDGxQnfNs8MycMbhatC/o4OFZkVc6+EH
+Dc6Zl1R3IvjEIULHfm1MYeyEP+mL47BQ0Q48hIrAJOKCQt/TV9j3EmP/DMO6KQP0DeT/zUXdgWl
eINfbQK20a2EzhGhf8Bon+znxWZ0IN73gMLshIjSby59/6ybv7oUspUGNcmDWcYsDWMyWibGezWH
nGrnpLN4e8Adq33K7WWthDTCwzytUR5tRPtLNaXgsMZMsf1LVpZPwSNamYwHraGq3SY0CWQxlrc2
t+F8HeaepNhfDLJKJduA/2J0XRflY8h9r3bP9SEz5yAOUoPq2rlaVYg4zHeCKov9b4lFcRRlZpVY
NGOazjCcuSIQGWKOqvwSg0mcB/hfPbR5fdDKs5ShhB282GNa8wRUGt3bZ3aL2WYmnp4nTaSRY103
O2QoJN4L/VwxXbi9YBA/tVnWi/Z0ipGjE3E/k8gE/A5OY85QilKy4vVI5ga7ylrjQen96oeJbjQf
XhpdjP2J/nTofN5x9MLzdFf+eC/7ICGcoo+mYbyJ+yOpi9qLVQBqmofKV5Oc3BxfZgr8XH2JwYpk
Qynb2BTKb1hQNrX/XA2XdReBuavESomqq80EkjgcV5+1oJs7SZ4RpzIuNxYMBcS0yVaFYtOtwR7e
1ky0NvXS3ueC4YqaDH2C0QJeTKL3N/6UDfusHTAmkIhJGGJLAXZMEeeAuHGo6G9mtRNrxemjNJD4
4E2uqaaS76jsiw77DahaS+N1OFuU1i/AlcmvbiNGyKF4rGFBcy4DuRWQpjq0fk1WxI0OxrHRMQhu
LFJJaolVRwDnp4BSjXqcfHji9/6qm2sg6PEUOOd1ShbOTqb5OPeDhEM4tsLADCrXSHSDDD8oX1pA
brp3k9ZpKqSmewDSluz+Bl761oxedlA3/3E+sZFrS+JC0fxztRgRW/ewoMwlZe7qsDXQqteHwlHU
XF5DrdVW3ylFR2CXwkEFMEwy/FLzvxzDy8EABuswQA7oOvPQM+xeWNAKCyEEdXu4b4FtZNWvdGV0
fnZR213vTGX5252LVAproc7IHjmnPirWBWrz18gDkmLHz/sIGW9mHgwml88UyIXvB3WQKcYnP32R
6j0s8/TfnYpUnZHGuir8frffPKOSmssRihQ7lhkPK4Uft/DnInOPvvVmpN0XJrSCTktGPcRjli5x
mU15XS6DZwfJlt7tzbmSocffbRqGHaaeIEgc12zSDAooQTjufIuh/U2VdNYy6EXWY6WzAwPmvgzM
IE0OhkWTOm5UKL4lmL5wwobW2Wsj6UjLGMwJyLHWeu6aJD6XNIOoQYFv9HArrSMP1Q7gHfZMsMFl
tPr1M0jRxPtd03dsQpWLi73TasG5JSY8rc1YoHCS4/eaigdHZJzzzVB+6XfzIZru2BGfA6faO1vV
fHjof6DU0pQYT2JCinTYdt3AQaZxp6V5Mobw4yX8yRSp2B/SFP1WZspCgwRr1FIcBWTpG2XoJTYk
JvGrujeqRAkmjiBUuDml3sUzQS7aKTv2kmJ6hfh8k97s3naoCTFKca013KJoUCB2tnqq15x2QOvQ
Kp40+Wdptj2MCepVlkQ47wHC2TT4ezUDtAsSySfVAtIEbZFcljJB80TKdqhkCOJm1BP9z35UCL/q
lSG6vNKoUCmYm/PtGnri0t+4ZOY0Idom0p5z8QG72nI0m2CoqwonvsFYyvy94odykmSlN7udgTCC
pagB7bLjrr2HcYo6ny3Y1Tz+XApfglUieUKojSAIiFyarnehF46mteXW6b26Ia17Od8lXFPV0nkw
Afaq0tMAKO4VwW6FHHY0uZiyV6ARwnfbfeRK/e9Vn6VPr3n+ponz17sox1o2KnDJxlYHf2V/wRNg
eFI96C4klJ6WcdKjXy8jJGL7nd/q0QlHNeoD+mtxYy/kRsE47KNLpqQ/hej5hN/IlrYZ2h6GroLs
YariFEOqmKZhRgglfcSTIQ1irY6ct03wjgLhk6+w1W+JvznLEPiqAHwjDOo9vKCqTfQCgaLl7WLg
LP65rycWlSYbnQvu6oQuwSUPn5QcvGyhZtOplU9XWrYUPmQQhDjj1us8uByWmo9Ha2H316C4qxKv
4pYPfMBpqjncfUezQrSClOnOS1vPYwlCma8qjwcNgfKrNMEE5jUCeS8XoTR6WBOBr4BBlPmx6tJv
RbNzIdPXwt1e6OJfcX0kCrageCKerd+uH5XeBlpyPHs95wchRDxICaQ1XYAkOoa5FehwARZ6VW7h
iPTlRJ2vOAMWVx65opsmMqnrxSm6BCpQgMeSof0UJhjrWoaCEREcWofgHK4o7lRlKi8FUAhSd5RY
Rt87kG69pR7xQYAhKPWdDugMmQo+prT7JbXM3H79VTBSAs+ZcGRuzVlR/XjxtNHDDUH6QZtHoL6c
9XoMCVTb77eQBbmZEgHXcOiGJ5hDB6po5qxfTE4XvzGE2+2TL4OoRJRtsxHQbdt/nm7oBqZ501Ab
mbs93Htj7dUmseoRhMyMIwFP7akrk8a513rR+UWynan31JGOQ/qtTh3vBxMD5CXLq5FczKGZAlFu
QiNVLuA1RnYcsYB4eZ23PGBj99AqLcHv2IewD3tX9a+I7zNSIoITtzpljvSO7YfIM0o2fOfChs0w
Q75/anPoJjEkbBvzmx7ylaxcVp79i0pYCFL24judGay4h+JwI3Jm3G9Ip1HenL7wTpy3eBSu9zPY
rIT7oCXZKJ8tBFQcSYDnNo6MsfbXbIJaKeyK2cqOnURlxuk3IWwJxDYLa5RUSV3avxYhRRrBzYw1
8WEUbJGNdwnOlLieTcGPHrbMutMrQLExJMn1tZe5QvUvcGviH6iaOABtt3y3S5HXlkFsdLRKtXyx
/vqiLtXDx0XaNGoL1VLVcWcGSb261209REnOwjC1MUHJJYWZ0y9jMCFA1W0pM8ZOBLbpwy6/ADEF
TvTsxDcQ+iyVZ+zxwlbVXmMLkfDTu8bsNV9Mo1sAMXgn6Xxr1FXtAJMfh986oCfEi/EYhK4qzOji
8UgzdCCdbDGBLApzsuGDqw2ypJi+h7seDlnbDNr26xo9MJUj2aFWF+GVWI8d2nbegUB+C+w7iqtd
lxyFlfTJDOq9iTA+sf+7MlEcfd5VBd1vnga9F5U8QdOlCMP0hOCzBPSbKXQlhHtB5XgKCtaQ2Pzc
Plb+b3OGTzUqlFbBoKhDAi9jMj4qM2OObSn61zEYTd15VAPR6vQgQdk0AwTQ1rjKbUoANUS9kSrw
8v4ybQkW5Q2J77+XeIQhuulP8E3JmrwiPpPngZfnHH43LOOX7DWHXkjdtbANLq301jlZhzXzPyV4
swE3Mhf1OtF2hPCtTpGq3saP/P948BPI2pNVYGF68SfnNDK7K3I3VggIwpcINdzLK6Ap4hqofqfL
OpobhuFYLlDjsarLdUQ6N49CanBJmwjhFna4JH+HodhoFPevjcZ/iim66DykE3UYHxF5hBQdiE59
EoxcT0jLxouR8R9sKj1zhmXSCmw5iRkmAsfgZQVAMW3I7tSI1lvdqfYcjj65rDaMaYf9I1Pv+zez
JWIJZw1gPFVlqTOG7Pp6DcNf86kvkMCmMZ3i9rrCPEm8N9MxakBsldnRIiULjYV39TbdxEQnBOft
XkeSDKqD5lDOKvfsuc5RKpWjh+PY9ei8ijGUHGp78dKzImZNF8iRgUAA0ot7sDlVRrsrSzbyPywJ
Ay/YWHaDOtJaeidvAUDr+OhaSy1BsNGSVfnTqQYupn4MEUc16jsKIBpjb4VPv3WyaXUhXKeUCA9F
KYhwSX+fChDVDsPp9tkFl0akVp6x/nqaqdqaASwOYA3JF29Tg/72ezRx9XsT8iEiF8VX7O6a06G9
BqKk74EREjexMHZIAIOSfm/98wXSG96HbLSD9NaXfzC3G3jU83DYXWp+Dm3zaCzMgGFLjZ414qGn
VfB03dph9Z7/3zRn8+1Ech784HtqofWl8tMUGYay+P7xW2hP3OmQN2B7GmzPcJej22Qmb8OPbD9P
VX7h09K7/QewUi/P+OLT7YrCHamgCocQb9B60iGJWDk2WQx2EZIdEepLmARORPwySES4Th9tMojK
3SjfSGQjrn6jPrUg9My3MlxyC3egTwbqmk9DSvcAwtQR1XYG2AZWfOyWn93sJ8vHdT4LVnlcBvN2
QcgRCho7A/N8j00X07RzHw0q6N/SE5aeWqsnVEAXya9ZLBMK6NlzKgmBTO8R75PKqkhfInX1PCOn
KeGcTBVPqqEQsxURZWW1kyPOaoMvH+OGmaG4RTcboR/ep+1b4hWHrb/ZsmEWAiB3QIUCgsL7Kfzk
auOscykPVCzH5cOXJNkoS8Z98Avwt1PpRQhtb2mADQuCHQXiE+y0AJK/L2VcOWWOR1/BuKhwUGsi
mAK60yFE7tUeo3yovEhywz943s5OYFaZnwBY95Z2E67X/XMnRez/Do9xa70FZSV07k2OFYi3zQOI
ARNR2j2XC/Ks9K6jmJiMxhOPg0aO9tYmx6dpNvt/ANk2R7wmmNwuA4yKY+55wqCLSaon25MCffu3
NyP5n3gShKcBnYCZSa2EBU2GY4fadFJXRVzxblRP6o1ebrIeE7xiIhB6tDVR4rrTqmtR3Kq4PZlb
ontdtb66L+w77pUPD6yWjznxYOBsgcRIHJb9A2dfHtn+lA2pLMzGQjyB2Zj64pTGpDtwLdW7z02w
mkWsoRsRq+GSR2eTjyryVkuOETM3hyg4NEzPvNm6wqehHS4SPIVvVOHKvX1W1GjiwgytnDK4RiBo
6ubtdJkrVOc1DQtkJdBCL9X4f2F3eI0WWcgq/m+l2AKXXZKdh/nHF9QHxhmTFeehmipIagIqDEQM
AXg6V4qKRIf1/fvbLnIqrquBRVYqwRtq1BSntYOf+eGX9kRh8DVyDP8dfRt7641cLHv/cIzgA2jm
2MyRlcnphzSyeEV8Iyv4hU4nCgNorcQPUNlGUF3cGYDKAkM3zcZ1lyn2xf29euxQ+lFY8QC7azqi
Vzw3bRX/MREy+/RyABZ0cTvdP9OO6mM0Jw7KCxfYSAFnk8q/ijvPzk/MVqPGYfMUsYMZXYUbj95G
A69ow58pazjXtzCYkmpHhta7rrTdop0DkqwfgyeVVWABhFXzH8iUDmP/cLxWdLE5BvKUeLNvWaAn
rJA5zZU35y4UIKaVbHkjIJXIBieF+9aAVx9QBEjFQxxRGt6mP50CbWoNSMehp6EIHtnlwDyJB5ia
zPdjDLJK14/kYkxiDUNsj+UxxlZU9iBY/s31IQ4p8dH12kYLxOx3EcyxDghzU8Nwss1Qn0HMunRw
/6pYiKOKWcO56cpVdcU2tlJkZq8QWC57enPvZNXRSNgzRE0FkkvOFS+SOi5HthFD+VTn72K45EDw
PzHXGd/NSX4BgcCYQW40mhf4R6P9V4ROzxSzIZiJEAuC31KD53SjAXtHHNRblYH67Dpcw+IwWPA5
xyVVIvbJkZR2lc34MWupyG6ExO6E7ZX42Cxe6ip+Xtv3V5HsoWdqKQrxkE7LcCiUvVx6Qd/t9Qgi
YHvbY5bIJpNUuaC+KeekL0gPtB3aRovnT/MAr0FkzTU3QzfXyQW7NwLv2+UdHMw9uY5fEtbHm3p4
zV8Nk7kbicxTaxFzUwTfxV43F7CzaODqe7ENToqse5HCwCwEMfFXOrMZPXGmAw8ZW+SBrpzBJM+4
c6lI8hRo9zMoKUEZCkMo8xojatyxUJ3pbyZM8Q0OagP49pnDbxyfwuDnQEADcIQ+wKTTiKsWExLA
BHadiYgDPNndgRO3h3mQqePe7Rz5UHjVGVrJjNldqXP59VmwOoCPRoKCvSiuIh29CghE6Glr+Bv8
l+kryR/TrQINfgl9ouBhWJ2LdAutJd+VzZgMCQA6mynBy++Pd4YpvRww8kdwRQE0EqGlG+iIOMTP
2VTFFr63C3RSYXvi2AlAa/z8q/tTOUoEwTmHZs2UnpEe4PFI8AO4P+okJPMn1n+S4MnGBo0ZErsg
siBLusEQ2i+GRPnF3eQONEFPQFbkvSIXoMhxGE6zlSNloEF5g2ty7M2FBr5TCmFR6ZLDH1e3o4pB
7uRNQjcLx9fHvXm49ptg0USGbMTO3bNVN+kF2GQeQ2awWvUC+q1FdxOIu+aH8JvtbKxISu91T1X0
xz0YsL0pF9Eg0z9kfT0x9P3L/WLGsJbsDoVot+xZ8utHLzZvmETFhJ4rAgW+UAysHMYYDg+rKwQG
ycU6wgpqcllrmSJmnpfBG+APD9GQQnvxZs6NlvzAZ/lFS4grmonQtpA83m3S4fu8k+vtJgVbnC6g
vA47BU68cA1ipYQJm5kkUPGF6bQyO8E0XKj/5ob853F0Jq7RdiiGunaW9zav5B/JYDsSyPzrXHkV
0uUkEN57lom6Ccf9Bw1vxYyvdOQ9X0l6pqvgo9gowjuF/rCOrWj4Wmvgub6+4VJAyP6ZHS+Iz6r0
VexVLLLts+4lSCZL5V5DbsWZc+SSrK9QipK5KqF+yEy6WqOzpehYqU8+5zTh36SDBau1VxSBr973
jn13IFEAc41t/G5vYNABoIJi5Zkfc4mnmfKMxsdfHVfTHjexjXDGKZdAuhqFuoZNKwB33j0rEBes
OPNSlFSf0Kx0a+oCc3WNGQQCPVMQSKIj4SyAVIvOr8Xx56Spqg1wDnQ4iT9lfep1F8FNb25Gw60+
CeRqsUkvP60a7sogHw0aDtqw3SLSHBngKAtKg3S2SeDEbIYdhu+gwkU5esBVU2xnO3OfpmZQlhhA
O2kDebmBfhXHlRJA2mel5zGCEyKWSuaXKLlMOvkk+cdH+Pl/mwSWBuFdvovNI3voWEGOPhFYoTHT
HxEmw8+iejvZ/D+cY4xXpVCLn8eRiQidvPW3KQuXBPHqdhF5/sIcDIfcightMCTwTkoqTQepGlfK
NMnnDUBpXM272gzsqgtiSW04ALzQwFP3XzqL8Gh6FDKQK/CFjlzeNERpbBvzfxt9VbdNLoG/BDE1
IUrivrkZoYOGc6NURZ+6ADGAJr0iSEeb0aAQlUcavLIeqHKGJLGQIBhkVFjlx3l0UGN3fR6oJFcj
SHGiSXWQmcY04MGbDKsaTwUCBU2B27nsjsXXNbHr5Vm05UCXH7ml0FQN9y2WtPy/lRuShfKbudHQ
I3dTH9kx15KaksA1ecnmQYYOcLiQawMtH0xN31WcgEtFzAWO8Y3WO8iINiE2TJ9sYvD8NqzptdyU
zr08niMj2OnTKE7Bx3ISw+Br7i0hG/yICOMFK+2zXha0tOB/k4dB7ZLyRC93Naz4mo8v6EsL7zKT
mUnGUOkM46sbB7irmJNwnJ189E3YHdR/gwuQs/tl7Fe+0KwSuGjHEMP51zvCuvQLUZi2INgHP9/g
atJPl57xhhzWkyxdJAdJUFX6YHBFS/hk0wszJknIJlYFocwEQXXL0q77JM+jqBI2oOZw3G29F1sA
9QfwtoQy3nyB62/bvhCHhbWCLNwAJB19+mCiVldHS2C2CTIFYO08h0HnQbRZtdz3pJ/UtfOu+J+M
+t+rqOKpOWALv3D5l00ZhHpjM4RyjBMRAXO7xxyGFwmkqeF/qj5axVh8P4aZmfkmQo74KYRFt8Kb
m08fOQMqZygClGuqlBslnhonOsYTkPzC7PAphwupPprvCBXSI8rha9Y+lyzTZdltRHmANhLy81Eb
kwwoO+6Jc7nqS6O6Xyo8kR2BMxviVcizPF3ItAC9nf8mwAcEaiDAptHr/7CvX/7mEbcewrDBP+rx
hf9qXnhmY1rfTYXZFPcG4oKLeAUYKvh5t5GeV3R0IXIMKI69tJVxFQlPqa3qJEOplnK/v0ffsYCv
68ZLKOSDdQLUbV9wlsiQI6j1yHeJl+Trqet7zq+TZ0hixLd71uoOzXxaDUJfLgMANBlZczPhKsZK
VQQE3c6/QBblqRWorgtne6QIlfBrxqKeaFfqV3RsDGXr+Fth1REdpPa9wtEEuRVuL59LLKeIDcgw
j8VjEhkTCnzDu08T1r8rVD4wkwG4Fg6euRkcDr73e/MIs0GUttk0683eVnsANgNIhE5L0EVUghnk
KbLm9wpRNya4T4Uo2Aasb78N0WhTh8Mn7OvtMnEEQxJDCo4/+CnXcael56LrqJDqFIPBSOpL5IS8
YHGPJbWGlMUPeQueOWDOh0QK/WCYoF1zuoZ3814ZTlOCIQaeQa2bgB6MGeIvwbpijqV3Kfe3LPWb
eFDhYGlOJTIOUofCvmEuefRSnIWnVWu+YEWT1oVNlVeKrKEkRIRjFOMNRjpe3IvHjPWeYRhzsSWR
NFGG2Ae+WvjoN2SeiLvLQdT6EJ7H4IYqSm6gYZr21mVf0eQYIB/T63arr6GlpDtvfapv8GuwVE49
DOc6b9TF/VOy/ThnsY5S7MvcU9nsoG61jCUU8NBOJp5nmp7kAflAGcYofyucLTtC7KvOt7EvCmXZ
RLEv6/HabvJbHMMRUvnmnnRr9G/x0bOtcTbPWvCl9wWx6i9dFQ/x6cRbCSyl2csKdLU4WGQcBOi0
4xQqqgvwSw7YrkCgRHtdVl2He9qkRaqx6RyRDZ3Fi6j3u77VSBMo7WC1G6sbqFanEntH/FYaZhnl
Eua1cPJaapbFCbuVjROLTTjf+Ih3B6sVokgJWNhh4eAv8eFKy+as7b1/sPvm6zQRyzW0ire3sFbZ
Kiy/SJDgajU+7HKEojsKE1qeOx/7fMOfq+4HPc2tQN/9GdJaX8GO/6Ob+qLRyU0vxtyX3Cr4OuPO
izfU5cFV65+Uriw15jrChYytNSibKSJjjVXi2Yl9EqvNLaru6Mw08DtfiPV+HvFMekr8M9j3i8lU
GH674szIWGi7S2i/+O/A0Dk5n4d+ZSS+25PHrTdzNfjF9V07s+dF8WoU3mr9X2ZT1uadn1PBeVIK
6dV/yhnT605yS2kDVS+Z/52fDPa7+jy7i/IzYreUo8b9A3646BSjH+tGBWm/wEBNDKy+Scc0P68M
ILNL4m9J0mchEl6Kf9cXcr/NmqenkWyUTqx4p3Ey/tK5jvUHt40uyQuTSvdPSPK+44X8jzPgjs7S
UwNGfV863RecpRUyn7uq8DCmO2xeI96aBcvaUGuSrLzW9SQCo0L/sHND/BGiKdCIT93sTm73cwtq
XnSmpgm25iX9U0OOz+R11zcp+sDR1hyJVZo1Y1AOkinK4cwA7az+WyXtKsw/9RUAQD4OVEQunfBt
Yy+uJr+g8wsuJiwp6YcrDjr2vTC88kxDc/V3QLhWdsQSDvUTNni3uMQ5Na7UnCMaDEj8ltfE3jMd
6uOWPdd/tVSf/h+2EN5anR2H7Wi+nEEW+cty+P3LPk05Me+UrEhTGpTbHk/QXtp9t1wWbqmVyDnW
qVqVNkkIXRxiGkiBcctSnpuh9b7W82STL7Zf2qR9slDHHjjdtmX2LKW0kaRT0fprppBIKo7ncAXE
Z3DMZG3qHEA+ll0HeTskvohgJojO53QbFKRfp38NPW6weezm4VU7ANVtxP1lJh/B+XEL2ONZva/l
7qzs+TzSBfkpdpEw5F6CjTS3ATaep10glULZfkzn15hg6VxpbvshQcnlBg4DVneoaAcKt8OFtEhF
YRYQIu1E/dsNu7wI3ICtPtUH7zpNSLLe8d8USQs6RRY+VpzWAOKAUDQQl0u4O0HiJaIAfmKF5eMT
fJuMRC8EotVldWw+rBQEqBFxRbs5LTyvSHeLM9AfFOUJiKuQvfz8yYLY24UzspZsWU8jwXYWYDJG
0DcArXgD029O1zUN+isjr1hm6DF1t5Cz7dsjc2ah4fQ/2fh8jzgZQsde97cBx/FpeUo4OGoo6l+n
JnrAsGzBTnHG6BGGQgJTVy1bWAiGrCJ0sNfPs62vdKKNh86UVtr/FXc2yQIG95NGNGpm2888fv+L
3b9ZPdoQr3jRentwj9tgDl360ECqd6jCpj5Hk+5ctC37tgYDIM62/8luxIaDiiajDgUGE2I63j+C
4pqRZ4QrdJMdCKG4XTrkLycGivy/zcDukyClV8Lrfs/Ta2AkfWcxNMU/MifBhnCDISqHui4BnRQG
ntX4Zme8tqHlpYbh40Qq3FLwdEP6gsjn5+nsNgSKvuSLowjggRIPic1tX5yV3zSIFkeRy4JnANcW
vmWZ3BVta1Qg+maNnWWWhL3aEEun5nt8HHI50p0kgFLcFeBswo9fSj/phoxrigkKQuHnpBWr7/5I
FpdqyHDzbfF1c7Uhjkk8yHe/fd18mBbF3wTc+MyK/sVYlwzeC6Y11ABR7K82nS1qxs/ljHiyqRZ/
lZm6g6JWsLpHjSjca8wHJ7KD7bbiaFlt+fXfgpdPm6qiXUd4qJ5S3vVWEAElqixW1K6i6Xip2wz6
O0Xc40hH/3jN/8OPV+5KPd/Y8PqKDaWI4wg1YeaXXINg0XQh/f83a1B8alfQdBxOPtTTHJu1cZ5o
h6Ie5rNiqV2WSq6jS9tYPIFCocofz8mrWsVsZhJIwlJbYaV1Mn0vhXcul04G34y1OkjKtd5DLz1c
CvekffPndv7KbjVqtDgOLgfdkodNhupSy0h/KxQyVyNipi/y+atHUoKwx5udK56zZ6yJyY1YG0Ae
0yBgpzH2PjhcIv2vW45QNdG2sGGKCK53vRe6ETIzsASb7tppDmmlpW/Jw8WhSEJvnba6XvA7hNSp
zFbb1qogpboDk2edbOcsjxJY59V97nE2AKt9gt4i8qS7e7sPjb+l4msrRJWcXBADMH8E7oukceRA
RDluRDfwjJm8cwvcfey1/NOaHj3MjPoJ8i3t5+0tXIU6raiKWNmPQA1gfpx+uWdTg46J8U8hdNMj
unCPdvhSUNOHqHCZP0pyl0TE6hBXo0alcVN/bWddAilHYUZNJVruILgboUGGnbiJGGVDZUjvqeCv
DIunKKkRazU4bAXD4L5NnKwsOcSZEVNgZMUh85BN5k3vWIQeJPlqJexl5XVwJf2T+BMaS7lOJH8D
jEJIoMwEwS59XwmRt1rnf9YF0wx0UG+ccseeb8bhub9Z+ekpe3RV7urbYUJEQJZYSpevqqO/T5go
LgpgLulJKXzrChl7HxnhMyUelYPTc49/avfTaXRWBxh5/6J9afrfUp9zOacRw06oN4oHo41Ir+Vm
5OPBVJY21bxvabbtte8HMeU/1XqG553rLqjnpkbk2Wq4eke4AvdIOPe0oQxYe2popJmsc89J1+nj
d5zj2UMOfBI4rrWF8HoFtCq2w3+gg+CtJc3+xBmaZf8NwGKgXe9saBICj0xHHDXXg1FwPHNBRpps
uD4wo5Mk+FMgD+/I24+BqELmE+uCATqhNYjw/CWIiNxSYFabuQ56+gAvo3sdFlTpxKWVSninvx9j
Cnqrws2N0jwyq1qUZY1cE0Gamd4PVJelHwDVR3lJWSFbmqK0bwQEDFuakJVkJJ4hPvMUAOSKR5ob
yGUThpxp3RJKggQ8pOoI0UnTghNuTGxldDMzRQmrf3WVEcmf00Gwcf7fofah2GC1KDj/dAr6cwFg
xD6ThR39HmfilNLbxE+64FilfnScZ1g+7K5EKmkqVvXPoVdItR7zQwzxoZuf4/yJMLpHvj9W7wAf
1OiQQ3xdm5ADGUVyUWFm2Z1PxD3cLgK1UUif/Lad8aY0WrjVsYxVZnLCMbtOmkhd286B9ke62i9L
9H9+r7sDI+28rhorsnwCXsX3+EETm+tlR2fdkOUsNvNunz4w5F8U4PL+s4z/AFBHl+1VE8ci4wu/
X7+oCePnpq/oYoo6E4bMcYHNICXxJjMkIPWfWtOIoHM4u3IfxPrv/sNQ12+l+ZvvnBLabj5c2bYf
7v+Jm/lbCkqb+cuuajmGOewUx/5uTIGya1XgOsJgudGk+QCKO8bGfeCi/1o52V/1bIGbx4IWMHAA
q1H7//+o3eUw3dKmEGQYc3LZdUA5iCCo5EQzOYI8nlasVLlGAIETWQA15P1b6eNU8x+n4EB2vK0R
JkLHK2ixB0bDqDMidbfCGA3c2elkC6Cz1qOz9GVVepe6e59exma/xqQK2xoNb9/EjWoN7a2EbghE
magSMZnIRZGjCq+nigJQGeUi6SmpmPepjEmAlBt3VUvcI1EOzmgIvpqSZQSkP4xke1qGClNQ7gXx
hcxdNBgSSTwCzCo4J6xcQDSTEc5uz/Py2yXXBgEniE3rccmkj/5cJmsRklCx/p1rMF7jZCJnTbUN
SGKk6Rdk6qgHcSgOIhjcUKvSaXPfKunvMXqdrznAV5O9TYsmfYEfzWgRyR03uFMnlMZceyXvDTy6
LYzkedCDKZc8Ox4o6yLiW9u/5HaIsXcIb/2+fFb89hcV3TvmOKtZnlC/h9RgoDUJLez6Nw4ifpAD
lrXHyOjVds9SnS52a585UPVNa+eBt5dgGXX4Vurbo9shrw0oCBRr9Mmi4QD1LJgH32pqaotEAOHa
FjKT/BX6ntkQLP0lYk5uo+1UfzMryEEV6IKszkuPUA/Z2MrGMUilRdKP6GMMKw/XuzfPhChBQacQ
vy+rH+fS8tsT5Gcp4uovpuzkfw0o2OL/VVImjDK+yYTD/LKvXLhgIOiNStMquTGyu0dblbrHT+Ca
3cMUdVSezrF/g7aRxApo1sbsdTt6R++UDv5ymoDK7XR+M6vvgHybC8enBuailJ1ZQqb2xA8ijvmZ
3kZ4/rWAJQVAGXyIfoNT/3/9Rhf0RcIDBDW8/OZ7aGn63CyABzR45UNjnLd5c9xMckEx+s+dczVp
uRdKHoP8F2/wZB8eqoQ4goKN3YMSEJBOuSfF/VUHf37290X3SYltT+0mUgNzqqr+3NZ6k6FT1Zf+
tcUnUZUo8Pt4l08y2Z7HfO65rfcE8iABmVSkP4mNL4xqOMZxjt91oIHfE0DbYvIJvNckX8u5SnU7
Ya4r14xgjl9abrCN3jYM2Z8A/00HG6BwbZ22pe6moJP89Y0D2mJBCe2dSEH1vTG/jNEFWxCEXJBZ
zX6Vi9MxYIHeZFV1TB6gccrBtoV1txkdFZaO8Zb9jnYN/Zvo+MUF1MgQNklU3sV+suELlbQWpPD3
dELtCo3ZktBL1w8D6mDu3CEGR+0Owd4crQc48YMq1ReChhcwPOzY34j1dtY01ZdY9UzQR9yALD7M
HRCs6Hi+/k4NQSdhAm5tqcr124HnratcIvzcRJBCjkceT+69GUm4CCjoP75EekqYSrouGf+gU+If
Uj8/X/dvELDqQMmL3g3tf0ahOGHYLEzsqP29mnggm4kah+qHawBXMmPw4gu7UC7mrAtS0qeR7xT5
XMigqUpGvjSZQkTTt4Ht9sxNKPLz7UjfAOJbNcDwV3oBwHGlIbsPWpuTLjtyabW5bcyEG1OK5oob
CORqM7HpWv8ZrVqSKhjEAnpoIN9RSTOnT8icHEwOz0jCpTnynAOiy7xF2Pb5zqHQ+aO/6KKYeUK9
7WJQfiF/Mjv88TpojupKy/I8t/OeZR9L8Kh4qp4AtAFYWKomp367jBRJoNIoGdVl5wDmjEaWQYZ/
2IZF76+rUkLVgdm8LQEXBOimUoJSHGJ59+fFNkdsnA5ckQHCTmIkSrcpMKj1xvf5hMEao66+L8U+
HqCwSww7gO/1nF9NHHhs3a6sXMd3gKKNJr5m7mTcQOenTD44X2yKZe7rsItPOzW5C4ZCJ/O0+lC2
OK5k4DRi9S8qDKoK36EGGDtcD4mX2rNQ8Wo1vFRXNEml4OFhKcPj/UfX8wiMZISRpGSUeqr+uSmg
0b8yv4UKFuZPonFv/y41fOf7qQvM+FDYN5DuLFYKvZU4NBicRlUtj3FA5lG9tWBUzt9ZpsS4FPcO
BomZio+JXMUalt06dufLLYTObjhDKzVOEYlvOICW0Em3GitFWeEH+r3nE39Y8F+BkAmeEuE8amr7
mB75VB85nVBHPZoS9P5MxqKLg1giaKGv7wc6yJq/oO1sNdRFmKT9bof0ynMls4s6xKNOuObr9Ph8
0AOWjOpXpAvp/uGY/UXAY5SztxIETSQc3HXaE/y2+XeBhp8fb9Wi4qgk2xIbb5+AaKlyNML0oOMi
VGxs3WjyQ6GEn+Gb6mSs+G3tx/on7E/JzI/BmzbHYCltzJ9fGO3sZx77NzkOi/ziJVPMt+K6qIhj
Ty+d+MoT3jmIfjzjEfRBCtqzPLiANp+0IjJ7mcSgwC5WdAsu/VK3CZW8vP8p0AKVXPA+sAznvRrt
sRyug4l+DuBaD+2CilSFdsJdLLHj0tydOtj7mgaXgbHKuXiTOY1cSIdWmDRqOrW5x/BL6PNONbiX
D9aKEz8ZUMluV0gxX1wCJ/500z0SxrAcXoJBbvCdUfKx3oKo3miaMSJhI2Khi+daOa7N/CI8D9b1
zRpHKuSgZg0dAKt0J1SQPPFi5WUQWCYoZJaPIjyJMG+CSkznXEheQd7UhBhb+YKdMo7ME+XAsm4l
Qj5cccm0H3R1f+CbCxFXKYfC32YRRX287U2Rbe7hUqimGhVLnnWHdrQxKQAyy454UbxANhRmcjYi
zNvIePpFbk8+0I3PR05uKSIzJR+9PYqRXR8ZLDCOWItp/rMCRFxHZ48E9tji9OnFuJRDm4X5TM+o
JJCjZIdzzg3RBpJhaakemYN24GjuRcTZba1khTHV/AI/UtHatYo0OAV3ZZfmE0BNIIA3VfLZP8No
y8BSBfXLTgZ646DLkzwphFKRHb40Gc9emquvO54OEhLN+GOvQcWikF5SOBatvF9wkPE4KobZ2vXz
mNwDK2rQIMHJ2emJpm2GU1euv821RJ4FDmrGoxwRtRThZcg5QwY66aol8UZvToQdkimD0v3u7OT3
K75PzzV2wGGQcoDRIhqiNBeWrj2tHrFW9NdDEVd7KqcyVcy1kiF+ZjNnmhbhkJZXKIejRrVTD4cq
P9VG1BqkNNlyPS8X+pMsBMDobQGcnD1ZSpJc/gIT0Xp7CjzNWpovnc89rKOypbUoNjixmldbgwL1
BK/CoXTppQUHSUIArfDD0hrAwFGsv8tIJ1M6FeeOwDpvABZmh+36mcGJc3yQhO0fapDCE6OuNUD3
7wuwMrO9o5jyoohAL84+DPzRA8ts2xd/QP/ZYWnmTwQ15UrznApVZsN0V+VGkkwphGgfUcwJVVFH
MpXT7NsS+pMBbSjZODMAZZ4CCsvhr1dEdFODwfk4aE1bW2GkwFKevV8zPoEKQL6u+J48fDcSjly8
AACVpB0enY/rJMq1Kc5P5Z7fnToMHEfJi9EqoBuhPVLFVGobQKCv1AjSJvARZepBLGows4wJ657W
hjUpXgTzurLHdtaBnZN3IYv1WuBTyooQop7NKcOVluZZJBNPuUo2/zAgaOiERHV03GX9gCJalgV3
++/ChnfrGQMYTk59XxmWdgijLUwSEPz+l6KG6EHhRtls3FvJs/4XBwlpnQ/cbUytTaWPpR/DXTPQ
PDJKg8K9+NaHL38o1n0n+M3sJnLfAFIGB+ITSPP1y6jJmzQLl+4hB641K0X9BJe98cunDU8SMYYe
nPV+qIjNTN8HD9UQf5uU9ttafN5x36T80UcH5E6ANvcVZzesOayY+9GzPqr6JfmS+mzNN3+oZ2iZ
lGogu+EF8DJz2f9h8JFH2mX/nl8xI2r6sKY/3FUbzLyiQ52aKAj2h68S88rABduRC1KZ2FZ40ugI
EMBmNtgqWk5B1TZorQYllSD1bX45Z5qGu5gdxH9wI/IEWVC/0ndhV2jFsYln10unk5CnBxGEf2iH
1qpI8BWXLwT0NjItcVR6Pc7Ae8bqc0nhy7FtFUeiXZqzc9fzBPxV90hoGgcw5zcxgojxJ8SLw4c1
VExVTep99IM81GDseZ3ftdgwesIXQwFdQ154XxfNwv2UIYnsrdDBhPmCrjUJF8h5BbSE6/fm0hqp
a3Ej9OXz/g46/bHVNqpn7VBCeZ12v3xQi6Zx2l7KwLv0Vs6ZCtQYETW2XVmQh2ulPJV0Qt2pQ9zv
ONrZx2jMAvCiH5QBisOp/XFA04b+JGuejbVp/QEXko1vaTIHiI/fnQSBiLe736I0WO7uy9xHacW3
vSkF+2J65AF4hoGMRe/HmH+8r1VvPWHzN614ah3p0Oe7hcG4e6B7G34xvnIdcq6/D7O2T03XK/1N
Yn+4HK+tDsP4Xk7iWWWuvLQiSCMHt5L42DwCQqbLW4LvVpEwSE9J3WpdJOgOSFIPb8qfWWS3N539
pLjfMNargU2uqHbUf1aQac9ugdoFLjNKB1w2PKp7pk9oXT6XcvPOYgdT762oUOrBitW2IGDph43i
ptXreV/aW/YdjfEaSNLKNEyOgIoHpC7Z8gli/0g0m67FKj9rPfJVvoRgl0M9sKuGv+mw8v59RiWE
lMkoA38gCfbCwTxi3SXKmnDqe9ixcr76r+y7rQcW8is58p6Jz4j+qfoL1WCkg0jbSW2yVyOYJYCw
gwY8hJ6ewEFtial1mZgtV/jjwJlknUf4QWh88FOEz/cWNM8eGzhLmAqAgrYUiMpDNn+eovFF6SUA
piiowJxoPGekXPKxB9RCJcQYVEDVv9D/FlHnFsUIxKR5rPn2Tu6tiQzbSIfuRT2PVwvcINM7KL51
6e4pzJktn+8fn2HdospNzyBybIX2QuqkqzgI64DoQh9QQi08iXKFxzbht9E1pFnXYlGxniIZ6cDY
x8o59ZV5edDTe+Z9zRP4vJInioQ5CzOhNBjBLXcHgKxTqYTdagOO0WMCV1pDQ8aG/GY45m7liKrV
U3WSH0XE4xsbraXBcNO5/mxJFOP67UOHKvXA3W6D7XdtJEklO4x8A3rKAshb1hvI8ySvKQ0HOnKN
qOX6jQfRJiLwXlfSZg2P0mDBLU2UlG4zrj1LXnpvKB0/47gpwxEji/SeJf2LZ7jN8kwUpLYvfHjm
pkGqg3aJcq8K5bVYwURRD4zHUO00ejdCpMk9BQSyEIMxyi5aRznM4Gy27Iz8KSIAQEXRtI4COr/y
X4ey+F9Cw+an122BqMV/qcp9OPW0CLhm621+6CThVx/7CkK9eII6wLcpm3XMu0nakS/hIuF2nYS8
qGDH2n9meTK1RKAi03FtYUrfoyjziQVMxMdmTeMwl4BYz8SJK112D6S1DYQyKeRrEuW7FGpOcjKN
y+oYjPVBZ/IvBsDsSWo5P3W7vldUTpWHgG1pSfsbJxXIeVVI6NG/kuoFsJNUwh5t7NUttn03KXke
taFaNSZkjbkUfhb2yraw4rrDzMGgI0nzfix+24t8qLituBDDqImegW8ucLK8UC/n1PGBu9qA4jD2
tNnWA/Gk3qS2b1gR2paq4rKfKLe04l0KUDwN/q0BCvQk9171fz8lsSSwZiBkvxsRX/9nZBzenkEZ
m/LDe4K6lxL6Ua3kyuwnlKnHF55HRxdGbYASu14pXHaqiDnhNkwyUcUxB58BzU+xb0hA3mSYO7yT
FUS/UbTI4tohlIEzzIF1NHWRj/aXO/RlmVQpLxhLKYoenG2eXkeJA6URMEpiQHcD4x8wdH2JOGer
rTcqGn01DDCJX4fisjvClw0Z/Z8uwWSo8+Z/7P+ofW7redVa9oMczc1TQgUorZqZea7L5K3oOgdc
VHHXbn1syu6Z0vO2QS506FwE8lDMi1Rn2lE3LrDH8n3C9yKeqs4eHQjRxkbvV9biv5gOAT5isvhI
fRj1D9dRTExt2oUsMPr9dh4ryAvSBTTiSOULbz2KYmTzZ9JF1PqOIZFga087mHZJ32/noxgacogJ
GucVK3IZSTcJC9FnPygxUyjwA2b3p9rrhuJU3HpYg2fDBi9Ai9mFz4iw4IKuuJCpSKOh+liyJ5lB
HnhsfFPcITPJZIMKzkqeVo9JoriocfxAgUE6z8pd0Dd13G94bogG+lUV6y48U65gCISMZEbn5dYb
QxjKD/lGU0/PyHq3FUerI0kOYPRWAqf7bmA14xvKcCFQPd8xIvvOFakuyp6JJ3DTyGzsTaW3+n2F
KdCJ8ORluwqPiCbAGQyWVZHQxtt3zpDkiRAWpo5krMTy24u+ubkfwlgxOKAlRLoU+FHvi6nYuvOV
U4YFUOyApMTAf1x30DLVyEskPN4fJaI8XlignzdPBvvZkz9CuVQ2EBf2XESyGA4YZizwUz1Ufe44
oExP4OJL8ppMUXaajXAV6JzzVbfGh28yy0QPdkIQOqJzjnTTDVfP3Dak2lkCYiAZlHABu1FAldX4
TD4GLoNyhJ8qWTmZ6r3vx6zfGjoPVNWvM3b13JUy/+cMotWnHuliJuUtgYhgoCqpMkFXc0LV8RNZ
BbPV/zDeSdyFIufvzhBJpbdZjN2pwd5DMTN5ooKoTsxSCmhPoAZvpntcf3vHmInZbH+lO0eCGTlg
IG2RL6rCquB8Kj12o5eUMTUg95QUkd2OS6cm4AgtsAtkvykm/PCHQETmarpXlBQ6WkdOv3RsL98t
qgtMQw6AovN4g2U1HL3s+H4jr5IZASEA8suz2mge+L2OM+jxWwhlBgaNg9rFocFwIp4k1+ldRkpr
cef1Z0AduZvAyPiJhM1gOP2fmoE4j31kvsiQ1ePjQWALHV2pImM2OZnOvJHsu/kLwx20T1exVSgQ
V2LQca1IXFcBW/rcq58zLOQf0zAbIJjE9iGLELX9D/jawjJNvhr2LziG/rg0nf6RHN3WHPneTGK/
etWbhLtCF/fvY1OU9K6R/kqzTz3geHbpyb2uGAEBIV7mAKev1JyfRM6zL2ZEdnW0v6PdL4//PkI2
KEWAhSH8q2+tFb6F4ndKxkf0wcJq4vInq2Qy11RcohwrePFk2k3vjd3aiBEGBZ1a+RtHpV/1vnkx
goQ5Y3Moh7X+rLJmDc7ZxJB1H44+5XOoBye1Vp26qquMwPSP8DDnWAK1jQirUVBGIrszKP4zfSaH
2y0w31A/O6rIaOzVUiIgTlF6Ux5uNp5Y/ceDikbG2VS/uOQonHdhWe/M2ETj+B9tzelv5M/H85YT
UO64nOdAqRJtRGk8wZAOkMAL/CDTxbCRdcdaUPrNDsHm2Ry04ejzz/D2euWVnGW756WidgraEfwh
irnlFQHL72i5koUtbmoa+Po1nkYPm3zfOaPXcWfD8b1Iby3M9KZ1FXVuxfZiSQe980I1xQFpcgH9
BHRzTkLQKjikmXeF9nzcdpFMzK798mcYpE/mbS9bIxl4eviqel/KMXi7QkvgUsrAMtWB79hR8UqC
8pHNJiNZobM5Oj/S60Bu6na9XyE9TezQdGN9cqqwX2LRatLtW5ZHHzAlrlZCB/aKC4pOr5R+wzhw
10+ht0kHBR1HAqr8eC2tpLkBtJJZZ+m3GX8Ji9iH7EdyYuwDqCOjlkgJIAL4LSo6g9DewEx2EW1L
TDzesm9WjUMXPcwLKgs4rYYD6zYr2c76I2dNx8ekegTFD/cJVEk2crY7EIeZhucMILeRG6ttw/Pj
wHwBadKFBuGKRayM/8F4lmctXQpUXodyN1EVkkvbEqYr/iOcP96Ggu5fCY1xwoASlwbmigrytJV0
ec6uPTjXgF4jCCF0P2jvvlUSwh+upFP5cgBRMUBSmLXFRQ9o148udKoQYL+YnBnV5MYl/QU0Lq0c
5V814PKHxCP+PjPtvSZK3LQ5vqnkZke1mJBswZ00i3U/+r5BCULom/fSjpp9q+XA6CH9gvidwg4V
raYZVBlf/n/4Ros1HDlnzjfHJOdAnaQaAjnVMr/Ugqciic1sc862Oz9R0LjO2sUEgaZX/CF8laNu
sdUR8ci8P2FjECVdUWXcJ0HAllpJgRgqHxvU/uFefbmgE/MlqPT16ADoIHGbx71iiiK++V5EgQi2
IN1CfshkW1rWQHSAsmhf7tgFMfE96RYcRwwtbQumk9oDSYc7QvC+kyuDSuMyU9mwm6iISy0gIZlm
Rl2JN+XamrAl+Ns6UU6xqhSID7/C/g2h8gjIqSVTS/2uHuLSJn5HNv9wrkE1sguaqVTxFVJkC84r
e7alV8VdZmOpn7qmV7zouCvmB05YhN5VW5/RptDE4to+vj72vZbv2RsfXI+FEvkXooXmhCLNgrat
exViDtTXABi6MMTk91lmFfkzY7Qbk6HAoCgbtdYxz2EwV8Apkwi+7MUrH2pnHuZO1Brm9plL5kYT
XfWPhJd1o4Lcr96VRmOWfr4btBOuiRLv+secYA2Q1AH5S8knSL61AEcJPRf8dVj+H/AydiJ8l0Ln
0KSDfhjp+Wp+Mu3FR5FHqrkP9OvDf5VtbNjikttliGyIMJCAoJSi71z7+KRxn7U0Tz+w2KOhpnRf
4XVjP4heiou6IT8DwZQDjXD3rWPdodceNGa4ciTOdFjb7d1WvcpCx8vHkX6bQq5/t8oAIGZUZKSd
/1jjqzvqtWbVTp9X7LdIYZUJXmnioZXMLjVepJg5pIVXSpDR13wnFKHvuzFAZD3v9iLxWyOo4GFq
ynDqC6hnY99phx7GLs8zlqZSd46QNuo7qnvtHm5v3rD/Fx0XEECPIFEmoQGTyyibSzfP5gOfBBrr
+AUl34izp+2ZtE4Oo4eBJ9OLjZEZbpraKS2my57Ff04sDVc6REh6SQVNAKr29B4F5tP3/Ytxp71N
+Y+Jc2nW98PLIwc8dpDR1ZfF+FxVGmOeyLFBMzDSjnc3tV0QhBAKONJ3TX+S1JRvq6qgS66xugtW
iXk2QPyQCL/duThTyHaE2ITzFxw33lxdxD+zcEwuZLHMjan5h68404I1SFgPxsdKbVKFBCM4fHZT
P+lQj1nZZPqOge6H11LIsXoyfl/oBu+OpVPVciMcfBZxuwYVxQ2KPz9RRWIJ48etkO/MvUCivruu
ZkABlxZVAqlCUJP/XA7f7391cueL+4BZMHvveMckW3XU5l85r27qoaQLz4jKtf8Z3n1yDLW1CXrN
EPB9nHudElZ5Yt4EDpxdFfL9T1OzPEzCQEAOvX4zRdEFTf7RdIQbbQeASDq7SAGJFyyajlwaQi7W
fIkJG/ogm7zMQbTrx7w1dZxQo0qbBIdmP9d3GwKLeXfYQxBN02+N800jWbePJvtv9vpWN06y4n60
Vx5i5nHF6mLkHZH02mx5S6t+gIwOAtDTZpFz3hfgy6iPTOQ4O8QM5WvFOJnEMq30svjSuDz5NIN6
lssuHa3JBaIgOAfL1o/nowPkC2PQSBxm7Mavfgn63dIHUMFUBxmAT5o8CBeBQ7bUz849iEaKJlOs
OAPjODLdO4czgJ4Fc43dMQ8Eluuwv5Hgq8HgxkIpxAh5nxnlXoRJn7jxYZtMx9JQdWY2H/bHqO2O
b+RhjLztBCRQYhjMNv4iwhVVoQdDEA2sqeAEYADHFVliIAWY+wlyVb6TW6tNeqbHDtXekYVQXpNH
MaBySV34QUVdyvBIZdkKJiCYax2qon4ZTcWJ00KgC7EfLeqeaLsEDup3mxk9wkW+0oxZF0yPIRQU
fTccpez69ulmv2mNNhR9yliTno7d6edRzgSk6R2mnGRoIRU21LBlD0yj/CORUuetYMSJD2VfSHit
88QvhhVkoWjiEYwr+V77STo+BvejHPiz2Nty8+EO8ZVtK/wdj5gIB2HkyLDw15mi4cIi9MFX936+
jiRILSisk67TLSFTZdGMckIAYuAtlcEF4W+HEwD24K+6u2gkUAZ2PB0zT3Ufewu/Wk0I6pQU7Mj3
qe6TpY1eA4nvCePnRWJbJ56ecd1UwHTq4lW+QePFJ7NkjuGGJIfM2qMPl3owF3voJOVIqG7vr1mT
ME1/qE2d6DqBoZHFQiW0IGZEvbPx8IAKVH7cySRNtgSQ1VAZjMq+KOx/K8sBJtJ2hqN7/mcVJYnz
elLe1LbgAXy0LxgDbpYAYIPCke+jIdm+EuFh63dl54TQDJnilItsUxYMwQYbQ79j0cnlYXeBG06c
ABd9pyt4URKBm8cpcUqYmbx2MFcwMbqv/Lv+vlJUEWW9MvTZ3KCiTLjMp6NHWqNdQx0wxZ1SJ4Vk
WOE7L2B53yXQYHt7ZvKcRm5tHYaSkaid2Glh3lXuEUv8vYn2akK67wD9sm4w80hkZyNvXTQNOdfk
xfb6ftRnMnpzkH5nNvCy2nFiWuQtEt9NswiUl9INMkBwMkWvzhfhP++GYAPfP/iBg1GE6oaraQYI
Kpy7DkrWUaNUa9GJbep0u22TegNM7R/Yw/Qjc/GcjogYNigdFQBFv16elEuSmqHpYZ/T5+EQl5z1
gOf6igxl2NkoZQ8fPKQFytgf6g2xjNagCK533NYLRlZNIUI9aJv3ITRCVPaI3OOO5wouwPgq2oha
EZMtTp8Vl2B/813GGGsm4lLGWkFykfuSe678w+KjsiSnFyiyZK1AZJ042s19Thka89D0tluvV97V
+ikzpBoZeIIKskkQXb7N8kl1X9Nlzcr2JcPhkGxBY5/9fA+avJwHDCNPG/A4RT8bsBVOkPeDnf3W
my+LO9b7et4jFo7bl88smntolVyF2HpCoxf986O5RTVVi3Z0kdXUOfOProUKg5a/gRaTeWH1R4rP
macSLOX0kV8M2yj65fl7oMcMdLXf3HyXPnf16Jf7K7e9RKXsmM0b8qcsxUlQ72sv0lll1aQAIIZS
cjQ9nfPV8VJWMuvPHs8j+n0HQBAFLgmHusYdCnbrBhjzU6gPs3kKlzBS1QNWgTRTkkHrdUFQPXcd
UIHDJpPR86WxPA5aaFK7bwdM90sHKExK2PKFZabzToMUUzX/CUO61rKWElkfFYIbn1LgcCO8O69z
hO9xsN4zIFom1iBW1qyqydwxh3msm/pr3uQHhbHeRJ/nvW06D6sRNhhwItdB7cn9HHazmHZ39uWe
d+xT/scf7srlbPWgJkxcU2jpUb1ehVxjWQhEAm+6FPswaXRdDllscVppirrE0szKRmwMDyso873J
nMqEIaRDz7bWiQcZm78O4WuULfksJnVxe2NIClJVP8ng4RA3GYAdRvvIZgFu9BhyLwyOikuRhbhm
+oywigRPD1uCS+6bSh9bjOeRoEGGQOXfAZD29QvNS59z3lhW+0yL11ZMDmhgU398FmA/p2Yv8ONe
Z26djf0q6xChcMkxzcKfgm52rMvFgAfVh7UTa8Ov/slWwVUdwhuDTuJlxxc+Muq3kVn1/4QghgvS
2g4fhpIbcpK1gZF8CDl7lCRu3xCTqaJVyDP8T2XIrGFRv8QVTFEpLHtMjze3NPZMRfHSpDzSLagI
zKDHlGJvDYuFw1gXaTZj9XnZat3X1QEok+OOHS7ox1bcNuwpN34Ez+KGrB23zFy/96oE8kpnamgW
RxMEdLL4Gh+r8LqV7fi7ZPHO4+I/iR1SxbDTw8vLka5DpCBKs/EXCKIO5KwbpBox8UAUgpo9kfIQ
j+Hw21Lh+MXkuNr1aPbYG7TgQjfHAbXCBLVyaMmvMK+sVUdiSLj4lGbc7KtrnFZ+ZCPVdxZG5W9f
++rD2EqQewa7Jf0kkz14Zhbkjqf0RyoemUdMG2R7onEV1uoE0Lktt3Z1Mx4kz4lECzBROimPDHHN
s60WUE4ktN4GBZGPCgpmWW35GoO2WD1kYU4Swa9Z2J3ZToblWselbB6yQhnIP9yXO5+UgRmcLWfg
HPF4j4/Wge8VOUeOJvv4ihSpkOJSgbFN299PJnQk75a2vo1ds18ioqaREqg077OQr6P2ubVtyz07
VBRqXJlVj+sJaaPJExtwFbFlpXYcafBzRyFeRWYS/gXm3Bv8gTtzuXk/z4w3LCLhXZR8g34qsmtN
mTGNvTUiB8/i1ieet1Dovi7mItRlZrZLzom0idUTrIW2Pd1vtqVhSdEvgcrfVkD2LoK5ytf1tvi8
iT0zSdL/USO4usf/JeXb2sR9PszIiqf0XWdIqOBkQAedeqJ+5D+f0oWQDeZj0GK99K+dYRJRYCtR
yCOLFTJa5iLtT1n4U2LDzDptmL4ToyvrJxxrXRiqyx/NznVbTh1VCBE2H2zcNOaoBOYUpQ0cxpCq
n6x/Y1L/FLHsAi2tytAAROnZQK3UTOLS7pi98GhyYIwkLn1PSNYUw2d7Vf8SA3tXG6Bdj/XnyaHV
a1R75RmNbNSRrMw/auZ9SH4F6m7WgAf9cCPdAkGMiAZ9qUx06ub17ARC7+AsSgLnmMNFvLYelRyA
9By1SpIhgOSk+ycctM9r+mMATjlNUZfzx1QOcOxuXK9n7wm3Mtms6tstHJFBIwt3T5LRwt/xTBk3
i+O+PnuoZ2GRXl9kwZgnSiRX+P0Xb7OVGABLhYytNbuJdEV3nhtMblhy59QrofMvDBnhO08EJqA1
xHFd2FmAAto+5AichnMd9D9HexyPvvO66SY5Kpaql5IMZ/jXCPnQeSK29evWJn/j+CGtlw4VwEpd
C/qMhxKL3svPK1sd+G8J0ujtgeIAhXhcAtrwIjcTBsFpDGogE8GW2if/xWoGIjJ3R8MHVapx7kZN
fAJwfJDdLp6+c+CQS5sk9/4vSKY69yo/UqTAQ6xrzdoqU6ZIzeU8hvRbrENB3cZFydHJk+ylZYgZ
uYIKL/sADCBfF6jdFvDrgrP8DGMPZcxqD2xz1ooMqS54ZOEysvoYEgwGefI0r4FkpMpckEcraCof
NN5ldSuqXt17f9EzhSUieizIdLAsLncKqNUqYv3V1sBgnCQeFLSfa1aXrx/J5PBJKEhzNMfzUO34
+Wia4XLKvFD4gjS4F7qY/OUKK5duNu6+gzvQwqXbntQBZZl6OzodhZcpJaDrgxK53qV9FuRDzP56
dooFE2pw+UURRHYKLG6awDuME6Q7A5zmJ8TxelSTCXRfpjGwI2MheQYNnYKGFfv3gZXirDrYJOg1
KuuLbyY+8IyHcQzSeDg4cq4bWPlZFjm33/l6GFe6bTc2LvjlbpXpcp9U6J3MAXSpOx80fhUTNMe2
r7CaWYxxPZdK+A3wAYL/ixLoUcC8fkHvNHXnooyMeFHsmOyARGyFmJ0AogFeHu+u/yokm1H6Up8i
P0FHCoWY0zFIjRCyksZ5SIDxDCtiGUCZMNFrLg7OC5A8ZPwWbDRBbFvOGzjrvjZueVK5psCo2+s6
VJaQRaHFqKFdzXPVI+3LuSws9c5fF8INu4/x74T0DlaZRgdtL3dkmY+fK0W5Xh3Y4OqRuAKDLYFf
r9pLnatRrFVg551pphdu1GI70ae4ybR7XgzJYm9XQtNiStwqz6hTTRrMgXHO4/MmUwF1dArxi6gS
nz69PSJ1HW3np9gk+Q6NWcnV7pR/c6a+1W8d2LUUWrZOWhPLhdYczOYwC+f3OPPWp3Dyov3ywjPb
vliYv0j1nZxi1cERfEyhZzK83wpynqFs/EZlpJKjD1HU/HOYnYVztfgsISrEckIleN6lBVkjWxgm
9luhdwWZ3q4qR9GECLBuDT2Cn3wkaAWWnfblGIA/fOgelTlideU84gNAmwoDag/s9aacvz9AOFbS
CzIKjSvZkpmI0FTKBHHCxLQ+gYkyAIUzZ3YKZ8COuqd6bF8BI4YaB8ojuoTQNO2FOHCnDLT0InVr
ehJrY9XLR16kb5xm6RT/LIfjsNwxOyr8UXfBdS+Voun5si26xGT7uVKvr/pqz7skXCbbZ6OF0RUH
dF4Jo47safavn6Ni6Db/Jr0bzE6gFOzbRnjiBHqSgPmAwocJsi/C4pI1xWVIbMOAVOBz0/9/ccxq
tEUl4/2eTYrHR/RzPfXKK5DxCT3m9usbTrNFMtX+Sm69Xm3BjH8wFISxCaoDRs7BH/R2z4RegYeu
7bpmTWE0lKbDp/oWtgQ6xhLazaVXf8H4edt0rxrOg1BbGWnZ3wWcH84A0DHdZwj7R5oLNCL8m0SV
sS+IcICvPCldI6r9yJdDxen9jchplaVJWW5ao0+D6lhU+oFTuG+teD8PdAHDvIGRmMouHohnnFcm
47FRGS84oinmcrMyVATmLiNDpiuVYZphLouPpHNC9Qquu/2aihZ6hO5aEhhH2hygApk9bbUTHlsF
3QQ9f3Pk5l0vUeIHPyMPVWTSMAwl+s/6613aUM6+6vyS4CVUzFFxXwcwLP+UsP0MgeNUGviHvJce
bkgC729apZhQ/xNsrq1yqx84UfjlGmuGgjyR9Ay8rUlyUbTLOUDcUPf+QTvtOl3Xk/2gb3MiSK0D
wRu/b5D/mxVxJI/iIXPTgBvbjNn3vYZQ5xMK1ceGfyuUusczme7InR6+JMQqG96TTrPd5qSi2T2B
k9Im7o9+3vaE51e+guEWEriXlrhvOaxRAWp4fq7mn1X4Dw1lPmjN5+yD2J+bslah8hEFjRB2Es2B
HwvsY1n4WR+dgzEa0EknLQ+mpO7cFfy6hrn7z7sc++RD/shpms/xSWOXFHYq33JOf+v/jutR3RIm
CJhbdB3u6aSGtUb8SQc/Aj3NBBM5BslL0kHX1Ozj6qUIiON6UqRygF2RmgVNFNF2GvjgG62qJtAE
OMeUxse+KymJqh4g9utyjfyC9YdE2DBWveczdq4DlaE+tdjF+VWGVo5xyLQlwI+XNRY0x7Ks994E
EbwHBOc3kSuvrfTNLtTdlkXqrYdJghCONGi8luK6ggUB32s7QQIagrTFNV9XXpvJLXEubZFP8LrA
HSGPkQJvAZ+OnWCuZSU9qV/EO++mEI0fU6LDlyXZuiAb4t4Xs5EKYQcKcYP9I/LbZYlU7AMPiNFU
hwWN1e/JjZcci/Y34S1xBqm/FbVVJYYNFA2J98brjwhpD7zly5eL33qRLlbbF/Z2q/3iK7TSjmKI
5j22u860m7nhj9n4oM+ukuwJoBKFTUY5u6diJd4dv9Inqvf0l1MJpnfyehPHL6JkTZzSGiGdwJCI
wNnIJtV9DBhMDhluSj8ay4AD+KnoQRENPKWTKW4RfxMUpH92PDPVz4a9JeO2vhPt5ASvJLWUFNwo
taXXY+AP0ifJGs7Xk6fDqPEoM9dUfIKTC49A+dzCSZWhbMeuVbv4Afp1Zqyd8ZRg+Zn9NMXpOkrK
hg1GAHdsWVbJ5qWL6z32CquPowQUjhxBUQOmotNv4mXVYc5vIzeiqoNC94LetairtpMWfIAgAks4
woh3Zx2OmmbVuQ2Ri47C2Y7ohfK1TPKstbK6iaUmlMVSoapgW7smyGdOLWAb5KVIr4qDg3VyM0Og
dhWRdSYNgYAGTxF2ABbN7BXgktB46gF13J27wXhxI6/XvOHc2zBNKc9dxl3Eq7W4loWFltZY/7MG
MtAnzaz/w7tIWo1LyHLCpzNypeHK4hSA/O2hknkcNYeBN3ZbxT7XZGhnyiRJszIDYoVv4MqzKMsE
i5KooM2/j5o7pVho/Jn23T7Q7Zcy1CQVvK1HLABG1ozPgjwme079IemLgTSzE2FWiGX3bUfvcf6s
dfzap0JppNZn2qLXFa1ORUjHqQ7uTBvZSv3BXCyeN9QQh0/V6hiyand7moHe5zI1qQ45P9UNvn0U
aCsyFYhe3LkRvk8UBWcoVKGlSsxCKfq2g5DfMfzRU2lidZFaiUNH7tvQhmCNclfpVvjc6io23x+W
X8BYxZdnACeU2dyjkieYHPUezcPIQxsjMvBEsynVDIPDd4IVSi6JpgVermyUK5XIGOu2Eh4Za1xR
fcLMf9aq8pPlTwm8rkyq9bw7RXC9NTfU9TG62F8AzvVmTu724waZlssYy5Tixa9jG65MfQQA0UDl
A6fHwzGB/qsV/gwVBGwL61OzmZBhKwAZTT+TiUiq0K1lmUBuXCV4yFN5CjnMZka6wJVea6eeqNZP
KqFQOvyIRagKp0BuZF1Rkn77w0I/E0u02hwZtX9IocNDJ2GDz5KECcgodd2MuL0/C8P2d8wwV7GS
CEMNZyDHoIZF4FS5lHMyTYxkCNcpOy4gtjxXR8rzN6NNLdjznK23TucGcuHeeSPCnDc/ambjKgum
aEr3FjUYijDGOn8HJIlF9pJdPPvEwj7NC41EnfKiA59RVXr5OrSIKJritKrJO3gUMHOZgnKC2Xlc
XAyRCpU9RxoKWReHQJujh20QANQe7NWDfWz9Ufvr0up0TfxeJZtUUpceBlyIW2uX3Qht5PzxEfGr
CIQ/wR5l9KjIVDsuUL83vuNwJY2YKgIoGrtAjRXtDwa/zAzNRm7yslDlhcYM+PeEhV4+Rsf8sc65
0/9qzh8RXImroGKOi/Orr9a6fTQQ6hUxvBQHQogFpcQ7Jh3C+oyoq1U0eMc5wtfSgRMtl85aaWNB
a2g/NyXpit6fn/mS5GujUUqeYC8KC8k2TSMXJsQu1rha+jeD0tz3OJkfkQ4ypp3WeEAzlyHOyWCV
Jki++TsuQADcK3AT/Q9O59qc74JM9vohIikbBiVduGo5KiOB2v6uEogRjryAKMo03PKsLrbtxWD+
B3ftDoyO0pSf6l4IWnY6xs8b1251IyKfIJzxXKuOWUIsbxLDQPY7p8DYq1ADdlOhb7Wx+Mf10dQ+
YwkMKpCG9U6dDFk43V3PMYQ0u58bBuRUlIMUMsMGG/RR2Q4KYiXpFm8VObHGk63W04x/OESGD7Aa
Hr5OqcV8OgYFIzKmQbAQtAMfldfIWCqCmulpeoyzFMjo0C/aSK2uSY8WK+tDCtFHoHma3PwxmHVh
xKOWPP9uq+j4JdIIKtQolKa5DHX2ArBwRVV1Q2n1qah5gooSTUnWWGzD9v0/scAk4jwnVs19a9kF
z5rAuGqJqbQu5jwvapMRpw+Nug6KlqD+VDVdH9MIRkH2t/78aE6wqs42aASOyO8J3xA90Y2N7nty
PRisQDXM5Yy4/BuomCuJ7YfQcE6T9Y6wFJ/g/jW9pw2oXuqc7DoUR4ZKWwX9Qg2BmKkDO0ePht6h
eJIHqr4Th6Pu1lJRQwFTR55h05uQaXgYBF7irwQc74sT/gjtLqcI80ubqtsT0HihRVQ0w276RRRa
eELPMyz/fZk/w2g0Ac0XW3k438k0+W3WPzyTl/Akztp0TkYUBrXlpWLYXUm/wqhEHprMFnb6XRXo
BbothEapM2HT+J8v4EV1pO45t13SmvNiGWPEPZoU5XVxV8MvTNc4fQ7bfgf+gRrKswhqxj95Ahws
ar+43fnXJh9UiLpw5MuZL26BWYmkZ+j2naK/tqqrOQoQnEUe0TZSFcHXTkZcKdJqu4uNq+Y1YWLa
ti0yWuZEJj/QWWMUvhKCQSDf1InnLPsVg7ihSzigQ4GyWLschfKLMCDmQMwmHaQTahklhIAyBpt1
lckprI9nKWV4Z6nLFLbAtn7rfze5Q7AGsRhYQWZ4/4aJOZupSV4E+IQyu6fixflLZ4xGcQP0kM7J
XMU6Yl7I4Kd6TlUj3uMD7qcMdFT1Ouj2e7lABNJaH8baL6u+EuK608Ajy423FKjp3AXJzR3Hx185
GOHJzTn3cw0JTqs0I7XU7zlsVUkBsksNCwrmOQecNgJqfD4oIoJ2A4jrk9p9g2takzkmopY/RrTF
HssUDmJQRqtawI5uFBhEQ+7XmcoC412iOZGmQI20o9lKUxqBA+o5+/D3cbdXUM5SP1CEKcK7ob5H
ue8WfrbnfcQAPQgieIrizyelIk8ZVeoujTY7OneGIY5z7AY9AsZVW4kL/uvlWfBMxgdu+AsOIw48
WCGsWjh6OMsPSvBUA4Sc/7x6ANs09ah9kP8OihU1Z3HBK+xUXnWF56ix6mhgeDfwnxoNU6e+TbcY
fsOGB+VjJEMMs5Uedu7ZyDvrfCYkgAG40GZT84St9YacIg52RoI6AymWRtX7RmqTjeWawh1pp2E/
SMHOy/0ANw9m/yK1KH3xHW20ntaWU3lmhq6NUOfM2N3RCSG5rcX/Em49ezGJnyqrVNyTp5KvMbR0
xZ+P7v0f2gPLNRoL1ttG8XXh/kPdA6L8JdPG1FBXfExDYwARUIcvCchHx5ypePqEcDJ4ZiedlCiE
cLxkZ0Z6/RBKiL6IAGVDb2Oo4ysCWbxqv2xBG96AyB7O2CYI7tXQ/Tcr/5V+bpcvvEidGaS7Pgtc
kBxL1BLMKYorrr7/KlQ3WODf15VsPzjgEXekGukuyhjo/nIs52WzwcZUftgifL8uTRL0QAYpKyUu
rcooySvnclotQETN9J/GzQm+gWgqPp5AxoBR0oDzqnbH2MkbqORocN/hN4mhMvRnqnDnvtilHAC0
XKBo2w2j0CEu48bkEAqrutOQWclAZ21bsITq2EqrEJ9akFs2iQE+osAC0h6OdWTXtJbU+MqhClqe
nE7wKAm/vk4h2ooIcCFpEBs+QFbidrzIF/Y0VoihlGK/gEYFyi2LPGaSzH+snOep+iDq7eyfkIwX
zR/nKluinF3DTM5O9m0Pv+uuo7QfBT6IpLADfZM5dTHIMADgsjopFwNVZOWZSxsNjNXmAcHa2mjD
uZE2E8rY+T65kBXaSKWjlPBc+uHJ2Ca8mOT8oAIjaUXc9IGVLLWT/3IxvW9upu7CE/nMT7SrfMBW
sQ8WfF+kSnMLvNc2WrYnC4s4LpkaDP8kdPPF8UoCsisUO6i1ykz5PFZ5cUvEAqhJfWJBIZcXHIx5
HhAHHEqVELgt/Sp+Ow/6NW4eltdXPLtnHWvvurJlam3O3lGVVASkoKHXfo84o4Ov46n3dSQzcD54
Fwamzhl8T6o5H4W/poAJI8/EWl+O/QsKg7y7FJwHNbklGpWAmg35mcuOWKfbkDGjDXbELD00q3qN
+9ncWRwvTVARc0iaGuIp4Nf5pjYsOiU5qBwrBreP0WlWOhqPWvEcH0hSGXlqaIRMfybQWOZ9UOg8
KN6BX7L0BuTiWx3xRurh5mG9aLxh0Q5LcMdS4CwYE+kVb+/B0zVBDkOttRk0X0HL5gw/zY3TSx8T
5vnPMsydQvXgd/ocaXcFzbSTr0j+jeR1kL53FGux/YIdavG8iHqtmsI2DuRDEn+Lvq71M+tXza8v
EwAiItBtOqVG4aNtrk73FFtWa/oPJSY8K3Y69u83CryOUvHBKwa2iiHyaETQikgN/NSH/NauiNRB
Ho26gt0o2xrB1bEOKYvEZ0lJSBEfM9kJEtxPj1QmhzV8vvUz7SDOkv7D11BWaL+nQ5pz5Fbvf0f5
Uf1oub3GsCjAxZLkt4GcN4w7XI6zeDH7YDSnGZ/MmxsTQDGbah0DAJZmMCin3ylNo1Cg5tvdt3Vn
DQrFEoxQ9JJlutYxo9uzyzjw2IcwcfQSZTZroxacJrs4yyb0W8iulSvJ0jGQuDjmGbG15WLoz726
1ql4oFLjhrBvlMVL2jad4v+NUoREDZpHJNiTWhSHYcQucIWX0GBu2kU4BtfC8Wkg3+JY2RT9n3kW
1oq6+Vr4nS/Qfml8gwpt212JeDYh4HWPYhB16sw3VvGpTqzrQTVcnmxx4h/lzHimmXV0p0FX3mLU
pErs1W91G5Av/ugujVN6JoL+wWLVfgsBKN+vN4/zBgnDGE4r/vBTYQTFAdyIFeBuSRvnQjAcfxtu
pSTpFA6O7pDWbpNLVYMTV4D7oHpF1LF9lz3zEKum2TBIo/C+bRF3Y8RQRRSzJ+yYQe5AtT9NDuch
CTDbPtU1gqimnvUHi9WgLsQPnNobw807h50TcqRUnI2PPICFQuw5cqeNVaPy/jTXFOtJK4f0dqdF
yrt6m3fm8SvvTKznQaqzj79RaP01GAGZKfbHvdpq+0CkTNxaVmJKNvuR642iDIZojo9xPUhgdx5Z
QFao1/vdcVvqzJkbuvhncMVHaEClHs3vVwVdxLjtisPRPEl1N8kre9grfgG7xLUoKPQWz0oS8fTg
6RU1MtN1+AETyrmGawa0YOE5WCwHMnqRBFWS592xngU+LHLIYxrhWr6J6j6cg/0FfNCgSSmYsuXj
K7v6jmqK0Gx6RAfEB4h43Vp2DPME2/+lId+XU4/EhFizDNoIfOHXu+IiG0ObZ1SDFNzKvAhZe6c5
7PwJscwAdk5tSnX8NSOAJc5I7Pd6+0WmgSuxs5IuJYGqT6W1knI+mVsXlCe3D4bhpHIlEMVlxK+m
EcFyWw33rNBS0AVDFyxWII4PmpTdmYOjHs+RF6ScBY2qS3a984qM1iuCxR3HbErNkoVTHzial64G
fQR1huW6VBlONVLdz4Rm3dn1utKN/EP22OYEn+b3izfLk0i0DVSEiSC8mB6geFbuh2QFWVzetyJ8
E0Vvp8JZ6vPe3jhuxsFBXn9tGwFr+LFDJJuT+IOf3D2LCHhnfV/PadD6VVD8KXgN1qhQPTHcA3ba
T/DDkTSOININlEo6obLVvLOi435VG0lj1JkWDN9rh3x8Mix0QK3EsZoGP1bnmxUMwTHBz8Z7XggJ
Xf+nwwmn4UNtpXQM8SzUBqTrtw8eMVRJgMgP26YH3D5Hdp6EGNtY+iuWKTVUN/DtZQW/whtxnLCo
g12+XGrk7TODlEesGYTXzR0CltQKCif6vAw5F6lxxm4q8nno1Y/JCa3tM54joc3vovM3OlqXBRrw
CM2+2IklfEK9Hdf6Y7duvn14HYjfRTqfpAqMS5MYDfIXbEDWAuS1pL39TZSK88EP6RmJUWIdfAmF
yDCOTbishuSbSv7YPShN+qj++vKsdQkvIqq7YJbnNsUfOHtgVB2fHTULzQ+arZmCco6uN7MFy39D
46sqsNLWvbS+EQPveg3iTbNvW8ChlRClzrB2VH/T/1c/lX6J3FND0MrHNnAPsuzB6tP1MeGRpPoJ
LDV6wR8XHVoeJYFQyN+0EIIFGeHAcz2/Op7REst+EpSFV3Dx5mAuEmSm6bKR25tGx5AlAAC8rHqd
OWrcWHZBT1KTouHZqeDe1HRM9DD2myYEmdcP1LLYVFe654+cJ0QPK1G6dtSoBBPDLPhW8ZmhyNx0
0Da3IQFDUkZWLZSXbkq79JB7llxldB8VS2ctCEXL80VcwiCeL8XT0oY9nJfa9HMCLPuajj3sS/vr
VfXcV4ek4sHzyrYVupAtJkk+tvRkMtPeEKVMGiGdhxU2pUnbSAL6GBamCQLQPzt9YsNNOj/ST3x7
nNOjXrUNCnvpySOjzf+DsUvp2KZnOeVMzTPF4dany9R2bRomyzGa4z+6RS3oqOAMyuiMBahVmkHH
95xuX4zGTWbU40NsOKHDyzp57xaazjdHWOekSRkpH255WYanDwYVhOBPdBVERfdOn+V6ZJTs4qIk
QRP788C02amZxeJ58B6QISwp3H755kJujsxO0636kegrbbxjLFXVqf01+hwiOys1p4ScJkjnIeWl
91UtgSNhN3/Um/f6WRBKPqXgZdc0rGMEUmlRgv+9lT0frmKuXZkiWcIrHt6mmvH4G5z1H58gPbfR
XVNuAo/x1UGTykNukzstuPZ7RVxPqatTEo+qwF04edKdcy5xcx5+i6dS9c6Uoqo4t2px6TnRvOdL
jcDOAEZSHAsJwaDy9XyxmiCAmcMg1EnsrSVKIGYYe+GH+5/NtIdsqsT4vuNiEk3TzUuJrU3Htas5
YGC8tVpb7FVncVDcHBePqIBKPqi0z5l7Z0LeQnCwbs2oIb4yYqugbPmPHwiKwveeKPp1F1sp78+H
v8pqWX3WlRrpRjGQZGa0ZjTvaSxiQ84o0MEkLllmPBZRfyMYGJqTastdDIe7AE850XZj6Aa06t/r
ecSGXCReKRHhJv0on8SGehS3CK3J2sqhheFZxzK82y8kMqyJO0RKwIggLtZo7cJYDjQOchXraQLt
vDP3Wkm1hUxJemmHBmmHRhRr8UueBW8SSB3ZVZa4dgt+ZE/z7kHKianExzZmBtAJ3059AcuBVhth
0BZrOudQsOi+TX2BIUF/5yfpi4OizzQ22A4t6sepyTK8uftrdDEId+wr8QdzvwVufRyMr5GG2Os/
g0DrZCCVLHWXBKlL2ytoDImoaQ2FlNZoMe1ErlmWeyQ9Zbmt5ugrqV0DPH3QoSFjPjY0VZ3PITyu
TGlBZlqIoqvTmTMaI/+P4kkAx4CQVkHgDx4mo7L7iMTtRhb/d205YIiFge3WUv9LUhZzncBQLMyf
lkEhhUqJU/q/FezsawdUK/JjY/jkkIk8LMmYxoIxZ0mO3HZVHRoNRNrCIrZVTr/hLAs9Tqvwi/Bf
qr726XcSRygZjkBYiDSGx+TiP+wV9zlVnSK06cESeHIocCGjm+rEk8o7ahbhDNPxREJVnIi6pQUc
u3x4eIaNVusaPQJf/JOUI8FKCDtcs2onxgImROAHQXyTGBuMGg4JqyKf3z8g9P6ilbxcUbXQsjFE
19pt6hel08BLGNgwUGuxNALJgK517z3rJ5Y3Hl2mpZj1u94l+Vby68Gm1BKn7WhkuAjJKc9E78Ry
ZQO1Id2409WQBBFaTQw/RbBGXze0sflgFP5o120opbPVDsoGLjSHxtQz0rV8/LxOQiQoyY2iSp6p
/JauVQRi+4JDivnthXcRuB+UIpTQqGlsoeeeTct5O2AE7BrZMa3REK+wLvxNwlXbiJ0pDa6gN+nP
DYap+YFH4UnamiNfDxV4ksZoTtonaDDA/1t4xVUWEM8WrUMVmlUM18OdOhkSNs8ZSnx4kVjSJ49J
yI9He8NiuyA05Pfp9Um+GMeBBSTGhGO77hZHQ842fV/4PS1FGLTyW5zcJOt7Ix9vIVgl1R+aBr8c
Eswe5gu+PUdHf2FgeWeLyF5F14SCopZKY7fI84Jrf5Nq1iHvYreqvQLAesVHidmQgyAwwW4OEULC
BMjj9JBe9lFfrZvvGtByV8LRwVDTFVsT/no4hIP0R0QvUiXagcKL3sb8U8FSg6j/ZsH70GYEfoZm
qa8eMhUQ3nQonXHdOA0eRJSDsjHO6T9CgmJEslfREFEHWY1G9UfI+BP829PJkyApOPNy7Q139UPw
BBgwOfUXzFBwX4+OR5JAaL/7f7nhqwmQTrHJ9PgLSC0KoVrIjfn9CYvIypsigjbcBwhbwaFEaPMa
gpW68iny1HuvFA4sxJ6qTwATmCaLetxRIdMllc+J3hN3MPimV4eZ3dSwn3N73XBvlwzIqbg5/AjD
so7zUIGt9xifun6m7DSlBLL+FVWok5Q7D+kZwK2o/c6CaX1nMtd06e/UtgNF2cDPyad3cT379vkB
jCXdePrxuomrHKFkQfR+AKzcoV2A6DmG37mRlV9mLC5q3Zr6EbK73rBikhxrZEgDJ/26AYAEoE3E
V5GDVn7U230cxW+MZYhnOyHbH12nqJ+LdUtWhyh47on6HQw5EtZDmM7CnbRZ/FjyKX+WV3Sfj5w3
lm4UssqalYgapf2Bm2Sj6qIjxuJ3pCf2HNReItqrh0Y7xtwJZnKVFnj1RYL/MAEJu951t0i+msg+
8eKAhsDqDjXUU0rtDVYR/mN7kFLpDN04GDWVeAFziSMXQ48n0JnW6+U751l1pVX4Wks0TrnwXB6U
MY8iOzXGHFYBONE8AdOtdYDdPzC/eY0P844c7icaYHUFOZntNXys8sKU9V/IWSO5tKZ1fdZrXTL1
npJGyLOg7KrSwq7jmMzFDuSmqeiFf4WaUK4RNhjJJg6thLYuII1fqyLtlV3ENbpBufLHkKhbM4z/
vAer2R0fq/N6EfJefnvyT2wTSyzI8PD9apDckSbkHNTRD5+jZwH1LFqjGk52ath2/5PkrJKYcyEz
iHciGwRK75NSKRDvEVfgOsHxi+M016/UsuVDwzGXa8ch+3k5/B/HahYBeD+qDJXDcxSRNFHr5vB0
NaaWglrTJr4LD0xx3Qb1015h2oH7rev+cevQE3I4F8b4+yM2h+TtP5Q38lwbS6sof1kZl78LQAzZ
CyT/iwVqJ6OJuNrH9TmFzj8mOHhH9KM8aqeTt6/dMwdPItni7a/BXY8fTmFQaEMWyJDvxPC/YPj8
BZWnHOIdYdF+YdPVVX+M4ofufyInGUIcz6D3CnzTNcDjOEogX5WEurF3shvu3NnH0iFk0uuwm1B6
PJeRmpFhc4ey0JXg9Ffv39n5SyeI7rD+jL+cmMurJJO/vTuexSi37AqNdzq5wZC8XkClrcSg7CLM
OybLAxJKq3OlUzbHePGmwHDoFIESyIvYREIvtRbORBwEo4C43k7OlOK8LTPfxGk5V6B6RYFdD1Cl
uiPibtgSKSgW06FldRaOGqtlMFKaFHmWa0aOKUz5QYoYAuiC0dixVcmVUee2HTseL9yC1+i6hWtv
QyHwoKW8e64tHJgtvbSEMyYGZUtVePwIJNgw4BB30HvqhUm35shWrLC3w0UAeJWfeBWzV4gD8wtx
/r8RKBqj6R4XrYGEJ7395QeMI0vlBtp8HRWc2LwbqYST4s9cwEmjSnV7DOFfNMqO+9pBJaq4P5ne
PBTMQ99lt2zywDv8BNihX0glxbjF7i3BrEwdWRe1q5rTWNaPjZFHJkavC8Kv06/4wTKGyGldtxR6
PENchDdWkMUxH7pR7GYvvBBvYC3iNpUHIbE9EIefpjsTnnSiOBl0Qhh1plap+kVdWxmwz5PZhcNt
Oqmik4tB/hpDnqgSjqJ3kHwldlmdiP6XtoZmVJ5Y3mkeCOTA05slR+THX2SwHriNUUe9/civlpXl
NQr4wLL70/fSJ2WBEPY/Ezy+ZMAarz8SWMRSegbyMYQE7jnaocNGxsI/fqBCTp33ryJCEiftIudN
e9amaQdwL9sxG3j3BYJkqX60hwuFsdy/uNlxLo/j3Zzz/i3xIF++0NHVA68++qLVA9sNVHvC3M9X
sqi5KPi+QklGEx61gLs2Pr42YjccA/pN80Q/+F3tfFxMKKitxtULa8AYRBKdYaybobbhbeL772N1
ybCZBBxbxthFNAgt6qDrR4gRSTwJWXI3Y1jj5xXprtpPtX5Hzrdob7EFLGgFtSHTH08BkKq6dPQx
xgwbBqiVH3wSohdFq6lFLhvGZstqBomkTZQwgjLhscpQ94krWMn5b2BB1Sb+8EFBiHSb37xzWMJR
Xp/pu4PtqmuWETKuyCmSokErUdDswrcw9SaMEx1ztsdruwWMiV0mwW7PHBpQ39a+pzNe2IfYoyc2
LFHLTbSd5nCQu1/mRmnNI/45HhL6tV/prHgz9qJsQ0dhAbna/EqCkzXxuvbcX2yVnb3PLCrB8PFo
SG2gFCWrUk00Bu6Tm0K4KcUdTWD00oEacAaAlSmiwYk1ETidK1d61X/1Cv4afshU3FUpG7b5R7nq
DpeJg3weJ3qqVqUtpZ9uI6kLad60mMbv/wmZEHFQElQkR4/RfwLTB4CrlZPqFpVEr7r8UVzijQk5
FQ+mYMMx+jrGFID5VtHeZGGuGgCCCav/owHtot05aNpPfKxiTEkLN8YZjmkZNBq0Iiq1xcmtPp0Y
HJqpZblE5MN8LuM6y9xUk5YdiQZe1CQHaS4EAAHY6AYNV/ScsdI1tS9p73sSSoGIAJryJbQUyUt7
IX1oRbfijXkCJfLAsS2DuLEzBlvUz7HrJrQ0qv+6rEj5GgIRtwmPYvdvlulkPRcvL+qmC6VM2GxW
vNjjSpbP8N0JM8D1KJLXchcs9nvU3FCzek/QvYSLWaKhe4tlohv4ukYDPbOHe+urC25yH4+BFT+X
thBZ8GgoHxTBmth1+QyscuYGfXBoMsfd4IyeBsdpfbSTV+rKWvQlAx3YVDOu/l50cKcwPUjvvjDq
Qu6K6bVNyPEP1PuKRgTuLp8nTMZhlrmdYfj51fP1PsmrSc++IyCu6O+sNSI0N/HrNpPcArQMtYSZ
sflBZqC9aNwv2kBwZwFbjnIi46seGB1Xoob5D1CUebV1gQjFYXTm8/fimPRA482bUZ8jgzBk7jSx
CiioP7GBhvp1kYG1jA56OoUbYkQOGv9oySHGI++p8Ry10pFHzODFFXq+1Mwy9GgNXFIheCzfTX8c
Wz2xK707Pk8w0JXN9fMK7VMczYajHANYeEVZhG91Ex11MEzRSL6y8JzkoAMURaaZWyKtdUdMdeTk
8tUZ5Iqr9PbOZQxkOkQnpMr+lDLGy+UWp8UgLswEjSUKAaS7RpJSx8Lq+nrEYH2u15uLo6fMtNcm
n3l3hoPmmHdRESWYHuID/gHMruZzYSLqIxQoyKnsLzrHf5tuqgRZkw/B1R+GKjSz+3QmJi0HyzFg
mJXyrfQPMnM0m+3p59aOfP4T63TS8EPSRc0Frqnkx9FPaTS8DCVhWboMsfCRqJYYgW66nJNYFLb/
O5I6XCXa52eW10IM+ybs9WFOpf5dfQxtY3HKrOUqBpQSwN4OrnV9YntS7NsF4XjhVWRZD3A2iqbA
zhraDKc/ggKTE8O+edE2v3nIjZ2gEb9dzKoIn2b71x2UqRBWWfdefB3noff5hiVU+HhROwzJMrK5
32/UR/5gUnwcvYXu7aZ7QdAeu1VeNa0y+DX6b9Cl2y5XhLJebuedcV8nwJuzSz+SDcpYslX6PJZJ
EET04HJ+PyaS3W57iQZXN3kEZiBAI9Qzz1AkI5iNEmghAVNpjFueG35QsM9l5CY/Bpf21fUUoWQw
5tHPsoJdkedkq0cKIh4dIwhw5kxHDhTgFKfTM+W2JeP1sVoBtEV3D4unUsty72mWHNFqYTMy4XMe
S7JCcNxPnt0jXJYbQwtowpgF98c7XMRWhfYxNcrRuAQsKizqkBuvlAPMsLJ5nzQs/e19uDsm9og+
dJOh0qw/CqyX/3DJjIzSMI2LcwDjfKoSC1IrYdyq2oNfC4jo5ZfuH3N1C4OayIowkkO08CHJlj8C
TwZGX1cLX8ZhhZKC7eLtndB6XpxHoJEtKKlSp1btC3Npm0XjfKzhYK1aYU5K1IReweGsXX+BE9qQ
vbFsGB4bI9Y85V0mmkltRuR3alfu0rBInewbP88mQ7Fk10JJZHhISMkXH+VrfcBpwdZ1/RjU7t4O
rXIC43SeLR3Umkkgpj9GAcjFwnX3Ny5RI74ACR3G8om43iZ+NGfO/4T+J27N5QmSquJEEf403w7i
g7wmw3813/3uafoPP6sk/U+A7G0o+sCSFhxfGvgpt+c8+xzwJecrq8elN8grv9V+JvD31VS2horu
0NaH7XAegqVRqs/tSnr+wUxVvcSlZTtA13LP6iFs3qZfwOr2G4qq2l/NnvxrcTHxDpThJzMLwVNA
bGa4DBgupT4AOTRoU3CzfHB5C76UzB3xWwdMemS+Q5kRjiNMLTo7jsJscPh9wt6b5t/LKD87e/D/
SR0qypdiXBoh8MGu/Mal4BAARQR67lvQQlKuZsJc9OyCdCJlh6cGQPF6yipD78op05mjvmLF4MGD
8f+8x24sj4ikyI68O/Z252TzE6/5jpYiXew8iOvwT0l5Ocl7D8tkDOCwt1j5VJosWt5jOQV3TtSS
eeSl2Dn8XBZ9QPpBqRtjXwm748TSWb914HlD++Oo7VZPChdH0gNHfyosr2tCsfNRHi7J7RV0Kf82
Yg9HJjd1jzacvmISCCXbKA83+snyMS7P6CugpF9jSTZZQvSjESTkBrD+HgJUO+R8YNYNjMyASs7e
HBLc+qqc/nxDYr0+z7QhTbcEC5ybbvKCuu+Rr3XATRyTkz6Uf/KKpPimt/6cPdnla6bD5/rQ0fP7
/o2Ln+J2bwGWyvJWEpnASLJFeHbG3NtxjxkUG0XnPSxSmVCBOPY5XrhuuXrPPhds4xlh+t4Au+xE
KnmMC2oqoeUFHoqXJSH4pB2rEoJIEeIC5l5PgtiKy1KzGDP4OlwCQUeu1tPfJkHm7q/cNViwTcKJ
geyGSn7XvdZr8GQaZhhqpKkmsqHe9D+KGCjWjeyEdorZN37oFmXIr/uM9Ak2EOyQhDD8eAo1k3Eb
hZjgzFO8L9fP7HldAR8n8lSSp5iajFHbG06NQ6DimAlWeaEbLYpMyJV/BUXAScy7n1Iz3k+I3157
OnQPWrUO3dXXO5/MzVRyu5Pfo5xgHAa1qR3Pygf2SteQ0JMhYXPgek3IACpfEs1XH9yfriDMv+ii
MuF9P2wuDwbbYnfjS1EqPyzW9RHAVYnObKn8UakvZZ73PfkrfjrzHkdl1+iEmZJR3+DDL3AS7LwR
lUb6QoPehR1NY2UsBvsc4aSA8syKKTp7HCmlbJcHNY3BlsnRomGOZjaxxuDV8rxGWIDkfErWgv7R
5XY6bQYKMUxTtSCHjKftEPv7joT9c5XWSCTy30LI1iuX3e41tiWl2jlM0sLol+RngCEAu4NVjJDA
FJnuThhdA5CSDF82oH+TzeHhni6LCCHeD2AMOQk4+GWaXPjLZFluXI9P7AtjIHKXFyd0YW+52jSf
8HpRVOnHxed1n+19KcFiyL0dE2/8iA0PESjOWKhBiweBBGcxn1Ie217bR2JwrirATwW+N//I71qY
Ae8eXicWaNd4tlkd63xZNxSZzMP8TXG7CJdcBDcbrsNUxyZdjdzFJia/CqzLPZ3dyUbcLkhf50yb
t0OiSzf98Xp/khxXi2soJC9s2AL1Y6LMeFhpQw4l7whWSbo527yyV41EZXAioPNJPDhhIrxd7J7D
yDOp0YEAAP/oiESjLTg5LyIpVo3CtaiZDPeNDKJuocAAG2C5NupmIhQLpeNYGCxQUqdbidqChxsE
aT7WgVaKUMmeCSa/iDBvasU8zCqKnCrJhv0FQpmamRLxzbsN2mF5UtqTMz5cGVcDQLZ8c7jF8ikC
DdsAGTfvZkdU6ylIWnxB4/t4qs7CjuF3TgP4BKgCXcWovyCieUeHF9N07zLThv05rRrwKnk4haRR
rYT6yL9c2Iouw7JSvu/WN8Lcz9arfiYU63lM9BHZZmAmapHc68+x6QPFYzW7/y5wYHwnHpqYDRr+
9Khm7hpRy9n843tYCIxSvneIvCueBlp5HYBsZnIxVuHaNE9wDiXksW+rF4YrWun4zDX7x/c1pwxA
5w/YJmeNDPaKEIfeY1jFe9pAL6EBX6kOqL3zAsPRtVptLFprNydPSo09rLdTK+oUZ+0xeuU19rmW
+1asc44tRPg77nRyzDp/b/f/4izcfLnOPmj5E+5whPx11mSTVE2T0LK8NqFBNC8rbY2H6IfT28zc
vCdWMG2miABjpmamFQF1zK3RuGdg5Zqo8UW+OJVCCUzxmaZpoCv6+STPKvpqCIA9wru2JH5WpGX6
VCIichpZVTNF98jnWjEVx9ghYCgjJ5ioclVd1lGIUWc00cTWKqnMHMQzpRf9y2+4+E8YaGKkaWeD
or83igxZY9WeqRVWm1l2rVvSRDDlKNjg2G11slYNsDs0Md79rj6Yqc/So8dGFpWRf8t3WPAZjeYj
Hp0y5wLgj/Y0U0HXT9H5bNYpCK9zBT3Nfb/8hSjE8rwCq7U2cSThDvawfBJfZJWpORzxSz0Ws9gA
xwU2DrIm9j1+TL/IHqRpmVzHtWY9qzrx/WNWfWxJb4qvwtJ7qcystW3ctcUerzuQFXCw16ifrBWI
RK1+Ej54EC5qD7fVhy6Ol3PNXGA4w9shZLY1xqvLe7fKMA90VOYN294PlEK/Eoclf9PYy+/6zaCQ
vIAx1MkvtzaKxt0soL2l39XxQQuOAzi5NFWcD9+q++DwHfvuzDgx662bIZd1sLRS0PUfgGpCuirA
32QzWn6g3kbtjYqxZPQ+wLOCchSFHcmWkfhHx+3OF/X8O1WNH3a5jFjV5X0ld7EOFQklZoykUdCk
vU39Jd2Zu8QKIALLEyME/p1fCuGWSBKv1vGWvywij22sgr/eZgxAy/Cclaf2j/NiOcDOkKQ2P8nD
xCUChVpHWlrdkA0Dv6BpxQKRPiCCbiMu53MCCwpsCcy+qZu/XAOZ9M2iOobrQLkcQNvPfD+o3uWt
lsoqpXBtrMC7JgYD/LmylfMgcLa6gljcPZaVjqV+pCDl4G65qdN43RKgDzeYHWmHlhUUFEt7ppRy
B0B0dig7ulI10kGVCDJX59Gc6d7BrX/pvLLsyUswu+yxtBrMKtLeggYwCThUQiMx+a/xW+tY+1Nf
BfHlvJZH3Rb04zLPvZEMjmj/bh7s7lRKSxj3IBQkXcj2TUEMZd1XV0PdhxWR9GK4vZwY5dMxgrz1
Id1zJbKceZmM2cXDR27l51xxuAopRCcxZOgP/NcwVQPh7IX8I3ff3+sCtxxjjx66joCXHOVJy6P2
LTqenBwrGNSlUhYtcYCOz10Gqs2FRcjhi3+SwAXR4Vk9RjefdbnumNy1ALMkxui4f6JjChmmofHh
g4UZUvhUJy42el7B0kla78wDlW2Qk8RMyuVH5M5cC/L16qJ97U7qYJq8FpzK4xgeeCcOfJMCJn5u
vryrTd6HlJGdxDHl94cnQWvPgUiYhRYoA3y9kgrYWM0CSixHjlUS+unCWeZhjkAeBeIUJbQeBVZ+
4UiRM6ePBbDs9ROj4D5mr2d7WriT9PpUIyjJnG4JrNuSZ8R11p1eYWGYeNgJ64e3cf9T0w/LQV8s
MacCccCRYLBWJBnlgxZFEwe6WOwxfNeVJDqIpOWjICMAaXFUQX1P6Hih6mL0Vf2M3orisHGV/0Na
S5Vpd8DKf10h3DBNYI0y686mEDEvG2cB24b4J4K0TBBmTUCUCdmJGv4yuD3ZeXxFZtN3QlZ7FL3c
0ydcrTNCy7YhFd3hyxk3h+jaWNT5zu2u9AHqcQ3XDMQNuA8wNTxSxnFgjvRmoOLdy+B8TXr38iZI
lClaNUQTqzy9+SXZtQofjiZ9Qdvm/e8Qd/3WSfmktI+3Hr3UUgws20f32Mh00Th7kOqHD9Awg/jp
Va/eOOL/CO/fxYFGbOG8L/guhKyVS9s/ZNERutFcrB2rtMRaEpNEJn8E3ZS01PrurFk+1ydQf3DE
5akrlKDTOsIavfTQj/iIqX6UXUPT8I3beCxgcr5ubKQc8NSCsOoxW4z8eSx5Mmj7FqtEOT9Xs6Ym
8xyJrvHOQ43IFscQZqaUvLEbchEIuz1WnbC4nTv8zMAH86oludNYyK9MtEZiUJ+BtQ3I/cakbsaN
Hagw15CaBkcLb/3vhhX3pXSDoSxf4wT7FcYZzPJsQGoiBuYQ6+yy+bXvu53doBMC8+qU+oygxDNz
3AB3KiWMmithyheC6iI7xqcR9A9lSzwGcdROslmobWXVtcNbUM0Z4FRz0lbBho3i/k4etx04bAig
SNYig7A/htOwacMvyGZonL5G33sgADIfNDlMq7W/GtcyihE46HAbCbB3Me1pBqdDHS+8pziqLjmy
s0ikwOZtYQFyHwsPDTGIFb5wH2qM726/8IUnN0v84wr0k/c59/gO3lmJA2FyytN7ZF5eeacrYrPT
c5woqF+baFBg2LVzZgDJNbdmjfzJo4wd3Le0dH1XzGc3eXrFnk6yKmqk9QrSJqQ6pbWtxaRT68tO
TIsqhSADVEtpPx1iR2n1qMUZa/nPGTVGVVoNzOIPNaVuZrROI/mJhc/YSq4MA/omR8QtR87/vjBg
LwOQj+UnaoTeXefx2Z1u003gHjMkm5RG5CQQ4WAwHNuelc5Pb/MB2j1RsoLdsLQmjadMSEUEhZuX
W+QM78WIIypXN4RiMlw0OZYPHKnHkti51GaIK+BXPFWtQtEHendra2X7TmLw1GEej18j7nKP7k6i
e12BSxKRnrfdpb9b3UgspDZARTvOhDtj3e0hT7k2s3LZlw2ZdjUCcWn3t4fJ6mo5fR4VodQSRJz3
sEZmlwzY777HpE9zPF/xCtXRsITMPRWx8miL1isDiLN572e42gHAf4Dqsv7qQSimSL/PlVKDIrPW
FPpB35qUW/Nm0g9c8eIw9ajQaIh1o44clo+YuLhxtQkeVCkj9CD45gkQREkCAnC5sREJhLGdYhC9
osLiyl1ohFGpV3PMSnrFGGG7pP2PmWW4LHBPNMuBFG+9jWT8zda5NkfYvxq+pT6RZ2wvA28UpCh3
IR3O3q64nBfDZn3nm8NKdLkKvHLnrMlcp8+/x5XSv0ja9a6+vPGfDaacpieZ1PicZMHdGYN/rcmJ
Z+dGrjwqtTYLgaOZ2hfLezrTt0RqlhksQtQCU48CYGzTUWLwSmjfiDakTdX50WMhQ0bdPmNrfZQz
hiZ9Wm6auVZ9eCJMQTLQys+MnFwZlcwvO2pDd3qKLq69dSQg2xtJe+M4If8WHDHqlE640pHZl0Rc
itgn2MJEz3I0oD7PC28g3XmK4RvLgi/v4YK+SnQYKX2GEDSvnwB7mMY3hzXs2lydTClXYOLjRduQ
XcSWP9LP/LbFOfGRlJxrmp/jj0tclsX+LtglTrWrjUMmGHMcUoLvAQmjeSVG/9VALM85A9ZQd4GF
k+EGFX4aEsM9Nl/xjcoUn1j0kR1upUs//M04Y9yF4YMWWTWzHawwAWkmjVI7fiLjXKE2RoqA6uSf
+Cg/0Vimx29ctHqB2mg+8PvfRxfzHEQhv7r0Y9WV5c1eZ9pkQQskplxofLw9Lpv70HSRG89JjrU/
5ahVf5TNJw9yxwHodQBxe3+1wm+ZDkBu6YMUAt9qNGWdSsTMn0hQi8qYY4nRo+MxdR+/aoobABAb
yfAJ07ffNCwh47QAVJn42YlebuTZjTVHtDyIuEqm9/LgQ3fWBOt4waP4IDWZ1+4ziB6vE6Av0z2D
rcuqh2QMqfprisDJ/wlZ3QnrmRicxes/WxPTfb4KJlNLya578VJV0P+7VYtuQsEqwOud8arU490g
9TIn9lhPHbLBPgFNDOtsjFmiJQBzPBLMfxaRWXP2isQLQ8HYfjch5xPDxyGlmOGS59O73pqoG9W2
PHBNX22g70BOQ3XYBDlEW330Mrftghlbys7mtDjy7hW2pWL06VrX79z6uhXJs5P24OSTPJjV2ehN
/Oq5fPekLx0QOe2nr9Aoy4S3vkTD/x9XR9aP5Z8SqMMr8LUqEmsFaWnHcVR/KRbevL4hQcbQflwR
fgVM7u+ZBuUCIn/h92AxdoWySX3GWWfYAWQ1Q/5TbDFFQ70zZZ++6vENequ7q22ldiK03eCRI6/G
ga8RUyj+i++ZtK7aEcAfT+XY/GHP1+5AQuTHgXYLbOapNmCD7o0UacX+gFhmC/ZF96F0cFnCXE8c
O8uphVIcVfb5JAKRSU3jgwjLm3Lt8CqT5rbv1rcc2DrP3TjWCmws2+W0VNVgxdwNnRyakncAV2YV
iTuo4uGRONuuOS++ENm9nb44ggefqqNxRV5l3pW38eZcVOHKVocLBEDhl5k1Nm5bjXTx8yK95vAT
LZOobAMkzne6tP84K+CO3Vodl/0bSvONJPvdgmB40qiCaIOjJcwIGNFVWiz9q0fRtA1zKcyNgRc+
KdPKevmechH85myeBQ19Jv34YQc3YuS+6SAXWFXENWE6U6Vxan9BZk8xb1DrX7eFpNp7WhHIsbLP
n9NiVkP6hZ+/kNLKNIvXXDODT3axzz+/T921IAS0rGBXL0YXniJMq1Nb47MySUze8t+Ij5n/Cci5
5lbNXG23nqEYct/eTq9GWPlbNVsI+44D/7S7t9rYTLew2aZ15fh7/UjAt1gH96effu30mRmPOHQV
GDZDwSc8qYCI6M9fhVfVckZNRMb+saCqafUJ5iz4OaZec9BwBYLJtfB4Q355jhq28/degtsQA54A
qCueGoBkHRT29rkBx4FBe5Af7d4JJLdatEoHD+qLulScV8p+2jCgpEQ2ZmPQFAGmlARHRvtZcfih
Ynfd+i8i5vE/kHu+vVgo51z6etbZuysA+8QX/HfXhNZvHBdkvLPy8XMfcuw4xBUjaqGFJhtkYTDa
rtXYg+CxLPSxUlE2WF1sVZGNzdivaN1uT/jkj+O+oLBi546U+/jdM5nADoVzpfiKztd4mKrnb94Y
5R/Py02HdNpPClsmTZoAzdbbB2RYdx793EU4AgcLE4diw+eGhFcJ3yNfB0Y1kP+PUfO8pcOqKMqq
GaFepFQiuSyjm3hXvV0d+RquHUnu7RFVpoQygiBXP/LFwtYG9vLIRC8km2pxI5L5gOyavgtD3io7
Mxnkny/BkqsV7S8BnN0tbdwYkGYJyANvraZ/NhUqhWDexJ5L1r1TEqhJhF43npVzxoMHcQSUMILu
zATYoh6SuGxD/Bu9BoLZob0YWZYhRRGbJQcM0k87V+NMLv1OdMQa1R6NNbcA+a3WdjINqBnix/xr
jXv8zRQbOzcN+chZJqaeYZtXy1ExmRKC3uLZquJTS7zkKwwGjChHV41lwIzOEtg/vyfcnfsxoFeW
yLQor1Oq0YOZymCBez8qgb1Cg0m5GL1Jo5ptFX7cf3o5LmzZcL/TW8aThOBEgdEMjGvFQW4/x8oM
/h54ccIFWadFF65rSzVcg399kOICggUr1LOcRPMiX2EwrOaRrIX8NVrZamWV1Ut9jCw024WDnnLk
+7Xhg5SXg+SX7RVZiIynIQqFrm/2WTOkd5ILla9D6bI+8VXnlrnyF1yiFF1asKPtvbXenx0pxGTe
t/pZxUuTPDP8qpaoXXILa2za/Tavf6vMj0YDatp5BqT9HjP8VLQxt6Ngi1F6SbbUUvCBSz/VzJBb
Bt1sQv/jKRvnnpvhUhLn95KNGpRL9NilTA5qukooPsVH4Z7gqODFdza7UEV+R9CTLSWky+LP80MS
6UFVkdGCi5SqP5UjvYFqJMs2wLVrNVkcXOqyfkAGiz806xtwLxUZAU6G5Bv8FQ0S88NhtvDN/iIL
UDee9O3bv+zTyry8MDTGV92IjhfUTXBe7h++IoH0Lq16Lr3Ey/Y/juO147XPx3521an73unUdf45
35EN4TpjUpVi0UXu69qYF6AQFQwSGNPc5e/mywTGNVR7rVmC4Ym5Q4a8CyTmuGZ6eAPNo0EIh/J0
3A2ZzadsKxz3mWJ4IitntwBLsuc09sjD+RJ/J9CpBczJJnTcrtlnBGal28+yz2yWrde7HECyBFGA
oWYjtNhqfdB3mbRV/5lZFvIQD17HacN4AWKlg4pPVBmLZxI8cvvjhEk/LpUg/SPGZWrD/GjsWr+r
bsS/S0gWkG83Gf/27TG/cGozgAtwUaf5FgP0s1+Lg3/vd6sMbusp4M8Az/EzJnMfsAAXQDvfdzvo
hpd35lUWjmg6R5RFGHWq5iBRKqrEJjMK0ez1HBLAj2JkbFY5tG2y+JEFjoSvJzPFUVsg+My1EZfb
UbHRuIGBUNBu9oFKQO+5xgFndW2umSyvKkMyU2iX1d+C8778zPx0WbdTLmOM+2WG51kA9itrHjet
IjNdTtao4Gyd6h5FjQQfUnLj4Rew8zK1sZYiDcjfrOf6Uxb+71dkaz7SbGEEFc2gMgLywf850OwE
ihgXeqR1GYsR1EnulqfuOZlIPiBVoMsLrC9xUbAliOeiXbj7q75dsufmCDgmLGlt+bA6816GT5aT
Fel2l2TCVdtIFgm04rjLh9f5DFoEAXvJlCBTS+JtBu0tQpmB8sCoBMF00eWDZ/XfYZe0ZJSefLcs
//TLN74RYhXnH0KNrgLe2laSljqpEa+U8wSHeNmOQ2EjluAqtclSdKG+mvfPSp/Za+Dydc24bZBZ
jRELsrVZggTVUnZ+AdBrLj83R9ByJjhwnd6thwFpOa/UpOWEGQIofMY5fn21/f/4nm8eOpufu542
pk9RyClb2xk2jQ2haWEChH+fEGyE1ELjBYiELag9q7onZhRUnYBypNs9OYiuK5Kmg90tjDrS3ujN
kV+SXC1/W1SB/a82GT02iOskP6dG6DI2bNfi0qIqC+PHTFU2GbB9lwdcUCNaywf1GeUJyCNtCMih
Y0CI/w1SVKMYGOHz0MSJOshlEAGElOBnpfbLbZcfI7YLb43+xpj6MkYacJdQpj6a83s6GVHk4p7r
ynU3hD5KSYlyvI3hM/HTb1RMsLFSUdu0sfQWwH3eI0jEe6ra+bu0qsnMfHNwOqGI3VS5R2DYYGA1
UV5r649P9tIIJmWYnaDEl9WvaQQW6d6F4juRsWa8sEZFcO5PEHblo+/gYmFWaVBAOdjicWR9QEHG
vzOL4G0nfmVnYTMbkiPVbBcRGImnnmtYOsq0cg0CZznrbPDgxcu2pH4z/HPiYroXEklv0yVblmEH
YytOWIcPjPTqbRtyRJok+eQSfa/nu+AVozjYRnvdegAC6CRnc9MgeGMZgOjx78/ps6QJ7YyTiO/O
BIxxG17pFTFMa5VRz/s7fte2HEn6EV685ZYrTnn2wmXH9LirY/VT3g/3dYY9+fqJPGBLOXBoduvH
w30KIijVJbu8b5DrL/5S9BPoNbB/c+3BLrBMuZFasUzvl4Fw0i5+qgz2x6Ua3KdAvjDJRUhy4qhJ
oJjSOJ4bCwUWZ7WrX4gY/wtFcF+ND/xVmsBbpJtXCGgoSuO/T9ZriP7Ua/4V9IXTVSLb5eeCZfpQ
mU1CWCWuNhhHE6FR807VmR8hTcy8BulhmwZDkZTbLplXoL3OXaiCvgmezHBpiaxf8jx62i+n0xdU
CF4dYk7sdskw6kqT7wzoIENk8u+kavfi/8excug3YPLmE+0IxpbsTycHKmg1vjdjcwtXg4nEGYUS
zlSZFz+QIV7XhptjIHJw/N/f3HzZmj685oiclsAN/2eLVW5YAe56M33YQ6UY03vAlLgNDathKynr
KDiPmdz6GZpc86RkTTTWMf+H9Zd4W6uGLRdiyO60sSChBRAt3Hq/F4esMSiyHW2aGR5Sfn0dd+a0
j5ZWO5vxn5zgyUoWFRKrZaqQ9hZ983XlMeO6R/Bq9lIsxIGc6aoHQILLOUwmw72ynWo2bfneEf4H
FPxLRyU6QkHja+AKT0fxYJywkeCQU7GfGIwnCsgg8cWn4Ll/W+ZsFCCzB2kB0PrCoCD+5OA13G1f
854gEaV8Dc7hv3PbkudA+fyr3X0fP3EOt0ByhUw5aHjRX0voCHitxaQn6Qga0WsTsgnKv41dbaj8
8LZ//5GpprucMmnshqC1sR0HEEyfeRJiG28gdtZVkQKnNS7LSjsO/0VZtjH3ZW89UOFpT8hrmzd2
4yx9teYkrSK7NDucTA/TpAfjagQpikDa16kM71wDyswRIN0IvodqAWfLWIWtf2/mgS2YAgPBxJbA
LqNFErjAJjuQA48ZrNgtTxDSDsIqQYTwO6Ph+0Y0KNOQaaXx+7oD7EXwEeCQFySsaceyK3g+gox3
XlClEWEFtmf8Vst1hRameU8HNns9QQNMuJEoZB3oiUo2WrRsNMLq+E10ZHZsPD1qjSG7meb3QqLt
tA4bG9eZJ0d8J6zl1gPNS0os6/8k28GS2TnhmVqzhowjO/gXCwvevlsbC63FoL/HdrGJwK4PJdSM
2tt32yjpRxxx4+uU/d1wAM8mHBOB07QuL4VttpawPWJCif1sTeFgHYHQnQqEReLfPI0xy69C9XKr
LoX/B8um6/ylHpq+lFZeq3PT1llXJ8nqvTSppacdfGUpyt5tDi9t43hTPS0wnnP4PMBAffN487F1
NdtxCaXZN24EPJuajiHH/WJs+dQs6DE0ZaNH4fuX0aseRotaZQ6OXfwcyMPSMJ9kYcO9pGMpVWRT
WE+5oI9N/rsD7yDa2AitrjbDyj8oAZaQ9v0aEe/Rinb7yUXwXlGvsVLE4de9wh0CcFeMDTLHiqO1
cYSqOZ+C5Wb0YTSPpnMWHMuLZQH7jzFKUklaoJqE9ae2K7XnkYALVHzjVQBS0r+bzEFAeciR4gAH
OqZPuU9sAH44N9nZ7yF1IeSG7OT3rNq9/NREe8/GwhY4opPl8p+ceC6yUCoiSH2sG34zMZyk9UKz
sCjicdLynyL6/7z3MSE9Q8WjNi9Vpc2cpT3EmpUkG+BQ1xONURnUQNhptSe5PKktA6NDppGayUu/
OYL8LsYYD/rC5G+sFjeZ7svsipCxL5aGjXd+2pmwQ6qd7m8aJwHPJPABgIVEyxyidoQ0+IK1gikk
Wm63iYsODCGiW6JpmZrhdPXsRTMnojYXTuZEvPbZzvGikbrbD3vckzEyh3z+wng40mc+y43bNzab
/zvDtj7i0vYyF4oLKHmZjoZjDZyErfjCFDtk7EBWF/yoJgXZQfm1dMkLDx8G1bDV2u8B+EF2+zJN
X9qb8O94otMQkMWayVlJmKm2qSK9cIA7ZIa94Zh8wWeRkPnI09CtXDdhakJZJq5ITa2vutkSYiud
H4QxgLV9NU1HUVGB+tV+TVaO6hkN976AbEi+nyc2gIsU7Ce4fHxRGzqLfZDvjnhmwpAQgkMKsfbl
hUCbNEDa/v3o83ojN7kJBO/PYHtI7/rQd60naooZDAfPReNeUlvQMEUTtDqud07vM8BORFrj3XrH
jBWa0W3tap/kBKAhANXJmWSITQcjgQUSumGUbWS0VRrWKiZCgq4YFNvPWvssMGbXyG+S9GFwO4WF
/fHA9BnAKW6Pe0qZbHLOC8dUpNfJPTs2X9I6P8SbbACKqAcnN9Sg18iyPspiTVySTnG8PvtIarkC
m7HlBMOAf6V6ifR9vOzyEGZLgTK/zHpGlVc8kY4AWafB1SXSZxUKyuXCioVpcH1KJy88SCggIGsg
E0X32YiD/RUhAJQvDP4FMyjr+j0DdB/TTJAjD1m+GPuRRqM/5P9ZVeG15S4NsHHCL76g5uhBOJsD
jzEKq1v9mzMB3YYRIO9w71yXBBzpcapuwTr/dWV+cVthJgs0JBKKb4D8n+wulqNEXIJporLaBp/G
+pHF6E/nlLZw2PjNhn8I/nUaL8eKDxGatd5lreLYRL2v0sVS/keQenRQTkOKICXWMe8PqlaPtAHt
lT1FG8+5rUvFAzEXFdImthgYfwNmc/zt0xgBcBVg27Thixv/mRGvHQQjlTZctEVrRS/TJoevNd5S
YKMYiAt63vSZIHICkHAubfi851d9zytYTCpYK/CU4iPZOS1CGYDYLsL2QFGjaKleEq7ITZANDmXW
T5hJCUArNG5wYcltmnZ+uJMbd30UntPnJqpFqlAMM45CoTrrSalU5VHWmrZYyrckPqOcLPYerkWX
eeGHqehyeXqpfXTSo9ILS1kInsmLJS8Bip6E83TX71R3SK98PjSXk3Mbk43O8lrX69TcTiER4SBa
jlImzWloMLDkLL5Mv5du1EqUvjEBP+zjLpYJfOuudoaULwPcTMmqZBXxDSbD93mKnclA+Hxqc5Ft
fHplqC9AWk3EH/0lG+Ntrk5xfiSIrvsj5CEFntFzDiFVDreFTzy6Mgd/vAimqyCxG+UNrxoWQ3CY
SrhnP916/pjjwuKMBO1IkQwB7kUphbDJZntCCPYqfQZg5WE4sFPV9NjYqSiLNpI2y4fZ/n0DO0gb
LlPMvpDmMYRdNLMWB3utB/KY8AYT9zjPFJce3pw/Pi2DeJLQ1omtce5Zx3bMlUW2Mz4PI2znKwxa
Y3S3vdtpgEVTQ23nejiGYuKjp4QBVv05pwrOkEsguB+T2FZO6UgE3b6+F1ehTn/YxRFgM/Gu0ddH
VQT7NakVgD5B0+TQEDm3UfmbN7YvrATS4Xm90r4taLrLwq7kivxElvKwWd9S2Ri/VVc/Qv053SjT
SVcTGe+VWTMIwuy8K5Yad3lGXMSzH/QXkTZZ6/cWGjPS9+KRE39ci93Lb9fIQx3YcXCwmaQpGH/u
dqyMQEo9mezOjTm56yFIY4ppngMje+g50y6jKuAslenu8xH+xlgbutfU9b0nXtkshTFRRvsWmClg
pg3auRDAzOjBUwXZPoFlJ/S1BctozE9MxPfhGzd2iOCA/AJN5iNKiJrkQg6tfUiqoZon1ctM1eK3
3CsUj+ZaOEU/0a0iZD7YTAH4h5f7Kxcnrmk8W/zr0yCL15PB8EfaNZFGrRwHHCTXlkCFogmcQaVv
9BpH2H58GnaLZZtMdtAC+RDwC9Wjj47hubmPnor0NAlUm8OdBBGepZEeDu+1Nh3MCgI0YL6s+ga6
h+Y3yCmd3R9Kbzx1kraFMTCxuFBMfBvkF5HawRJWoSstnlDxKTgOJsEWk3NCM8P3IseKArd3Hzcl
8xzqe4p+KLoIuLJipMdWuYHKIgh1bJa1FPZN1SDaM+uXQQaQAJq1rENSrkxHf5st834kQvuFWCBN
W0cBjh263f4Sp8GvZBbqf6omVlrLWc6np+b71RVwYCiMfqRfXaLPivVIGYETY0LGEiYLOPOCLubD
WQekc4N2KxHYChrHn/hfYPY3Jd+REF1NOk/xxhH7vYiJPH90WWiZrcyaRUvnhMwVVo3UIEDm8CPJ
plZECvwthMoTKwd8ZGlEX17bH6EMUYKtbs1jzO0CWwj4gVO/4p8etVJMVH+LzA2+dOoQexC/xlqn
IjU3b5B4E2Zs9tZ6GpwUjUUr4qp3CHkxcgMqSqHBQiqBzHfbzX1Sjeb0IXM3xAd16HCmu66j1tnz
HC97zFMdbImZ4D4WKOAcFcDweJaQ806xd5Dorw5ZadvBfHfvzFbvqfsJ5cO4MT42pxBIq5YHypWB
b2qqJCB7qaOFuQUs5qo76QoiTZTFhrAcuDCiWlZ9X1464Abj51aL5aGZpNQWxwbOSiAPoG8gA8wT
2LE9m231LdtqNSO2+76EgvyaXkyspGr3NZAyBLYUlRDbCGe78JCxPC+JRIUBN/RV65P6XVSw84Pm
YXfC/DnZfPSXjqvpwKuBEawhHvEdWmp+Z2M36YTIgweBFEfVf9hWyiqS+ZqtFlNLZR+vOjCyouaM
z5DvbqEBTo+N3HdVUd5WW/0HpltUpcKvY9ZphPdhddNRSijvYXnvUKy8DB9QtNmgSeH9HCdkUc2h
kAwIbD9X/63fWSZBzK+QkRlrLRbvL972z7z8n126Yv010mOSLWpTSYq8agls9dLkaaOglaxtwKxv
SUuaYL7u2saU/xE0fmUuBV89CxrCuXEo0oaNgEa6DF1l6rIpGCA7jqfJ6f4G7YKzmMaLR3x0mODT
B9bP/7uYVRQIWGBrTAwgCKWEQxe7z69h1Llg6wb0bP7lZ5A02j9vmZkHSNjuLTncmEo01g3Uu7O7
I9dqktZEruazUfFgkQuWG2dTT5P9VLnvsoArCJc292LlLFFt4t1c/kT9MN1/5QJumvqB9SOZjVn3
a3dEqIg+/Uqb1EkC8eMRmkt5V7SZ8s8U3UAxpRY0b4aS8Jd8+ZTjjV6o97vO/KMZxtaHP9gTzJhH
TLw3UIyyCA+mA/Jw2/rMUxKLzNkaQ9oIMT3ftb+dt/bhqeAuVqEej3X/l9pJz7WucAqzpJFIATz4
ekqE7o9nOWyTEhdo0rVSBnhjS+ws/RFLwm+ScML7p6cpBNddlUEOC6HDrQWsYXwfwLDUvDVm2vzn
n3G6+DpRQeN5H9S3mdURZ0guLha71IZ93j7DEARNYuEyseH8fQ1CBdxrlfOfEpdoBBFe+K2udU+X
ctuaXvf63aYmjhPKubPOVJPfMYVIa1/PgWJ7TOOhzS7Ubg8S3lGbZLbvWLO2hjCvNkUn00pGbZlA
N82OfdjNyyNLHaE7Kvvup12O3746sAcS02MuAcDsdiqYfvq6bfs5xSQGciCc8WpsTLtOEBMXUTnw
rXvFXWGwuT9N2UyGJEHWxwUVZRB2ootN6kktwwOlNas6pYuMG0uO4HpbAgwEIAdLv5gCNzvEz5n8
w9WMefRNlNc9GMbL+T+fRAGEMz9G2cWRNydIQ+Egb8WSQZN8qAa8ah1PlpCufM3CjJcZiElvqxbp
uesDJ4kfnXzhmibD8gkmKDQ4fgwjZxf4HNqF5JW5TNCyY8i0bw1vp7qmFyI4Qz77jw2TSUCOBWC8
q/VnPEqVcRz26LaFVww+1Sbgf4kqPj6x+HUAvCw6p8ESZj19Z2MdiDRta87mwNkbw3orqPN219Q/
ppodTnTQyY261GPmj5V52ug7cMwGmP3AZ0NzXyWivYMovEKul+sDi1SAjDJJ0p9bu6TX5vWQ6U74
H2Ke/inCt/L1wsRNH120/LK/4p9c/PffnBb6/q30XwJXz0FAxVRK37gevtB91J+gMDudm5C21m8P
eqk90mU7CdBlypB0IQOA7vq6F9KGM7x4oVLQ6BYAQFLyqL4w1V7/rg4SJDhx/p2Fopt8ddjX4qNM
bvYuPqrCQUo8KpW4vgi7GL4yQcMgNnzjUZeqIN8DWzl/5IlY+ZZ1vJgt64Q4ByJOQqwd5b8KcRdi
vg/AKhySakKedGG1oxO3Rmr3DSjQ7kFhtrJsVH2GbjFhA+ZTFK+dlkX8q2CmHDLEppHnJ5ckHFPP
+UAhli/1BRTZCICkwBNkEsVtK7xj6lkKlQ88E+MoaVNC6R2AFseN3S2kF09UKHvPvalfPTeAbD+4
bjuXpaC3FZuEVh0s426D08CtBvLNGxDVNn+1L/lx8jd4m6yY6ukMmWqcG4Mam7XiiR7EGFslxotH
18nQxJHXr5qk6SaHpvKm+DkPvs8riABwlT9O7X07B2cFKq/kjD15gKLOf0PTT4/JCWQ0yFQCjsw0
GT69SbzmW5i3JqD4kcOeMDfTCFnzUeZ4Lgdv7VK4lUKBiiW+tw9GfT8otnd2rHzE6mOgvRT/5JBY
H3JbWSdOywuYqZ6t11tvILXBpqjeYf/VTrp/HkTXhDKasr8xtOR+50bK7Cvi+LqStW2H+WBFpE9t
hZ6v0aiqCTB0UKa8D4mWve8rhu3iOaHm9Nh5jvS8xayukQAV94GVaQz+j++CVF35qc0H7G7mHzYV
HX1lcR7LVMVXsOakqnbCxenfwcf4fZAKZbP07GpUpfaAhZ4p1IKW8NPgO9XlnYUzGMk/TnU0FqLx
bdiFwKDROVOF/ihNUZZBBqGvCr192LKKX25ohENFgejYdoKohfVn4eX1UiAYyTI33Hdcl3VzZ7Qp
+9mJzO7opfIkCR1WcTjgzYIxEH/wDaJDc9wjwFzc46kDQcK31ofL0TlDHC+02ha5qLkUO+ic8MvH
1EA/skwZIRWMlPsBNL1hFcxgVM4VHGKt7cYHwAuYBygyc1JDY+ry7WMZK8GgvQlxwta+1y4cf4Pk
Fg6nU0O8ORZCfVW/X7WI4KCJbiN6nif3f4gubh6XRsdEW+QUH1txgcYGgQlEQoEwpxpNX/SPqNF4
Xl0lmQofdUpBu3iBtJkXs2U8jT8sW1wAyhWOH2U5OsDWC9JeeFDvtBMTBvkHyjTjBC+wCXDtF1Kn
5rTQ74chIy2W6ABILaYRtmcQYO9f7ucg1NrYWss3dxETuB4bnBTNIc9F3A8bGp8s/YZeveUvgD/q
pG+yzU84JjdNo1hLztUlThSReKM0N8a901b7ru/gPtc/g5T6NofDeI8Tqxff8MvCSQ2hbPBWc3Y1
GhiG+frn0G3qGphgJ8iO46kN/4W4GmY2Q5NkJOh9FOwOUKv5DCrXDROA5Q5kKURbvpuplYZ9L7H4
I/Fm490jgjFrofIkUd6X6sRssvENE4hLma5fW7LiJfAjk02Uo61eYnzP1ZKfYAIIyMxJb79xWL5F
4XYrFJI4QdsDn8zUzPhCt5WTe225GtFyy8wceEuQOEnzZqPQcG/HSkzIbX63+NYnAnsW3NRp2OnZ
Li9ni1l4CnDIJsdJ9ietzcMdM45lXL3vGkz5uLxeujjhjHKApdnn05eyRAb2MA46EDtH9l4RCBVZ
VD9EEvZRxUWrvUJReyWOv35QSLBZynOrWtvGhyjEoAzNi04OGA313vX6V+nijrXAmXgCFcu+A4P5
wZsFvcJyexeok4lPXFEdHKSyLIbyUPpuM3Edv7mp++xNRKXP3TAiI8rqVOox8yOCyuZeIVStTR0g
n6nTV/CDSBhoNrSU7EgDM7rk4Bo9badBLZbYh/HH0gpkr8OBUSiqMHGMlm0JO1HW3RliLUJmexFp
i9QAhn1ckElxoYiEZ/IGn5YNaVueutDk5riS8Lnhm6dY2WRlXRIUXo0Q5yWKdmQJ8tGDancgxEPR
AkICp6y7+y9gvh94jyQWuxAf4SKAllxYLz4QxSsei8hXvoIHtAvjs71g2mCW+fswk8UNW4kc3jJo
98w+E8pdwZuuk3/qSDMW3qjbiDEZZGpSVg8O4AQuRRKVKVGBl1cUMOk/yOIjGACXv4rh+jz7TbuW
Fl+p65nR4tbrRglT27nE/2rydk7ptSDXe0ZHjreYfx7aPsjrRC1MAUEp+FZ9KTAN4QwduOir9hJv
BssaQn0S2eSuqlZF7UnwKptNSdcQ2tPZ223/JiAvvzlx5+jZI6yECPqpRavVw4umQigxaCIb2VoJ
idvz6M2f25eAEyV0/3rPgcAgKa9e4lh/csX876QBg60t6yOAnuYthiHGLAHpJdPmpJYwNamuyF9C
dHQK2vlgbr18hHOW1H4YC9WnH0b+GFBJXeCDY2Ro/e/IQeI4QsIdFxb4/VwDZB6ABc3lmIg4tShf
yi0bg1CGHigov+7qNGe6yhQrxImz7ExgmWKEqvRMA3ms2sR2AWB+YPsnx+O+A++LU1Pd3GgHp/Ot
OUYbl8JInXcj2E0jE4JsUaiPt2cJbV1uJQFldIVB0R5A7TsDE94Bf6gvsB2CkdmrCJ26vU6zloF3
+0yqte75HyKLRN+HnA5ysRYXTcwWtOeK7AaD/6SC/0HmDT2Pu3GXqaPApg4P9dBBdvkjpmd90SO2
Uc/22lkdQem/IBdniq4DqCfjWIsNHep5uGFNOs7KYbbxsauG1vTWkrAoi0WaAqlpJ0VgQUhKkdIt
N/YIavblfW3NbCCL0fLFqc8JKYV/+FXZC+SSEC79Rrq9cSah5G8nSUdnTQfa6mTf9rZJxKQ2YiGX
BWTH/HEvAK83ZfK7dshyFkaBjKzLOn6VJcnhT9CqYQOgk7qp5hwwTK/ssSlvjknE5c3JKIVnmUS2
kOr4PqY5q0v8AXJHKTHUD5Lb1U3tuo/1RQGNQ08SP+MuUMF8gGOMGyVAvmMYDLQhte/nkRcQ4XFA
/Buc4hVziTGM65CAfjHkjbP86AHmj5AKoLiAaS5a5TdBBQbOfVkAYiOHuelbS0A07IYObd+7uCGp
pK/Uzs7AJuLghS4WWc0sPA3SgVcBnDRL+kBu/Tgty1qffqK7IeLM8VkKnzjDyeILLIZFS1IRqMkO
abymOY5dvvHksU64EdnOc7E7IdNd9yJOzJNKIQW/2cE9JXhGPTg4p98zh05pYsOaRedJrvTTQlUI
Xzskq7h/pHJOXju0ElW4ch8zMdRHw5EY8esCq+VM48mF1FW3kf/ybbBu1LrXah/Trj0JKmCHw2PH
hkwcwn8sGYy2h/o4mR+/ga1CNhSgZmo3uVkvt5qrAjLCFCOEwZyC0jbhrrDxUogWIXz2j7m6Hp6q
Gc5GBpFwgKYXFZjl6YoTcfw751Cd5NJ6tvWUg1bmWPYeLSJP2Ufy/mamq1ZgVXqbntDS6Camwho0
Aghp3H7vCQ8ptKGwgNHuXoDTXaenNaXYxdGzGSEkhWCdhdzf5Th6PS+A9skf8j2weNLMsypyv1un
C+LuAjBhckdMO8WriNKc0UYfGdbYz6xKTduwI1L5DZq799jd5unAIQLSKX3jkftyQkYoud97VnVz
JTW1TIslFfSTS59JXJFePzAdsrZGoUETIP80dHIfQSvo7g5BZ3kesd3bSVqvqwBps2e/vVTtXth6
jgXKGaP4+eTcd4NKTG5MS/1Fj34X3Xf4xsO/SE8IyZIguqR4Y5nLnCaf9v3wJDtgF3qC0BDzxk1i
jRbx8REsmrGQfxYcwTQsjONGSCVAo23+jCvPgbPy45UCWqlxcnLNCUJ1O9N46GTWLHQiq1Mm7XGv
qZ2i2UO8kH+Bg7KEi1tQ+zZlLUGZgu5dqIg2aZ65VmNuZyLHPs/lKrbNg5FtuctAPA2DEiypn9NR
s4xt8hnn14FAY2eHkvRetyd2qQdGB4mvLev5nY71IAp4d+jI9ZHYnGGnp5VjFeRAgPiO2GEVGuAc
J268rLeIiUwyf8uISFaRiPv3BmlNPcxvK5tZ7rnQ1QvpD+tPzpwxv1c6lgHt7me6szkNOVb/D4wd
xm1Cdb/rEF9RNwU3M76T4ykPNMIMmSa1/IPui2fLLm/u9BqcTtoXi2KfyiBNzCdZ8E8KhZ4oEJQm
n+4ti8e9RMletHUfBSkOzRS4PqquNWaURj8UTqUYNhQAEEMTAYPr+phtL0dKfARYuo/WyzjV219D
l9PTFTdUQCYFvRNQHcWCilJa3jYRBQTEPK9lSsA3vA1kAAXwPby8WkT+ymQh5RP+HitmCSBbrCkh
lpoTOrvFTlSqtKaatU/vcglXDXWcrXhjw9vVG9+JZc1YT49qYGmGiBXKxHhCk6hLfx3j+zu0tp+F
ThqELvY60OqP5GBnXgUoHIPq238a/mvlN0p7VZPAi/UJt4AkRcE3xkpBvJqBfPbyxm8z60BJKFwQ
4XDqAy+XGuL+BoAy4QYfgkTEwZ1ufXdIEAhAgJ39sGfog5ePFNx64vFGWNzG8VPYQ8mDQlctAeXy
tdSEd61tJVsCYLiw0K7ZRUIQUKR8rdysUr2tzrfmq/5j/QQfsyuV6bVY/Es8uFYFkxcGHwKwIG3H
RrXAh552Jmj0sn/voYI3gmMx0a2KCBalLvAKkQv0vf/keLRtBV0TBZmq+E5AELiQZaC4HgTbS9Ua
4heaat73D4dOkQ5J4odHPmeug9R7dMH4KeUOrmPMZT6mOPeWal93MiL/pyvIHCQXENHSJ72Se6ki
Apc1VDK8Ii0uZMtfV9gOaYfnfXocAgizu4VsSEejVsCCzl/7vVHgYTV6gJDYuXyFRV8uStpv2/zk
Sa0rU8OZG77KtQdpGTePhgmGx3KWkGB00Vw0ADa1G8W9nwiTnMjjhr/e++CGGS+D1pcBfHaXq/KS
Tmm6bD26jkqU/RAixUij/oEjbksDVhXBB4IbNkbAOqs0zGEXkVGpRPB2Cjgu46rH+UxnBZ9YD4Nt
9KXjTrkr4A70zjvQkYStPxFkZ2aZWCifkps80J4uXyy8d170QXRsRLWbbnXxnbzlVKyHQiXae2jn
qVUPg2l5OT2EbmhtUu1hWH3fC6B6vdQtYdyYB7zFqBWAKWkzIeyrh9Yp8ZVzzXmuX0p5gdsPQJQo
xX7LfHKQFabpBCYDDBnmP6WC65mOf+Eaz00UYuhO6J3OnN4N4kvzGKefu+e3q+yFmq+W3ttYh4ky
6FzaD2FTLPiRKV/IkW7gMKYZs9m0MJwkm5iBwjq/X2nNSd+pMTYFavP+6p01ob9f/p5YnJRF9KCZ
d3v6+0y2xIDJ8YtTvizTOeXFQxui2cr9F7rSQKT0RWNSUsV8rgtuwLHKxL/OMKZF5RxCxKtYW0WC
3SwL7nfUCjCtEx6U7pVx5rXoPUrg8mjHoksncqq0mDkMNFE2c29AlfQaUfGrt+Z+5n0VRpS22piU
lm7Mg+TLUjyqb09cb5GzmfURbkWqou+QJLZxI5Ln8cblHdOSqbJ8buq/XWjUzLmOVUb7dGt7mcqB
92XrFwQx5FQq0p8NO1frLhWjbuf7v64za8xwKkEsLGq6zHXOGxcXYzXxfZgWHd69abZEBEfM5sK0
nAlvdOQ1JP4GFdYYTYWlkEYW0v7C6cGhlTDQ2vDakqEIBZ79ycMnSKAW+Vgg1FDzJNXrTuOrGZhp
5x5OHOegcSjO7f9Glml+vSAIIojaNde6LLVUC6cjif156oNVlkhqdSWOnKuV9IJmvT8FGPFqC116
oOWot6pm54NmCZNfC5q/SLvN8V11gQHssuXzuDzFTViElpYwYGtH6KUPe9ewuAjpTbs05+lWgWFg
HompZ43aujneIjCEyZcV1H90Fwq6JRUDt9h7QwHuTKrqaBzk5I7neTyOMfhW8C4sje7200XifZiz
q0je02NqqsRQNGWlq5rF3xTR9ROen12GKBRWMw3lMXfi5qNU/fLIQcIO0BHLWMsBz+74UZW7durL
3KdZKT5wCxn5qvfU0ihFyCgZp7smXS81XrZsKEp6PA458b8tVRKiDU4LGcm69znupNODYx2Z4/gb
5T9IIW+ybKP2HjbDPO0iFH2PT5R0H0MeOSoCQCBgJvccsh0JnPZjcHFwWmQq+70fiys9uK42zCZ9
VtpTTYxO+AU5Sn6kUEJVN5HpzDlcAwgMt3rElmH0pjiMKiaSB3lGgkKchnW0LGrUgmpxKG+10ii6
p/VChI2u8ZAlow58rPzhLTLnlgUq/FdzDS3Sc5+4xwWsJjmauqgQ9Gpijr30Q/CyoV6cxJOLvSq8
tvk6kmk8P0aGMZlco13PagtrupvhwwM8DIAALeWs/DxhAVLccaj+s1k7IQpQXDG8g3IDYaHj6Gy0
epthXZv/T4VnOJoaODaOUdctiASzyj4q2iwBzr0eDulCXBieWuWG+wwWWzHA+QDAtYdpl0ek+su5
nt8I33Z3cQlaxYWXGvi5D+pKDL9pALCDqTXrR8huRGJZG95iW9BZo+FSqBEDRa0OE9VCvDL8YIFe
d2AwvZS8LhiEPr2U+hMS2/nZt1gol8IgxJZRkt2mgQgWHzGfUX8r20RrFMPlQzErU1Uh8XzGwPxy
f7uZLnZT6Ayrl4fCDte/aa6aqfRe/zf7Cm1znnWMoNHC06MzhnDEpBSMpmgdd6WP/qibz7wOq0ia
oLPN33TgUIhDVWx1a+FLzubEmg1IRXxD35ALNk29L6Gy67KJsJioxiPyywTxFuIx6BixtDZHApsB
KjFZWZlwKSGOhiT2gcHFgJRKu7u6o/Hf2y2jPJTQdnUKwxd2LvYLAdrvoSC1jjnqIFucqhBvVKWA
AFXH+8AGwDIC3RKBIAF7uxwRdyIzh6rTeNzj0gkNVgXyIh5kZ50bKWgNPbRo45Tf8yUR4YgfXUtG
xgGi0Va+PdHeY94V1O0lZD+Mx8gY/X2nVEe1hnseZADYQZpKESlM9Q/BCMWiXNQwu7iDQ798Vqrt
DUFCdyW053jmwBu9NPZZaUtNU+6zI2r5vRiHdbQvsqyBImbZuECm6jSd9OFYzowHtHkNs/OE1emf
yldmUcb/QdrEQsBPMld+X+cUXqX+15f9bF8Z/EPRPuPodwOImSHF7c76KzRIuaZdRfoWuVJLkSYK
xqQfo1yErYIJC9buHQRhZjelz1mcZhtGjrRxW/ZiPOPfLod1Lf89TMDik+uinmAzo4TMC9Pag5iu
MGS1OZbzbmtWiO1vhf6tFlC9si9z5IrTSrMrzQYDuJgZWQJoUU14HYOKrS62CleCjIMHrlKw7mm4
RXwCGIKes3AMr0jIVV15whII5hDQuPaRYuDHELcnjAAfe3ec6kT6RoMBewP8f62i0hxSo3Eoit8M
75+zxPw4ud0vxyMlKkFQVayB02mujzz49h8n5ABeITKg6Iyobx6qK0bhihRpEvsdkxl2bKaOnj+C
mIq8Lpw5NP+GU4TQ5Ktt8uQ3OQInjrcNPD9U4vh4xQSAXcKQSOyOcTphqbXYfOhewdn30WWhIYcr
CCrPbNCr3gj49P6W8U+7jLcx84FbUJq4cQ0WIzn0qlELkq7yYAYrzT8tm0HGS5K5lgzciGUs/PIp
ZZUcgcyJS+25dum7+O5GIaFO0ZO2A91kBZzUTYS1VQ6K9+B7asEj1oHErvar3uTBsk4yNEGfIpUQ
rw7VcaWXIGh/AEAzBUS39OZc1HAyzPhQ0QjrsYruwTFmUbheKtu5XJ6d039KM0aNW9MxLdL2sFrr
brfOp715K7ohwfRmLU57ZiLxrDz3g89QjVGBOGh/PrXatFmU34UE/f7KZLKtDJjNKrBTpvna10nj
b0OR92MvTTidZ3J+olInt6Jz8AhU1H/ZtNCrHXyIM8r780dCI83lEXFDAR54sBzJGOgSz34yRUj+
cSg1WPm2Ygnk+f6IQuG+FC5h1Q6ef5O6gs9IZ5ShlGk9T9bnAb+DJkzyFV0Sx8/CyBYIC1nLLTRn
exCaB4LKSx3Kq5NbnEx5SOMvCiKm0X44+NshkcjXDa1unqQnbmvqs5KK8VEaYB+QLb+pFNU3je8n
J5SU1F9CHAtXKsKJtu+Bce1qXp2+ihYydQkpirgMI/NFkGT1CUxAiKVMCDJcslDeGV9cLBCaD0Wl
x6Dk4Bi/gnph5CkFiaESedImMXCBhL+9SqG9SOxyQ0k0sD2tPJQpWaW5yAPV6MI4ivN1mu5cfg2K
J4brkbPgLZfQp1xUUe9Vfwg/ZGJCDeXVOlHZQS1kJbCw+6TIq2dAbmvTFg5xzl+6UhV8EFhWGKAE
6NmiQFnf0Lv6jauleKDy67JTlabc21+gU5k4Byb9dU/pPBnyE+PHcDVQWOj20Qry21FvqK5QjLwj
H8vFtVZXHduS/Njy+/CHFWq9x/4ewPwQfykNltRJFgDswQpMQXvk870Qr1c9DIYOuUysiEh5hGL9
tchz64Plj8Pq8UJw+qB6ai8suuraxZVFHr3vfBuzRMX8puJ52jmRrud9wQNryJxQf3QWoY+xd4cS
gAIOyHEYagDZzHRQveTM8+TTMcBhHh3lvMSH7iXxJags1qa4pCwkSRkXZvMF8A91HWkF5C21e525
MnkVDNyGN5Z1pyEMDUrLRrD5MbyPZUn/mcfH/aqj0V7INg0zh52Co6Uy3YVn7cfhFCnl8ABq44FP
k8PuRbxWZMfx2uyQulHGoUrg0/g2ml1f6e67f6+AnNBcBCZoNuBEbuPgDEKf47RL2ohl/h64Bq/j
o5PtiL+nlkftf7R2AJVWzGIoM1jPROkkEvkSc4ldAX1G9SRUuU0mu7tbN504e/VdbVUqHORgHJbe
p05FKRiXZSGfn6GtwJKUaIoOaPjVVV7GuakWF/lXDXqBDvR+ndoNXSkPSuFVeF3HhkElaDeqOtyg
d1KfHLRc3Qz9A8HEWG4w1iWoZzFRPK78ZqpxEklDVJkgQwCG0/9zq1JIhRUjyzD5//+RXFplNUhG
IhdPZAtD+kj0yV3RrcLq5DQl4347qcJSb2h1fk6Wwq9Fnuqji2zre73s7EA4s72IM9xm75Qvb6Oi
VdctmXSX5+G919DDITB1oYZmtvBwUSrJFO+0uorDN49tSohwyQJjwYknZlnBcQp1wxpxi9Vhb9lf
wHFvJHLGAUMUL8g17Cb74ar3QG8qZNDRW6SIxhu8IRhq3foqlRbmR9s6zMjPE4f6XIDGfR9R1+/2
w6lHHx9rI9OidquK7JFQeXYCTXn0eD2Gu7afbh4f+E0pm8qJo2JQYZUhlQIZ7Er+tGVH50CjYUkf
izgt9gJU8RQjmoWxiti5YqZqLhcr0abuoCDesJ76oE9GqOx3PazXGdebu1RbvCl8cMg0r8jc0Aaf
wT0Vmko/ey7eFHPdb7F0iJFNy8QwefXFzWdinwhJnfLZOYgFubdGxBnoeWyDWMqHFvnyNHfHFmGj
T/GEGPtaBKPALDgEMG6qJcZdwAZWKRClOX+nJcmzIzKb5MaXYze9AWqqnSqwHczSeaQh719LV98V
JBdsFUH2BkSdhqjxyrcl1OuMynQvYcea561BgOekGoBNGNPSVJJT1TOlhhjrvbev5mKloNkv6KpJ
W2PoE4vC+wNS7pqGpOsIzxN7qy/a/IN1qCe60JiawxOh67Kk6lpgZ90HL5SXPPFqDi/lYesQX8tr
gMWzLRFn8W2xK5QrrLlSame9U3w2/YWGi3gjHSlmq3e2+cL7/A3oSsnQgkzJUV9Oap2KSX3MFYxp
T38BRFbkxghEgJ/Y1bld9o51TV7ZzdXrfPA/S4V6GDLI+BcaloPm1E2XyY6us+K/eflsJkWtKSdB
aMqggVkTjLR5V0h/Uab6M05Nzw7MCtTMbkEbS6BwjTkwnzlj5tH+IkF5ReFrMP8VGdXR5S1NWGKz
GQz5DNDoywONkRBOFUuB0yQhCAJ7XtbwH2qJLU841p8uZsL9w2KqBNE9kvhD3ms8Kd/8pcqAmEJZ
NCoQlUI+fHf315rjZsNihjg0LKoYrllVyz6qxGXckmIQUiOaHq7lZkZgJfJULnuYB2DCZfkuWl99
9UO8tyObTmBDxpivf39dTKhVKASi1uqKMarFmPZKgPo4w9KJtfxHWnwShWL4Dx8VlON011fRMZnR
cLF/ot1e5GZftI10gKDOu8B3uRwPe4Q+sPFFwzah0UTmzCOn9wvC0qjp8Qoq4BtuXGABeYqI8zkG
wrtLYbYp2zFurN+39k3k+whGXdkG3MiO5jLVef2hO97Z9PZ4n2tAUp78Xn7uHZ1sTabL9i+j6+FO
jqm3vg1HWnz8wztsiGn/hDmvzKxgwmky+LpwOKMJoGz0JSIgnyoAbSlOGIdoSaJeKfZSfHgM4C+n
7EssN0oV7D5a81PG2UIJV5r/yuURYwJOTD1xVUXcIkXuKJwFPZUEkf4p+dUibekhQh5zk0tQn/be
gk78xkskcn8H51ayQeMrCYKS96TYpDmT4SnFkTPnhsjO5FckbtHRQw00wwH7z/+g0JLrhuiv2y4A
xWw4A00CwpabS+NeKOyJXF/JmpyXIdPZdeSkNJmJLWJ2FGt1oi+TPb8Dsc0mdNkonBdGWtLJqCDN
bohjtMTNlRVpgLZFylk8p+Dy1gXZD1lMVkhle4JrQyYz6qgsM0xwZfXiknftHLO+8esRo21gRKpE
PbGHuJCR0hwG0qdXv+Vcevj65YtwJxF55FAXy1warILCZN6Q5gpKIjWsRuzE7lxLeMR2mxv9/yBT
N+fMA3eJQ8XQuNdKmR5cKTsqU1bH39ZdSNX0NSZqduKZkNRL4c03r1mozcPeQdxyGqu/ke/Yhptu
xc/1NxYiLZjewoBmguXaiNn7cu7j1vbHVsLjV5Q0N022lBFWWVF1HrylOdulMz1jIftDtYuLDk+f
8Fur95bJZWKy6FatxZuj+Qg4b6TsrIc7mw/7Pvny34ESnT20hN7PHhvaqd4QepkO3MU052zYZSck
+eC2HFl5wMuPPjjjyL7rX21ccp0kAbvgJDeNMHg5CCHyd55B69J1tyYuPrnCXzeXjis/PxNHOk8E
sxst7quy6qfbnWOAePk2mp8zHyIR+jEJW2eTrTWUG/G9W7j3ZC7E7YEEyUQE8waaN8tbOEYviIv9
OavSg4ENz+jlREDZXapAnO6Sw5eTHb72uaVwQlUe1vcacrZqLfNSYXnSWAGmSmi23iSq4ccpgdef
/oLl9cHSYUZeLpST5BeNnt0a42xGMOUmZx4AiC4QblZN75g6Nj5SbZuTMPpYYnMWPhF+GwtsGyG0
72G6WnuI3DhahAR7Lny9nsp3zWqnyS2IM0ETQD88Vi/gtYdmpndF8RLbl0NaFsGcwQV5gVB+J28r
dw9jRw22I3cjdqtPjoqtfOSqAFsddNVgM/yau1+uQBW6CJuRs6MP7N2uXgKGqwOVbkP+1P9eGQ8V
FgHBcuyNPKNIM3e/S52dwbtcZYm872oNbDVLXhEpfzUjQhNzGfQMT5hWeA2qu+2sQEMssWHAHGLZ
HtiSnYILgiz1xFP3wVAzzt/tKaAI+Q3VgMKTYYgT9/+s1EcnBv/GR6STTbjMZeUZ/g+qwV3t0VK7
Tu8VStb7hs9Skhb+KWfW44qnH5y1wg9svUBS6OuWPDkh8xE0E0aY1Gqq1fuHno5YdNSnFe49vaBC
1GTjouq2qpSzOqxbF3eArAqhv+3v+yebWbo/WH0aOxZYHvJuyjngKFKr1Jndbb7M/d0GsU8dkIDd
Gm/UXxdJF1qLaur7RcYYZnWoGEYBg+RF1VpNdusmV+DSSbxllkn29l9mKOxjo5Vbksz7K6eRUQZW
yof4R7u9eItuKYNpFd8wdY3hGUlphu7bzEblF2+1fa135du74e3ybETPwA2sSDLXDtXUnXlBJDwX
8X9bCrdas2ksJ1tiU146TFJLu9plZNs+Z9zMOKcX12o8SUkNq4QfiVSTSVTGejBCMROO1rQcaA9k
t4INpRZ4ho8Qn1d8AmVriYAPSuHYIVzBKeVbDfomQChlPJN3Yy5EuNNvY9spjXlveJXjBl82U4f2
R6d6pkS695l0ZYFjHokprc0+J/0n7Hhq28wBpgUlbwDvQjHBm+KypH6P8At81ZGu9zG4J7Qxe8Nb
wxKRszFrPflT99/mx7NX4YQNw2JJD1s602OizerVh1X1PGisdPm51jhRBjrl7JXXN5Xr7Jvgy2+x
40QZzAsg/gtfB0zwezF4tXC2j454Mzoy++Zd2kRcoeF+rA9qXDw/ffKnBEzr0PO2h1kJd22/gKfc
b55Onpbim9X+xGelQ/xjiuE/zli8mcszVv9qHWuzPyHArCTqHM3dKme40FyVvWBL/GkPA/q0sh8f
Olg2PYuuRsvSj97blOr1ALAzrppekJzIUGkZRKKG6u6m4WKympapGu+cLpmY6wE376VaRdL0Ljbi
PkqLP4tdmXR9+nzwX2CAzHRHGHUdm3i00nAfApZLAdR11LMHFqdSshIkD8kuXEBnF0XVJF7GDN/6
cnt2cFE1nUDEp7IGWHuFl4g2vcu+MCItHHDzzR8oK3waI8XBTrZC6EUPoIiagXLnblvwv8uT/+em
z60EZ9Xm22w4OXnKLAwlHq52+/8uBxkpkGFqi+3ojc8LD7MKvrN7h6PC0uFgTpWxrOBG2GuBJWZM
shFbvYf+XGWZ7TGNhYDqeEwH4Uny5weLuowWkG5CQi1jNQNssv+HZsExHVNp5x3qRdQHOWWkK4rA
FCFI5FQiqlfzN4AxlvmmraSQR69bBbx+6Ch1ElODTQQNKTfXltp7LKd6rQyLnMJ7kEmcyyXiV/vm
520uOh/TxzVEwdUO2Cpti6YWkLTg6x8SCw+vV2LUe8r5gEzv3uYwjPlg5XizBugYJUJO9zS3z/OK
4dZKQEQp3SdhPV9XKjs4x9NOtH1GQXoFS5daa7b7B1UPFjvKbTA3Wc2S7eGS+0u+aXd6kgCPyn7t
s8Od1HLogtW70+Jt/xNyznsh2nmspKZAI99AkvGQwGlg6j21XWEMNz1zmhtNPO80H2n5TF86ydoE
Mj1ly1+nrc7bhGmVmoYye2Vpatrluu87J8IE+UE9JcEO3yy1m6su4IE+4iuDWPG1zwPvPeM6ngp5
pfwDLvheQsD84Pmv9NWMiWbdZBZS8dZ3BnoLo1TPLff38QcdvEmFkva6L2tzUt3h9nur4ykmJeG+
nxX75dt77es9Au4JchL6SUOoEBJo+tEgF+TxBKXt5iGLMzbcKWUyyYqjCK9+udcLqxQPlInyo85r
rA+AF5NUUGYz4lv0vJuimTbRMOcfOFwAvmWTy58YSl8Vf2HcUkS8ZlGxCVIS6Wfmsx8q1itLU3Tf
rN4aK9A1/DaVk8h+0JBFJYCL5HK5HSj2Kh2Taz7U8IETQSw68sxzxmJa5SKd4quM+I3uQwIeL1PD
G7K0WhVf0CvrrZvujQVEqGVIB3Io+zZY7BjdrOUX29mMBrJHVomT4KnmNZerjWzwwSLlHnQq/jKu
tWSrPHai7yfXN7bMOnqTszVKTA6s+0CAw8I66kXt4dff4ZWy49xY2WOtv7vCwK+QpUpEXaM/ldb5
F/ygEOYxQEVy/CsT5n1I75jYzfSuh8sOTOL/lIi/a0hOSBqzyYyCwxq2yh32x+EmABA+oIvrquUd
9TbRT3tniuQMugk0ARmz0pkg2pA7ar4SqJ4iZVQNJ7kfV6UBgCDLgs5uB3eLC6si1M976d4xovZJ
Zex4yBgRKT/xdNa+Ykcjumt5ljojTHB4BH+GzDJ6MnRJ6hS+6PYx5nRPYkdhGkvygGe+Qd7kkOaK
xtkl3/lwpV1wVYRUeEqsK/x7upDN8LFOUmsEyr2Q/7o9zXDtFpCdAVkkxDmWTdajogAyEqICK6ca
9MUyCSu7WlbQvNcQfYa1e1XAlIFjrp6CnH7mUKYXrQxkahZw9Xinm/wrL+a5bRcmBKVkyq6TDHUR
21a030sHg2JdExJe54TOxqxKSs051QoiAr7Z9vsF8PXTZvHDiYPhDo6wd0/L+PKuQsj9QMCdN9jz
HAX8S3oEThyfeJE/FwOq2+JWsax3REHX2hXE3jAPRy8f4UmEiDWwtLlQrMNLA83dZoCDic/rddyT
Xi3Wdp1Vg/S9c1bOgD+h8xlOX67qN3qavzbzqUjFC9N2LEaoZDkTPY8fl+tlVJ/DdIj9nZkSezF3
5v6wR28Xdows+C5l7DZpWak4v/U+/w5PrfcNccB3O8NlWmWGpJgzizPy/kB1aK0axCV6V9dnCOcU
ZuhWlhZhkyOnqEiJOD2CJgslVlolsURjHlmR10SeS3Y2i1/oLZhPn+YB2hrsplAfULuVSnFZLZXu
SQfyqxqsmJ/8E/tFujSUwicOl775EPXOjUPrEm4cdXP7yb9GplVs9QXr11awLarNEjgyqmVCGxQF
jubxRHqePPZMBKz6xs+huj1n87O3fqA36vqyigxGZkCXMqGK3ayXlEVZmOlYf3QUOSmaob9hR5PS
l7K5kz3QW3kp+E+MBiXs96OA4PcBUMkaiPGR0ICQKR2WbezWwkkFKe4jGgiF/vVitnMTueyBvYJj
qKWObX2bzH7J+RZ2AFboun1oNjugnNX0mmcgJoTROntq/2V/FA59Qja8opFFkogAeLTRF0L2Q2nR
4QElXIMnZMvb14jvRES38/tV6KsB0N+Ogt+xAPC2hogpklbeJq4j0Guz5EjTXmrK0ekN/KeMFNEQ
CyJBlCF+tdVAuotObGjCFv8L37gf/XofgL4jnkH+kcKdZGE0Db43iFMkYQkp64N9cbNmmqXqupcp
dwjZCmj7VhJzO5ivNJcTnsjk/oQFEDIxsaW80p69Nev19AGGCzxGwOKmxBysQHGw5ieh/A3XLqcc
b5q+2lQ+OEYWFV2fxdL99GOA00jyyizzecHLsv1FYku+ZhC7+NNlZcxl0hQyiP0f8G9/JVs8wD7j
fDMqUhs/jWXsugfNRQHCiFPBTLBSGx7Zd6QFtpnnxdRb71g0Bg1nnJu4ZUWdJOp+nLRc3V3kyhSE
iY6aT4rINStvmDg4Wp9ddS7F3Yrk9W1FtOvjpL3vd0VnBvQy4rWv8C4+AZwWNuqwY6Y1zQy+psrN
HrGkbv1ChDwWUaNv+wLWRUyW62l1II58U/bmnmpvRIFSSLjVUZ3ZBi9FEdjeNryATAliT4puLcZq
tjy+83uWrjf3GD7kqiE4AGGi3g1x6dtlS+2Cj9mXM7XdchJHreZl7hAbg7piu84PlR66dCERGWzj
68JohmfKZoPmQnzNfCAPAbj5wRGtzXNiE02VZAxqZmOgXe8SqMszcO7r0KoKyOoULyOMmMPlR5ih
OqBfXrWDN81PZ0x2LsuLfNbNY0iSd8lPqiiZ/imkOgeL+FB+P7LipJrnJJNBM1TbCD74Donr5JRe
N8eoyYH2iZOcCoVaqsfOl5ynHm/nG6TyKZ4fhpN9XAdgUfhB+oG04KQrGSy3iwA+1yNZPI/qa0jq
v6km78JBLZj533zK93xrB8tlRNzSk0HPFL83Bltz6zgSKdjEKAHImi0nkRCgzNmDZfOMqkNocqZP
UHjEUtsZG7Exn+4sovcLdnIJSRmrEqDQW6E0IxA3GHKH2EN2yKcViOyIK1StzJ2hbbxRLbQ59a25
zit06tWnR7gfhMmIwqrRzKL/SpdeEum5rt4G8pu7WEpYGasWAXPKvErv6I+ZR9esYXu5s8a4hCj6
Zv1pR0vn3+kZ5K4XDfXTPE/qVkX9xf9O94yqwGFUD56bEf/Szo7GPXBk/+qZmwHRPYGHvU8kZgoa
zBUWgRhr8ZPKuL43mXHHXOwcF4Xa6kV1C84OgyMYXjfQe5/7aFceR4M7k1/XXPlqAAKdBf/wUp2s
RAbaNBliOFbXC37RQ+e4LO0+Gegl0yNqgQco9Ri3IESQA91TEaO+Xxab+iBvDYEBsGAcIZ/WpBw7
yqp/7sKHlzjnX0XdqgrmOK3GBLjT6Mq4LKq3RGODir+EM8ehbbQcYtIi7x1NctdkjOKhVvjculAf
/Bh+HeCokLQb7SxxgToM/J1BYBs0m4XRCs4d5DbcKpNNweknhCLHa8xX2G3iSdYKfZ/UWIcYulcg
bCnfx74Q6+ld7dFEczdSOgZZpCV5VtA3H9c8TycOXsewBMMGaIVToi1mbOEs7Fb/9ybZRV0FJ9xN
4oQLtnIm+q48aLK2JLu20BqBJTf4qxbUv+wl1d3EPS3Mb1TyKDU2W64L5ULmT0c94FTSgNgloFBG
i+NIPx+fmnlX+3VCu3Wqp3mS/2CAw8H2iA9nFD491VMAUTrEx6nyaV94HCTGFrdbj/ClWiQp6ZAX
EZpzto/A8uYyXQLTjcvKqQTmvKPcl+wD9kqf62HgkbH/p+40Zqs9i1VLRFiFT6gcMLSop0HUckl/
lWpdfPLZ+Ep3FgXHeHYXkTNGhMstgxH5vXhsTn58UDgu+YXl8I64cA+ybXgSATQAmYmckcmhUEhW
ssz7J++VglI4hgKOxfz2NNaOH0FHrlKoWDw8ArPJpbKeHSSS9GLO4gZnrx/q5EuzVMy+KlFpVWlL
galg/9gUGDcWTvf+0npzfbOYrnlRpLHE5eY6cSn/u3fFK6W6ky+OqhNp2KQDe4jKZeCnE51y8IiU
4QHOkRs3rgsZRdj9xGa9uXsumWPsgytYVroDhjjLKnVCrMOCbaGKBBxztv8gwtwPzlYCXc0Kdyio
2Lpdbrva7t3sfIjfUegMvE52GLLMi8JH5LnIFWuQP09GsSPop6BIbloJ+4ERcJnCOEcfxBbQnZEE
dZinm2nMz5/HjYpA0zSMLqyILq3FsxIQSCnIv1ddMGxmWjfN6gKElrNJI88fxZ/FRPsgm3KoQl/D
SRD7W/V/+b5uWV50U5QMAyYKank6YcJ+HbibH4x4Kb62M3XGCAV7DIM6lIpAs34boj7flbwZd39J
mSlvKC0dzO4q30+jWdQRnCaMFxEeLOBsIChAsldTBjmuEr513aIrng6AH0/gA7XTm9Qw0ft+e93D
Eou/B+iDvuPoXj0BQ6CuePxCmiB5m1Z4T1GFqgty+JMMA4UFx7Jx7SL2N83mY4221ApinATxEV7O
OYD/ixQ07dBaqPXXWeKdcAzMGQfX7DMsVlZ6ExZIMnBETfF280pGNoPjqoRVIY/FV5O5OW6UvFGl
jjxtAHjefrtCOZQ3qaFn0otOWSiHZ2ewbkKBda+CW1IrwMQD36WlXLafM9I9YsPSnML/yKbXrVLf
aFHW+ZW9935F+ML4zFi3fiKp2MKHDOvJXgKGgrQbTlKVEsthZxyiqidgAV1wMPBgR9D95kx61kLl
Mq5NifClrOpS9f1FaOG1pJe5bcMCJuHAXla7KIDJQmAjPzP1kp+8bQwcTF8bK68xQQq7tWdznkRo
QfdqNGEcwplvq+19JzIUwBcBMjinUfvjPwce6KPTRkiebMRA0PTQcswYNPZIcZmGGxTzKVw651ne
fPeqjnKbw5Bs5zqRw8QM4W63hLNyqQkMdaegNizsiUDTvWfj3Q2KCxi3DDfNv3BxFVZXkVj6cTCG
M490t0d2PuZG8j7cwxBXScpOWrTDml+LKRhposMXFG2Hd+pBU/z+KPeJ7d3TpHTno68fEshaAbjX
F1h5qz568shIRJ0EK7cT/1qNfcyHrwqXBVyHtjhU8fFx0RTxUHPbX2isTmIx7zR6n73a1iwF5c/i
7Jg9EL4OJb50aKVcx1PU8SmK6uKW06shYeGkORvBgTel094/TqSmzo6jyq7iSmxg0Y37dzjMRL8+
2ahemrcK16DkMyivwW5XMrU9w746KM3oqpRIdrdZ9MDMiW3aiCYi8ya0mtra5oSa3wNUUzaBX9o9
Xz6oJ0+N1z8tHVMwRsXhb41nD7qkomt+U0fSvaSIafXOIie8r1b95FSXjVE8xKbK2g71bsKxlChw
rVIfCTtxsAcclNWnXcyEox/YsJyXPb9CJ7KA9RlclqKZJVGgdBUR1NE885rBJqyh615exue5tKQg
Wj14uzdOwoCHx4QjULLtCARlFjyVn+rn0BQNcOEtYanNfQD4yxAdaY/nASOiIgoS+39+5PCIsbBA
i4r/i1ngUo8bbuF53O8vPN6JAcuZf3TBCw8dNT403IQqPsptp8MciyC90gqBcOYKOcLQzIZwTtKJ
cXAF+ilNPCK1ZWIVAS1CWojNE1EZCeySruU/ZyIbIBo2p2N8tpxIHWfyI1Rq78ajnCQYnAFt/wL0
UkSLfFf6eXaMO1ZOBLThNmajbbm9fdaT/PBfCUJsGPE0Mr6Q741CMMOqO7e0qpEbDValRucGyAEu
qge+8q11GfvGBz8Qrrv5FvNCF1jZJ18/bhnMBCgYZJ0vezXcEtAue+VvrGefD3aMDNtyEdz4WEsX
h269GkOKqvrBQBPKw3N5+bhC88MEu8pPuhdE6Jy5TzGY1ukPFdZSRYgbCTaWPsydq0mVTPPTIYpw
kxmsYUEMsX20RETAKW+Mcw+m3G8rDtGA+NG4kXjCmkIV0fVkpB0VsYjJZ8cedV81fyJvrD0POgxu
38EVmSmwg92FIy4zwlpsFUw511S6wwS6oOAb+Lj1gqiQFP+HQ+F+LTowxiLsSlId+fdGSYn0JCCS
axB2k6wWnPZdvonnZjPpnm5RCGxMem9X9lc75yYslmwJDxYERLBIdjOCPwqtfaGxnFV/Y8ERu+8S
Y8VBT10pZts4NtCMRtaOKWqo5g/IHUARXxvqqJPy0dvv+k7J56IHSr0vittFvbMrNsEqfEiscONS
HwuurNevBAWrpmePKumO67swRASj4ON5GlxthxNFOb1ZFpQnuOKSKi4i/Ol6CUtSVyKUqSIdHBmS
me1+7IRqRB+wwDdYvsziidNnXS63xmo/9oxJ4jQLrVVscLlQiT/yw7h21vK+SaTeMSRG/0eUYhXv
ffAN44dkP1iIRuQ9IhVI5bqKwSufSSXE4GhiGgg4PNd2dWMXBtqDCxsEqEcxdjNafb3qyrK/il/5
MOGase3kwM4lUUAzl/P+jhrQsSS7lYjgCjZmvCHJGPlAF+D86lBF1oGDkFvHGEXFQrE+hynJ74gw
6n7FnYHZu6UH5RsexA4LlQT6wH98q3O1O11a2AMqrz6bH6W5x1KcnUhVna2l7vWUN6tZfN/pnuAm
clqoSopwKY/b0PgMA/GXd9sZsRI5CBPmf6QgvGBZHJixl9EPo22RwE92frurC+w9UIcqhyVGSOEd
TVPXlxOqWDCAnbNQc4+eQCJXaUs79H74WVmeomhcx7Q++jUEYCbWXAjFALFqVn0RD1dxYcuzL6G+
IM0j0Ypz+7wAnR7ZshsbKy7IsHzFgHTM3/syRm2fjoWIvTkglKS1AOktoM+0YvdYrpQf99I5Auqv
Q6ERYK5Ahl4X91F15riqtJyjl69fPIqpRaDeS2Q8BfI00j+Pn+IzwdG6umdS5Wyny4FcQsUX1wi7
dwgg0EXoP51O9QQ+1NQeQqUknN1gycsIh90j524s7ho/qTYIfHBeToZt/+3Dz3fvXxxgEb1+xztn
135TGIkNHUfBpjPdW5z/dbPY4c8F4QHJdz0fXm7Lqgvm4yP/SzsyZ8oAWtzq0+3qt2mKoDYSaVnN
wzZ2furVo5cxmbXT3STWTNnkHiDsobUdhLPoiL+hoFPX+MXRtHh60N1Uy4I02dHmAcXW85qf4J5t
dGbr4J3BSRN72C39XIRQPwhNS1kLpYYIw2L/TekWVFILUGjHtICk/B+jPbJEX5pFcVgR38G91s/s
9cadYKZkL6WmtBSd/4+CcIP/t9swwcISXhkDE5acj4rPQkgVtcDl9pOBongtRLiAXECedi5ppLXr
Y7a8FB5U8wq5L3IGssYu9J7hzrjYPqosFo6UllC31hBrq5uoSngtj/dB8VVMFQ7xyC+VCF9w7CRd
qHjE+FZHV0yRry1RZSmSTXMRn8S2JAb86WGWb0xMwYrL6snpw31f5cwgenzXwct/TBu7oo23JE7w
ReGt9hjskqKYigXThHJoJ3y6m5z5II3JtNtC9MKbCqpG1Podkm73m1QFHpjk4Go9Vip8aILxx/r+
9ewT1WTqWzGyxoMDnBQpuKQpjwXa0ZiGxxzJS636CBd8k8cZ0/9F/SYkGzb9ogXzcsQF9IdN+KAT
PZAF7srmlVv1ogm81E80M9u5ncnb0UwSJbca/HxqT9JR/pSUjSBeSqLQXDaLYaTEkLmIwPCFBiQH
s5AdF15HI7AbTSHlzADqsMiO8fkulrRUrpBi8C8k/i7lHhhzhn+HK7ymyL95FuZBUzyoaVgSeFJV
EcQFxoqz2oiYgZGD7bB7BHICid9JwS88R99KP+5dZyTUNEucqXXCHlC28FdcQJmQBTigdNfAQar+
RH3xnArVo8mDpLJomGn3l3MHUnaoSJdiaPIarZq0pdiuSlbyB0aGULyXkDpCk/uanmZkkF4WUcJA
S2EF+TetSWmOzu9rXDuT01BeRGS9nvd1q/VmXrZQDoaQ8MVfaUmTcyATeo1mxOd8jgDgU6qgi+g9
fLgtosS62FqNkauEVsHzuuAqHTKaFfzIRrCRbYjXIY7pRP6x1VXwvnLln8MYXr3SCZDVYq3yhUvF
zpP0E8jKTu4LJEvDBjIlogWPUXqrYP2jTDXRpKmmAsvoBv1UpGUSV58+o5vCiQxhsQr6pDhP19yf
lZDS2Vkq39bJ5rTVcd4uxJqwIazTVrRAz7yGWOkvobUhZcFzR4iLoRccS8mJwJU4dVka5CuhLuTI
j746BiLPqGNOTyQrplJ0VJfVI7Zk7phqJfwcs8PahZy8l5jKTrWpwi7yRAHQlvWbrGESSw8e+Z1z
OpnvNHuD+duQKG5HErb+mfezDGTh5362zZju1wB64Oa0NyWYifkhThzRXPBkLR90Hlh5AFbXZl9l
bpnf3LhrLOSSl7KLwuS1LtlW2/l+xR81bpEahDMVq9lXuQRAbhc1IVgkSt+T8BgNkjXGjS/59yhZ
7CICdMCQFZSjSXkBF3w0iJ5UTeWD+GgDac05Xokn4g8TDO3RCq47g0fzVhLU9wdjC4k45bzr24UN
HJAcqJImculSeTs2u++/THIyUiK2U6j3GXROGA1aYvcHlBwQW8umbguQEjUDtn9ZqUdYwMVIBwu6
eRp/7YosK8CmUp9krQQK2fXFXE8GPpb2pgcUwRld0UnXeZU/DiHh/+1KyL+I3vZyqXh5TrCa+KXk
b+Zyexh1GyV4fnt1FD9yf3PRfjGGHHW+469RSdM/yUnPMh902S8ffrXakJBD2y16DssRvuGTAliZ
JTYrtwokT+WY6OJF/h/myZ5fPo8BC9EvZ/16PQM3w3WNVz7oxduACA9uE50AuHc+abYi4ivlooQb
vdZ8hr0rYQf7TrnsWhUwZkdVCCtJCQFYuDNsfCd0tW9eRG5RkjHoDj9mgjLhar/a91MJAw4Ovrt4
VyYoY2fa49vUMk9T7kTFqHlgYq/ZAs8sSWhu1tNmyxMoSs5TJZkh37c6nbVWSHpqEdC+q19tfv4Q
sQKq2ssh1Y9ry3OKt+bAouXO6gZcmrzsbuigeTDo12altTs+pb28UC6xmhtTUyfKT0RgBw8pp/QP
ihGegDPoFmEppb4y1gnHvkWoesbf6IU7WgxPZooamafClO37GjVjR1XUBdJKN/fG3fOqBdKEvibX
R0x1Y5MK7kk61HhdHPzNVVE7OtOfOiCp+ozg8YUTRgEncCylqlMoTd1Y1pwns9m0q2nWiNbJGnYR
78wtID1fmHeRk8492LyuJOeViIcPd4oa0NKJE6P6TCAbPrX3E9TCKzjkEPMKo/N9QolG38owlgpX
rLDaXLQesP0klrr5fEYdtvWklm16PTquXdN1m1LOWPMkTPmizqbaE9YRH4wPBnA8Ce8aVg2NmKpK
JGWvL3QNLnCbZ1OsjSII94i1nB6IHXWy7fTZ7KtlIwSBJwufAzg0LuibqO+3IZnhi2GlUH9M/PcG
v9kcKlAO0CwnO33LdqLqfNf6vvn4de8CEuppP6NT0syT/BR4SUB6qEMuAuptNyiv/TPkXmGyqL6b
K+R+/vWayE+ETnK5ECwBVDteID+VzE6vlLHbS0FDvedCffS+qK3pyP7/fcrGjsrUi1pxeMlek8X2
1Vs8FEG/Ty9q9Bfl5L3NyObvejx8Sjp6LBhOXuX263kDYaAq/9o4OyNy1Z0MXJAH5p6NCFKnhweo
Pv7YDA9BMTs9NGdqCvRYsdv/LA4B7HPxKYRxjHWAJ/azWNVO+Tg9cmzcR9RpYYIDqrlVrVZ/ptx7
F28xPmXbiCAVdf1r/PozBpdbKg+PjUsVjCOEUTiGv146J/EqJ9CpFNn7DV/YUkNIkwXcP0ROaV9G
T2/rIn5SMT4l2BtLLJmILQ/23NHoGKI7NnOiGFjfdnw/c+Xukxi1ONYaaht7LkgqePD+ohBwMOMf
zm8MZ56LofcEqeRLdjvwHaKKoWfYDlfPnb0E7cEBYCspNWp9fduz1pyZX5t73TQ86tEaUJ+ghSF8
xJHDGMyZLGThlnYXIgwBCiBY5ZowVNlWNyjifNL9bJiZOw3eXxptTrtnj8EJNUNRjvCu97CY44m5
fhijISi5Vkm0aBstiNNO+37BbJQWPcCK37MOBbUgHhjPFDhROAtlRF+XCz1WNuOHl6UFmBfR2EGf
pjyIAIyr0E1z02WjzVs6wc/XhyE6VdQZMVG2nOIVPuNqAGY5bcBEFua/fL3pZTOcLp+GiQgqvqzT
6F+BzpR1hmdsrMLFE4vxv9WKUhqXi7d5dXZj3KZeliZ3LplU3oMVaOgRUTdjk5QJxh5EzFdIrJZh
Z7bmGKTBWmGlpRVrKwmzxJxyLGVzUb4jiuOmiE7lwSEd26QMwU3RMjPP7tEoIoGQ1ilRhAFuSkv3
R7yspyoyWFB+9QR7Qt698HUw7CRcYmvt6x3YiBreYq0pGJFJDLJ4n6WbwisBkK/RCkyZpazr03x5
1MMI5V/OUcFQjvJODFhRrh8MBR0asKo1Ef8UpH22eyW/FV9iT/eWe6SAMwuR6EUWQo5uCSlKeZTS
U+YK1Bm2cjaOnXsotQhwvjNWEJ3OPs8dSmqMhUOnfaPVtXhvUt8YSSnvTnTcZZncah/HncYxMlkK
WnFsUMv64I0endfDklfKnhxPzQ6f3aMzDhskzKynYdXMJ73xeiphhD+ItvvXFZGvlfA6n24MoWTR
LlY/ZNkx7zFSuT0XZF4QpcNbOvghsXcCUIDT3yqT8NRnoNn6Niq6PrICDWmfuP5c2bX05ZG4m0dt
5WtrIlCW5WsWYV+Yz8lGOpgJi3qR0yeklpNXqz2dFDgfC2TbUFBMAQbUqzTeooGDOFE1perLJi6W
cAg/y8hig4vXJW7iM0xWmQWrBg0Nn8KWsF0nuglj+RfqzHVw5KtNlbOZnTxry5F/zCkcuXp4ZdEq
OKR/BSOUc1zt9p1HeRYHZF1BF9hrFjztJIjmlib2iBNnsVtK3eEZOmO4+BM9Hc1MdiZjQpyHYrp1
2T+Jy3T15Sgb+I04tSpwFn2DTTcw/Dq+lCroXaGrxTgrzdrdnmNQ768xEiDPDHd/gVIU9Y1CnyG1
e2cwmKE51HDICsudOAgwgT2woIM/qtjOW/7pdc7ACxUo9G/h5R9J3h4m22mn0LFHK+SSiJhHJosO
lrSRD5fSicO9t1eoTDTCmvaPM5hu+PwFkT3oAmOK4dcmhUNwk3LxIJc8nnB+K83h/KX4Hjr8P9DA
LKgtuirH3esWkS0xb8lqIi8gXYC4oCqDknS1vHTuBdS8uq2paHYo5pAawJJzHWQcnE9Qaz/jDooN
6UNaESrd4XTMnUYKsFkoiJeA/Kb/CZE9izqL+uGFJyXel6HvtliK2+u44XeWXEaKLULn9InY6trq
plpDBO/94M83wiNLBzANkAUQrgCdjVI4sukUInjjITnENQ0goPTwZtQnJw5gmYLpiFbimrWcQ7Ln
Q7VUX36ahd9t4NEWgEI/pZV8jqoXtbmhc9amMy54MNIh2MFypRDO21D72mw75YmeBPfGlPfHGTzQ
GwEENSsKtVvhnk1gT6QAQNYN7NVH1kzsTt16DxyFxQCXU1RR/BmS6DalUpolvdUB4MAB3Is9KMBM
Dosf+mcCSi1sBcP4/taO4AyPV33jnIBKbMuqX+HtY4ZGambz6P6CUAN7h1aFF9U+XpVKEG16Icta
PKqsCUO6iaMTBrt4RzZBuY2j1SaL3clehgxK1K3clN+YAZIC8iiI+5wFuV4Hy+mvZF5a29wsS5Xu
ArGa+5E/4Zrmpk05FEJ9qfiQOB1fUCDgjIp3ycW+pg/4iOH1tEH8XgxHS5/zvW16zsCNVC3jkKtT
kBLRIT9HSslHzgXjQlPnMEXVFuPTqii2sbmxMfneEkgZe+Jr2PFSSq/qSppL5Rn6tSPhzStxJ2OF
kq7prPz0cl+t1O8Nv2lfcJFviouWYXRAfYGA9/a1ozdFd/rfzCJTh72TCHGZACW4DtDg6wquHj2/
iEic+YaiOOKqmd5oZm7Xey2oPS6bqw0IyNjLS2Y7owJTUWzCizZq6temeRuN7YONxAg3x/EH6pG5
vtr/Evjt8xkm7I8l6nFQZEt9UI0npPgC3JCpJRvgwEEnL26B7ea18+8iC3lUl7QPw9EOnmkRcyQa
eMst6Y5XJ2CFI2ULLcdgs2PyLVK3xFsnHcE1dxSkSVUDoBsuAHmNwcEOUx39kANFDGtYH1fLxF79
igZdhm+LYzzk9O0+s6fTEsTkCPIDeg35OW+L6DS2asA6Nws9Jxozrc+yRO5BHoIxCnsJOKMRFKup
XSgqKe2H5rbyRB0dEFBKftYJp8/x96qzjzFlQlkjcGcZyq6Kc+8u+LWE3MYUTSCoI8R2b2CcMLqT
EkxW26f1Zr7eAvjqvLFgD6k9fLP+NnWd/h+15KNdkKMI5TIKTMmYHZggYVY8pCKNwsfHPxibYyUt
EV1f1ILTQ5E6G3JHmqDnNti348POTg8eFLZYiv04DynYr28jtvPT6k9eH3ym/5vn1S7tYXu2e9xm
hBzUrehZOfKFywKP54ztIvCwpCUsFnAno+zKRHMQHzt78ZxI21j92fjS4rAgHU//3PREiYEtpYPb
GUXCPjIPdZaf1qMkmWZpsycomkgK8Z0zkJWdfZzU1erXY7V8HlTq5l9yxs3oKBXDox2IgBT2HN99
IcDDzXvQPsjxggBE7J1hfOKtDu06il8Qbaoj6lCZFjFe0GVmnEJ0U6TFat02m6h+Tuo1rpb8m8Rd
got/Lp//znZxUFKRiXgG3zbGG+xFcL5vjgxuP7CqAjAysjDGjr0GR4RNYR5SNJX31I3YQ2UKapvS
wZhowq7TEEDWDk9vPQouWOnOWXi0KkgxmaHFqQwNUoPvDPhOP/GGTv5rigb7exrq9vfhPuxY3Fef
XFqH6H+64HqF/olq+FNwNseAFBivU6GWBeQY3FXvULcxZlY8ecCWUzIq8ouUUyLrgxTuzzE/mfZ9
HC/NeqeMIC6qs4pW7YcSAP6yI+5ByxeWNryMMfJKQ97hUQrQefDfBsfgTKygmu0ceDw34YhgiYNz
ucLI4FrshoY4PyKvWr6OCWE6LZmv7SCDllZXNc9ZLiDqZZAYxOSJhFWzSMn7b5cqjUtnC0Y7cnrQ
/kY1yy7L8Q6g0lO7Pwy7XbOV6W9fSoX9U62WYIXsJFQCkuLzjozYzCyfJ4UooCM6ssDtIUF8X+pd
TnCvUOuEh8PZmGwkRTfEkzUrn3iG90FQwAzfQGUL/316w9rbmImZzmt1cJCWbNRvTsbZ+VUHhw0Z
nTtSgLUkOUWpXjVpWGWiS/xPLAfxLZAQJic7NayRMx0r/UnGRihk3vjOrWSF4wUGDwCZaFO+PYXm
/hEiF4qOvheVL2niN8/9pZQmoV1uuOrxqf87m+vbdaHsc4mjOyxvDr5RCsJCQDgo7NtLHS3fxx+r
42TUUvrRvpkDyFGhct9yNaVmkfc9gRHPqDsARF6g63XzSMHJk5gT8CceKdalNJXFmH+Ve2rbVFe9
QpNMNvnsH6k4eNi10jTGZd3E4SnYmEu7QK3bWYL0qBYT3m2E7603nga73RshJHwPww5u4Td52VMv
s0oo8w/6aK4pac38PfjyCcs4BAYY2CglfoBb2V/8DrmaQyGopjvB887d9hXHxH0KPCVkZ3KOCs+R
cI02QYIG4pF6WrMLGFqp4jaUVJptuCYRR22ICLXpGCM4kJpQcz1C6dNb7m768i0H/Ffg/Dp0VpTe
Es9MvAER2yyk4v4WpE3WEZgzOHG6uUv/MCce1b8CEif54mKlbSdby73xmlx/VkGQE5lDJ7HdUmpQ
ozrzsKcyhYDRMMba3M7/lBik+tDubkTWlyh0cWaIMEgsILFO3MI6/bZwsXUGn1SyRhDoU9wx/dWd
wxzPSTO6BiDEyscRrqyO6SLvNcRNkPlNRdOf4yQ4HTmY3ee+K53KIWKKZY6bkE+JXlMctVEmp1MR
us1iHqP6JPanomvRB8cr7mTpEJ2J1LNt7B1Wbwf4VijAbYplUZ9OktezB0dkU7YNO4vcXczjXAs3
6xPkoRmeqq831kfRNPiyiCt7zEX5cyV7jyStuA7jfBis1v5ZVsK6k30QUFsT69d2efpLAB9a6FgP
BMxJR6DrqoVq5yv364taquM6b6hQM/vFs+8rOIxZQ9SkSbyujMzFoVuHk6ho2rCddGA+Nkpb79Qo
gAx43Gnzg2CM6/HN3cUA/bDsIcxxa2OdFnpAPDyYwcxtdV+OYb8fdGKLrlFEhNm5NSUvpvZnWn1o
osySgAV5Op3KFeGnyN+goxWMSjbqPA1N9sjfU1xVU1iyj1gEvXe0fwQNLRsNp78UmvXAW1ZGHQVW
YNF+yZdBM8wCdRTVlOHeqUDNbRswK+Ty/urNk7IWOkZUI9czWms4r63RF2q5ncP8eNV0yY9i9hgk
P+IPiPytIP2HHtLYoHXfNBGKdPy4LVA7rC6axNi+z2kwRr0+lhDzMGIizpeN5wnigDI+O4WdJoTg
HYPoTewSuzQYLlsWQaDsWhN8RIgUiv7mgUpTBaGNGYhdyBtFzU0pgd006qQ2sNBCbsE4WWx24eCn
UfrH2Xb8rv9iyppCPIpG9y0Ec2LTemwOfkOOP5mOUVqtEnvIAURdYxVJaGycdKAsZQKFwnZzEE0y
BE9wfl5P2iarzVSNkXydHVwnbm72IDy6yOD1bcJ225+lxgjKWWpIM7/Qc9uhyyzF8xlHWlT1QUPp
Yhs+0+B2p0mhyUnrb5hI7wUHspg1vl4YjM0mqjazjiw2qAf+ymfuvSEFXsr9pUfhRd83kmCEU3yU
IzE3vYCXalqXOWZvy9Ex5yAeJ1v74nuoKom0NH01q7h+7EIxl+BurxrEaF46gLg4Xezx7QV8Ax3M
HTL4z+our0H1tHMiIjog27uPPdwHrjY2+nmVMwCnnPOw/5SeSpHzbAN1YuafBu2Fot4GQ4yEUpyx
sn9I43VGQGH/Wg6UsChOBFkkuCVH9xdD4hVSsPDzf8yrw8ZJ4rAdJYGBQKHe5tZh9zZhZsTiP77v
NfR9B4r8YR+bJ2Qn4hTKNOueOPtQ0dtTAnPsntJs6aFtIPMvPgnLPhJXEXUPYE3/kVdbj/hkNA6U
jguphBBbPzERAVcLGuZhxwgu+VOx7+lfvyRtc3D9t40MzkKgItUCc2MoXsK9lK2VkgkV5Ujgr7RL
gNyj7PV+OekZ73uuEqxUBGXAJeo7UEm0Td7QHZhEGtrJoRrMKu5TrrLHVc25+ZVyQkdWkrXG6Cr4
/xRLLZVtVhax64B/pEUaLAk7ymBPwbdhZfIDDnMHTR0LU63uoSi4npsscUa0aONW0xhxNHAWg106
QOuIzOvbf+AMo58ujw04MU696YO3ZvxbrCDAHrcivRfze5hHLrhMoQRMPq5b7bAMQuJWbDK3lPXk
VMS/uWXpyndQqmzKDyn6grvEq6SpkYgoOkMqn+Y17O2U7MAbPGZK8C7gqET5vzmhaHIXBN/xKOMW
5BYJ7lQBquZiZoy02qSNTglYN+TuNDzDtkCDweD85tw1NE2TaAb7oj+VZ1+knwNUN1cH+ldY1LzM
p/nuSDxNtA+BNZYaKhnCE/och9tJg7yl3F3umf6vOi11yl0BgegxnOvmt26/Kj3QJufGGXab8uye
XIfeG41NXiVQTv3XPDvS/3LFQr7pJtBqJTpNJR1F56+/4ny3NtBnUbDsbdcpEQuv6koB7FYV34E3
nQE+97o+j/0f2VDp0RPKFT6Kgmwg8rtLRBg48wVpBhaY+YEuF4mjQpg6TvtojX+iBTE8FAHGZDrb
PYuqaQERHuLyFw2clQuB/4D7oeHlRPcDp4m7GIMmwQSVWpMSZzH3k7leZqTFNGBrEB8q81lIZj4f
NH5CImmLK2fQYj5nzCzvwOATcbwBaqYm1xHcvOq4R4KUcDeVowd5aAfzezOpENpYfkl1eeRZgp2R
JsLiOiDwtZaCYvVdLPx7SF2t0jZL7+1ATFj3YRmc9Z5Nx/aIXjvSJ3duAOGjbT0DUZXJgdovBqSa
ala7ICdrgf3EtnNAO7sH4MSHwszgU2NmmT4O3bqviNBmh8ZMQCEBF34K3FZgBFKpxxtuPU2e0fU1
DRYpqoGYa7MMzoFEz05hiwhwpax6YMxa5Z95RvwFVudqr84mbOoaa+ty46ESx405aIXj5Qvt6pQc
qaoc2hM1DOqNKNAsOLC3rG5e9gNZm0DJOH8ZOVBnFwxY+CQ6CBXzE9sfU51pQOXVyE4mvL/Mkh1q
Tw0WpRlL1qdor46YGQAMkrEUqYemK0wnAF4r4P0HNE4eeJQZ4m5K2TzGcFp4huyU8WVQhaC7L+zi
wb/i+nTot7MhRYeWuEpijbCMmegP7GLOaVy17M3qdlOQSE8Ln81H7IVn2hGyFNImzHo60T/wbmS1
jC5HghZUl3GKR0F3R1lttDBTl7qMwQ+K77etfU+EQpYnEe6/y9UAHMP/0aXqUm21geQ8cAdryMY1
5LYJBaKkMN3i+AWXI39fi9iGotffizCEc2B78c9VC2U8s5SPTLh6uIQmXs0dv7Thdo7CzbcnLcST
w09MiFXDepEseMbBIZR9Ff2TcyF/a4MeCkkd3B/WkFe/ybYpvIvU7q4h6wE20Vms/b36yXo5GXDg
Ba9AIbljTgB+8L79gY5/LtCiWlaVjhiWz57NWhSv4rsUWOc2l0VFvnROcI6siN8dM2N9IoFdOuGu
eij9UHuxEmb2r1qH4mRjQnA84Rkz9E3vy5BqH9UQfzM2weJIrRdKWcvnfw4o5rF+jR/2USdjIqcQ
lHUUpeTlWnQ+pOOR/kaQe9kCsl3v4mHbKpidW9dYB73dkW023r3WG0LDFLvGNarjPFVjGn1Q8xjF
8DTLuxJTDQNyhR5jnVSpY5XagF8+ZTVsIABRp2FYC5jeOHD1iDJ0oSoBtiD/vQPbSW4v+HPB/CXy
EDBEHAMeQL/AweUbOPAIgrBY1TzN0t+xKV1cXwpETncNUUqFE3I7T4RHP6z1yzd2ff9Ni1A+uler
YugjCZi0n1vgIJeRjdoUogtPzBvpWXoNTPVofm5OQZDOiJnpcYUsr+f8BRQB1yQgGS5P7tDyQrSz
Z0ptIoqzJ+fohK6yTFlRYrE1+tU4qmaPAiiwlmm0UywpMOp+LgtmiTHYmzlaaRyEGmuGotvhUhyT
gvN5qbYNdZa0c3aH8iTIpzpEMelWjBZxeCekJE25/eOk8yIRt6ls8WzxAwIufwtka+Tyw7jICn2J
wp02WrAkAohGalBtW+nS3gydKhM2qJp3loQgXV+zFdlyxE/mC3+87IXcT5kyQ9Xwbp+04VPshIRf
zicEdw2iPgiOOl8hCAlOwhOXwaY8jqUJZt/UhYvK5zDmDxhb/a0oaY7sbhWoSvuSdDD5sjUmv5od
K+TS8ZNEH1BcMul1pbfv2IZIr+rYPbSKwQphKRA1yOYnMHonUEDqUeVKXBZWP598TfpQt0nzxQaq
ML9n1Rmt9FDtVX3+yrh89iW3uXFUWoRLDvmcCVBGvZQb7Dnvq6XGj0Z7Ml/zgWN06z3K8ybCtysE
jrPqcb2fHa7EMIN/ZmNiJL5xFLG27oufdNjjF7b029UPDo0XII7SivENIeL+4qsjpY4DLsKGKhr3
FU9p4sRG8d0nKR7fSHvwJ/yO/lfpc8CVtwPL1VswodJrt529iBx97OzMA/tA2tRWx3/MqGpY9Vjz
wrwIosQuuZMbn7jLD6XaireZpaneds3ekgja33sofxfO8FAKRxFYPDUbfKsJ6uD0D38zZ8Q9SBW2
EEyAPt/IQVwNPEeMCOWc2JglYRKPkaLxh8NfiyBQi64oQdKE+/WENE2B4NtrTKeS9bJVbzj+hyAd
Zt5lN+YC91ynGTMH69XVWwGZK/wD8rZBPxnL/jhorMi5Okrbm0F2OWYuEkykxcC0SIGqPqD+K0JA
R9w/OMFnJoxlkkSPmUV3J4hDbGuCeWe6hTFV+U9GXQCwMymkacMWUMCjBXt59CIpBFB8BwCNP350
7DGnNHY5mhufJiFvvlS8BjFXdUBZbJU1cIVbBOO0kyMbl6thR6T+VRIp3IpY+jr0Tux5ucjzgY4Z
qbDxgSuqDR2UAfzKssEqDVJgcoheP7CmmuNFp6tC7EO9sNexZqeLRVMJN1Nkd67XPy+juCriujQh
fRWuSylTObESNUVXEHx0FWbK6HXg67lBZImektM/yxIjkDhOYT0N022X4dlYCTyzTxf2ir6pHo32
rl5lzRQDjFORv/b8Ij5YG+scmRNetpQmdyG2wVFk9mp1eCHRuWHmpiQwexKbz3HLeurp9CtbzAkc
fSaQXjNUvI3UljBfE+RYOqvOSIOVKestXF/bKLCIyqf0DV05uWk+UXGj2+loi33x1uaGhJbwlu/1
ZURanuFqGwTmGq0asy3c6UhuwJLxrq2SdlMhdhsnMIyN4YpFdzq4a3CwKRwxZISSBdog8ytDnL8Z
DwcG0N89lZY+q7qJygBnmxTEIaYvAiWMDXT9NKm+P3FF82vQyO6t02oNUXQJRa11hKdBGCUO97HC
xP4YXX19301KyCfh04Ngdyq/3XzsFFDwKTKb+1BTRoc/yNE1YpPyVeNn3P3RSd8FVTTp1XPF8mwR
e43sFL0sLFwV8wMtiCNSC5ND4Ng1fc1zkmw7+7GNbAn1MZ9ui5tmj+TdZdJuXk9+Ha+N6yWE6jTo
u3ZyZHvx/VCrQmlYbB5A2uqWQp4GOXQXql5DGn0wl7HyjqeCOsswucqtcRSA9N/Om0OIpQl/tuW0
4/9RyoTT54tTS95B2837fgap/L5cvu2xcm9w+WcXCIKEGpb9Elhq2EHKsJ3/TZpCCRcmVXw8omWL
LDhzG7ThFs7wNv+4/RdQQsn++xYKjwQtewCu3eGFp0RFscyL91wo1Z+KKvnDUHeRUvyye9iEMJNo
+TAjmSo2tbJNXC4xQSN8O0rjzKdi74NVCazolKo7SCuHlcoxZdx2q4ik3r7nuPGlFVF3LgHb6iaS
veM52ljffkVgLpf4vqSmPy7VI20GWdztTtejA5tMVK0xURjpkFkKaCZrswOeX9rqXNpqNBCUf8Hs
rO2LTV/6h+Ko3QKNjZ0ofajNyLJyXx0IE5wVUY5gbH6pUWxExS4CdOAjFkcPOms7TFJZs/ETAEv3
839pSLicwnjZJ7FHkxh1uNPyw6bxi0sfYISefoRrieo8UkG9qBbL1f2K8depkkESftBieXaR9Q6e
giXKMHgIeFICcDAHsOWuZG+5DizPXHj2PtopGkAuj9PPmt/xgr+53jhcSdiLs6UxA662NWirn3K8
VepK7HNJeZa84uPdo/dg8xBHAuRfMfu01I1fFL85HT3/ovmKRiRwEsw/eDXiDlq25GYMPOb+kd2E
5IODoSL6vjCMVH3EZntnGiTNu3CkOBw6ZNDJegzi/ErxpMRUyl/QXB4V0ZsddOWJUri/i57Msui5
SeQhYf/ZFF8XqS2/qDsKr0v8SmSr4O5fBbyW7LPU8CEBb3SUYmJ4rjdR/A14TIWniqgo/JFYVKyU
77XipX4cIznDNGyRm1QAXbvVLqEhp4wWG4GOQSILQykAw9M8pUKN4cB4LynndZdCy7UNo1px1yyB
66yTrHKHcvyE18YYJl7otmbfHAnHwVC40sAahgG2RUEFiEoy9Y01jputMcJHdBE8yWPdzpWn3qRq
SpsJadFcJYi9kehQSm1Yb77eWuwbMmq1IJfc+jf9JI6gdr+EIYWRIaSeDKWOqktJBHWAzjzwS6ct
AgYWJzvYqFOGY+XYATHLNYDRqq4482Aa7aSIg9Nitpn0AOWrwQWuDCh4CR5ywOO0ZVwPvL+j0fPl
zCwEiMDjCI9aP+sNcXsHNQwc2DOpyU54uNvQJURmNFN8DLc4o6BwQi49ZD/t/8qnKKq1S+ZVbxJq
luNzyFTURLhRAArl6h/pjLAjqyT7NU8i0EDIhq/p8CBnrVkHWxq3zAvB+a+T+w/ziqq2hbb1KueC
s4CF++S55MhBLkgLyP3lFa9FEC9v0z0RoxSVqPwrVQB/z8xWL2umfl1N5He4DYpJ1dMtKXgClKnc
jDTWkqEy464JZI240rvxAfPdTgPQt57lnYUcdA/+F8HHYG5bXLLCI+W+s0U0n5dcza+kO3HV8GKk
SqSGW+CF1qUldveQAokG1ct2arOWV5oCXzLIs7lilqTI2acFQROtRsys3L66hoZPS3Uwt6Abkut0
4PFt7WVhCdN3iuv0jwHDIHVv271y2z8Elsx1QMlDPhnp7wgsBnWaiIGZ0CHYDvA6h5wB9G18hEQO
PVUKYaE1j8WB53m17igGts1RZhXgqCvRB3HZsbbNSgeV3WXNjav6gehvkBEd3z5xNplko8sGuix0
S7c/+nrsoshcMlFtlAYA3xAp+lA45dOuxjY2NMHD8GYioDC+wrhWlebVMW4q0ZaOG+jIwap5QKKX
ZCBxR3KxLzHCmxgzQOONFiTQjkFPHuoacye4SIuqne0HsALCTOENeeL5uzzOhu/m4nRv3xd9zCKL
X2bQKNIivFWmqWyg9RGBonzjmZowkOa/x2gUIBSO67P9KONgZNXlib6xFm7qZvyOVs7rXGVNiD11
NocJBeGuzZvJMbgmJzFevwqPNJvzfpxKohBeHrm8rM5Yva+8aEGQScgUa7iAEp8bk02gCl5WOjLs
YRj/y95MZrTNb1zbT2T5O78IwuO4j58Rie6yhuZfzkNft3xFqpZUwpOWw1SoshTJO/VRUWVDQaez
HJF06LAyseEuCdJXpqgM9Spmh65Kk72ShBkumoLOaWDP4o0Yaplmb0I8Pj547bOWlo4WsBzEYaQ/
p6SV8veMxGdNJXlZhUxBf08UCc+z30QNQoUzT9IRF5zO15l4PcHNUzLwSRBwPCqvLk1xCXFipqJv
npTN/DI34tg+9iTKRnx5e3mJTJHx4x/RGZvHZcjMybLfwlL3YQvRTnoLG2NmaQTUSyXaUAMUnXa2
9ClLfBTNH1U1OuRCL52Uqw11Bq83KDPSHeZZWNu9dApYqrl53a18dGmqwDV7uS2mhwnbq9/1ZbQN
uItbZ77g/toK7tn02UfCN2YE5chWfCLy8BTIzU9/rjaBME6SnLX6W+rcnJqhEEMbz7RuxvwTVHUP
MBCutC3RiCI+Kh2dsQ44cw/IfbzpzXF6sO4NonME9g4UzbmZzVBWqXoVS20TSe0EG7TRFa5+nv9y
88xoXjGinNtMYux0WbWlrXCCO24bOIwrvMoQt8MfMwpSmVALnPlRkkSu2EdUXqRsD4qFSMcDAOq4
v/q1anzT5wSAsANOHukYnE/JqNUtcnmXvVmJIrPk3rP3WHupFL3Q4fiUwHfysltc27CqxJSlO+3a
3jE8EqMqSgZUN41hevpMaZ5FYUKeZzSoRDfJWsLP0NF78Radg9vIa8OXbMg1R4NQDvyzKpLbV+us
j4oSb+64HahJ1j5T2/5l8i4Dm3Pk2Qme4BieKWpU2RsUQmT230Q6IoCzfzuWzeQfBxo8dsBKyPLs
+TQa/Gc+H79mPaEwnihaORPVUZTKcYDvdUwKw9ImiOUrps54K0FlQgFTZ7PSM1BzNRWYHrNBTWh1
Go0kJUXMsy/E21ZoKfOqGs3zsTLtZl9VLxW4xeuQbUiPNzHYsIl3v4xROVIu1C6noLOg+HgDCNiP
U0qc90yxr6e24qyidG0WTQePXTJQ5bBIzknybYrTtrWkJMezk+D3mzW8/nYV4QDp55OLA4ws1686
OrdZ8bgMNo7VTovnRmFh+AWGY7ykX/LNw19evoDxNMNJQ0t+C7UG30lhDrlX2CMCOM+XBaV/hHuC
CmrzlASGA22WTb0qe8kQzMa+dmuAc1JKPeFI5m+HG4XhSrc7Ru6GGw+CNrhwF0/efkGtmG1hfgGL
1qBRNfff7dA/UMxfIr9xOmcYrr29cNS6GY3DwQjjW1LFsRfXL8+w5YILFHypZd0FbUWADGupbsdO
bjLHPWp2n4TRQ+ZFjRMSo8EScrcKgQsrw7YDvX2rTrsQ7tcigrtsjXrNkcZqjTakf0N1XuvsgEWn
HU2mIFdYPWYaI2TEVNfvJcvQ5Ng7utXN7A0qPYiDLkziilnYmqzrGZiborEr/1OSnoMTGLaNo4ZH
LmIUoc+cO1DEsy7Vdb0IUKlIp/SlqoblaU3NdR9haYIJqP5LC1vdax47MsW5aOlFuaDReuTbu/DA
makmPmfla0f7STmskZlrAXjNVPM5YQPNbNsfuEjpjbgGDNnQddgx8XPbMdSrRsJ3ExHo/5AspyX8
1G5Nv/CVS2jhwBvJpug0ccZ9JWZ66X7GMO6sX263vchkz8kjNEb+UEw8rGDGWBxeZTBg05mlf99t
uwY+MssdxoNEFHXKpTpTVdGmMP9c1Db/WhiBkAh4r1oaqkneGZ3DlXkyXrWZlNNkKD562+N0rL0N
IJpYMsNqifGBKA6wk+pEr6aCTJg3g9x/Tt2tHx/UMBEMtHXsaXbtgUYHZgF7+kzwG6YSadHfPr0S
ISz9dvW46knBl5DOBKK7gMGu9L19m+h9aD+F9y7h+Z3lfk9vS9PMFWmGaJLfXwBp2ekZBZ3lwXtO
0qE0uHyOAtRNYX74hCOZbysFAfjmFVMOKNJGhgSCCtrsF5DGWFnDn9oxiooRO4QqxePU+uZLHJR6
6Lh0Ftm0C18WEzh4hRYmM49KS8gCk1oCCiqRwxZTI4ka3STI2IyJ/hU5+6qVyGMPkpDldddIPsGL
PTtLv7QHLDT3ZLboL0uJH933uNAQQ013QZdORnGaAWcYHuHMhB3cZ6Rda5rHN/rJmH3l1q6gtA9W
c7TT2/FTCY87qSxk9X2VkN6rsoDXKdg3NUVU3wwC9K7oTG4gbNvXwojgHbrgOm5fedYM/Ox/+6bT
iIy3tRNNLLhjnD9Kjd83rbQbEK9C6gU0aDwBDPx6nPvEXClkjzm34t4J0jT4aKs8SJcDH9GTDGs2
IwtWNo2YMdbSt4CL6k+ugNPhgadFop0S8wSlu6mjvCeS097fIghv/CegsqCiMZtosTh2XvG01FqW
FqNVjzBERmmqueUdP7sGxzcWBh+spi4ez+2XPzAcqbO7wbsBi9KN/6yan9xZv0pYRnxhKP8Y6b7q
U3gcyEjxAnQ1BLbYMrnQN9hZuRvYAqT9QbwhIyAxGPW7bpM6NfR3b0ULrHIWwkD35xwXri3i7GMA
rdAumbw3ra3p8NpZayOZaNsDzk6z7+pFJI7Sd40lfSVaVfvrlIZOu7a27hNadQULDACbp/6lAUmT
p9ODfzucZyPDyT/c0qMrc7V/pseUfbekbsuufJLKSbWPn3FJ09C52ClCsC7q/T1TOS+kJarCj9Ag
akJ1T6CsaFHJIMpa/eAHUReRr+M2opdBPQSVRw9qLBt4RVMl+ErS/OGFSRAEEZ/9LlOemi0Slu/K
+3VOPWYqt6PduNq6Lm26EQ+n6XZmSCV2KUC100abt3A/RKu+4sy+Fr7ZxMqtYkCtYi8vAMhrVK3U
JEZxnA+esbr/wGr3NA7CaBx9ANZUKwWdAqb34caxTcNsVWpWrcBwF/QHlZdBoTPuEjB1kgHtrElk
W7QWzamh2h+KO6JKSK3vCgnR2UL91JKhroc84xSOUkmmMH/YasWNSd8Ofx0PsxCW/TDbRehLY7KH
XjUxG2HzJgGSIy3cLrvEMvclQFp06wXGL4LZF8XLCvjQankntr5FX10TDF3wnpaZ1vqcfr5lF4jl
LAV4D/SEKKhlmk/wpdF+geTMWhhRC6EEFzkSDAJmzmZwSeB+iZjyoeKolaoDSR1DBPCtapguGw4L
TxF1EXfMl3t8ihYrLTMRIWURrv4ak9oqG6ReqAUwNKyT1Kng+6xj2Ti04RdZ+168ddo1pufzEqZh
M9Uwt7ziVCVY8PAea/NI8amv5O3IxjRn3VwWxio7HxSmQ1A6CyeZM+SJrSFdoDmoBNrKbJwWiLzG
NvjA3/2JQ8YuN0JRvqGHm5KdQq1iydQuAA81uvoC7mfy25JtWjqPOoj6EW2i7HeWjMBs1JtzF5SR
9jX/SHloms7Cc78EzKIuAFfh/vzWgT7fmAV1Zwxvc8VvLYyxdi/6TEe/BLjzXv4atK5zzMJOO7n7
9ETvPrXcjJfQeF32AodP+/j1Ih2PpX40MElAPco+x8laLg8XBFnI0EqYMmZb3Jzh6Zt2iV73T4f+
l4GwRquscqCs6/24S+YGtbq1V5bsU7+LIYACBr+hzUCchyiaR8owDy9gihPO3EYnTAxCstYNjb8a
qC48OD8lhyvwW0FGNlsUMRIVH0ZQ1+KOwpOVGTpIlD/Yyn86mwB4E+LbwqrDW+MJ2ukFp7wb5AeQ
ec/i2RfklHOL3+A3D7yMVXQHiupk0iOBQaFRXtchjyJoLd94i0XZqu7Et/LbcZRcI9I+qCbzvtzG
THv/2YOTAMeFW/VIBwozyI8sFvl8pkLSD1eVereEjm1+Zwz+ei6WzKJ0XvkOKFOtBMEDxFSq7Ldm
nF/KPhfKX3ZUADAWr3UGMxckaXQA/AMK0qALO9CfII94HgFbDk3ZWss2P/5d4kK4GjQlC+BqbbZl
e9YV/MUGCnbyf86ENQmWaBu09xRyXLCUa7qLvRFyURFRU5ymS4uoSFRzOnzN/zRuA9hVvbb3kuz1
4b0+OexknvtSmSBT3S6XeJR9D2ZS6YeQizCTIi0OjSWWGNnXPKuDR6mTydMM144JHZECrT0UGqJC
kvXqxpKeeZDl8SuVvYW4vAxKzeYCTkRprjEh0CF0mJjZpg6mvDs5DmJbWY32x2bj1ivc2GhMXt52
6Pa6CMhlBNmUyltXN99yevTTMiY8V1rovcXoaNg7eK31/ba0EqgrvCsJEALwLbg2MM0IxFxkTL5Y
92XQd5eM6oCtxYG0YNF2oWg6DxGrQIqG5MfENN81OByjnXLoIQrSIVuyG6vRKBSWfu587sre+D/9
zcgQ2oqaWheCC3uY0x7Wex5sc6m9SoHGEdjtrtq0l083Q2k7IcwTZ1DAXgqrOqJGXJY2tJZVG/qb
+GAXoWtkhCGFer62/skFFOgMYSY3eL4G8NqbP0XRNh7j8RbiR70okar2NUwoZKBZYJ/Vuiw+C++5
ASGZHcSXdFsL9JrZ7Clzp9A68G/Pp3eBVIWOXmaRK0UnQKZFcWp54Qzwwj6SkA0bu0sxqC9Rmz4G
uChKvDlhshTLzEirttRmQnQoQH3BceU2Mz2M8krDc+vURx4NgA4m928xplHWOeHO9mIZlM7+Dbpa
RfE0Yv2Jn2yXWDy1Ib7p9ePOf9T6U2jFS+DWfui8CD+yPo7zx6xcDBuml1nGbFE5X0qAUuoFBwcV
1bHTdRLMyCM5nULR1OHYDIAfCPzjs4jTFqUZgzKFXFxykZe3xN+X1awLfQa3QIoDVCrfd3VfIMwt
h6fn7EaKMn7KeqvP/JdV7/e6GObQCxLWKjV4WHaPBY7CMMRyV7mSP0Q4l+GW5rShFxl4NlSqdPjg
vBev5vRnBHw1nTCoRQgWab2BCB2kNV8uSxmPGIWsqcuWCiWWHRqNipQPrQvEctaeuELsxjG/sx9+
VDLJDC98pCqa0fgczl/eAWlZ6kxHM47V/fX0kygs/DkLthSejDa0A4berhjYE/eTSvGDRx2HHoSw
Ifki5zQ2Y4PIKJGii+QwihLqi0FqldmJIZyaESvSFbPIBrBl/m8KBumSS2+EB8PQfuFzZ0CHhbio
sqvSouF8yJqP8FXRmi5BSd4DYlZQwetv68qUFVd0TkC5AotQIkNPFP94Xujzgl/kbk3rC/hSOw2f
AR13UNSnwEDYL4s0X9xRtWUar2P66uUnx+uqSCCjZu/bLnyjDBY5HCYh2n+k4+ZuMdEAj31b5FKZ
m+jCeiYvjgYuJ8TuLQrJnYKKieOZfmXAd67Evwf+NQK7RNsJ5lwxZgzwudd2QjpSks5bMfS5ZIco
vthBAGbpk24Vy+VYQe7dXr0pqDc5k1gSx+qHJk3oVHIkl8P+tIfJ2yEA5u5S31QCfVuPSTTf+XA3
eO7rXQVAkfDia+Ugyz+G4FI62n33eOu9PSwl+rcV5h1wBiYeelAjGfAiUoAO9yTCSuQ5m/yfPXgJ
qwUyXyB1HJ00zjdyg7SX5BUnM+L2jj+LNW83GXThq7cCiz3W1XXghQThYOLTL9+mHs4a3oyYIJyY
/FL3L9xVDcft30cqLYDooIbY4Ieh+kV+Al/Rsq7MHdfkfJ4jIjZUzDZ+YADGrwsFsJBGsuS1BV55
q80QqNhg9x4XZUX6kZGpvK1EakOg72gCfFsid3RZ94/aileMmkxMx37bZ9qjNODlR6WOgNETussk
ub5gIANTeHDIrM+GgsV758OPJZghBSbHqB7xOTySSuQSahHs/ieaW2+wSd9MN9KY7xnjfU5kyQT2
kpW15TywiYzgbPjkjO17Ndo9UfOW7R1aDsR9VUAV6TV8b64TI2zGrjT0hi7lrj8hkr58mkQ/P/lb
NdGAIYyK5V5AFZJzUXVOitTKsl24HflT30A/ZfS4CDHIDNGXM0az1sczqSWD/tLiS2j1rUkVqrjC
kTCkjGg5WK50S01v2mPrEu1hi75mufHPNe+kYTZi9yopN5gvAa10NfuDe4QwYpSWajzrGmjVqN6R
wVqUnPWMQ9oEUW4s33/S3Dhsfo15YOJsOcsArbN8TVkyFbwN3iK77aIaoN34PnewXuEM+X8AyJ+5
jHdoNwnQ80TFYGr89uyXNDVJhfQNn77VkzZ2BS666VM0w6cNHottmVj4phBIOfAwJa2HSVGa2HFQ
35miD3KBD/YSvC3OPkp/NvMkviaFkxzZw4xMmW1xwLCKuNqP6fOEvQE6m+SZKeQMpzhlgW6axrm/
X3ck4Jj+nBrA701sIOLhz0UhQHWhAX6ejymdqIHiA/vsTkL2x+DGAxRAZdYKB4QjXoXm5luGgZl3
FOzcfH+K9ECPR4yyIjourpMm+FzYpA1RcD7qIn9ous4mP/cCGvuEdpM9dYUvtpV9vF5ldCYvqRMj
AY1phvbJBEhocFVE6WBW1m12MqMpZYA/LP7zJpV70jyIweDJugo/cr3OYrog9l1cxsTIQYMrGMG4
AbaZfQL0ob/z8DEqIbcXR2cYXMNMzdocT0TM/77+2lQbZosBIB9WFoTcA1+mo0KfqdfIBDMFR9p0
8Pp5Tlix+PSQ7Fie9CX9EVLLctM9FnwMhSJTX6X6tGtyYc7PLOcv1n886nx3mpltTFqLNHd63ji+
cvFpDi9bzaED8MfhAcmNobyOJgewDbqoE8n1sMovLqRUtGXrLEdq8Phv3ZTuX4lKCy55b91HNUGo
P7Ou5Q2nI+Dg1Y7/y15lnfcVpH7Fh57Rl2xH1nZbShBpwYttboJvnCF9b767lW7sFgixGYveTGKU
u/i2U91dpiX2VFYI5Vda4oYuKgVIjtPeGXMCFVjtBQiDr1MfEsdNmam6/xs1Hm7hwu7nz5GOG6hn
C+BHCH9uyqZMEHwAT1r8lecBE2BXCM37vQUN6hjDNf5o7q+jPHqVQ+CfaczTGAxH6Fihuk8CCcP1
4eIWNoVnqa6f713iAxBprZV+NS65vg3nwtp7mGrZ5ZTPvzU4HHvhQf/QqQ/0DljFQcARe/RQSyq3
3P2xb7UpzjlDBOZEYcXQeBtTVF/bcxRsGY4MqRdD/bbjKp5C0lTN4vPYUj5OUR0jvcUc6mqPrtAo
LAYyVQuK1YQ0+lZBMwMZ+IrcFQIhHift/UXMHo6tHZRAwfrWc4BnnJTBMO14ZjDmQK80HVJ13XBJ
nHslfZcD04xBi+sDhh2TVq+dVYT0SFJdTZL4G4NWRUqCdEUgKawqJKLURl/bj/qYVNW3rDPVKWzG
U6MUSSqD+Yrx4w+D6a8I+kr4G3Rf8NcMku8398ISLgrOtwcfHv0VLXQuIn7ToBJyl7qU/FdwmXlp
rO48A/0piLgiXPck0rTntfyPpBhRsUtzQ/06EX1ROpA8kTZGkMK+cDwC+lOp8Z/ke0FGImgDTX/P
uv2kq+lxXXVdcyb+xgoKSP4JC0h1DwOYiHQ7cLMpQyvOApfI/8TFdBFO89AqMJLzjYVszcSeFMSN
tSwM2RNCpbdvsse08hj/98Z+oAjZO0HKW5NfLYvD6eAt7ZjWkMs6EtHRT7Freyhtc3XELbHw44QD
0kIYjfw/pULbeMRR98EzRc2ygv7zO8MVBTTECZs7Tb0tWMGVPnobKE04AdnQwhYHzZhmdr6DPv+7
MSVrmb7TnDAPx5KtOqzA6iCfffS9/SC4P5LOTRQpvclnL4on6Y4yN+yvYalb5FhQpMc9f6N8T0v+
giLotbANMCs2gbQuPYiwqkhfUvwULErsRqWIQ5LNZ6LqZFRL/Wz7Ap1A/5hFbsKamApPMnCi3ZkN
iA9k57D2A44LQiPfB4IM5pgHCFEUpG8Aghtmswj60FsBGITvr7s8HV6vUEof+zNnTa+PS3CvgDiw
G8X9i5krHUIZhOSql+1YsmGryQt1vCwK1ZRqofMYNMdTVuDZ76X/SmJXQbsT3o/122gljE3bcvrn
vjnL81duIc6wJjD6nrVS4VfFR+XJZwddJrEl3haS33u9Rf0PWBoDFVpTYFGW6+3/PjKVe7RIZy4m
HmVmc0xTzwqOqbpUDuH/DxegOPt7qRuoJsawGdPN5rjIHjgJOsqWePOfpaK50GjHQAcjbG0UWqeD
4pWUcE+V2fOXMYy0AVFJJ0VFJoOulFAqgpTky3raSaB9nXDlkfB7P7zdVyyAv2F4Xc5waM4FtCrz
2qNvm0hwZJCtmezUJI6qpbsr9CMgCglpb6TyE7fc4AmeYOcyEQcqY5jIUFE6DTItoYSr16e6qttA
z+lLfDYLGUqAmPNZ1wDQSh5k7DIc0W5gG5iMvggs0e0HE1/ZEXonnm33zwiJIBGkCTiWKD6cm6B3
lGOL+/ZrBBGT1MICeto7W3MzJukGpqA0FZd+UG8clvp9QVieo1uR8GvCKOPa4ebBjXoCHalfnnVt
tl0ZZZ+hl8le0e0mRjpLVkr5Au9MLPES1TPwzHmZgrz1hwebHNdWs9efYlJGItxFMykY953dVfAy
0UVaZQMXtbAeX60fRHgZzFW9K1Qytyrzto9h2w4AKMdGXCk37eh4jA/dcwxjo8fYqkopiOjOjDRP
Z7tH6Sb6+wwRWLmuT/MgNqxbVfRDPwKv1+qoq10z4AcZ/kmj9b4W10PB6QYU9+DSVholi56rvIfe
Mi0epn5f1FmTcpPQHJ7XRqwOYmBQVAp0Z4zoyLPUE/n3uxuWLt+QgLCIohMbLT3IE6qriBuykXN9
WKdStOaZAXOYNxp5FcEPm4bG/40/7r0yAIsMBA2SCjZ1hfVBfJLJYguXkmZa5VoSGtS9zmzCNmPX
MRe3l9Wuj5d1x8LmYAXEbJh2kzLzqP42oNWXUdCR0vG28eZ1Qndj/bbbsjaL1VxsOxvZamH2wjOv
9kW5ohoSGCG7bVog6YGZ7ex2cq7wpYtVduGpR3jhrgjFcWjf7E1Dd2oOH3WuOu5wA6dGt6p5yg7+
cJlK7obmgLz6YJdGbT6cEl2QZo3VZJWTXF4i0aBj0qG+D0gu2L26IgWd9EBgSrdImD09cARbuT2Z
e7XTuW7OgKzELJOXmtZESPsRVAvEdGWjB1AQm7uW1Clpd93aicWarWOj9hVhmOng9eB9KEDelSe5
Dl2TtWEtQAvUWlH/URgZzOvlBSgKHLckmchP3iVhtpeuA2FVVFOHAvE/q4DOZtmOD0P4KHVWQEkw
tzGDLqpQEuV3ef/L2KHYMSWQkjAHOjddkyOH+5sumYlyABQe/STlocc+Xg+RS5cJWfL4/N8bOV4Y
NaLrwD+oWXiA0TLgXixPMmTbuVneHuEgzqlFBY76S9RcAw713BgBitlHddLYvfFoSgVPrdZBrEVE
R4Fv+KQr4wGzsmqppD7OiURTGQc6Y0y1i/J/T4C88EQRAnfVJJX1YEfWp/KbcmggpNocgXaN11Ff
r6S4YIjUSaYq4zFqT8gjxppBxK0x5d52QWo/J+Ge6/sOdkfmNXE46J+1ziuk7CxA9n07f4t64Bo3
Mn/KbNA+U9dcA9+rHPKggJjha9bVW/F8dgakMiJ2Xndx5I8+8mcCle+BFI3Lq35wkC3lAh8N6n57
FWCIyDFigOVfYjd8abZFJylS8/5ruR+418C51KOGN2TurVXMCjJm5xoiTLEbUCc++PqaIgScTcOW
biyc5SuFznAATzmsYYfYWCqtCZ0JIl7M6+ah7nQqz8AWJAWs0gKr7UQeLpOZwO2qaTyRR1enOVxR
YC4RC+kGK0sPHhavL+KpWNwh0aGfSZ7vTdvmtEp9BxrG7cU4989RadW5+En1ATfyka86ydF0VMIJ
bb0bDyWmtQMGFtmKjCj9KSnLrvvjOOguy5d1TeiLT7Q+IYaolEIuP7PraDCvts4xKJl0L5IUrpVj
ANYulAyyeyT0S6kdfNQvmh9Nq6sn2qfga3GzAsaoHmAZ4uKJ44xCIMvhCtBvdXAIFm2Ei03FTQ95
n4f6Bj01smii44bBjn1gFRlaa4g40vADTJ7TMic++O0UOpCAbCuhUQZRUUV3aYzUeuMDiZJL8qFi
xI+uCAChVtGseBckiotdXc99IOnuK4sdNUtKo7wodZ7jUjUrnS1pYnBDqlIjuxI1k3OSGoClUtOy
jYB3HpQmvENtt3xWvQ1SWUsjDjjq5v9Cqft5law/tYD/EnttMIyKZyqCWyXbQuX1Xh6Rjvbu7xAo
rz5PRY+8s79NqDNugYjBTVzMZee0fk9bPUg/V+cDY52ceBfrY+c0jUcV6jh052Ig3zgFOXFeJnLO
zEbd7lS924uq8aeeQql/riLis70ajuPnhLJFoUgxGDSG6uKL01yBleqv6rCaWTZSlc2TiTG3tnBs
zp+LVlGcKiUMH9vPcpVVHgvTdORl2VlSlFj+YGJs7wScEJO5005xePsmIui2TAq6mHY6OUuTId1X
2kofnjPcy9ZJkWtjfZm0m5e7MdJiJGilU1ITYjKRgR4+Ja80sqgz4Vk2ZEABELLMdDez9GBrm0gn
L0+LvC633Nn/M2cmx0Y08exgrfFw7QrdAZS8pvN8Zn7STXGCyoN+2uWSnaG5tiajKur5PCUz7kkY
dXoJjJwJRtmCyNTGC37qrM8gRdy+hDEnZ4oE89uF+O4dcJfhO/PwatuJ3xzTpZuOGdTjDiWnSXzi
ahO00ORRqwUwaoYVtyJJJ2h9qVez7IdqjUaoexc+AQXK1MAOwhreEXRxCGOhhC8cPCqFolJmN8mq
KZDgSFizeKvZpZzMi26GqQDucK5sfQVuQMktkjQiP9xnQ3G5hRpe6JYDvATXPyVaAqLGx9tzuk6d
NYB9+OreEl8Rv/WKZ6pJPRejEHEOqADmbhq5oKqg+FVV8kz3z2DgOhLM70sxGF4vT3251+jf5J8h
hPXpzEei0ZHjJtFYpwsmFOz55oCVOX547oTEIK8UPH/owXeUkY/r6MMxzaxZHIjCEfIXumn98rKi
56hxgnuxRIcZU5eTF0uhSyq+wyDCIvkkpzLjnnsz1qW611NIu76+54I98oJyFowXVPHQQJsQC9iM
ebUf0YhtBOzYiQ8x7knwnijzOIX5YmNT4PzTF0Uiyyhcov+tGaZ+ZWhmMOJ+AN3rqWFpn0UF66dn
Qzk/aK10tH0Lw9sLFZZ1hlsrwWgXLd8Quv93bC3TkduyZMbfMxda7Y32AfyCf4/K/FXzQ+nS5Mhj
3tgffwTH7X7qmMmTMi5hqps+2SWIJZ5VgcRf3KaqIT1ZhSq33V9JnWw77E7VNPfEUOoNNB4Htpmn
KYVh8bF4ag06aRuVIRqH54lCIcMY7lm3ce3t/WOX2SMfYm0vIgkDHQWz/fa0+JLmZQRYX9TjNTZb
B75hCWswy8UZPwo6CYb0zIfx3o+CXmIn+h9wja/TlD0VUSAJrcVPQZdmyCuDMQUfSIqUVhDqphJX
Vpy6d72unKzJHJ1Fcg4XsxAjAMiVV5jmkARIYx5M9Q/UmyS/JuWpw0pq7N6d1hzOjwhxnpVHmTUf
sdiPYlMA7fAnYkvZka4hrActLIRiTUqgiTLgECehAFX6Af93BV5qngTBngYYBncxiqSeay5trlw3
XwPae3TC5H5/Ime8qn7MdeF5KlAlyDkHD6+W2rMIgdx4sJweE262BhkUdoxeV34Etd1j7IN4XTkI
4dl8RylZa0wzB/2E+vLnxL6SGAZxZbn5MyWiz04enPrFMnq9BjbAmk+N9fcUAwCaolwAia1hN8ee
OevE+QF9H0R2ol7ikGXtYjbWfow7pP+rsjQuDPwbYVpi+yvRUTtPKKF/yPVtYz3bdrEApXa+su8r
CyagAmGXsxYjZ45H4E6yDo/bpbvBzw7hCPs/+cNz51emWLCgFlSar8lllalgVqljMsffUj25hvNd
gpsHMXgYMIco2iwB6WxIhLVzn6PvWuLcwyN3d9WcAGPISKDGniubYohFJazLxfC9YGIpAYlwS5if
Mx93xvqX4XCYYAL+RDR1FwFJR1ufp8kWgGJm9YQB7hzlH9E8k97MuL1MsxqJyItXPw/zG2ZvMxSw
UaayS4Orgbd/1LjvqWCrYZ0FxFusUA+zGl8TUOro83i1S0Q4cErSA4JfdEmkpocBAsuxC7K4veJU
kr6C8DFhDJfXqhsLF6FDNi+quPVfjCGkNETShS2PLIfo36m1LJwEAHpFkW7dSAN8VzTV5i/mQ5oN
LQNa3oDonHlTVWOZgrs8HbggP97mHnK/sqJuY9kbEuIqcNvIHDcYrb+9jqp+d0IRdLsHDDgPb06i
bqz450kuAzmG3A1dfHChqPMcQKxPG2cvv4Ba0O5u6/LaNNWe7uyxfIYH17V09tZGnArOwiftW8I4
0JUZA7XieJUJ47pDUqis8u9zn+1SZTwS75mOQsD/qza3hg0xO0Tmi+Bn49jeR7k9be9WOwa/829u
+zondCXJAJYxrtuIlT4/jLV+zeNvhJu9JfFMO3X4xHWGtFjcqWT5PCpAjUWGhRuLrBGGsjplqtBu
N3jMp++unxfLV0pM+kdCXn0DwoMuz4CigM8Ws7R+/8gIAMXT5sCEd2zggf26aQJU3xMOXHcwUZ+n
l4WlcycAYyFSAqxrsbYnhy20smtenagPQqI5RxetuLS5WoBFCofNkcVzOMYtDKGyGXuqzBlppP6O
pM7NiM2VfNbBT+l+EtaM0211bAw9Np+JW5SouHzwZHga4x8BOSaPfWeCY2MBIU6Ti2XgBu3Kyn3P
G8vy/efPmvb9zKTV5HHUKzYu/8CT6EACeH/NqCOJUMTwkrlnIYjkVwS0tMZadOnYNlHXTJG9oqSA
CslsiXQBgn17ZYbmUxYvsA6zhtqtbmYGSvwkTLwFG3daaquhjddUslg48cn5axW1XluEGeVNAupu
BCKNDWxd30KV3ZdlsQlOcX4wWbIHe4l5MldyRr23VYNZYZbSkXZkVPA2CtUUHxJ6FdU5ycFcR7i3
LPN83XO+Sq5UUNO+OxV7Kep3+vp0uJiMOiPcsfMuvU7Jlw3gbAMJv0CkZXGlmBSE4O0x2qS7ACSW
d3z8kBMAezybQwbUKfgzOWnQNxjXDh20Ar8A5F9dEDoy79kF7sHWaI5rtJGyfVl3p3BPUwwX4hUO
FgfXvUrW3tQ0sFU1u9JOnimeGN9c3myTwndPhzOKtS6setQri2LIv4OA5Mo5SB+P37zPrV4mqs7d
VTXzTwumRdshADLCB/9phGPiVII373vWXZU9jBh36znsJeTrv816dWg1QyphvmlvsolS5g6i8lhT
7fZ0Lw8J49dmtPr6GXy/t24ICpFsX7SSY4yThaNjQt4PW9Uk0Cy9ETNLsmfUNks3X20FTGtQij77
jTg0cVsWURyY3K+7SJbCB+pOADpTSwOHs4CilCyMCDb6mEf2xobORVl7BkiYOGnmH+EVm4bPqdly
f9uYQl2UxNrncjvr6YPQjIbXNj6HbtXAs8eRnxsmKX0xa9AMYCKaJMfGr6dUH34D4UCQgFKVDA7m
6kJscfnOO/SfIZBhm+wIkEpj5fUh0rWqIof1aMwly0bCeXt0hMaa71Pgtwo3Fc6JjKvHVMezlsl7
CLtuHZHL5lPdADLO9ltj67c4l3GSTA4zhm2bxjLC1xbiGzLjxCEGrS1vOvL70POJWnTGR6CGmOZd
otPXGIaIN/TutpEegO2YvUoLS7HZ54bAGhKW7cLe4dhlKuH4+gET5mbY2GfIJbNBi3iiSkFlv0ms
x3wu3Tx5BT9C7jETAy55S/UTo8RlDpj1zmP+d3BXaK2nib1AMSmXOl8mIQGW2zY1RYEag0wglNwg
NGlXRtOhGY+jMP6en1FIO4cdEwf+XyofI16izRjSlLWoZIl1fXGboE+XL7VEqN23vsfhwbw/BRWg
Wv9IZkJ/ACiiLiUad43RmJCPV1cx/4oogzHWw+mAjYInBZUkfVUPmUdZUwjYfmGwePjDGm9m1iul
EvjG+50wGedq6qhiys2BWN54Jm+UIRViKmnN2DZGmajPClU9CjY7gC65HA/m4PmqRK+y/x/NCre/
gJN/Bcfn2J94fwpDX/9hbQp4tzrE5HYep0u2XNKmIoC1DCoJQraAlbxe1Pb2MgQB5toiN7oKAYuo
1IN5fAM7ic66I0fBzJ74mY6YmMe285aA+kPT2VNbQcorUMU2Vc/bucWBwrjv75eAVxMJWzWbkbNN
+7NUCDf0vAHe9o7pShDerAR8RP1XcQNp1Q4gNWem4XxxiQ5euSg8UnWf/xKQz2odnHxPQR4Q6RHr
QB/cYifLeQQflb/KBgkLGWd77GrtkWDgnapN2Wjzv+3G1yf/UX8lc660NmxYwhLav1Y6yaIAaTu2
ailYDkygwc6S/wci8TcWbuRn3v+vvZwGhIkLc3Jzr+ZEs3/P5J/jQkJ+iTPuVUQ3laivaVc+LCAR
zNB86j+Jj0yWNXZA/HazdoO4BJAOvmskVQ44Tx6rq7o2p/z7TEv869lkafG1tshUFuSY2TTB1/n/
rmZzpCyOrBqX3TF+eOtl5WDfFovsKIHH7/y9hZmp1I0ebads6aRWOgGo1BMWTPTcCR1+JOQm3tFz
dtq9O7hFENlnBQdgPAIu6tA4nKuKRaQF4J/qzdPC+/LYMJISUZWaPmI2w7xe/KkNRKpUq4GINwuS
iqnEDPrC49SyJBeooTiFYAwjjItcB5S+oLzgdXSddLU1YnVWkC+eL/RSWuObKMskO6eGhmqbAuHs
m9NwY2seDCSBYeELfI7FQGclPpiCcU63tRQHpyHHWRLTj59nU/vivsqRCTMIO3UDGS42bu8P2NMj
9TeYqLjQuhD8mF6QohlI6eQVPeNSaJ78bm0jvFJalopquKHxyEMDAggTD0MGk/62lrd459PTdaH8
S4yue0zWDnUp2D0PJFNJxGz+fXG9c6FNYmiLU7haLlPP8PSBqb+6tZ6nPJNDQ4KmgrsF5SLPwcgD
MrPR0JelBYsnE5N84Ush15uG4Uii6dYl84SZqbbpfFBSg6/+Oc+gOykGciym6r1traHLiBks+5MK
rTNWTS3VOsanRts+Y/iTEq6jySrQLiA34eFbPvOA+aOFNOkiSgYOZfaBC2xg2dp8QSdgaOXcy+DI
MCKnFHpWzLuajIr92z8b47S1W91KqmbLYVgYCybFEFCZ/bPKBQMN25tzAyn4GHhOuPEPXSFH19LG
bdSGBqHVN2FBmfYfQchkvQpNL95vbh0ouus2JWCzT50z4pu18muh4YQP4qZeORqYIqiRYRz4emV4
O/TaLExwmT1XXXs5KCrXQwqls3fiHiiPhFHbOPVZfsGBscQeWh/L2NrdCvkZyBpzj+hp+nUikh+A
7F6l1KcBVbK7zLjWAYN4AVvsRQQCqklWETxJlLjM7cvkeqRXu0oC/gjnWPqW9tN15bVKIUqXGNkM
30CTRTajRVazB+QuShtGQgzM3N8pKb8T4NvvWqCWlxoJ+rQklAtP8FiHihGRpOnnnxPoy4mTd5Y1
e+3Ab7PLOyK2yD/4s4iY1njyzT2NcPo7jOhwkykC16N4SA6ZltZbpeMETrQbKe0ddxTca2mm4MqL
JH/sVgxqRZp2pfoRbB6vRJVKuua9Ahcj5a9O/AB/Chx+cGi3Jk6c4sb2zQ7g1CZawNfb8qPf5D46
MuTXYuHAXklV3/fUFdEeZ4yHxueH6kjCr+cerSQdQXm+i9tqTfRcs2CqSBB6V8CU3+vX22AWKlHK
fjdtVRR/6r5Zih4sd9zVXCkeKyQD9oSTeCp3xatJZny37x06Zatg9osrjgRQpjNzYlOZoqhl4qak
jTCqE9gbc2gzME3dSMBXwHP7PSQz36owTcbOGiFH7YEE4vAVJGh7btpq9qKFMBP/4Qeq1xhI9T2C
p5+RkR2mrI+Joy3FycyIecOnKsLQvpkQyXIKwnLuTEP60u9cE0D0fAbR3FSaEsTtrNt6b/szAWJp
BbGxD/JpmPXW3fvtMXGG2NHFH/HQYs1ayRxzff4q+l4TjbYbB5DnsHbcJXnaheLkoFDh7WGtXVLE
woARpsYC+CjU3WoIBT6u69X2viv/kfPeeFuI2PobnrxzynoWVQXPAjwDyFRdAGFTXMBCX7Z34bL/
X78wecbne3QkWvRogm1GBPXRxhAD4cYafNN7ggiD2+1xfWJYGvNEijvYUgWrWA5oUew0ovDTFCvS
DDJtawWtJhKoDEIBbg0iQ97tNBw9xV1tXExEQn6ajQ6hdSmfy9QMYD125N0TL+QKoTEE1+mx9UBt
jgXtVVOPpUBI9mdHE9VqYs3lOeZ6HjdAw59UlcPnqU4s0qP/hTYyBz2bubCT4Jg8S8I9LzqRfX+U
KedwwroBXUc56XFtG4I9IjaZpyXFlymBWpf61U5A70v9BqdcelDZpCv9KoaHDAgeVeCrGIVp/+q9
nzv0hIA1U/1yov1Yn9+kaD1hUwRfZaxW0Naotv0Z01bA+VXj3bdOyNGj+NiMbYFkZWz62wFT+RaQ
gAjPviNxbQT+xgOShFNNUDQFcvkORY91ksiNNXh992gNHddYgCBPKBRDohuRysvJnXIwBbuwiiSy
pLVnwS6x0t78oX6MzP0qKOBUUPznw8Kg62tm0jaMlMjH82f3FhKnNLxReiIMDO9d6S2X48XlVL/a
xZOtrLradR2w040MMW/OJdttHnvRxU2ab2KwuOePLC9yx81X1scmmLCKQ6q2QYyn5LxbrVv49fDw
9WKLKZWEjPmdqaQuIhjYtFLPHRwM6lcHuMGyyR/VGf2+lgTN6xkI1fWBabJ8a8MkZ1+gQrUEhFC4
x0xB/UqNQrOZOPcOGxv7BV3+X+3P5goa9+b0Bos1JlhRhhlozWhWs8r/pM+81kwgfZn7jTX0PVcN
KQucx5dofhQy4oWSZHz5+NfqcedYkcQs5Fme+X4hrkxAMqFUfQKP3qPgee5xR2T0VDeEk2veqSuT
qEjjaP2qSP9q0vMY+/LEBVUqTnKaCLv6lMDdUVTRcBnbm+TCuQf6Xej9AH6XEC5SXC7tWwMjFXxl
e5UnscUFQENXsL+1XDLu+RdOIpcq90Uu7DsNRU4lWqWS7htg5Dt5Vf/saYyeUGsdKnrxYxtFx3KG
uQs1k/i3P/j7Q5VF5BbYpB1gX5xYL69/ZRcbBUKoe7Sxz+Te6Iy+Nlg/0cBntmfgfLfL2vxPbkwA
OTwNB+/BQFqXsC3fTJaT82n3Tqh6U099wZN0xbxxqrIVJxJz+qn84HxrEh11PXfFaCWbesAookp4
ztEqSwj4cjoIrt3mi8IUP7FZPdEzNXgskpUuzNvMVyP+3lZqXtlbVEYmEj8UJFECJGuzDLk4dDWo
EkGKjZVSspNB+vD848nk05ARaCULpKJoYgi4ysDwiHDTx47mgOmoCHdyhQ/uL9SJudJYfS30CeC9
NNvbKZEdxIzPrAtTpwv3zCMf0YErJt15OaF8OBwVyJOlo1xLi41fpNO2eQTKEl/vSFdOcvbjnNf+
nSvvemZnmUs98SjJslug3pZ8waAGG9RhNNNUJlBzot+QN+YM3zRpuYzUi+xkCJODCoOtD4KbF1Cd
Yyujbt8lbB/DCA9c4AGjC5V56wt6kO5g+7oVL0fi/lH0UcS/P6la4QJFvx4boMIRL2N+buuown1c
DugLOzmH7sozqkYs+r2yR+edl0G8xjRq/L9U65te5zihAI4R47lOiiifit5+Wps3ia+ZEPzdkWeq
SMUZ1ifA78QECZvovGDp8kqmsxodcTgKmorV7kXXRw4z6O+NUDFZWCCOTeYclVUJR5I6EHdt832s
ndOKtXhPb8L+5QX0KJ7MJjQ3Ney9yXB8gEj27ZWf3LaZ5a2vViF0PURiElM1Qn31+H142sBBsQRQ
cS1LQG0qEGo0nN2FGrOcHcwPVSpyLTs0FDNrWyNSOPpY11gbAnX1yNFyKWkKUfNwHhcxYdEKIRb7
G2ZqRuIXXWoUhhH76CM5+uJJac2Kjp/pN7s89yqt++TK/mgq94TtCLsccOzp8o2ktrdHoNIHZJ7U
6jdpx+fmc8cZzKH7kWxfnBHQaSinviamdMp3JlXBoC3xNMLTyC5EzzKWSt/f0gro4TqXAiCMoQa3
bHkBR6+X3yy8wzqozqkJN5m/gtDKPI3Z76/ct6gwe87L6tug5NELXwDa31QPvumzYj03S0UVhnmN
e/Xmftvxj8fm8pRzV41iWr4Brmm8fSRhhDxrcXv/VU5eYkyMysp4G2/XNzaeR2UF4Hr/run3e5/W
Q/p6N+/WlNgFMrqFpHdqNf8hZPQyXAanL1yFXg5IlIM7kKDK35RmdLWpsyBIm1FuWoDYXLH90DML
cLU6rNFkZdsPUPPODqv/iUZWGlumOnTceBaPazsCJywyoZy3kPCJyun8jWeR3joy33HosNsv3Mlf
5AGcn3+YZiLwUzqIYBhPzmTu2JqcOhBkO481+bh5VzMEPgO0aglGzrL6f78sEiqKRdptj2zlYjKM
hXCVrYucedEmKd1djZhsYnZnpPbJxGS35iiGtYsjtsZTnuQVkl7x61fQ4bRSFgT9QPN+8hkq3SQP
2RVAkLXdstuzKzepvAL6F9HsvE7EpVz5BlY4aTmh2TlCoa3FJK6QAW+OrdIwghUygafRsGweK1iJ
RfcDi07kxaM3fdJrhi9El8MHt6ySM9qVkzVXoZpi3WfpFIzfnh6aLgHy88aCBRnpBdG7MVBpZgfG
Sl7yEMHkdGNdLJKMhNFDzE7gelIx46q8Q9PhcOOI2sFYXEEVTlypx0Vh7/i5Cgczo04jy6PzMtHI
EjhnrhYSsU4fecYIBbPmZcx/mq4dKfZ40KiKh2+hp/gmu3JcwUDeSEmj6ZLC0p2VbOzyNjQaGryn
F1wZlxE0dKY86GpBWw2VSV9IQRzEfTNF3dRYdgliDrK14UblHp6j9C5Z3pgnTYqHLFDpxmIzt3nD
IdQYQJRT7MC7U0t5uWVl4VIPivsNcpgUSxPvQaWnb1J5bCqmPFoMqXxP0nNf8IzQI7YcMPtD4Apn
OFVPkW0BxlL9TLLQTKTzC3qaiAr4S5XBWwaXNy29Z3DDeEFuT0LwwctkQbs9IKmci/44GterD7rj
NFX4038D5yHYXpYJMYvYW8SQTJa7fUTUoxFDZM2v+mSyk2pdm19jLuT6cCwErDWD/0dFt/J57CaQ
gQ5SZ0pvvp4sck65Tic7W7/kNwVZwxlkOfORteBZID+371Le5mBJIuOw3pCul6nXkdZvfzlKtZfe
iXlNFJwQBrqPfrQeXGTRDXhp+fUG797btNf6LuFuBPkGWdFoVats7259hX9o/Io4Hvh7luJoC2yZ
qCJLP5i9g8NEY6vRXkz7MJUyG88ANoG+spxxo9uuCMS/oXKfqhVZdvSktiGfS2RDwdo0JX/TugEm
6vQwko4UnM4yfT/8TfPRmqd6Tjs8AFgbJ93EMymykE4IgtyXwPI5wmnWWzsIoOCILLDEJsINiOgw
PsQFoXN9mJQu5eH4uaFSE0IJueIXv7X7OObzP06mT5xB+y3RgdxAXgJQWSKq1PG74NqKIbHr0fom
5jPgiGfhbXJtZzUgd1ZAzMHm6GCnVvXEdmLdyc9AgefdHlvpEA51BPYwYZrapzzgknKryBVDjIDN
2mGHP6CZdc2Nsby17r+u/flrlOgfEMiik5SPHXo+T9Zkq6POgpvimVXJDlvGciwaFl/6fa/qrXxl
h8nAEin1Fg6XBy2evDQrG+gF/icydjRbDNOt2VpRswSNv4cH0qr8L0Vjf0fhmMyoLGN70LSRaWtT
oVoyEy+LdF4ERXJj4owNLKSJoPaSDDcj+0A3UddnqhXY0SIMKCAAx6V53xQVLqEGFSDF9Id+duhR
zaBeOi3cLKSn5hBAKwK7xUVAtWs8Svm6q6UZCFMRHtRuxXOeBU4KtTEnHZuQjQ7yU938zx9GBZ2k
rdM4QHx0uj//uiQ/Qx8Mq5acs0Ac9dZH0iotWCHKQSF+w7/gx8zB6tuNhUzi/xR2/mgUAFZKAGhQ
yn6MSEgUjbserXOfvNx1jyBhfvX8GQZMovhvVVFDuyyDT0lbY9Ul6tEdfZa6kHpTygRR/IO5gBUh
FSJF5b+TBYCFwMrlqWoNzgAiJ+7shh3aO9tNEHYWWqFNSPDM7rrU0eYwy3MmXqMDR6+16jtYwWPb
AoRNn0JujKbOtoQHeL012gvhBYd3BYnZaUQb3YOeGUh5CFnbuaMHPC7gGUhyDqwMAjWljaa8cC9d
obTgcs+R1OGjvg0bLtqCovz+dgOYdU1OIEdKlTafVGzWZ8pPE3Q15mq1Il6P6WcoH8ohvWaAx0UK
NtGGKhEoGdhtSmADqaEBy0sKTQ9rgHqY12Wi/mkgZUWSAm3m/gxuPnEmoB1/P7g1t/kW/PidDnTl
RnhS6b6Gs5qW8m/+AwAeFaeabO5lNzXYNa1y+v6e6PuKJiLyQp/sy39X0WfqrvkC1Ywwb+7nvWBK
8zeBn8cwAQseaip9BWV6Dx/38wgbVjXOtTaFcaZ/eU1TCB4w1DjIWnLsajgrUXIUZBe4XUXYq8Ek
v7KcLrhkxqTohze1zmkLhWtV/tmNWDwWPIxCyCCQOJXBU5b3i7aDairp3Tzg+YTV3qm3kFEPUDgz
lyAaoJhdh6cOIoBmkIBrNLV6GxEDhnp88db641utOTPS4fch7Wel8+805VUB3ND+5tkFCSCUk0in
5zS0RXX/6Y0+z19ajQezN9adETBMBAiGb1FVd7wYJK1sEDQMCpBbLGK1GQifJUFrw2sI1snDVfMt
+pMZ1YD7RxG2ZfMwJGCUIILirhAbSuEm+Gp7dH2eProZhiWny2O2z7MBoLwQ7X0CDRHgk5/rGzwo
q8ikUq9xxeG6s2kLTEKWV9PdenEG3Cag2zQYgb3R6yvm/xygtoIz/Mj/LWIDLf6nyFsO5Z/cj1tB
RBFtr80ScIssY7L+tDyIICoAPSIN8q0IgI3BbY7sdkbY4me9VEiaMK6wamL3rImeZ/wbeH1nZScs
bIdJc7zMF4ES9CbYsfnLNSi9QAK0iRttEe/TYmrjuwdPy7ykcx2oBHxJsnWR+6WTKYd9PVtc5NL0
P7kKG+iHbALWTYhp3tNlRe4LLAigOc45wGfZMg01kWYvoWeHyqCT2VPcOvTGn5tGDVfHNpmO9486
rezlFb7CG328/O2uArUjyVzAfv+0Y1Bia08gC7f+gh+BXQuNOqDssDE+jb+xrAv+t+FL1RhHOcga
+SXOwq+INC6MV6sO0vBU4LxO94OXIq+02EOjGeyuiXNj6iN7T/vgCdrJhB2t0RZtkJshPH8XxWrl
ON+ouxwJrI3+E3w1ALn3aAfJrphw5t8wDd9kQjn0PJnK59QO01EXH9KmDtzxc/DYKOebkdosY9de
dadm+gds7M2sJtfTlvb9B+Av28dJooRmo0C1+bVjdykWozpYtvRR2NNLeax0hUqBaYhVbSCGEzkH
WX+2S5tfeXSQc/d7VPiDVib0zYNSMNTteEa4EJc0VhVPDqUPIWPDpCSftZUxTNtDEsvGy4RBBPHk
4YDqhfYbPV9bywnnSVNvK19i3nIt9oFXQkxT21T4RrXx5oYMDMBOlJTq7q/KR9Ecid9GBnn7uu5D
eQv8PwArpsgFkDwaiXMTNBOtbwbwq0V2CZ3KACh/CroCPrH7q44pqOiUkwkS8J+lDIKUAqqMZYMk
jIha3y+8InylS6NHwbogLJlEQd/bIYW60ROdHUIDvMxa+H/hTHBOyzVy4iGaQk71PmHcA+10pbWu
sRHSpvAorNg+eP4T6Rgk3/YBT+v7FveVXHWFNrmT6SYXjW+JBZHXir+rwCeCiL0jwIp3Euv1b/ZH
8qEhaaD+aXYPDhp19FBpCvrYdPsZQmkQujPeNhRnDeaXHQo4ZN2n7Cof2A9nVX9iwTHJz//zAT6n
DEfO3nS1Y8Ogg8STVNscVdbQivtVJi1Z2ffggCU1uIxhqn98eq+YcoovvYTsW3dIdsYZpeW5I7Fb
DVReCffpsomOqiZNep9wsFpOiVXlfew2rLqNM1N07IBpgzml/jB2tNS6rvme0SzTwyHXlGHUu/c0
Ey2Iqmp+Sd40k/4j2kMsLTOtB//lpKeHNU0Bm57VYeb/x6zDBYtCLJOrCGZe0xtp7Q5wny+FMuGE
GuYhzikyeLgsrGoMIO59Toqz6r3oM9G9x8c2BBvfJMGEuRY2BDBDCrcC4Ud0BwqZKmRBbadeWtq5
dP92c4lnFHqiVfn6GMu5HuPFZEvyDlLtsVbtP7zln9d3R4lkZn/FFZ4LWCJFS3PE6FxlKCfPAxNx
paCTU5ae+HZRZG58QvZsIYDM5WzQZFWxgN0gZk3xtOIuDMgHIPi5Z4S3yDpo1mtuF+ycOk8a4gpa
ufT85rDAsadKyq8xGwgfci7ehHZmQIYddGhw+T4h8pplSMPilj0EVCxQdC7/bROQaoyRNMLYz5xK
QBGrdpooFmmhA7LJdjtqkSsiZK1loXrVuD2sJT4HwRR0qhIpruOTIehlbMrsZYp74gxKhuzW8P+F
6uqwnry1LKXQiUIYJEtbVd8qXpCWQF/C6+nqfPvexB6gb6x9GF+1n/CBo0IwWwXOiaprOfNYqhjf
1dk6mc3dE6nyTqwLg1mt5OHr0rYmhQ9PqiAqOKqNsltruwfmIjdMg5F4jh3W/ASlJvXGS8Zy2w5Y
GWOeh9fe/dfVd4TfOxV14o4CVEU7yIahyyoDgUQvIEvK473bnY6OBt/2RchLsTP92RjtIPYT08Km
fiOIGaqzD9N/4FSgPiJV7x7OPz5ISlqm/+XaQAP9Uw61LKhv2MpDucd+R16vkrec/2AUJDBa93n3
hVHTVODBr6ukbBghmjRXjikCguBsiCqX2oObRpJSKOWrKlMxT8WySVsJj80LBrI7e+B4x65ExZ1v
BRJZRbdm+XP8603v32p6NMQHQ3l3E+IQAwvFyzJtqXGzwM5zJJNojhKkj5/w7cYqJOT/WzB9++we
k9LKyPuuxthxjZ8IyAICsF/eXLlABVjxsXYWXLCuD/38xMJM+5f+nB2Yks2wy2mY4QkbpdlIMuez
6k4Ik3Lv8VZjdcS1QHYIj2E8942LKUf5BPPCSt3YyDvB86HJEOksBWS5t870t171mF/HFBtHUMzd
C8xlFRHtGekgnOQIOinXz88ilq4KWQ1E879hCX3E89JjWRxyl3pGU4Wq375zhmTm1srSDdINS3N4
Q3FlCpuaiZ/wqLH33m5m3+5lKfBXXBKN+mniGL60J6OY+CTjqIPfqAOSEZ54OQ69groPAOkLJrW8
0obMNnpJHEMvQKSWX1a6LXjyNBp9gjA8jPoQs4x7wQw53l2CHejBFiffK3mIumJ8vIHil3SB5eck
1Kc9lpjJLy0gLgEBl9QtSROM9GX7ZXir8RvcOTJ5Hq+1wNUSzHRPehVjImi7M4dLhN9yh/CiS4ZB
H2NauR/m3rfhJWYYfP/YFJaLpeM/MdofUtGaQ/H6fQ0Rie7lD3lvUiy4IKcBbB4Ke5hxxUaMRUKG
os/JAzVF6ugrChLKKChY24yqzXT3y7pUv+jEDJSEFjemxnDfysN+yl3Y0eH0IoQKAjUT8NMxQwaE
TIO/UJqfDKcldZLbbcWcu7kBVOrZojswg5DPRBN5x3jYqE2Lxa3c6fZ4hoKq9Scw88/Ka1BwMpwM
VhPpic/NwcEr71bAMt/R+z5NOFuO6YvMqJ16gOSMgWeN1YbE/UlJJI9VE46j2nlL4W/mwP459gJy
8nFVCZqDSGE3T89azrpXTp9ubDNh7/ycempi7G/v53T2eiw/QNsKx+EgqtWIPok/By9ly+kSkS4h
GcutTnAQ5Omeu6j3uCKsN8h6qfN8SpszCYheDK+vSjcuVvvQHz56DViGlc5sUxwCRUcOtOyCQM19
T7TDoUOiXQU1oqN+li+m+wiUCDEWMNIADeGvWKeIOWzi2yGTyDdys9VcDO+nPXWHrEmhy7weW7nD
S5eQ3HCP/OGm0tYSM5lID3EBzhzDfYx3CgKIDWHelmJg9Bmtnf2bHTb9wv9K3vC3Fit8kwE7jpOL
tmxPvjU+++WxnSUJhHQui0ENvg532pffsGYaw9fVN/AmEXOpYnPouL+1GmWcuTIcgXaPOfpMQrcl
TIEmZuD5+25xkJm3oAEhe0dDVjVaXj8mQgVecKF8LpOOBuBO4t1u1V7R2Ke7zrmKfGBHdH4hFZjS
C6UP10DAINCfW9FdqXaMb9qNNt3bIXc9qze4K9CznwYyn1mN8DDoJEWpttVcmKlMLxfDy+J2L+hr
bI/xtHv4hyBcjODJAfLTNIC/8dw7bvOB7NhOGR5ucy/YG/CtHA+QagyZqwebtezAYUMJb/csN4Qf
hHFTySttcHApNYcfnpSH8twQgvt7/mpa5dEC5tywloyR+aoZQeXxESEltIhWBXfnZE1hje+S46ct
GbLsCdwFCMdRnjaCECi9V7Xa5wwvGXLekxkGSHbgO3sRMqxdWwWZ7vSBFleoGzkyGuGP9qcDYmSY
6ytH7j/gzKPlwEx4XNn57QuvnnKfgvEq7d8M9D+8g4oxXyg12XNXzVFkhpSiYXoVi3Gl1RZri6UD
+xDbsrHPwxB7z1Cgjnfut6KApO4UwIBokV3iljsJ2wiziqw9eVGgoFaHuZoUCvqbnywhvmiG1F/T
p5eNdAsNq7Bfx1tMcQSK+lcuJj8PQmLnIzbMVHyil5EW+J/6Vl5MPErk0zpZ9lwCQzIHkgDyNjZA
gDz8XuIPQlB4XmBh1q5bIEGILsw4aPoF98F7rrTaMBmhOMlARw0qvlZIgqgictvvGA+HFDEPu3Tp
SXelakQEZRYgEUx96krISJqHC+ejVnR4fYTCSA7AG51nwVX5nj1FR8HsqcH5Z31eD/jzO49zW40o
CPZqbKTEny+e0wul8wi1LZd5VwIMlFT1ZiVAoWZnNrSkqBy5MBrRxwpHcNd5jegi2aRI47ube12u
ZHfogLNIj02521Firw6ltfe7Q93nFkBeSVZBUQ4aKOgErV56O1Mm69Lh+mzod+jcFyeVjg5JZnmN
8mTwTNgEAEvKIZVbOWegxOon4ZDoHI87H9mVVfaDJKBMCzsuPo7nX8i7AfxaEjxs4qa/+7NTaZr5
j475Y4lwCBK9WPliy1lPD1rcbG4gjnsJWLxK4RsdB9udwR2K7v5hkLLDmbm6qkU3zveIqV3qZCNn
0fSYKYnBigNarVjdGMSUpeSxl/lXMTwDIBLQYUQ1F7DN9Ndb68DSLM6UA2U5AiDEtbJK933GX45g
oBOdNNoRVMZIHbUrCT+zZ+F33SQetkqJQsG+XoBZbLMgE+uca3WNnV3AXwIhUsf6ej6f1mGQJajG
ABEgqL2s3bXAABg88d0PUl6ObExLhcgnUdMRH0ADQA0v5A2qtGmq0wKCF6+Ho1t6nNYwEEjSzidr
YOMMAe9M71J3oX7j2F3xjA1krxSKUd0qnlHpFS2RTNMhhDw+73HfdUtUZ97ZbMIYC0y4A/wD1nG8
LV/bC1kXk6P/cw3ouBz86cnA/qJsTyOSpPyKDTnQMjjA998wjo8NN/QWKkvyVWyyKgdNQhzWzB5K
M9ZXYH5J4K9H8ZoRzwZbYLe44Fon5XKakWLJX2VqYELQFmzoKbvip4L3rjRozixEh1wbEc2qR1zd
0/NuDfC58vrBAkwfhZsHXsePSniyBteBOy5chwPgzKZwYils2FvRT4RzCUMjyxWdKAWaKrqmLuuy
Dka8zhiQPrdE3aIL9YOe3hyr08usd/IzwKWwtN4sP5VcrvR1EWiBK3aq1ljJoP1sNR4St0JH1nXz
dYyjkjU5S761SLN/tn9mGKqNZeYor8HKuLE2ZXQB+52jZHTq87OrhaeZT6HRqSym4Jj8s8xo7ya7
d7zfFTwNErbA7GXEdaqKQrzFn0P4ZIskzJdbX+t0A1y8FXOTfrPj8gOwxjqkXg55kecS+NSJDNW/
Yfu7Fhb12v9d1WY42ckiCAPEDFi29xcGOCdVxMkQJB/kxcnIWs+m9QtNRpn8Qyb8WYOvNbxv51kk
fBs/fnqaZBozHVMkkMAJHjRPRxc7qLIecXxbViB8tdiDV4m2l1F3dBuAHP3JuTIOM/x7p4guib5F
fuggtn2aZ6Hs3W6YJ3xP/VxmjGOuGGUVZIjDapXP/1pyir3rYO8STC6bLqgjT54RBljUIDeUnGep
iitVUupdyBq+G2YhNJ2dldTz72doum3+DrO7vxKhwoed9jFQr04HKG52fVb/x/YgYFFu03gftilO
Fx/q+rCK5Za3jdR1cCts2ZzqYzPJEIJreTzskByeo6jfMj6UJD6Tf6tZlJYQ423k77vlRrr7qWyz
WtNJ5w+gcnbrXXK337DLB5MnR2DUEBuvNdZ9MOSdeWo4Me8HaT69XClOu77eBOYcxH+qyorfy1/P
2kLBiCvRHneaBrqPAfYC1dy57t/mEdPQ6Xd3xkdhY3Xa95BdgHmgoZkNYaHflc9lc6gP5oQ2X71G
KkSgk8F3BJw3Ma4n8vetJU4fuXQwd3PK+rOPXNmNS69Fs2k7qBK7uxtTq+/GfBWjdwf2nuvRhLcz
bbkpdMuBvYrt10oJ+fh1OPj9ZCj7mmluwqQK5jtgwLb1ZoEln+74FjLZZkd7bbS/cBm1Qh5jpfG+
NLgyWX3vUl11UumQ96FWHZTRS6E3fl4LIhVp6AR912AUrIjrJ0OMz40n7//neK9/GyemqWOWjx0a
+gDZh+5rmcFlpWSGJjlGJWV3u7/jHQzF98PXmQzJZeBTOyVkaoqtdlgxgY0eIV5oYlq2U6Hq5DOI
JMTs4curGyoilpKTSxrlW35h1FfR8xrXga7WNnvE2rNUmbpjBHms2gvCoo8JdH4DP119z9vnSQSC
GQHaBwpLb24rx6UBtsGTAZP2VerLkiUYITo+YocGeACf5/+GNDaiZRxQfj2IvIYpxbPI07KffmtG
/Zw5Nm9WDq8j/G8fInVnduoy/mOeMEnW5fa3VrcTpyTxYE8aKSin2L2WH0sAlDLgbebHuroXMPH4
+Wf2jWISZkJWAkhMNYNMGqez7WEYHGE6no19g7nk/BzgMuJVReFznrf1Qio2k4yQAswRL9i/hb/5
5yrMTQdQ2dFJO2tnvhDhTloTueBETai+L0EOuQJkJuRoZzihf4OsOsViOf1Fw3P03Xvkpo10MkTF
sFsfXs/KvASek2HRQ6zbnpr6v2+hhLA89pVf1Ezf13mJ8qQ7BMVlf3oCizLFANIq9OKJCMm6sEkw
zCEecCsNEo0PaKHG/sFUTHU79az0wKukMc1q/i9p64hdZ1Zdu3UhToyH2HkVHB4CmfLFfPz/n77F
IbBiJDzzK1W4n8WdVhbW1RKxRDlLiGZqHR7qU/7JA0pLKD0DQJXLpil1ohj1H15whvczv+0/maLA
/vGLQWH3xs3ADlODqbJC+0e5rtC4xDmj56AW7yP9Ly+oiOjgXzV+QRJo+8PLLV2a1FEoOKl9dfHZ
+u0tdd8xLBSL0imvrRgqtlYX+qCGNHJDAXnwp0C6RzBeQUONR27jJLukGs4FfeMoj/YlMZmwqUxH
WAAmg6tLyE176R4g5dJpi8RCZgNKojVarSfj2c1//6FhGdTEYiPf0rkOOUquld+JfNoagZmKd/0s
ri0rdXt60veBW8u7CL8my7ZIXBxAD4O4aPhSRVjMM5Pvqf5LYbjxiamQ56a/ExTw79+II4HiZ7c7
HzSbtuew4fJHhRS95BpK4jqQqg70s3dgU+LUv4TFx+Nll++dxYrijybH+zxtv6XKaQT7rF65IRG3
T0WHmbuYb72LxVRVojLZ2PAUpp91KSSAZjUA2k4JpKXjs9mv5vkJPtZipGr23AGSUWzQ6H6cZYCW
P3HFRQPmJk+YOyXhpG/7BIfXJx3csocCf+NPYCKorslrosQ+EL/kj23C2YHPkzFzGdF3Al8EoqTT
BRbk9mmQxNXX+qF0j8y9PwLiA9lcGeUXZbSwSmfB+/5G6rfuD5kG2+YaKZoh4pJ6o2fCHuGybEV3
cCrusKjN2IPfURnTpYZ6fXFcus78XYEhmcC0KX8Wy4h5vPA1VQI6Ihp2nBqXY/klQ4Xn/Swl3Cxu
ksimMs7xNg5lI/WSwDtmGWqHVhUEen3p1l3e8I4dbRrLxGtO+QC3HaMKemSz93W20BwLJArCgdvr
DZYJ+i1Fkz1aca6RGnUdi7dGd8RxMKC4YRAJXd2RbljuJL6vjZkOVW2NLE2dN82f+hM5VYWY+b9w
wMp69Qv3hJiZxa7xbGttMxUBGmCnXsoQ3+iIZAWA7nnh+ubdK9exJTUQtfNe7ZcGjaUidoU9qBSB
dszPyEMGDpCArSKOLsZge1u/nCQe4ON7YST/1u6OFBr2m4699hTuI+xcxEsCAIgcWX1+FLSCf+hz
Ro3y5tKpjfhZfTuEicigd9Oq0ZNbCVSry+12vIHXnxZuL8kb8ZGafG7b0gR9nKdaoLoYRMIqcRKR
TSZFbnjl9EuRxfbgFctrWlaA1nH6a8NQxt7dcnuOrZgJuwj9mX4FzhtiCAPvDLabUTe0RraD0Pzu
gslYCpLUb2mivDDzCttpPw+OrhG6Ceq1f6XcRd80T1gJo21RyHZXI0GVO140ZIE3FK53AjUgaHUr
BQA8ekKBbfx4Lbk0W+CUx9536Qo8Vrno58WM5iIdpT7LhpSJvF26DBIti6pDTOFY8ATl51FrZjzm
W1PUYqJhzcrmvXPfUC8EEIPfBXDbK43ZXFpE5YrIPcBX+kiuZZto93BQSPdZ3OnwuB+qjUIDRN9a
WgrD+CUMAVfqp4TXXpvaka3FMWpUpYbjt4IZWLBNHfHBYJdLbJ3JYcjfQB6GpfjKzI+Gq11UqAfi
q7L7t57Dz1tvBYJxUj45uCj5SUp5HyESjawwgFFtgXNr55YbxxFGNb8r6r8O3cHNM0/OSeTUQrkS
eX1XdE2qUFN/+irAfzFXps1rgEGLS7rg/GVegZVGIlbejTD2buohYruArPKnNtW2Y5KvaI9at8d5
lU/1IKRfRzuvy5bNe8lBJhldCHwy1WO1UuzEoOpvZe+vjJfVUpRmp73LDVRdORVeyZVfRyYbwZgh
zecd+DXiSlKPtzT0hOuFQiY2tiEOzZ/jdfcjuxA9q9Kxd5A6wUDgbBI6azk4fX+5fsZ+46CYvEkh
suQL8dADZ3RLBqZE7jeDrylytWetKM5oLaJV7vHuwZAbpfgKjzb2Hv6hOtl5sWcUyQrnNZFFxE7I
rHy5wXJV/OuwZj/evqe73wLyoSKrknefrFMTzqgZWO//Qg22xcIIgOYq/3rHMQyL0+l/OJnVs9lE
J2/zYH14idTnzWFHhfJqUwuFOBlRGz2LsA9DlbDVF+XJls2XAY5F8336JZI7icvSKIl53obnWbk9
Yh9i98WzjcYPKDVlcOeVKqGZC5b+Sbt5ndp4IWGzXQyKS89lNff/HRWrqBqwNF0jMIO4R7cp8l16
Lq7JbodQMq2oIkrIXU8ThWZu6vULweRx3Fpcnc1pM5zqjtVgibsqLtJZiElOqz9DI+2CRKxL9nog
YFUDvgGdLSxA3BBWXBOSQQ1+cUshm76dLvu5IiE0Xc0n94EAm5syrmVyZWV0NoheQsZ7SgGh6e5K
oj6HGgv+jQ8HghO9Qjp1sZ/Vstj4QdJsWJA79exjrgAP9lOok5e3Cdl4rlzS9x3JhbOxtDORIFj2
dANIyqd1ZCnY+wkW6Gu9PEMZHzQ+jtxyTcmRTSfeae4gB+oUOBGuSbyePO3dYvHkh8PNofwOypKX
StgyNd7PWl0m2XAi9AsxoL5Ef1Dg1dBIs6Bri0KyGwypybqhK8gWSXL+8dTkjte7g+ydiynt1Pg1
9IPwi5+pijspB/7TLn5eib818I/z5QYOo2Jh3ZAiLAB/XyLj/BJt0fp8HKDJVWBgP++FBiXrHPKU
a4O3s93rvT+suZbjtcwdCUUyvypgcCf8XHK3njsIIw/dxBrBtIBzTKhZqiz9ph/q5ZfZeE4/8koz
KAGxi+B24d3Jgus4BiDtrrNOhldXSqbKgO3V5HUSROIExwgnxCrwuQs+OW+wIhQ9Yi/8yGMP8ZCz
FSNOlqDe35uaEmO73qQvA9Eo8cjj3TGvIYMRCrpoC8NPE4ptd0y7I+im5bRlm8omBUJXa2QXWdBa
d08h9Ii5PlrHOvZmyiItDYGhhRgAZNBAVmBiOF6l6CPosc61zY5/nT7EEAaoPC44tJSPGprpcAsx
RJWCoENGDtdwnqmHvoOp/c8DdHoAvn4JrzJJop/WboghfSDnxbUO8Rjk7ky9CrUGpc2q4VGM/z1G
B5xxnOG77JDwItsOI2VuCoxpLplBiFS0PW3kfXkc+TIDjX9r/GTV0LgHE1yMQjn/cF8ByM2J/xsh
l1WiSk76xFRXY15Y+O5ZbUiRHetkI5KnwOSvmiC6bHFGqmSyyyFd4CFHUSKKeJinrdcNjSsmHC2s
w/5HWIpy903KdrCVb5dmPHvlC/3lFoCLBK4PcV0DnmtloQb5yPhsQXMlJMB2ox1PKWExXHHcC9Yh
B0RqKvf9FUEzZIO0k/U6xJ3j7z8NoUf5gCx5pnefG/nX/YWtSqquKEZY/xfhLCRxpFNLjj+b0VWz
0+6q3zt0AEIOXGsB9qYvFDXulF+pZWj8ZcGsHy1GhfYr8+6kvlbdsH61ZMAC2f21VMRxwOk/a1EB
PQ1nD/MQWLEPQtP518a7Fdcfy5InBNjDZ+aeRLcAY6LNOmRVrQ+F/l7OIWZMIE03OKKuDo+r7+qS
XamXLT0DJ+w36JiPgA8t5pAAP2qiCTgoAenRGKuftl6jdWOW6fVd6dWUjoNnig94ZaULnPECQ5ea
MN4FD08UJ3FOJ60iSSzVMkxn0cHt9F8pDhemLH5XChC1YGvzcE1Q570/06Lqu3tm9FgcHSka6CnA
1Ry737lPndcO5zRAC4c2U5wLl8XpwKdVnmUK7ewLn68hUINS0V63MvrQ7c8e72aj9DIZXF4tAimD
f27QsICIz+diM+b3B7rNZq2GBck7GxtZAxW+OcrBQ3OgjKQjEQDoYnTBot8dPYEDwE9/J0chReyf
BnyR9v0AvXBj0+cOwVbfEVPEqlV+sz2/G1XQSKWDaMDlkLgCEouUtjuEyipyXreKusMrTpRYexAF
McdvUHRVY9PEFo5+eAkPZ1fIqfzGHuKv0MznoTeAIbUtJQG6ej9hX2hnhx1D3XVh+dbIiPc64Qp5
NG18OF2Pgkq3eILbOKQKMsLMj+pKuT7EkgC1blBRlXYv63LZ/hrbHJWwy/dIyBqqBRMEtXq36hfn
HkjS5d0FxKmV4vQhScza91L4EofMKsVllC3KIOyasA3L7pM4E4hfObrnADdvM98hkgCDJIWAkPmJ
1kBZun4BtSx8jk229fBAG2UUfm5I/v+a1YQ6vxBCPx3oRhPmVIcEUOUEtQwx0vEeXWbeEMZSG7ro
8kLXGzfvdNFbLK9ttq74/k20G3E4V7ambzygkOwdKAKdRkh8z+Hc73Uorb19Vdps/AHNxF0hm9K9
0O532gsGyCFurS2CatWKzhi/VNigqaCvVVCc3St16hV7/TIwhBf8/AY8tZQWTranoY74VfZnb09z
ESVB1qldA+jk3YTvYeV9AETL9i3ZIcQvpQirAyxR/+IunWB0crWmD0vFVjotKER+p9o1o28UTTSX
33cYxTGpuw3Qh7mtw5dqVNjCr1j7WDX801V5QJBvTS6JsCKIKTA9aNG+/uUNKiEBHUFLZqd289He
E1jCpUjrcN+SzrG2WIu5kRXFM6tRm2uvtdbn6wGsF67cXO8+BLA7BRRuSNoE9b6Vb/sbGZwD3xCC
43KDo1tnNSgN49gRm/3AcUPyHOP0dMxSmfz10CECk0IQ0wRvqJbS8yLun+xjnK4k0lwEXSXJqTJu
VmvwtOvsNui3QRaKa8PRYfCJFoUEDzUdAptwF20deiS1etL5Y8crIyDoFE5/mzx+IktbPKEPrpMU
N14ho9MNEgtcq2SSlTKJY2Z99w/x1i1bU0Ab584rrM1ShCrtSgj2Spwo0m7WKAp9q9As8QHY2wuV
6oKmPm+0AOlkAzR+7vEPXah8B0QSN/JdriCK9Y53XaT4Hl0kp1uDxMnmthB4ZBjboBjcIboQQv0F
RGD6V09XHqqtc6fF2GaaVvymF+PyoI+USDzOdy0x0PFsSDGHZj2SiKgFUqK8kH+qvhm8sSbJnLWI
f5Q1HSxR6phNQzferPZZspf5ej4K7s3HXIrfqhhzGKsmuMrqQzST/bWSdfeECWqG7j2zb/99kdPn
KJhxV/NZPbveIL4nuJhQnnng4YpuoQP6otNZpB7XcG4yQXsfHAKj1SkqbZ1JkpKOC49zIRmhtJWQ
BSPo8n3T0WEqSYQiRRDELX6+CzC36z7h60sJY/wGruVyknarKWLS6k932Oe+t46UTXsf+II/i/GO
Gs+4Uhae5t0WkpRon/lTk42c+oUgaT6+7Cwtuwg6DIlYfFcaVM9ZUzPKOari6NbTvZD+/U4xWgXm
uX5OrOV9c9hFQeW/otM9aRBJFOXootTzCuWW/CBbjX8GT0mkX4TnI82cBldrTSA7nlj/8RKonf6N
fjXjXYIVqSPm//KZWEkTaZK0Uum3j4cZCqnvSZfHgwA0d1fJ04cOgMOYV1vCh7Q63YCH0UfwIwav
Gojxh1toZ5ZUTBCaylEqMa0lAvjpAmZ+Ba+qIqpQMFaHzBxC93oSIQ7Dbqrij81TunF2Y0FTtztZ
DLU6sdXQOag+oqIjpVluRRQbwCLUB0wMawleVX/YockRvVyvW/TJezMIJPri5vPOfk7BoCAChy5r
CRmu3DHUKReOWgyp7EaD5QdC19f/5ixUiTxw0AcydzJkMNSNN69Ym8p8R/fpVRkEA6JAHjBr5zM9
EKybXHj4Bv7DoryHG25yelSY27C+J2/Bv9jp04x1KIj3g7ftABk2keWx8TC4YRzVWVk4LOeEfK1L
cd9pBr2Tr2PwJ16s4wbhPZr/mcjmcoSC8Vwfxq4Sv9IdxCtiqaB3pc7v/lCX6nVwZWo18JEpkabK
clRpXYf0y1NwIGTSFOJxE1dYHGaH/VCu2lc1VB4v/Zawy28SsVOBMhEksLYig9Zcc9bGhBDA/wPS
npE6/JVOBJyvaN3BQP9cfR/Dc2LVVPrX9KmOnUOJi3T8qurYlCsGVKu9Z0YV4O3I4yvD8UENvQov
99O40KP8aiqbWl5swxXwDepI3ve324UudLLiO6RJtKPDm0owgb14HnwrHI93clWqbnbabxSqwo53
0b1zPjjuCT7THRdURtCDUyV4h0XpGONpwrnk86sErZOBlKNLwr3u3OHByiaM5vBI1VT13tpMOiSP
C7QarSDKJI7B3CfRQ2dqL4A0xBFEuVBNteUQDkGBHy+7pw7Ojk/Cco+pqmraQhSTsJJtqeCvqB+N
bZ12Kek1TvvAr/WImjYQAbyE6/J9dtKfn0td1FOBR8mNX0ZZdc7yt3Lvm3E5+/Yi7kUQwcZ8oox3
b81/+nTFQmEFBscujNn14sZL1H2MqHJsrYNpEFduEzM/OMy4wmBydWlpcPvhRYQwURPrV621PJmw
t3MGxkbIVakazm2HPiqlFGawzUtbUYJFoychEo96hCCwcZMoFdXwUXh7Lsrlpl7rm3P14o2Mvi4H
5U5TbSO8x9KUic940f5pWj0O+QfO/HJpv1D8irsuWqC0UEW0XdUqc+QGzgZPuB4ZSXP9VJ4Ibxwr
ckLhHYIxXkvTjFwHADoopydMpkj/lisVjf5bXvqcKvUqhNFKUVhwfXWtuyagIWGTq6gdfjhFFReK
AW35bNEZcTILO0uTLHUMuCxq67bJxbWfFnwjFK4AW2NowlH3wPw+noUuLzO+9su2lWN02P6XWQaT
la8OzmjDjvKIizEABzrg9nrAH05Knn/u9cwtC8SaZs3f6tnvjOycNX0S65JiMnGwqVSvO0aOych+
v3sbkM1VWHZgJPvM+0lmD26bByb1VsLlBr512ynAfweD2OISgl/tLtp0IN0eaS0dMZbU66GvB+7L
mTXtLRTNB18j3yJHNaR2ToIuNKHCMaBRYDhJZ/+mx4X196CPDQNWXHfjHV8jDd7PYixonNmrYdU5
j/1AO95BiF7NBP5CRisI3XyCpen2HSaGGGpspUoF5C07Oe5kvLgQm0QnQiyfykXkRuzMw+0I9Bwk
Dp+iVRL9mrmrekG/AMjF7YSskRX30hnIdPRdvHIhxuruAd4p+cdRI/TflRTIFmukyjpEpt09wlk4
pr7iYGw0GD7qHpMzatmsrSaDzERuaV83uqKg0R4enNuAf2TpxfV6EA34NwyXx/pljKlK6PKfgMt7
a19frFrpqkdAXxip1fBIAQP14W6IbA/FdHY26Ru1/V/yKgGDLGp23p4viKlmveMP8rEEJFIrH5Nc
y0WxWSVolxjPvbk6CWWh9QsXO0oO7SaNcuNGNtnm3uonyHJ/2ocT2i6a799WhqUDypln2GJrGhnZ
47JgQPjU620+xRp1SKMynXuhhrWWv6Ms1jLwCz29fd25FObTmdaU4ShYj6oE5id/aLkfSRNGtkfB
DufS6ATdxuRmpWy/YrRwG9KKxfYdVT0KbcoA6mJWY5Sm5yhfd78dWyh5ygb1EQxzDtj6eaSncRIW
MV7eXxGJ/+Au9QoLzKdzV9MrOYrYLW3lW5us90xiZFeWKK12VbNlX0dyT2HYxLDO5OxnzpJdwEWd
L3HlNjz2/6VbHuIzT6alSzOkLo9RQz5AksCQ6cq8TUwm7lPdF4g1OIJicWtL4dnLV81UOP4C8qqJ
H45kOzlJPOZuidkccrYlRhuNoGJXZqQV0yq427sq7foMFLNeG38ef08x2c4tIziMUoB29wx36u6Z
dhk8K6S7hTP7jXUNLEZQbLGTPIYGNI6nbQTIC2JdOyI9xRufQV+mj1OTb9dUBRz/qrzDpB6kBilf
D0KzlSipYbBzTQKOurJBgNr8oSm+ZxKM8OYqWYHWU5JPyB+uCC6mw7ErjcgttBicrY0kNEWjPOFY
nbZX2g4fO7ClVa5ml1X87YV+XlAIq2V5VHuSB+s0Kt+scNdmK1I5zZxxbU7DYI+v2fOQAvc9MCK1
GUP63o6nGiw8JjP5q7wo0N83/lxsk0dWJwGQ7vmmEoA9SSyPegilpeHAiW23ByyjKNvI8SBw2CX3
F32Z9MNtyjfqees6FxQO+EFRcZ24jLWVQ83Z666rLDpSYC6RDsy2zKdsgki6xkvec4p//bR5BSDK
hG+0Vpy6b4/uQQaQKhDIPqOOAEt5MLHlOG6OvnGNK4TazWGZRflV5ZsORlJwXlsso/7jtsDOBNRm
sYybG3UIas6CltCACv0pOWHmWy6FN8ydGXZMW/6GD9mkEyhsdVGfXwCd51mj22pk5z2sxm04DFBf
e2BmOO0tlszpV5UzjEEQwd+Z2/AUBLeUH+x9EwOH4ptHCbDiE4p83bHpPrpXHGzY/BsCx/MFQuqd
GhaC9EZ0ywW+oADOHReqg3oU0VsYPk5Lo5rxKIj8uqMtDj6nr85fYnJg0yyITEvZjTArxwEfB9iC
cFv5PT20uIFmmH+L8L4mwLjmCZc+VhRwFZeh6mqAQq9Di4oD3bKiD/1QQuG065jDj83baWull7kN
6Vspvk+HEhowAMSIJ5YT0DqTI2AArnCIsVwnhJUKynicYPq37jvT/YKLzg+CaKAN2SbVjvKTKeFq
Lyz5LUYewTDuJ0hSB4IymrEyzzmP5xu5YihnbqsHqSny2TbOZPKPW9rCQPtfJwn2CX3YTM7UPmyG
BcRD46cNvJ278nB/VHL1Rc9FpAGnKaUBmMrOV5+VKXr78bzHnVmxMtHj9DdovatNgPiKkGXLnUaC
od/VmWVUT4j6VKR1Cy7yHsIHX87ioXhAYP4r+rEqj9gN3LuamILS+mkuzcmwj6aCF1wEIVU72xzg
6VOVwjKNf3qFKLLpX80ZJCuudsJdRFhzPzGtiUOEme1rFJmhUiaWgjElJuDJfWQ7VqkVDMpvVidl
qcg036zeXR97sQ2fQTsOilf8SHRlWY4Vq/SWuQH8d0rNWMsqgPsuo/uAko1ZDJM2XYUDRkAPfG0h
s8dem4BkF5AGUt12ZSKJTH43nOsQZUD9X8o7JvaxeMmfnmMcGII4wUff/uaWxcxOo4NHy9J0Bdk0
PYpGgT08oKegcrB8lfXnWrssBEuGxsQDJVKg5AixZ6lb9ulCGMV5oPooTENrZCd+/F7uBkYgqdaJ
mD0Js8qTu+utKXQdu0aRHfk0ETllvaLLqDH9/sZihzizUXHojqxTb/2naaX6mvqqjbk4GLHbF3AF
yKKu28/0jTBOP1DweMU6Ek/99AgzmRmOuEBJTLXFAHQPl4GwPNLc5Euwi9JD3MTbcgswlJiGh16a
Xt/Oge91uRW+pVfdf+O3Tz4b6qMIPvPTvwYxHZCa10Rszxmp6+usL/tvALQvHbIUlJFr+VQvTSmp
vMHtQejnk6t/8om5/oaI0riLfkhqjyfUX4XgF0ocQ/NqHSDlfYqBU3xB93eEpVdXNUNEgxJoX4/g
yQ2wEOHHGrxWNGLarxIXVsqCZeRwJ2Sa6Dm/b74i7Y+twD+mEVHELtORXETN6ex2SxaX7Sa70DXw
zi0fGkfzmI0fvBuunR/2XD/uYOwIoMqFMQsoVwKtLkOjkNIfVUkehdH062Cs16RLvvMBPPyUf0LS
yaO5oWf/lbf6JNPiFuWTHIMv4ElSZKU/8hC/bVE9OWCOhyWnw2DuZxTuRrWMCjRfLw4wesZmsdWN
LLaayMDX9qM7IGyJY5d4bB01PjCtz7+BjvMzoCEJqw4C0dVgzH34YJp+JoiCT1cTdkDF0sJQoBI6
n+MCcMEMjArYNcslifJyb/1N0FzwogBeH9tK9KWEP+fDysok4wA1h66Kp+hAzFqnBmdi8mP2eI9x
XABM3pO6McyYAL4suXVahMT8iS+1EDVAgwo20jaGumfDsikvrjrKixaJTrfTM1LFB+OHrIvtqgju
fOxF5FQ6UGfqMzINzKRsO6W3LAHXdkT8XCVZ23IU9gQTVmvaaX+1I75Jemsb6+x1WysIehnvhYNr
uDwNAJxKez+zv+wooSiAhIH4YlQF6/NmQHDi3J3WwD1pIxKrQmu9NZJOJYREEbtTNtiepjDcmRbd
whOJGVlF+DYN2nHgrurCDHjfaoCt0X1fd3JJZqK02/MDtdfA/iEG2LfaDoi/PXDjGcZ5KhGcRsgI
LkOtmM5Ap4MmiWH1SvNeQWLFQm+Nd2QPs4PQeQxRb1NpzlSSJrvS+WRVhk7t083NbyJBqVGcKbmA
y4am0/2i3c8KQSRjFjG+7DLE8il5tc2jeU/k63I/1tW0YUk+8LRalhHWzz1W4fHd3Iydm7KWl4Qm
EGqEfu5ejdfQdyfTujMrg3RHANKlECyXkn5F2vKh4ljL0cAq13sQr9GFNhAHszIb/15niUU107y3
e2ljsrtFGWnWEb8NkdMATAG/roHxfnxcJemyE9KJk3mIg9OlEzhcaWFTZGNzOtt1fwtAHz8KjDOW
X5Gnl0HIWWZRbRC6UZpJzPzJVNvXzpkDmC+ViZX87isNhKGzmNaHh3y/r2cA++coaEjHfgLYjTct
RITfB3RyQWFY/L94Fa2m0Vu1Wltv5KxlB3u7Iuc7WHhRjx/PqvN+y9NyO1hDaEaCzQfjdvlSLW7i
MDo6/XVOwt5k0dukYcNGH87lmhzklngS4dAoTIiEwzdpgL6PWmzA/rgJcPqRtU4x3EfAnDMOrD5Z
oKYFD2oqwcy2W00OTZCG1Nf8eKeHd6gbR5k/IJ0lMyarRc1AeH8fV2Pdfz/aG135grmOB6hsa2gw
+yRo1ivkXpme/KrSVh9Uf9BuPWkPLtR2eQSIGRoZyAHg2VUswHXJYAFs/QzGhrbFrHQdrJg8vCHD
IudIsdDwY3edMUXFKes0PO7agLYU16T3zLjXXfaQ0dfk7fjgdasBHYgF6XBL3o6rTBvkSIaTNWAr
t0soXVXCNLOWp1g7C4ecWlpY5pYEkesOdo36gK7K4gy1HYvva44Yb5pABctqv6IPQF9yJY1Nq4BM
39uIuQscVuYprmm5FB5fIQihnmhIe2/rBvOelyKL6N6W+JsiwL6iKj+kIZx5wj1p1hUvaosxecXv
Il1qx+YNfRjfstrKmPE4QJVy7HZx39dQR+hpH59tdltZow7cWTlYhZreRvIbkH9mGENGjc6iVj1O
vZrg7CmtaABtFCl0Fdo0X3GymsUqWhDAlZEMqZcyNYIOoQ5V01ZdtGZ8PHLVRwkmvPSqn26mgzka
FX/FsCT5885mo3XvZZK4Lf5Zbz3ekNzrHs1DRI2nduNBonq82zwj6Cgsd8FgAvE8b7nocK83mAkE
jx9yVL1Njicn13ftPjcIlymlvv+w7hxcPtP34mE5LpYZT7LoI+Wbh7smFXCkdOA86EisuUyUI8Jy
Da8BLOPuCOQixktiQUoVCOIVkBT6DQ31EyPCejvdhPkr8SgeHe3XKNXKxxqLmTkG9P5cdPxjAprY
Bg7bfoKF2cUr2B9ckQwfg4UPfrSvPsrCxQaoXfU+CoC7gResv81Sa5XcRtGHJprAgUfmBKGZr7yN
UKWilYC8mzjmZ5NT+GHaEaoqMpTENnsoZPUW29kV7wmBiQL+W608i/rcsuV0VVbte9zU3HdZb1by
DjXqmMeaPWZJxL5v8iuH3G8ZkJPU3g5mTeWkZ/5ypcOyXOsVRkN048XszIppn4I0UgaUIrH9l536
Z0IXRCS9RqfJOw1qZ7ZPpwRWn2QKI9/y6mTKfsW1L//yGIvs2rvARXozvfixX+7GDGdmDWvqaXwj
QOY95Q0GZaWOUFsGZw2R3MR3z05xSxD7zPaGApTvQVXI/Y5JNlPSL/KhRpCDYQNjwnoaPYCrposn
29RzkNg/ugebRUt6rmnFlv/zSYhybR+ub/FWGhSlo6puYYRQ8qqc7C5fBIUFlO8gKzyMTu+ytziB
7bO3uSskMTNLHFkN9GZT7em+p3PFeWrjhf62mj11me3Y69hWB4/STHad8mNJaUgGbUk9KiWKUi4b
vRC6D8YDwiJDTZ+BLs+hwyTSM7ersh2IsvSXs19lqOitiUef+P5qCMYDRQgPv+K4OX2vjFwylX8g
kdgZhmpfQ6menb18249jhXxaTLqShASHG7pZIwGOAzgdRD7AW0P+oDJwALt3z5HBWSWQYvULzdUm
VLmwPwQW5j1fgm+iBarpTiwaPfDztdLwHo6qAhCNhrZ910AJM6yZxAsrtooAgZLpBEfEgz7FXNhK
FiXaWfqo99NxLPEpAx/PmEIgTx88/YrnlukcXkiPwokf5WQQZCtfztqQe5sQ11+hUju+NJFdR0wp
I3MSf8zkCM8UJJIHqbmu9rCZNtMeVd/uMpv9VHk0RrKC70nxZSw7EkwRlaRh0Mrz7vOwvv03xcIq
FdwQU3C/13xucgP5Sgkss4Y21rC4fG9VHmqZanfwm53JZ6yR5xD+pHZIOC4PC0+mKqqyRpnowak7
hltSp65B/Vu3VC4qhXvvw49VT63Fx2D+ACoM0sJByB53LzCiPEAI3ecNmGSkbyRiwNgnVVwDMlal
J5MGfJOkbD405UGOUsm8r/KyhCV6g/SxY+5ijFhavynlfH9NBVciNqb5xXMDnSsX79oSGo4hxzu2
+tC7OsCpgGYM5IIk4aKurYEK2nZE+F/6LpF9Md1U1/9JxsIPiDaTUZg0KhRYcq1nN+JhLtSCv4Qb
gDqT55Jel1Sza8ZgEqT0rCDThTcIe1ZVf+NseW2LZUnSA0wBbq2kUCKJfTkmnLbTtf/Iap1wrmMn
EWWbNNX7aBiQgPkje+48GgyR0xGdXwSh497fyq9lJuxx9CApuR4jnGLwS1CwHNNgFRD7YdYLN/3Y
IWHrZoMptFg0/G92M3Aapvb1iR3GXIcg9PDVCUQ8VM7a0dnC1XLM8tjjKAHXxLTSnggRW0JciGBJ
uUmkiJOjUfiUW3n/G+Qeh2HyXmYbUaJ94zpC04ht5vfxM+yfoWvqz3aHBd5CD99zdOrFwoH6DLJg
v9NtwywuQFF9QbU4ztVrIS2A0nauzFdKz+VKd+ZaXkKRJ+SoaJoqNuw2RSLMRXzWS1JC9OqQMi/d
deUzAM4l2ao9O+ItmXQVv8rkcUPjzfuJN67K+g5amQtwe1ylz/6OxGDdW/4vEDnUuxnqxtEr7Cgw
0p36JRyj4vfkTAK2XXxZ4wFrXfjx1H57avlKxP2qmxiimcotfAHEZcL+M9SDvIObafxhLqPnQn6r
u3GSw1a+5/d/KSpQ9Up36pW53c/EAPjzamo9MVwSNfTdXbHlknlWpbHFOyNMSNpEcs0HElwq/ATI
1mh9x4eEX7LVvKdQLfzzCSatsTiBoO/Fj52oICKn1EXWqgGv5I1gs/J6V2k31nPLe4IdXdSBa78G
OKLs8XduQgqG83gHYJyMl6KJnktnJd6hxWMSkEpc4zhzjAZPAavlcfYDt/2vIebFGu88nZZxoqLE
KeUhVpvZcrn/lXjTkPr/ewV5E6Fsdo43UNtKG+GxRvSOgPc6YV32X8RTiqGuAUXMeW0t4/C6QZV+
CgEGbPTE1P5UuwBM+9MhkDB9H5XD4G9PZ3EdifjJ3ssUZk3Jdni2twToBFZSJR27vOixA+SfcVST
i2PKisXwA6Yl0up5IyBjnznNMG03Pf7Ay+d7scv6hh0zm+yO2kCwa9xMR43csiS6aBhBNs5EesqG
qcEyeVl1fBNxNa8JCNwuKb+WPIsPY+lo6BftidtR/HFt6NLYmxJyMh+nzHFht5IvB/3jrJzo2MZ3
gYcNR++CJaMbUO2blP9H9lT2rE3vKr8EeH2s/+qHY7aZr9Yx9xay6G/RLG1btBndrWkSQv50o2Rv
AiZkUFmopjmIpcq5dt4JvFD6WSdYjgZPzyU3YzGB6c1+WN/DbxO/isjDLwc+yHgDQLN8uWPU/mKw
jvgPMQ+mFmrb+WIkomGCK/qFe5ib1ay7WX22R64qCyyOBY8ZqiTam3K3QAJNF81aXj+t6VGqk7AB
8TJs3wtEhUyf3tai1nyoiXRqt8z7TNHkssCSMZg4yBVzJ4dFBcGsRP0XMJOBPtiNHd+OuieZvrDF
4vfYzzfo2rx0RYHh9op6p3YmFV2jEGDPkk/ScI2F3tiG9mzvlmwv12EQx0FzABgQwRYQNevmqsOQ
POL51q5vZ5TqaVwg4AcW3JlFmfOS49zHd8FQARkeBP8PcbFRvSCMUjixxptXATXaBfTfuqfIi0vM
NUbvI2XGrUq9nH+qNQh4uSG4pSyTflLxlq/UKduayBVpe+NjdJxV2jaXWXz0z0D0zTSmuhygeEam
L3XeQ1NiFs+D0NVDcj3/vMuvpopQAo9bdz8cbSPABrfOzukGVlozuLv4QaehkZuBfgTzT3ikbxXe
XrMVvJxYBdsYWoxVdZY03cmR6+HnezjzkDEheXCp9lHKpCkhcvk5wzWr+M67tX8d4w8tNiwbYB2u
K3Lb2PPPaA07d8B7FmGQaq9t1lC4PhCgsw0CO8hNLNl8TkLzmnlpHzG5Jp7LYAZhdtwe2KFaqu44
9wg56NWL1DiaQKX0UKHJj09iMrPXLxhmcdrc30q91OGxti7yVtB5Wq5chyAh+t3W1ZTOzE2gloFL
kMSgGI7qPai4fdcRoMTVDtgLC0F0vz8S55AjUqKFsGVNhfRDVl39IMbrp5IgrwD8lwbXmJ8XAm2c
e/CVnOHojLH+75MW/9q6D8l2juu0h8p8SM8+Rj5URPuhE8O3d4tVAM9NYyJokZtFAUryVvyjklqD
FJoedLSTdJUujc6WePcFlFkWKXrBqLErH4rS+KihuvShYrBSeSzzhwsC8PBavLMEq+8jAJDOMSnb
FdP+vI+AlHg9M5g7te5ESlWUMvxbIf1hbYUclSYX4F6aZh7/TQZH1ouFOygPBZnXL9bF4/1CJbUH
H6BDb8oVjQfvcHnl41bLv+24DtKI3pvCWI9thIe9H7T3SsVQP5VWxYXOCdDgCbVSSDDB0JkN40QD
vy5hNPYApgjtWd9ZAY5cw/MxTwi0d8QB2GAT8aS+sODlLdL7muh97kbVVrUgYja85g4AdFQwTB0N
Iuyikm/8/LP2koYBDMUhs3+p/9cc6Akj3rm7t/kHuAxQbpqAhm6H7ZKy746OoIeEg0gKh83D9Q38
EYCRjGoDzNYBJXblK7bAWEQC8RxbCOYQPWAGoL6NFXLe3Mghp9oRZNA09sg7SAbMy8y385u1yhEZ
54+h1+KcZ9zvIztcm/p8YuyOh9aS2noTlp7AfEp9rrdHOGnfmOAkFK1ASm9xU2rlCrFwZcN0tjHJ
svB01n+iGRMP5PlUNRmIq54IhKTDi6rHaXc/k3V4/NJ1VJwNuv4CPEhiVAnH/nf011W5djBUsY66
71hR2THbB6fN2txUejP7a5BqW7MnkeD9P7t43Vd4TKyVlQ3lbLuW01vWRaIuQn7iLXZljn0y6KOb
h2efKWKYbQ6VQFNMs7YSm44x5SwRT8XJJV0VVZ9VTt+TD8q0RYRy0+5RP/hrHQEoahKICKYeiEDV
fGLgQij/11aIbwifrrY06Dm3gFSgR7JCSh97goFS0QCKgQBZrHhlX2ee61mlm24co7J7aykyZ2Lq
C/LlsPOLiy+4M5oD4VgaGbXKAPTWnv+8lE2IHH9noslVsZ2iNEJSIuBo0sZLUqpwMTu+mmLdtkvB
RkvltelRwA1jota+yeSQ7qfjZJvPL7u/drWpIv0F7I2sw7IJjgLay20ArRSmJtHbmt9Ag2LvMC6M
q6bzCxFfpD5NmIi5H1nlbsdyDiEGHKdCv3K28mm0lqtgpN8UN+PlMoJkcH+b2hz5P1fLljq8TfC1
M+LsOIyUfaDjZGQKShd8F2S969NCwpf8B31RjUZ7CcPZN50Qbf/Rs2qrjYMSJsAAZCeatrntrUnY
7T/H6VPXf4ecor75/TKejn09vMCJv5oHvUfKL/XDDbmlaUUOATnQVhVJ17IS9BADm0fFQDbHz8Za
OgGd+S+SVQmNtZAB+yH429jbfF0XbJVAlBQ7QKuIpUf6YKx6g+dHXCBrvQEm2RFV7qkuwZS1VkRH
hOPPY7UNeKhUJDxW8Tf8vr+0Xc48TOJ4JDE4DKKxuX95uHHXcWnydNDk8K8zqLpUX9UJKY0wB1W8
EOSL7tGyvwbqMjRQ6wCaJCDJ74pI59wOvwOB+QVWDwzQ9Wzj58gK82ErrPRgal9G2UYl1AQhRkcq
mHJfi5WlFTNlgjav3eJbpUq+IGOKqfWIRZGU17mBfFHOwHWFPWpLCW2h2Rko4BOIdnzgDo4krfoV
dDfOaMxZSWRUn4Mx48jRZvy0DFMTYM3CwRAnq4YT0twfM1/14Lo6B6kP3Qa299SGUbEix9N97KdQ
YGbYsu+M1yrLVzRbQRMA/hco8Fi1nHOTW6tJIS1mjnbWCp5HyBQFTyODBiQJ2pvtb/e7aRPruzRk
hGhsj/kKAI1XbAKPlVzKbArzyT1t8QTn02lwV4MLdKptEbqbE6DD9o9vNHEr1DfTZaZWMNUaSq4G
BJ5rwEWXJTwnxjbX8MOX6ZZIZkkXZPSe6wzbH2IwwtV7aJbnO/Np3FHJ11TyYNbb+ErbO8QHBbuQ
zDEHrV3LNSYowLYXScpSrK7JzCpr8vydr4vJYsatHs27k71kgaYON8PfjpN5osXHXYzKONJTlXuz
kWU1fq341i4xu4RvvQzT34gRCldAtV4Cg8FsQy/p9yQBpwfDmuxXhFZ/ECWbnzD63MhgdMOfuelw
7DQho4J2zT6bXM00TkrsBStOxDcIsNB69xDD7010YTQMMSMpVfost44U6sFxOEoGI/r3Cf9Hgpnv
8liDE2R38BPzGLrh4ecjij4wyaSCsqBR3nwhyC0Nm5GZOJMKjO8eBOrvD5GJanLjX35qqnhZGCs+
zuTiL5vBWPezr5xBG8veTWp5YQ6Z2glCKR9Zx0iDTFG7l3/hGPMJpAfpCF1h7AhrwMjl4ORMJ2/p
BZBxZQdIf8846n4Oh+C7TUNZUf3MO4cwJk+nr5gMZ+oJ4cDgKktOJVQ3cPt/ydiq2IdSlaQKSee1
xYULEAqf4FhjNlFGCQGkVoRQ9iVd4cug6oLka8NKeJr2IX01EgKSVg0e4vlXHhze9oB8+3B43Xrc
Jp8U/+whq+1FgaPATrIciNAb+qXgrdQcijTu6CkZQgATEdA2A72WpHv/WWTt7J1vZ+3Fm/sd+8IG
vvb16VPcfnImWVSSqKXtcTzu32JUCXnBEpEz3eA4p+WY/z8w+VXBj61vleVUjng4DjorhDZlFKsk
MRh/KWxq+RspTjj2F3717eKvv8CCIwHTbMc1HBs48zZhAS0L1T2gKYRl95wurAOalIVa/4V04vwk
7qPwe3EUj9m+EON47tc2ykipx9z3NkmArhXnHtglhpfo2Wt2+57GC7fqBmKekIU5iHhLZW1EGjY2
R5ULlBB9z0g2wf3OXiAj4oTlrVgCG0RzaUE9OwDMT0cjr1vafbTTfsziVXoAvjLm/6pBsJnotCNm
tVGPRBjzjL7uCmKp8kqBapuOGNeXiEC5gmhhWuFEzOVGLSQAihYlIvsbKrIiSKkHb8facfFH4yIE
JCkEJU4Ql9JhTOi0GSEZPUY+smvtq2kGfnWUIorb+WBdI6LEvbxeeaK1CcMWyUv26qDt4QSu41Dz
mEbNYUjcse33P7U2kuBtnhOeA/+nQUi01Y8CL7ADw0h8EQ4Gr6XYbrtFeSyPYIVqDVfyQ/JjFGqh
/NL1x9lk6Wdf2YB0vFsOkdYiLy4JcGjMJkgPesQrGdC57FeVT/yecXxH8JecHBLcT/QMIA5Vqjki
mhFo93ZgDtHprGJCv6njz0BW0YjTPkqhig5g6cPIxWuwP2eoDQ0171SwRlASasCIgFlsnuo0/M4n
136FHziSwfezaz4cyZoSbBfSMQEN8upqRRwJaWLmEZxyfcJ6UtTWPkJLyykYt8iLv2hJa3Updin7
2ITK+9sZL0i76NVdNGIZiN6vJL4OwvG+JE9wifpq+Hkl28DZAu4JPDPuF9nhIApddjLv1e7+LG7x
y3qCr+wk8WE93L12+F52NkWc5lntDiyGAy6wYthN7JFBaBqurqhkKkGyT4Qu96aUeAsUTvIlC4+P
nz896BkHxRcQKC9wBPat7JZh+/FGNzvHtot1tPSg5C9zYhFJGlAYR6dQxtyZQHlOg7gDNx2ttgDd
4wVhFRh68taA7AXLDgtbGmwagzHCzDG+veXiahwxBIRlAHM1fWEnsYhacMUjsvGcnEXHVx2w090H
B3bgs5oPi3CDW45HMK1coxd/iDGw/UcP/wjVKmgZ3bhtfUigLNB2AKVac3YCrQsFfzCpySavVbPN
GQtylw6qbFM1NnhsIpu5oXlo+0AW8waq7b8dAZ1bsVCTiyZqXYEUsVn3TpFRzYhP7nMRkdDkApPo
YFzXGJft44gCKNtGexqwFCysGZuZ+iULfDvNThH6ne2Qn48klY8Qn9nxNulClT91kdjdgfHrlyJv
cA7G8WEid6KSURQIsxCTjRqMXmXJX0rNROZ3IrNqReCznRSKVFbJKoUTNnYyYmKwgUOmsSai7nsw
Q/LZHTGz0SVhacBCdRJ1+6YwhEyggCImEGEQu5msNgsnLwH8rfOvhEK3NgZCmUDM1NDRSSXYWM+s
j3VyajwnitcxouURlRDqegDeSNswQvU6xNJzcuHARz664u2ZF5/O5V+ih9G6f0M4WgriMxmWm6Ny
Dlt+rO8NwPN1TJs3rxxPrnUlmtRYdyNFM4d0gXydAdTyN1CRo9SNTm59t4x9v4fXWMknYP+49ljQ
Zt6ku1phjxA9X42k1z6Qi7Yze7YHowxTs/WtoSzAkY0sP68O8d54fgKHjKv0NOKPVOYVutg3He1x
7ZiTzu1+cx2jLGkrPIfJ8m/t6ZkyzA8BA0fm0248m0XwZba8eDYG1mxHorYj8Dv18u6Zku5r06lZ
L6DL+iJ+PKM0w3pZjUdwH4uL+JjMKkM+12N4ux0e4JzuKAxdZW3QAtg4TuaCCkSr0qu4J3d6K1Bt
7l8OL0pXz1B/AcNWxlvFu7oAYscc8Aq0uBtu468RBmszG3e2YTXR4rZyMwXw2WGBLVWq2roqENEC
hga3eHOhG3OCW+7jYYYjNfrDvkbenGzZPMCsjSJ/JfVpsgxOPzTl/dfsDuCsrTeB9a1owGJ/S9Zc
iY69B8CSUSTDXYMJgmdLDsuQdKTnYd5z0VtcX7di4znljQ0+WZ91puX1CCD54Z+ccI/qkx+3ZB10
Bbp42HbHMCUR31qDKvAlYAPc9FkmtpuiVMcqXP2espJlUvdET5rBqkEZXK3TThcCMOthTQ59DPhD
LiitlbeA5Q2EJb0XOewv1npwgOCRAQGX8IwiF5Hs6oT0LvXD8gpGvSoMDnujEzPjBgBahROelODz
PQB/uV1sI17aHX1FPp++Phn7y5PvdOU92OL7eh7beOUi7AuQ446HEj6mvJGSdpJIKJHbymkL9NZJ
htK5FSNrVmQtorIeJ3ouAculZdS5bdfoQ+AQ58Hn3ZPxz+ldxPj2nxTBuoIDbXT8TzRFoofTDNGW
HcL+6zVlwKzBKkMykYRmcUgGET4SZVuqNxZ3Ml/Kg7RLXJtmUJYiRVvXIcWQt28ae6hL+i3KaNQY
BvrmK7pWMJVame8S35UADlD8ixnctdpsxOqQ9TpbSlxLZOeWK+Veoh1awlxsJTYhDlaO8c27sevW
B/6bpsnqwSjrfk5Qd4ydUGEMROPSupNfwmT0VP0ArC4F99KgxaGEscZiPVfaid/bLx5s0nM4KBIv
VRwqy/y+ac0V3r32DW1WjEjklkDGLXOCiMeWx6D9sFd/3wXX0zfC3789oq8o7kLN63KA7cCYZmTS
aAjhsD8aL/Rpy7QwElwKFWAdkDMVHcrgi/cW0sfYuObTrwo3s6m5hCKAzNDK8MBtrBEKfv6VLJIj
5hdlIOsNmhri3s/ibZOk0pqG7XQOupxctuMIQbGmVQhdppK+oXZaPZLjT5Ivl+Is8RinFJ59UXzC
rNGQHjPfClV5d4ZVgd8NTSB0yxWBtJIH1xJzCOKi2SWuOT4eAzlSVKeTdhwXEnhRnZA/xjZDcz7j
PvD8vFwr9P4Oh6gcfd7JdteBms1mL+wL2SaYzsDFhcUMXc6PcXlYLMtjwdZzPcqmIff3WJujAcBo
zSIZ+bkx41kDWhPrRr9cu0RoJ+s/3Xsyoe63HCl8YhC8YlgFdaNaOw+rTRujQLGGNkzmgfEtgjeM
Grgj/bAo2WgbnSB/O7+m/DWeXgr+SPHRQqfH0H/heHMqOodDm6d4VmsPuDeCCkILhMaJ7pYJ7wqK
FehDG/XbjLtGdQPGdR8eitNRHN8EdCma7khMDsdZ8zHFC1qX347wruixDn7fo+rqskoC8cIgbc2p
B6ueu/B3a1LN9FaxbyULUDyLQxr+p0JwrhjqalUSlwDpn6k2wmGO+XoxKw8qqxwNFEeAJaMQFQ9g
D7dQbxoUKOwK1xuv6+ItkvFtzwPKgrL0DWsQAyR//qPFzp8cCQZlc2jupQ/UmP2ST3+KlR0/iMtE
CfrcMfDHp7xAfUg671gCc89TbDj9KRc/VWxid4SOtlg+REVFe8BFBgVyGsGr3FI6DJwXQNi2fqlU
o9A2yho8UOHrf15q+o8l5TaXNwbi5zChHJ1a6Iw1fasm9ILLTZAKY9ozUN6MSd6Ld7bxSdb+XjK9
qvQ6AMXUKuAUvOCkv9n5MRC6qHLm+HY6cWX3dXUdol05CtEDo6lSO33YaZ/6BScwDPmD0wEZ1fIV
h6YeQuoHbnL9Szhp0uXiDRN3HgSrWcu4FixBRQagdXwUZ5wOIfv5cFYpY6PWRxMvaoh8f0P5toaX
KgBKJYDu075UqLj3GHe05RoJak4uG8y4IZSNeoUPdeg/bDVassMrjhkwCe6io+Us+XZUYuEvIAnD
incbjc1mP4WuhUVouGuPYykTvOu8YSUVRRRGSRBeqeAYeFQ5NUcM5sm/wt+GDmyBvjf/mYOPtdg+
kNRq8Cz00QCWJle2R3bLitustOR1KP/qsS2OPQ63BJqSs3FuVdp46YGVy/GJR7eebu9DAbSzrBk+
RPv/F9lFWcC4jpy+9QGw0fNsq4VkVp9svRxb+lapUY39yrIrz68ibgMNA3JWyEtMjGymDyEzVzEd
PrSMANAtwfYuHiXyx3zh6NcMlGX+zH50QGiCD+LbcHc5IfCDut1BwODj5xJwX3qdaqfRUfbtEUTP
eXJsyTSPYKkrQ7tOvfXXC+Op4X0w/CfA6Zjm15678MrY+jxBSzVXWDIsL9+Q3cm9o3ziq0oVvDjW
7IMjlpDpefAWQT1y0lmISda1g2QabT7TlIxRHzEFIeqfgjBcLBhVmhXh4sGeVr/sqq2JP5K0oaoR
r8BWs9S8aSZBRJXFYrCQCJqsz1zZQV/ysvlpSClxGCXB1NXh4z6zVanS76ipA116KOpTIjRKHSTE
47uwkqayjKhhYZ5y8TokN8eoI6F5DGuBf8TQYLmJfyeLQOS8zKPtbEEekTwzB47/yRcohuTe14wU
u5qKRr8RTkhS3M0oObWu9rWvpJr0YG6PlDOUxtxzrw0AOMlFcyaTkgSReQ/oqqD9R1inR0fe/k6k
qUhCa/MU4sfpuBxQJ2iSCNxRKMcu3Gwgt7tFvLcA3dUsu+4Cgs/LXVOQHRCLE7ddoJud6MBYcgPY
HcX5W4eFnq9y5fiX6JbjQrA8UAYrEhxvvz3Q74kpcmGyZvxs7HADI29+vP4oKojnADdqRgmSaip5
aMyKJEUvu9xObiG/Iyp/hO3thiMEGgL5ZZ7WjqfBGbQDYC8beySKs3irIaipsOB6vuaZUBi60GJ1
Lll6kSnL7tc215txCABQpqnvXmHfwQLO1TXa3j1LZCd1jIWXmSrTB64dcENL/V3esJzC1wBLwHjp
lrmSvLycanR4wjBm3zSVBxvS6WMXlaPsS3lE6NbsIEjYcxag8pPTJQdw2z7j+uenHYpK7U8ZJKCD
iHS3ceYuZIf3aXZF61GnBW5i2lo5d/EHCQRugzYETKCYnr7wD7XYi/MK8/ZHKi0HQNfxbPKjkTGs
wJWWO8yrPfNWwD7dxRmaoBSw7OYn4jjpKh8/1h/QDpXNB8wFemga0rzDaImnnYKKKemyFK0evYRz
kATVd2mMm0+bLAoEvkxJrJLxY8afO53nVjVAMdwNRaxjAf/6DGfDIVyhVCEQkUgwH7aq2iNj1eLR
dLASZH9nR+3IL36TNUd48wVlb0gOC7OPEFIgKmSrgGTQ/834DitobPMga2XW0ev0S2SG6jIhJbDZ
lUbSttUeujdtw8wvBDrqp+vd+ybEBUILo517RWTqZkTVRH+9i+FWTwPVg6FPgO/sFFGNEJ7WTEFq
URjSuph51JjFbjjufF9euSliHr9dZKyGGH/viFR5qxmtLC2FNiS1OLJj4ebDKbObyU8011b3TNdC
JetHxT7SPXN56UR5cCpIs/DiLDcjBg48M37VoFaQW9Yzws5DJjtyymSk4wL8ie7ny30l0G4WaLA4
1qtcvQd/v9Sof+ojskekJGkoUEINHOigLGIMk/Z7yTUe8+9AwsF7LdY+QSL4dTQHWI0L9zfadJde
M6hY+ZEyhkSoKB6/lc8wr9IKgzy2RJgSv7izWnQjpypg22bwg8Ep/ajPMEuqU6qxNnT5ejywk1WD
9EPW12RiqdNhM1I/adDj8FZBS5JzcVQhC/tSGP8U6OKMO+OYucdg13DAKYArG7bRmIRxMUqutTsq
YTnl9NjZPMtid11v72QzpDbdQ+FcevlhC2gkMDe4+d5G6E4oDZO4GLYTlt9r0vW/Q9BNNREX2Uqf
E08ji4DwfVi0rC0ZcUZN8w1726dQSR1YLoYfmSTXTIUPINHbAHQfupFvX72+2LXkOOUIWXx50i8E
6YqkhDVsiGbty/gcXj0mk+spdw2a+tFXH33Qpe66rg+UE0IkoHdXaFxtT9MtIuQgo/wUoC7SPmwq
fScx5v+AthajfYIeHviYy2m5sYuk9KaCdDxWckMagi+p+zwe931Gu9th7lirAkBY8xdQN6uzu9Iy
XlA1osKejkya2PaHcaDeVx2x7cyFQ0S+VlbrN4Gu7ectJknjfFyEmxzF5eF5fkWS8Yuh/IbhAQTJ
Kh2CPOcZFXHwl13vLTD6iDINCcQjMFjKgVpYeWRbCIMDw6wN5XZZFgMmCK4HXls3rAMs2G+O60DC
lw03nkUqOeHKBmfp61x535cjSO89E/qPLW3FlALhSDKgNeaXIKXBxCZuY7DmqbH159ppPMFPV5RD
XGyR8VrEhGKfhuaqnZR5T2cBQmHYyugqv3I/tFoQ5J7ID/E7pKHsjAUY9UbxrIgJA1I+RVW6VYQn
cl95u042e6kbr9fpcrVjhUYaPv36+MEmjtPiPsO5r+FLTskQOYlmIiOyR/Mf19+u/EZ80FY7qLJD
eKvezsY30GHny/GCWMzj7Fn5ajvHg8LcwhBIjEdVbcl87Tgetn+DU8UnwtC7/PRgjCo8DWdkDgLO
iJT3PayJ9nuhPo8OE9hv5Fu+aFyPlRfTXK2ZGoNy+UkRTUrq9oCkeN6PSU+jY4wEM30MgxWKRfk2
yyae6FoXS4wX3kZhvXHDcRQcOFZzQVQABiSULVDbhwrpZpjecCURZG1emiJrIzxKp2yPDE43YKYN
TfQlgzWZVrcw3z7jDccc86oWZ3Kb8feaGVn69dPMhUTjdigzBSKz3Eg2fqeXo1u9u9BnzxjjPrIh
0lSTjeAcgKsT5DRhyVw4YDo7qwtxQa6653rJBSDNwZF7B5h+TdYbEJxssg1hVekRL2kvv5Gx9Bsw
K1CDkRje+ehTAy0eJbZVfioyzctxw2km9bcwwzPUTnydTRQ+eP9Z8J6WVs4mn993lk3ExRBb8GvC
1oW+a2ghpEnTegQyoNcuNbGQ4uYNOdfUAr7BiL7uQnO0Y7LvUHaZmtv1P0IUy0l8DZ06vWh04IDb
fDw3HdsMwbUtiypasuZFD74Kcp7qybI4XHAZsHu8/AvkJyukRjEAzfMRwiv7A+Bzp6CKMvJh/P2e
iVAt8b8cNd6JfB94NwegTuOKg08mxb/dVRohqQahHgiZRe+WIcgkWCdyFc+059hodlNVAEBHcsK+
XspyfoSzqRrXCfrXLCvHQoY3hqC2yQNY7yR45RZ49ddr+tGYNdmQWdcqCGVSTmiXYeNZusoTwGUU
6PS4Em6miHnj6uxVa3ncP/1tiFMyY9Ybp1EbX8LrxQ1+rG5jg7UI0l3Ug/n5VbnIxmXwX2BQRmHz
O/aMfmhpDTl3ckqRgNASmmm9etZfQeQ29JlAkcJ9lprd5GtM+il9nHOSvnDyYnNJ+uAXW4Kp3H7b
6PLXX7WDGpsBXAlCaCb85jB+NzJU4LBskWQkWUzNgh733BMcv2RKrYwVydc0y/XuFoEwX6rGlO21
J6xexD4kqhH+0VWuyRpeIhogmqYD78eC8CgZXWca71wq5aY8cEAhYjhnvVJS5fmVxEDHKdwuTtk9
VIgwKpkAEmJFjD2MjPP3Gl737HFC+gYDfjq86xPJbgG4NLsgkRJi89ykR71ZaYB6/Zs6DhcwRQyk
n5806RxBuofwnyMakaxGkBuZy56IwlTPkhUgqXHZAJiLVbNt2FKFRy0LtdmGgyi4QriG6mFZpnK3
IhTXrt3cnU/06xHLvvztFp2LG4OMO+OWPvAhNX6HDJTESRP/z6xRfAXjXMb6ysEFIKO3joIGi+ak
Ack169uOeNYIqeO9KZX7Nb8fStnStyYIcrnZCYoigLLVtc/MjiFrrfzil8khIqb9jB5YIaWS1srB
p+G1jZaNv22jYpPA70Q/gd1DpM9wS16+9FUZS9M/Bi4iTdy+sv1gh16/+KsmFtputjc3CMAAUGOD
4/Zx3yjQkKu+V4Ys8GA24vvMSctebbE3SYLEkyTNspKCxILyijR3QMMB4Ozclrt7niOKVQ8KddaD
3wllIZ/YydAjc4UKoNQmCtK9IZPaFMVG3j71ELj1ho9pogI3Mfyud7CbgXOfz5CELta6R8H4zIeb
LSl/Hzt/i2mA+CKp5ZH2Qrgm2UBqV1StU+zSK/PrYQ0HtrJwjbD4ZRI952FuVD9JboXVWzdIS4PB
FTmfE5lZo1+1h1YWDPtoaRLYkW4/T7iEwqSS8i2ClDXkI1mTPvsnSIVBJVxmonsTK1j9B5ZOorlz
c/WoK7scdBYFuTn6Fq65YNiEdYg+VsYbp/Gk66orcMqtum5+OH8PmMWEqbSzH72XbxNG86baQItC
vHM9kIQPO9T4S9xTrubz9BjbyiA3HkKyick/UKOJL3iTxlmIyrNux7Abs+OImAa6IkkJubtu+SnB
uaYJ9OIDlejgbAlH0Nvc4w9P2aGrDezDMKvxWgExmR77dFvSvIzWmUPJD8xxyD9iVMfz84iEG4fq
CFfOkY5TF9Q1Mnvug3sh8JfS2fQvEP6UGCEcOqeQoUJa/f03y2jRQIPxZ0ucHMNL62YwPKxMjTii
1MDsyftK6uwWxZ9SlKF77PiuZUsSf2s1WaKXy5An75EiRg4s/LvVaL7e6qugXMND6aTNSVBg4ZVh
6nJMJR7sfgYSZYzj/6t2GQIpw+d1OTUQry9ImhS2jLZXloNzBj/8uLnZIB4BR5k9oO2bg6LHpHcl
wbtR/Qkgnomb+YCOAaqEbByjOcicEk5NYzlZMow5tvSl+MsPqa3nMS1Cnxs6szElB7CRBibRhJ4i
XV7BwsevB0uMCGlnI5uJbkRgUo+Uz2h3Q2r2FDHoDopmzQNORMynHmY6D3R6+B13BbssY7NeMDnn
tSQ1wD3qlp5JLjWw3ZgIXTrhpg/D81ah5M166hBXTlOPiv8zWG3B5MGCYNl9eBdOD4118H92Lmio
mbKQArP39daqg+mzPxr5GPEhO3MScUN1+UVHKp7qouFq2G6Gf3eX6OqCceOuwpdy4/VrM9b3l7iC
yRf+MvU334KujFHQHb9H8yt1mVSjtZhehtrEJ+j3JWDOzTB1u77GCzJbq4iLrxKzWiExs0blsniL
bzRG2b/PncLqFK5qfuN77W5jU8hX8wt8gWAGVUBlKNrMS7WTeMEopIKeZYm9mSMFLBYuKGDyZ9oE
kN4vlaVu5mb6aDFacBtHd3Z21hiP1ELeabnUjokx8D/qwY3hB1wRgVBlPXivnvaKl7RqjpkKpH98
6zPcnithKvcN3FDIPHJ8T8K+ssTVqwhRLCOKKjIGlM4JqonWyIp/HSyg3Cclq7Hvwnx1YFP+KylY
gXhL9tbeesdnBNwPkZrybK1bMws41DOeYhxgqT7BUrn9vABeOYLwFUUV153e02ZHnZzxScDrt/xJ
E2p/eFt4ZCV2DyyjggnRGCzxC3cmGXTZY4cPUi5IFcDGBbBkC8o6hkj7wXE5o2VjKXf87kEzuhRR
zwzmYsQpv2RTXA6CMr4zJrdkzNt+EDbr9c44iANexA37X0BmjYB26kaYp30GNfxB23cpQheNbssM
Uz7pyxzuK0RqvwLaWT59xmst2WqYVyPfP2PkYMOoraCIO3C32btNegxzkv0mMCGWFVdDX4ry6qWh
+CYq+YCSYWgB4ggSWgFeBryQzMeY0ne2719/XUaPXrhkc7NqFvPNJy5B5YY4ScXq0cNFi4R1YI4g
E0MjjVmHH3O4DZAmyewXuv/mgev3/kmKCv4oHEmAGlIJzpOzZOtBmTYba1eT+oXW50BpjIg/c5qY
6T13HbuFnxQl37jWkCpq7drOnsnA7STv4pcG+7w3x1+lDoBzitvx53A/zTNnV2wgbaF+hLOZ4RUO
vOu7qSGYLv5KFnCJ3vtCwbXVzitjtqh/qbAVyLFnPB3qavoc+Be+GnCaTjnqQ+R+rEUrDJev/VWi
VBdF6PXdHkk/bQFhVZvvbW5qt+CWOVloz0XtCWt7yPFhAusUnusZ58pBSZ8B9Rw5/VBdtC90a15H
hLh4LVTVMNVk3wJG0BYUFr1vj28iu6hRp53J0ZbfrlAaUePD0VPEKxhS4K6ljKNBMgjHei8EtXq1
SaEEKGHsroIuF3f8ycLmaLEiHpumjWdB6hyu5GBhp7IW/doUfmELXPrn2fQEW21is+qGy54AeQqF
moIN6K6K+uLfklawxZ0dR4gbJ0jHtMLWL0SdM4ScikU8/rjUGiXyXbMKl9tUKJ5aIZpyDecrVRRW
JYQCQKQb9d4uKCt6q8GMnFF1RpIyIrloAoiy+7Zl2cW0Ln9ujBYUKa0XG9fbPCqpqvLdZAXY7dv6
KFWxupyvyS6Ao/EhQ/oBFOrsK+TTsYiEgbML6mzvJa5/hwox+I50TtiA5wIJ/QPrU5nSkj42l6/8
DmZ7hbI8PcTLrdynZuU5wXO4SfnFcBwxcm6btO8adOmBZcdDaEH12D27Rfk0IiegLNCkSxpd28eL
546iClkDfGclWyCM6cG2gzF0m61S3ofsbrkVqGM12GtFg6BlylObu+Hut8nKGxGQwdE7qkVz6xHE
3dpgHWiG7zAgShlRN0t8BZz9EsLIFlKbIONxOtZBD0NiahMASZD/DQSX7czlvinMORsvHaJNCWBF
3zw95GT59qftC6ctBEaTn7hjSlfyUWtS/YTgrJKlW/vRhtFhC8c/YeJJSLBHUvQNL2HmtfIztxhs
EpqN/No3B0TXoHu/4Ps3cMBhRZyHjqDb/cDbIrD+oFHnAtOTne1ruX/BELayB8YV1UierbIqiPG5
AxpHb5WMUfQPO/6TwOk+axh5tbHTaP9dwztHZuPg9/uqohqt3M+5reJ93ErKUND9Wddb+vyILsEd
2xyRwSBRgWd2izESvaUtiPE9Do3wrALqaXJXXXNd+nuXIl/urKzfhy2Y3kfwm8xVWtfngIUFAf1N
KSWV+LHqTGDR/+Rq8vt7J7h+0plponkc68Z8vebJOltrqWJ/d1iUj4gt2CwtEyq5OkrSeE+FC47X
1IIeuwiv7pEclnbybnU+7mPhEz0Egm/AbmzPebghNrBG7F9sS+NmerdLLLbIWXeOM+fuyJlFGkPV
YLV3lcVd3ubHnw7Px8Uh8qZxIrbpeE462Tgq5pdqva6AI8/pDiXgAyW+9tf83tsdkWP0MJQQ16fA
FTaKV5fD4tXMeK9nlE1yAEwpJgtToy2CmU9PCSfq7c4pKzbozFnYQ9Smf0tlsnbs9lVrU78N8yTi
zbyOUTRrZXsm9revF9zhReqjaEUENttXqmVNaKJeNUphCUNmWRkYM2YjgIUKIaMnFlpjXD9ZqsAn
NxMARMiBiVlnoaUlbhRw3NmdDluEswHjEGzmTuZ3O1xYGTZNPHXe3wF3krcCy/u4g/NvDzB8Xc75
IcHehOlffnnVkfUQ6KkLNHaznjFw+HkSxFsop7alFQiTgLuPeWe5DWqnDdTM7ANgmVswXP2MpjKD
9oAqRd5YI9LPydQ15nQ5RfU5BNF3oUjeTOXTMeATGQoQXxBF+E8aFI+erovpA4LxWH0/6ISm7fih
Qo+FCAzCfjhtEt/kLnof/0i8V3UzKoOborajxmB/u1Z1gL09lm56EFjiKpMSuCobE7v/r/IbJ7PT
UW/IXqX3v2kjnL2HPMZSLksnqzFho23agRHK8YmHbOi9o8xjXakc7sZMDIXwXuAvOfpK6XomR+1f
AhvwmP3KRjTwrOMCMhre3xQ7YLByw14cpKFSSSGfPRcsAxTkjfxhadyfYgamnGCTuQJCiCQrxEXA
7RVsulVDuAOXtKG3eExRu3690FGZCV1TSLHhHEmHXH8rQBP2gDk1SYwaESEsyhBnHml75BLCrCfH
Tz5cDepImYebP1Ub31B+K6dh278DensN7FVftZJhnbx0aqTP2bLTQzkxfWKxoIONrKns4oLeNcEB
U3Lar+E0frEhYpinklHVd5PmH0tkh0TDCPeYAJGNomqqYo3JicRvcWLDKYK4CucrIYpNuoRa8DAl
XKdNfIWlKiil0EAgwclnIuiog3/hfZRWEKpkjYnxc0Q2cPXGI16HgdCbM0ZgOnmmA36zR53Fo7Rj
JC9HgRQWP8jxADnloyIF7GhCuMREixBA76zFzQ7eBhDkvmWMYSHNm2O9YvjQWd8W1dWqyIo+rcA6
dROaE800w8XHWWhHoRAl5Ax50Jcd3gDwhCinrP+3OOEPEh70vUxE38tWYTUceTk6gEr8A2WqQy2f
a6fa5+qSmWKciasd0u5mu9bzJI49vqlWcHGatrDq9tfNtMrebZOw/sN/wMKmN9s1K2zrlUu2GTn0
DCj1WZiAC4N85YyVWoHRPLUCRfxTEV45UiYyot200MBHBuJUsYyBh2d05P0b54xgsknceydFFBbg
QKiMQzsYrz7gtdmIAgfEiWoRzy1io2HPdnPffCHqRmkgxAaS3TMIrmUsXX+bRwXjjr22RKS0/rwS
tIYVLYde4xrtdld9y5sEGs54i/nWamaYUXME7s4T1JBk/BqA78eDBkvDDo2Mh3HumYyIO7XAKv5g
MjMJd5GmhxHOBe45BjDRT9oXukcLD24lcQeBlAZNv1OMTxwjoacfDD+IKqJ/w+qd/uvk+wyFDDN4
/ifXoDJcd81i3bmVlRXl43Y6Tc594QBnNg/4P9GPlPFJB/AtEN95XMYIgA6B43e1MfqV5PA4BHzF
KERP/vrnyoKK9Wgu9qup2BxRwpevxMCwGkPwRKL2Y/tL25LMktJGKQ1ryEYi5hvWRIJAefzjFtsx
uhp9iXPhCNXpXsaveV4/YTVrdUZQFVP20MDLDbRYSi8UwqlnwwG+KwxOPirqNQLhLC5RDaNpEg8n
JUb7R5OE6/dBCpSpvZ6S+ZLklJFxfUDC8NAqrZ1j1+g5DnsXmyMchwipq2F1bZpg/M4fx2XAvWnZ
gT/yfg+ix4VsVImy8u0T8Mdka/qiVewufK9J43g8KwNejpIxqo8r8obGH1TqF6IxTOaTZ0dShhHk
zvAlWitoxAVzmaiXBRHMKF07Fyib97hZMyWTSF2BDmlmp8VYw9UafxM7Fdmi+H0uH4l3z9C07vXX
nSQItajuhT7jgvqZavvWM5i25OsSMtn0ckS7G/gQe8tsfyzI51TxQxzvjvmNLSnvNLw8vviOfjgx
SVSJ5TpxJgIFldvBd9mM8blPr5ZvB3K9mHkec8pCqBxqTIexhfH+y1/4/MOOshTSPZLIh+Ekn6nE
rR5uanBor5IWSH9TF93F/xpcznc8wJZc/PnPiLQpYYXNIiODYPhjJTmsW29zMgMsrNibul4QCFOe
RogwTKXWx2vpLVnHerxP7+PHU2abv3dy1LzN5afrjg3MFpaxbSMekeWQUFx73buBXGBn4apOvj5R
EwCU6+eYOTQ+wSoRPmuHTjEuIkVFdTACVrbpEXQoEQsLd9SC6S44T7w9bAuOg/K73g8HRYCXJHpD
jkOoiZbQmL+x1/fYRynKhfmSni+RebQk6OqMVVqtNOjjWuVBos+9TnTca/tj8GmdRSO7v9I9Sel/
LNRQRgtMcI7e+J29Iwe/VXWe0lV4YSD2G+CYaoEU7HDZ8xQ3MiSBTOpCz0GTXy3xmwBnAzBYQZAi
ZSm7gUXWfK1Cn/3X7CHdUU0x9eBYBKqjtxYq31UcVHnl3VPFrAAk4GPyP4YYE/MJwYHZ6RgzBnhp
VLJ5VcnbOFWXsE3kLB3UejQ8zCDW11X8fhzTluBYOAI3Xi+kPI4dqu4FT7DLUanPXKJHkUfv522l
5TzlKU01PTZpcX8s7c5mG6Nme/+NX02loGkexa8UImUNMWjDzG5hhtWXmc2uDASM8BaF+VR3dB4r
i2Qesu1VE4OJ5O3cCYdPZI69x4FUd12NuVWtc3GEyqeo0aaPKOTR+2v/JVA2qnE2vFKODWDQDf2k
Lq9j4bQU1k6tveeS2fmDPmNCzge5EiOD006hH8aGo5PPEDYLbieHYst71NaAYVcWERS7d6bpHGSY
04rMlc8cFMwRjbpey6IZGPCAQxHxiDnlfJp6Nn6IxwRejNAqXq/8XshUR3E+TCd8N0wqxkWG+euy
c+SqPT5Pe2PaQdKa5w80ItgZZ5nmK2GRDGSAtrVygJL9g4uHVW3W9F1TO5e5oDuX2xh1bqD/Xo7c
JY/yugqZQW73egHQZZdByhyO6p/F2xalh5U7vlOnVn2xgvrl2ea2J67YsJT1+VLsxCHhloRteljS
HiglkjUXIRf2zt968CpWjPRJ2d7QDoKRxtk2Td4ytTt/Uhr0hW28qZlD0JkuNeAbQ77EVYLr3glR
vxItVOAfCVmfi6c2JWxTpo+B7piJ4bb7xrId7UlwhH0SRIPRNiFfdtkrkS2VM+JROsCsCU8eQ5Jz
IHhXoD0CZxNwAyt5AGjTLF4RgQxZbL7Ht80e1O4nNk63erVHJtcbQZkTiCPrg5WBph/q3ogNMSyk
7vK3BsPntmG549odTZPrzaSgmrLM6zNuZOQibXA3VZJmKj86PyHaUShwVysAmFnT9R5HZ6IjH6Bu
7WRvtX/BKneVE8ZJLUfyzTALJhtGeR3xtZKS5kkbHDGizB+6erK9+7uUOkX/h7hmG+iXuvjbhGc4
YWnxC9UaxkFgypUVKerC/asPB0GIFKKB4a7eQD0+52oBe9qpMWwReUUyyTtJrefDtLTF3y2LWShg
YpsIpJ4LcRhO4lbbLfRwJnQLjQM3z3GtCPrMxwaKKubFtfy253FHAkwWsf+1aJKyUgBTI/O7ZXOq
O8LUBNOmEWkEmVM/kJGImm5ELK8yQSiHAigo51uXXW7Vrd0jroWvl+erj+j52RUjuATeqANHMzaN
/xYz4ZzidsKsWuNUa7G9VWy6LDmGw3MJ+kEEZ0q2QVvkWm8GLM8xZxrlwGyyKgnaJp4vBa8yyuqU
OD/y9bTzQtD54qKdIvgzuEvVCTT2KF9KR9vpX4dxkdA5uGFLb+ETOnZ0wYpN1l6bT4cJea2kagDD
QdPbJgG0JIyEx+ynrAN6UUtzR2KxHm5nB2KJVHY3lWnwCRK9wMcC17xTAk43sLdZ0cTgpMHJEPbu
7OB+Kfg3wl0WlzMaQBwQkxs0/f/mkB0sDvRMJf0j3hI5U8GMaQgwg+io1VzDm5Qcdha4tz8hWaTX
ZaQNfOMRx7ImVhGGwy5ohx76Qxtyj1kb5O+AfNA22UVkSiImI/cT3w79KG3Ba3xNbGJBeaA96Q6R
wFiDGxaOe7Im02UsG1VD1xcP8+vcXnIBPSZa6GCRIs6tsrajYw3jcR3wBWOoXO8ukpCFiY1TGt3C
HMKgGdr8KrGBKBRF5UnNZHKJzJePfGqo6QIoEK5+ZyH0j3LzwC1Taaf5CDCO/xAsjLdyAsteHRGc
RcujlxBzA04WE4ZkYapVTcPVQ5vt8ce/QevQBJx6U5t4kNDJV6IQTahA2hsw4sJ/REhDOd2a0fxm
EOcFhi/4+aTZ6HdNDaoo/GAblP3MEmzkDltCV+HGc2LekhPKoa3aHSMU/l6+lAJORNAi9wRIm129
DQGKTwPYCjyl0h2z584CrF1em3DoLHPhO5AQX6faxAWZuac8J7QhfJ3Ou2IfGE1ZAZRB+cNeqxem
b18w9QNpP4gD4SYvHc3RBZ15FIYhiD0bMBaR8XFi2zvSjFTm9t3Ab5bxyYJ1gGBHdWZjcSZhU2KO
+AElIG4nBYx3vsjctfKVPl5y3F9WdgP/hB7AEbN9wox8IVOmKcYEC4pVauolUgVa1uSkfqJf717A
ns+RU4iStQDBWmXa/nYeyvXtAaC5vaqm0YcUP9f/1DDH6loXpT6oKjVIveE6iTEzX3z2AspF9FAn
PPGUtu1IM8+MWqiS2Z/fisd1iUGn/wxzvO0IsqFORmFBAO0eZrBpTyk476b9UDL3t1IWrspu3VPh
F0GyGj38Vl2oBQJcLFlbr7hkqE1wDjCJRZdCRr3eO/sDehABZ1Cf0w4g55ubecl9+mOA2L6W/T4r
FwYXexEKJDFGsi1jtztthOXqgjEzUBVWTe/8/X+rzAoxUnFD6qIbzaahovEObeRP2BvI6Q5ZdBmh
yy3ATOHIrG70d4LTQdZI+y/UjrZ5EZE9odAEF+lnO0RhUCk0egZuNIcEOrKCjLE5E1t37pAE7RNK
POeQeZtJc2tCIoXpd51EFmqwvHWQVtUMTI2swDXRZxKPeSFBGnQPQfHKjv2whwW862jkmTwJ/HXH
XXMlBH441LkoKYkxoftdmJ4Wl/oGa4NYJplDkTvmAsEnkyxTXr19yD1FpG/vfycNIHMgEIVaGGdw
MQYeX3orF2uydCWOJptnE9eZvTphs9CLzAmtnCg34bfjZC8nRSaeviro/JM1pY9azTzDu7ogQHgc
6HUYd44hYG7Ka5z66akqsI8dMNzlovPra4abTL++VlDJIb/bdbkPTGbg/a/OAgjr4ONPpBjLlxXG
xRw8uSPDYJVZg0lnRCefuVQT4Uc7UM2Yl9znA09PDgPGaMKllHbAY72ySxReuYvk8xttS7jih7Qi
ovQuoi3loAkedaG3Jd9zRTjGJDg/ev9hOXJsp9YJUEA5BtMpklF5tI0mdmw5K54uehvA8XoyuIU0
bsayUJL9QQonsMpi9TPQmXTspiQkjyx41X9/aOx2yfwrd7LQCJyJwgT8VgGfuAqVjUqb2YJ9J9Ax
0wRXh8D85zBAbQIFywTuJxukTMacPrwNeeVnyZKVBaL663e8VGMOJJuHzmkTZEzMrbgB/1qKLQmY
VcE4LXqWqZGDSBgqIIeQQ+DSxG8g1QyMyTUZTun988aH15nkGwLgE2B0wCkVVcMDlpv7wjal/hxZ
GLR9D7RR3F+JOudC0OWlmUUM1fGPy2PQnK4MERn9MfjZuszADIHOcrfI7I9PrJny5M96PEWgcyB+
C2AXepO+PTWZg+s4t7OpLGP46kWGo0U5/HmaDsAiK8zORcbljMVh/5cAV+3K3NGUx2tgtmpbHYtf
ywoO4qtu2oIcOu/cxcq5k6v55NbRnKpqZT3Y+sYeRZaZxLFADX0WuF5tlJpFZcCAwAzSxgENYy7B
880jByb1LFGZiJBLoX5C/3osvQfSzPEKmRRwHVOFvIwsZ14Rz1u2fNWSIb5e8Tv9zS6yZAUvtolW
3DDHIZU88kECcj7ixvXApTjyLVkpwOfRjz83BFStBTWHv3o3zL99UV2555spysVQ65Xo9dW+KLvk
rtfYJUZ/UEHCQW4YJuLdXYMxMOOUv+e2BPwVWtBc26rF/vEsvdd/Ju202/gqWJeF65Grhsxwd7BE
qakVUeVnsEkBIOrB8qODpoCEqzR5WFWkGkWYqzwqYPjVZJx3oOmn/LrVLIgMPw7+k4wlxij0RxJT
o93iqlTgESEDGSc13mH+bvtiI9l6uK5SlpLhxaZWQshJB/zvE5eEJD40gtRpS35ZaTlbw91KlGF+
fkqOboR/A0jKm5J5XUJFJhp7DtRYyjF35UmRxWBdUC7xo5ysHS71vlzxnCtLh5vFddw3MyRWz1qZ
WeDXbigO4Z1/gT+5SoCaHbxdR/7vk4cBu/duS7MAulRAO2aZEKcENYxppEAAKUEdhPd1vmDDmCkr
BuT9ka9WrHG4TRjOQFIDHqvPihy8nNY9KFgBXQRS+32pAVxjBe4TPAc7QMX+TnSGD6kLaMN1Wm8w
SNQq1NAODfH4fGgIlJ8PQ9tmvRFiezNBzVxNyBDtsEMwlw5K5YzmxGKIg0mBwWA+uAqbcTqW5i0F
qXkABxxoPyTW9H45vdXAcvRQUmILi62njg5EW7ppKBg1P6w0yrlfsQ8LmJaC4t3Jh7yu1/MhOJ4f
S1Pi2RgNDKrMPis5THd5cr3Tx0W+pYjDHrj0usy5leodjGYgVdqaUjmcUBuPVAs0VK4vGTS/FJax
4egT7B7p4CYoypaFGnA7NSwNCcdaIz0xN14rAUzQasLFnNfestfhwIEurT/hKhglSZsCsNcqA6PD
n7VoaBXfXM6lDBWO4Q0tONZ5sKWNSl0pFa4uiKwbj34ewmcF+OOLiVMs/gBgRKKQCLpbWQJWA+gl
KA/2Y9lSigJCmltkjlHd3EhiPJxLOI5ABDRaiasvPXe+uhLDzx0X03UWfGfafRzaed08pdCAA7hd
EElolHpwHzJgJN/nbki8Yvh0W0RMgrz499Ha+T7EFK6wLtRjyfupxQu0gsQV3mwNkrnxrznZigV7
4ccbyfMZt4Ug4dQAJ8BEFtNeLGmH7V6C5iCIL/Ig+N0YKPrcBBO+tcfnLW4p6a7rf+3k8iG6Iyft
AG0OPZwuwM2VAeeP3yYVMQfoNlaObvk3s5U6/oG+DHGNMpWuwYIXmh0z1BwtNVjcHYSRPqwLYl5t
F7Zw1rkU/2LGV0WMVya7N9VLj+U32xEgP/3tdNgA5Q5KH/bkF2hHv894zrJMDql+HLsK8o9fNJ1o
1QkDZY+nW2UDBhE08Ak66aIxm33wkS+J46QKxd/lvd0KzStYZqdvyRGS5k9pzfI+jahhXYEH+MAA
KnYI37PxX6IEV6ykXlXHgUHivVJeK6KimK50zQu8Ls37O4JS/UaWhVLMQokb3vBMaNwzHK7xXWuD
CWuqIMqQIOR/ZZK06G8MBMlwmtZV7DJlJs2Q3St1jbvtLIngEy8GjYypXUY9y70ZmRaGuMFLorEF
cc695mvlNP050cTxVESdHZ3Uxc9B3OT4/3nitBLQdNoSVK9/Xgki4aJ4DM3D3bt4mE81a2HDwzsD
Z68XshXbBHtTWaP1I/P175UpuJTUpvBrRTlOEv7RBNHeL83BtaO+TzGEI1zx0NndhcuMZrLhoUPy
LFLZokY4QNjYjcK9f3z/jaOLEhKjH0WjxrpleqxTiWfYxPnnqDbnBBzTPgVFx9lj2xUsoQYSzBRv
yETVnjz31HqUyaEZUyu7lQxgIVLD3s/o+B6XtXRjXyKgOTJW20j3MlQMgJ01S5BQn2VcpzNoHeI5
4XJyEF2Li3m32rezomkR2uRQLhJnr0GaBIJEZuHM2tl9XVKT1WaFpeQg6DcaGVL7CWvG/w3ztWpC
rwlZnQu6g7Z3oR86mvMPgdyW5OZjpwwGS8Dj0MNp1TCqNl+VOS6DYn0+4oxO7s4tvvBbeW7Bgyih
fgK3zc8+PX37o8u+dphidcEcV0/ZydCrwYetLwkJiTrEF3oLtx/9u40TXlSTLHpMRJuqwhdbpcAX
jUMyvpTsZ5vlDyiWsKC1Df381nopWLghDipP39cLFGHINbGO9h6B4iVo/xSsoLaM+H2cQMFvvmad
wLc7CbZmSH5NEGJr/EAA3eFqZ6ExbmcVLz6qk2j99WFb8NYammI5OE2h47tjFgzqyziEJugKt1cn
ftLUdLUPcWNKjuxhJzCAxJHg5uYvNHL44PgRg7xaxhxH2V1UiimqgG0mSsKFDrH9gdttsqDwPkkZ
1bzAv+Jrl33LzDv+wR22KCnwmrCaHa5Y57bkO3+NDpSCwwU2Es7l2KEjAuPtbDJLpHkGTEMZbTRs
iT7LyPA6ckts7DrCsH+/AHs3aBEzYATCZ6H04+rm7bljI8ucDSF7+eOibuEZsaLAF2gxJ125F5V0
seeiZAU1WaMxomHQusEbmrxhUsxEa56WCmdOVLBapHbMQBZDZXX2wdXuDVSMW+P986Y8BUgwBxN0
9M4XgKJ/yYbyzIHHJ5mRemltMPHTjcM9pEJ6ng+/WEAQWj1b0l5pF2ubckFMxRRqkva8tBzX1+zu
xY55NhGIrkXQn0fa/DKGhA3bnWLF9q8Ks2TBv9TUw2Na6tVB5cbKrVpUA02c1G7z+BLDEs52VX8f
vrDQeGB6EyWyO2lYWiwqETz7fzoFvS+YsjIymzYwVbUe64Z/zIq2uePQiT1q+lCcUMAFq1QoOX8A
GLJURARQD7N69mNIa7OcYVtBU90Ztfane6PSpGRIMUS534mNVCPYy75Jkst6daovKAplYIm5LTPk
6JTStO1HdhS1RzAX4XMBAIAGEPnhSOpe6b+dosFvELlqA9UrtxBbg9N3RA4GcKRfsIt7So6HvF2S
zS+56FaH1SRGdxITeWh6wdCNNL4DTIq5+3/kNduxcBK8dObbpRddbojigLrWVFvExwlakEewIxG5
SALysSjrxt/53nQj3JWoq4oQ0uZMAlKM+TKg7g7HSIvTFWVmA+Q3t/6K01OA1mKY8awpSEmlYN7o
oWlddt/kouWBEo/eNMNSXPY02W0OAae+QwCEsfzfOQXm/0ZSpt6TMlfF/XLnumveQEG87+i8kJQd
KPMuu60C01d4GLzEvB5QEra9MHJYmZ3BLvEDgvAwjiBqoJPkAmGkB5sC1wWZ9387ksrNZAQQEEow
r9ExoB7sOZR016XPAQe1J0jbB41+1ppMqVQZqLzycx1NgrWTQt7R8yYNhxo2HNhgMWnYiyWtTJbv
6/8WT8ChduXRR468lGi4G47fIiuniOJB+Qs2+YHlCbDIZcyIP3ZgiFDxRQn0uMRsdkBwfzJdw0jy
FQA8UrE/JFKGUzjfHPuekaaCqXIq8Mnqlwoz/x6JN4/4qW7kF74RHXEschgVQunan5NFYMCye+rJ
+2Vso1gpjKr2/hQb/OtvldPh267jBvx9wC1qwhRK7zL0LlXo1t+rLVYKO3F6sw4KL2ZAog8q/uIe
NMSl4URBzDzZ9Djh2Fqxy8XdjJ4n3Y1fh5MNuHkygNDFKA2uiM0PmypL1mcd4UlDtsuP1qm3KamT
PzfxmmrSvJkIA3x3HDHQfW0XmUMz6nsUgTe6bOQdC3MrsiUErL1LB2cgcDO2OE2W/qvbuuwp3CVZ
bXbSnByEvGvTaYjQz0ITbq6Sc2AKt1tc1KtgPJStJ6RTtxYPDtIf64Kol1PO7T1y/tt1aJFq16Fu
of9Uab4GtKeOeaPVV49JvZZpPzi/EYJlJjttpOsuLeQMyeIGtSUaWcV4N/Tm9Ov/P7Aql/yFGkvq
385ilfR6OKYrhp/wrD5rAClUlWWWcIzJGQHdyOKbbBnLrcfAnvxERFu1iImVrXWxPUNFmiZufO/8
1+ZUy+c/VoulIViKt1+KXJdJayqQyHw1ZeLez/s1GJwWi+NUrMMtdhxghy+rg2FJ/pr2bwbo/Sor
m3aDXQ8euqO+QwhrA5VJ37jMHWR0ulDdCbrVnfTmn9Z9SOZ9sg/xW8wIsDx/mz8bGBzsf+ZnXHYE
TV6V79dijXNgMexwTHVWxEhkGuiwSc3cf+zcVV5bJTDk5CWzKdDWSM8Rt8ywLgYv54GJJSkSeb8C
wKYW7NpRJN19CLrCeTZNbgdQsj7cAW5+Z+EyOxP3vEoXGItVXBE1yBNqXyQ81J1Qnr26FY2G0Bw/
9CMb8FX7gTX2JWRSeBzBJ1J00pWtP01WeTF73OWATLKashoyzykkZaUGPPi1uO/LKJdJJdEcUssK
HEQdZavL0RA/BKL1zIOCpQuWebOS3Kobj0UFMIsPgJpiQrnwAIDaMGL69ZYwvcwCO8GPNe7b6xIr
rWSfNHsDklAzukHyNEanmBWSQUvl0aS8IqF5mEF5qk2Wo8b0F29fhp3oYTdLmATnZ8/hsNbsNDZL
SlnbfvbO+5lSazSjMoM27Pl2f1cxXtiDBA9HrhMz1M6OgwVjUwsQBORDfEBAfYE4jZW7Ki485JRs
kZhI14jLIB6LJ+ukypaqScd9h8Vgs67KwnOHwPWf3iHzGoPkpRquYL8V5WEYorEEXjb2nil2V9np
c1nW3ERItxdtBPD0UEwuZEuEyH8y++KuvWrS5kKrFjprTWgmgHV8Wz46Q3MWUXLcQ6TwD6Dlx2GL
dNGlFWOufLAEgrW29Nm8YYrEgUk+fOfQbxO0Dbwxgho057+/31H5gOeitQFNFTL5YauiD4n7GYiK
W8aRDqBWkolRH5k5B0lKwadu1f4TBB2QQmIuZ5JziyembQf7MVScPIu7c+COUDcM+YAkAzcXqMuL
EVbEQrIwm3CSNlNhJCZSY4WTelpF1m8p7TBftzSTn0hogrm9IuC/nE3sZraIipsGjyj0tGOotFnx
9qmCclsp+Kmby6ZRXnsQKw/SDZN70vy3GhpqWDkDNjmZAJ+z2qnQ/nTRp8+WYKnoQQnEpS6HBvs7
M2fJq2Dm5+SbMJeHFUMpx+JyGGWbl71cNCwHx4VHxvP979tR8Ro8qQBqLGIyPgZfmg6uRSCshkP8
V4k83RWaBrS2ZDjB5FAd2LkeLBiLrC8eecqG3hH22Pt1I+d42o5MuG4oHgOe7MMWNKx8QyycM8NO
ho12UqyndUuxAl4HH+Nvmy+Abivcz/e3prprSUWdoDpOPwO4cMghYAJBwWpG3Wgnjz6SM4bDQfvz
j0Yhf/EWdjELyHYXbieJSnf63+rvPvfF+nARX08ym9pO0I1qxhFGbZ5c7aHuqkhxdbs8Kvx0ETjG
QB+gPsXlh82jydFBow9QPL40a75TA2JjUVQf4Zo6/wdnmkKgzEQH/mPYva7ZM1bWm5a+L8ofqN95
aY+8tOkRl8K1qRBeUM7e0AS4xnxILcx77btBSLZxa4xxBmp7QKmoVvYGh7csb8/Wd1hizUnaDcBL
I5BjdZk10Xwerd5XAzR5tOlOUzry7eUKglc4EEDoM/nIkxsqmgJSvt8pFPOubZ2kOvmzGXIdqaT4
o6DrtDqA4JhAUnVGwBfFTsqjkEf96JLcRZVn0kkGUtJ0IFBHmno+frZF4T/GHU4zlYUfL6JUv0u1
Bi+PXFu9dSTqhdG8mJ1LNuijql/iVK+3QN2Rxinzc0EdR0XoPCUuggiYFLLz73UnuPRAK2eraoou
xtPhXLRQPiFxDWmNVbAMjz0W8H2fABTlx6sg701aLnBpuLofuLV0ix/PcmLxeiRU4MYux5AVwLE9
q6CZN0WmL5JMPpArOdctnOw9F9nsKu9iKVKy0+/Dvrzf/jwagq+cRkV2vAvDtyGaR9sk1hLAtvyM
wT5SVygbeuGqpeMCmDWll4/o77twAAgkrImoyoWv/eYY9SLignfzaXgbixQXYi618rKlu5yrcjNK
wRL0EXLDJmPGZgx7ypt9zx4izK2tFoRvtQrvK/1p4DyrigmIcELcqkGob+h1jQiKxDNLHy+t18Mz
bMfik6n8swbHwquHbJVdlHl2Wxw9qJiEnOJAJ0pf5dKI7uwneSQvHDdEhgm4lP3OwjzLvNVCnsn4
0Dd1grdPknt702qiJ3VMA8EqguPzt86Wwf8UgP2sy6jYwqVEFhbzPvcHzrmWHVmKokf7ayhzFGyw
JKK+AMdCBodY8qmTx7lluuDVPzm9kyroCEtM4rU37euh6pndRYM0hM88gga/vUjuRcTKl55qDs+I
d8CqSJbQDJDTXi3/88c2BND6wWGoO8tdlky8lscrIZT+ODWvhVd5QRINg3qHyJsB+eFOIy/cE7Eq
b0zzuaR+Ca2mFlNHU/IaQ0QwcSaFaJywpZB+fpuy3CjJ2QWhGvgv/CkghijPZxfp/+cuJL+vk75T
IKxWUS5DadScn7FZTGalneIO7bP5V0dNYvlj+O9uHT+ky0wJ5Jf0CWUa4kP3aVWLVtFW5Z6ysH95
ObryZsgCMvAp2lWhsUYIapwfbYr0UqXuJsLI/g+UsrZGHO02pt7az9L4nEBr4jyNF+lIfiUtQAxX
EQOsJI0qa07mzZpFc10fWoSEE8MUOivCxyOzd27SxDUBRddKY4gbre74AZKv+YCzmVmln020JxdI
ARe1bDxvWamnZz+sjR5F+seZDr2dVGO+gDOk4icxcb/z/kBDx3UxolTAqR9Hj0hb2++be9Q1xXX3
15YUYlY+wtLb/ybZd3uoXLy2WlmArC2FzoR7CHPJvAb3VFTAZKqNLeSauPtIFtvX2cUjUkyVK+5f
yVpNrtUdc4alKHGcBKXDLmE2XMa7+84NE86cXBdC9jYKD7+WRDPufLu8fzbhpRz7HtPkF/OrFd1l
f/aqZBButuQxTBqLdZRRhBMoAn7FZM4S2GZjkOPsjCfUYdw4qhGW0/AAqAS2GWd2cl5y8EvLULfH
M2cb1Z3DoI7xibeCH/4pMbgvpUIp+WkY8M+VPlX80qeyYjnK3DmGkn086WsYKk/191yKlXMnpzuZ
1XZWBSVNR3w4b/g+jyrf+VYg+p8FcUJxS+n2+P+I2W1V6Pq9w4DqT3dcWXpQaSxajkps3JJKktqT
n6bhSxvmF1qH1qJ7ouAyjldDRvXdLcFNW0kKTiLX05um1gGeZxiUUUiZaZHCWml/B+uy3ZZhbtej
sIoUpUm/pS/pZ7iADSqYdzOA/U+i5Dh+p0pxaFrTm6NXn9thOGhq18NHdAea1RbGLfBTqsq37twQ
r75xVyUdfm3UVT9yhpHQZAYfZTxkc8nvUPLvIkjI3TW0CcjTYEsou9JA25oYhA75RFFe7ZMRjdmu
k9REISpAY1EIEMEeDYZR9McydNuNxxa7hPQBpwYh66QL/4yen2yunMCAZAv/KkFC7nLqyt/3EJbg
sN6mdVUpsPjef1TlmMgAIjfOJ5lhp+gfI08svftrb2eMBdLkVttyTn8ng0rx8+e7ZsmPshv4DbrQ
4vbtiQM84EHP0okIzX0cFHexPjZFzldKiyzVdIBa2YUj7HupqknknXQ/FV72r1LZv4yMvRjzW+VV
cHFNChRrmIREEaWVjOaLEJ5VgOSKmYRDPmw7ahrzHk7REjWTOR7ZLk/EsfruJ0ZlHTpKMAKAusTA
wvEa9y6mcvjxp3b0qRkjkqPnYAr4EHxN8DUe937anMHyuKhR1yMiBkTPxEX/2OK929rLH881qGff
qf7UwsrOTq3Tqvrz5uWWOEJWwG+l7AjId7hNu8plHM5p0WsywnB+v0Q0cQF9EL3nwHo59s3s6ff6
P15QQscg+j59Cb6qc2oG+8wckjkzi/KRxEh500Kw0KkzYivFy9gunLuk8pCDvvbHhsrh5OFi5Of1
ZXi7DoHa4+hHsac5wdp+8M7AYEQeqhyEI4Cpv2+3DuHkBOQFJArgujQ2lBSXxPKzwb80/jEN8Qll
pwT/H45XmRCRDE6ifL55xYODJIjJJMlWWq7W+06J9CO6Z0cD8UK3W/SwYWB5jA0+MjT8GtbhJjjp
AKjE/yy0QVXJY2oNcCf0kvX7fpYnBiJFw69AVms31NA0F9HLQ8czdkMr+TbXUu0VTdfsbxvpk3yo
QgWtIvkIFcxypJFsyRmI3OLNf2Xl1Qz0OK8xCQzLn99mFkdY50wVvqHrj16gBIdVwVOI+jAcZgzZ
QKbNL22iJVmMG/s4OJrq+vkVlTatD92yTVKf2iGyfjBVNrahyLwsOsxED3yhPvuocsLsjArWQ1GC
8ucXQV9fnq8IpKd/Q6E2WHm3yHEu9Kva3QRrQvEI36gRMqPb5XXBzGPPZVCSEs0+7muiNIhPaWMJ
O5YNO7bEzPErksCO5xfHfhMub0LmZMbKyvF815u7GBXQ6mo0nKPm0vFSCf+i6uDW6er486QmcNEi
QQXyxPD5C/zkLPuAsEG+ldNaP0Q8RmcARqozIKSTMf8lXOdH917uiLMtUuEYNamkcPC1gskHOCnx
xAeRzaeV4J5Rz6+DxxrOwSAzUG0XQV6o1MOg1jQLSrq2zTArFb5BUu6RJM4j7X4A71RT73Hdy6lT
vGlSLW0cLZNW0NE/09ZcRILDUYRKYcv8gfyhswWF6OYvo0+t25dhBsynmDj1jIp76IhXzeNMjl5e
FNAzzwluqgQRF0+urbQSDOHwj/wQGvc1VPb2YgQ53v9Bd3DefZV3RY0QW2zVfqzJiYJsn3gderTT
f1Ul+BfeR7n0hjwjL6PyvwSNZk4kk4Tst6rYW+IVb0mJpEOEmFF/EJ5mjw7Ywr7L0DOn82/Zxkll
mUY4uiOoLXBdn82JgB5NR/YdbeY40z2ld/P5E5/oXyHsy0wLSEQLZP49w9872EkHNTmwYMDm1pyn
lglRxxy9UfQJBfzR5KqvtL65VgiLhUZNI4f76/VCNVKQzvtnQGwFHzG9Zrx5M0n2toNcHml7TD/p
rDmMZ41TyNL9DUnxok6gPPL1RhS5/Mu58vW/StztMaYYFkBS49zTmqulJYRld3/X5o1+ype0KW3x
hzwPgABvVHCIlzQcQxQfj8gPpHA09BijRTGrX4ehJrkKRIqHKUyGC85tnKBzzCFnkuRuorg7UyjM
ueDzNBQE0gx23rxzlZYv8Xt9dFpiBL5qmpCj+5SdP9XB2sQak6UgpEx+t6Vb3m4nUsP7EsOitS/s
WinqoFFGBDuYeS0wZXD4d8g2jlgLMmvxoQUfQSTcF33CeQn/4JKX4+PCUoehPHCrcXZh2nUDUJgZ
0HMR4uyEAeGsN7fAnldmYfTpdaqzXyMUjf5h09ATlPdwxdYlLuzNisjl8MjCpEsZY/F5+KUmxfj/
kiktCMRFp6JfwK0M6JkhNyXJNvjzm1d/QPyan2oz+KhDc5hexMxjkgV3kFA+7kCLaDHMcFTD30Ck
uaSCmwExp12czvoHsyqKbFeW8avHBiN7WRa/5u71kbHHpycOvr7ymqdO7qr05QxsACeoiHgYzQOm
bBJZtqUSQubcisHH7/TsFD0PX+kuEOBSGmaxHAAGan5rqmyeGZK/TQu0T8yqEVdRx0YnRYAQ/U7J
L/nGByBfUlIeOukHTw2VarygyTfj6v3DZLEBnAT2N4i5pC7H/t+YtwlhdGdTCKO1DUHCC5IhQB6Y
NfaA7L4y2jk6xT+3RRub+BYbyxMa0oTmaps2yOQvaRP7uiN3OBL17gidVA44uQFm7FXkj6Zi2UmE
6gP9VAkG9KAalMgdJdO3zf5aJGQNVfS6QLbe5UD8Fs0EB5Tt9kFSc9i19Ib3qkNo2U7XMmqVC8db
eSsI9NSD8OKQcOArsIl3ucZP/BqLGyOgQnCHVK4HR5YnHM44xw5+0bN0tXjki+Oi7CqRj+FhMGX7
zk8aGUuSy7Zevn5wTibq/iKOW1LVUoOHR96uKhvc6ZEqOInFowai7YfuHrCZGevVtbwPDaYYK9Rk
ivTIbqIGCqWVJ4EVtNwxwhObR8n/i3JYIV59vwlUSJR+Q+ksK6F2JwCNBLiFyP2qxYnwSoQCkrC/
nEWiArzanL71GH9N1k1dDoPxS43l8/Ay42Z4UK3VNCtPS7yf+t7h5+IRadBgf+dYPjds72OCpiHg
CgJUKbhZWDDogpFakouQ2YUfMkKI5Ipr/7LWAOFgxkyJC2BZL5+5IT2lGpyb61Y4tAXU/6o/pvT2
pjRgIGlqpUXTigmA05h4m5GBIGn3/MqfsNI5Xk3jsMh/3zqPKcLnMs9DbLHX9SQWPcqfG+yUZYLS
5GG+Sj0RlfVbsFXNxrw0IVw7uNPz1ZkbgQ2ylXri5leSSps8KeeG2GyF0Jdw1QVh/bUnsMz5jPbe
07kHUmCygtPXQsOB5YzDOmh12gB6Zf1evt/2rnzs0/3pMXcYgSXNvZZJxw1T/kUfQnFwXXHwnI/0
RFoKKW36gjo5OFQUY+n2U6SYbNxeb5IO3afuK+W4EZ1W99spCc1qRHhhryoAOgiZxd79dBK/sJKx
n3MTI37n0JPMkmkw/eFZkknPTOeFChRtFD4opyTqP+QdD/SEHDI87BujHNZx7YmoOWgpLO28enLw
Akop+h1teUrcw8Dzk/B8jq8cW4U5SYXaprcLh2Y1cDM0+pn98ibagCaF6WErIeoGerxKDJvpXSDn
AMDnXNf5M+//OYsXmeYNgiVoMT9d4aAoiE7iuN8/GkNMbFkAwSDIfa7reqae58CLho8CcGACLstZ
Us31Vv4D93zTFtHKiJ9WoVGTuG92nCad1CIDsrzF0lqUc7vJ8F0sGuAM4FpEwo0mwT4R/c4/JVez
CywhgNTpO16yRxFftGzZ0sHn+r5MBLRdaHMCjhS2VCqmh49EibEMn0eSTPNFp5s34Q63YUoZijoG
g/OLLAU2DHJapx6puOJE49J3WSiqokOUpA8KhvoHhDYVmsN6X2kNn5G7xn1e8b2AhbK3iHxwcnRq
VmuARyeT+wCZt6QeB/m5JUc2LWuHG6KxilSr0YX/D0RVu4uTeqqAFBKP9rEe22knVXkKYh8Wglyf
uiEs0iCijl2AafmVe6cjwqQumXQrg3DGbdvq+AVwmpEPy63OEsnTOo/2jJU2Knrq6SPXl4/Ik2mN
+Hpyjgiex8sxZdcMBBSth1jwusImnI5P/Ztjr2OIsi+ii2EuY2yD2pudNQvyuXE8wD31pJbN1NVV
k+0GLC/k/fZ422GzAg3c4TxSqmawW3xhtY34r64db/Z46HFuDscG/BSPKsswPIE4iRU5Nxme4boA
xtGH6oN3mRO+eKEPnolN47ToVPsYczLcCOUgivdRGrkqm5RAn2uZIAGytDgXfn9mMrPooVPLa090
yF48Z2qZBlxjDKeHe6EoaGDQENsvX1DSTJnN699CAj2BlZPKecXbv21kRDuJT49wogbDNm+72LQ7
UExqaoRHjNcgfrrFw8DJ7syAxiAEesmXLUDcttYqhyxgm6XxD25tNGpCtT06kJhI5wOK0kEHwq+O
X8sIDbRbbjoslSG8chlEF1JtetuD4wKbzLxdpwDnZlpalyUkqBB3f/sZacDuWkanphgkK5Ta1gqh
KauJ6k8PaqzcgDXA5Pu2RTVwvFUZeLcJ+QSA0BuUm/80y7E65IDoet+kBr7msGOkFr5b0A60qvvm
TX3u0UvHQ3KekQU4y+YZ+HEIZaMHmIkzJ55aD1jZuz9vQ+y8sPH4aQmDCiDVexBsdp/M3RkU6MSc
kxJghYS+cZP/eJY8Hq9G1lR/AQ7ZbWpFK+u2pxa32l7snPhKIW4dJecnTirmi0QoiRkZIqw79jnn
BY46q8hoI6JYsa5sQoIEHUYrwAkzbedWpSsC08k1l+M4D3I/FZdKEfN6oVnqCrWj32fM74iqtp70
TmOppzD+t5BRe99tLLa3Gg1tUXW+9LmCrguegDctP5WUjAegooXlMOyTKsrKEnFmoXRSVUM9/c69
TTvzWVq2/b9grKwcpDoN5/B0bVY7Bm2FJctz1KLfv8V3aTp6Wca2XNpVYbuGrzdACMpcI8d8zu6q
zvwg679Nt+FQ6fV820q7D9e+RRz/Iy2DJ519dsnbqgiyl8Ya60pdIUZbBjbiwAZSxlM+JXrL4RJS
Wg/ASR6gKKzOj+S329N1TtQVUGON+G79KbzPUDOASKH2Kxr/xOXPTYc9Ez1+VC3xy7AyHxS/hn37
L9NqvD0cYNTQtxXhpiqIUzgrfTGgqamAQ8JA+FlEk+SttZWSPLE5/gcaBmXJZCG7K1nXh/dGRLVw
GcWhic4MPdNuFY0HgEql6ASsMtWzVZ2JLYxd8RHoW0thjlD8cHovWrRa4ZclSCH40y5Qwg2JWSsQ
WVC7MAjJVZ3cyEZ6IVoWCmvyuTbpRN6Ahcguixqib94+ncCpVnEGh7jqEUhL09HjTDUkfV5rjeB/
KsgJkA1FUX7tFm8veECDCN7MZi0PyA9hIXwR465KJahUZ6pqHHp3XrNkAB4zzKy8ofzN8xuvlA9E
nlLk3pbfA+Ud6lTlgIBn1FdSoL3TUaOZJj/R74U9T8DYSpfgZwwXQkeB+9z1VFPk+cz+xPNTyEiM
0hj335urEwOW9Jy4lnz5kQZoJfsUtgFjbss143nPMOfVKcU5ChCu5Tj3o2Uegk1jxtUv98wVvxom
M+4xJVjprgLFODikfd42Dr6mQUZ0A/gap8dQWoN/uDw4W/q5I6nLaKLjtt1aco+D8RZjh8STSaY+
mbxEyzzf6QArw9JmrOvysMK0RizslkooZ82IcjtPdBHQ5Cx7uRZGla6zYdKvfFS5vdgp2fuSviTF
r77mG9hfab7hRNRLcI39fUm/58uH+CmS3ebl8U6oYLJqW9PIIWbL3YleOP9bozlDwlaCVRPunUnG
Ndst531SFaFi/UXLoABMdvlKx2FBnjkZJfEILXqYFg0gGKJwXVzfA70C52TdYvS5oApFIFr/s78y
B9zH3CtpRiRP+Ce6qzqp3R8in9Qc7Dx8ha0d1hoXZKMU1PZkMT7lPSSdaNEnsRSqowuBtkwiMtE6
YD9XXpiKtD677Wx9X+FsVzfbGbwZHKcU5AIiEer7HYDOe1ab7w2uKd8ZnYUQezwgtydfk41QYvqC
vQgFTKWRWcDMi4AFnfGsD10hLEKzg5j82geGvqUcCSo/wh1+LWQc3wcMiA8g0lbckWTZ2tK2q0fu
zzfi2tJxKScHOzN15VkqN/8HTxFquqgNV+nP+IpW2YpLDKigJm9nexicLS0pA60+l/GOMitSMBbK
dbxc6ZBTreKksk8+iZmK21QKCUW02dImaCZy4Gea0pTcJGyp1rM26HKFF8THxE7P+ujqKwi1F19l
DeYu+t7tZyD152giOdkSiyRxy0lNDRbnxgz8jNGiIhwxQHROkvzPjF2eR7YxgU+/KbjFVhejo7zm
/dZVt6/6og8JYSsD2AUoUW8cU9qYbvAjjDuq5PDLkN0eOJ7Q0zIsLX6/D2Q6cw+DhZO7bpp3Qc0x
X0t8MyDeGFbS8ik2adVEBU/CfBsaC7GpytvB2kVaOn8iVfKuhPMWxFWhZBbmKjqBXv7oMmf5Qteu
0SSXSvyKZChm5tf70F8+tjH0DUefKIsXfin58gEQ3tYpUwYE3fvJCQua9/nw/EOT6Qyd8tVeelj8
l8pr2wTnh/OXKsZzxJww1RiWIOeiQ2B2FyQ26sut5ofMWX+I3VyEoJhnOav56T9j9R8Js/BM1W6K
tzNMZo6uZtOoCo2Q+lffzSerBoS0LSMdpyYB4OFiDjIangOZrnf9njvbcZQ4miDpzn4Ki69IVw0P
xePgERWvT5tRBbT9V/9pCcbLpz3pBoITeu5iHBR7facZSKfdRSAcONLVUdwijn/v2uw2mRAaWq9N
Fx+5Z2chPnAbRcaQ3aklgOc2PhnisyFXcGvpT/IsmXzExWVCPBtWMY6TM+7Plt3/XvGYX/EBrs/5
9SbjgAU3JcFJp063n1+/q/4SwLlP5NyQQLRsdVjeIscytTAQPqEL4WxjJvH4lGT5WbMqCzxyTdJt
pKqv/W0lTsebvE/aiHieKY7Rgttp+lDkpX2GU0+jzwOVPPEPkZC1zygNxHqHEpMMobcwITUZjAeJ
2s4svfdOFPh0X+OW1a+pbqp7/Re4OYqxuPbHMfw+1e5GCODTb7Aus5mMDMYDTDHh8v32KtisGdBe
mnNuMuGXm3gAgHsvOZZ0ZKZmgTXJrPjen+Yvd3WG3X8wHFvs6U/mAP37HZlBb0JruJ/oIn3BihYW
f97Y/jHieqfjXJvMSHd+rfZtXParY9+wsrLtBwh9YZ/cBgtuo/e3K7PHQpSNMCHep2dxsqLTbJtU
ySDwdgBYvXqhcktxAX2mq41bw0EML4c3Gly0NUNdqfPLW0t7mbXGn0P0bR6uP9v0Au0eum/8kEGs
tp/Dfj539ncI5OSm3cjR3jxIuPgOWbWvJsgfgdH60TKLI4amIICBZbNjUUn/4Z4R5Fmfgkgo8d1Y
Gdq/pmmsg0n+l0PQrettKdSW2HaFpcMKzG2H3PL2qlIgFcTmHPfTVrugUMrn5sf/hDypEkDc968J
Dgvtel4AYkybQmGZwsDoC9IXK0hQa320eIEPiJM8b/YJGn4/QdNk2fZuT2knWN/dGYm5jODT4rCf
FMDKAEN0JvY92DSc9kIq4pcIz16gNmPtOnY/fs0AvAa8UF/2O7sbxNRMlGgF7HDw2q8jOwop6Toy
yDNlhT9Hc9kQrC3vCvDQELgTcx8ougBSe3Q/FB3IQBfGAjugOa/qB8Dm566MgfVob72T0ZaYMf10
+LP5kMEOCf5mlVCDTL/B/vmmd1TmaVG5PIsKlTXSZAJZ6yMkwlFKrgBeTHUxo3clwWLwO87qFnhD
cI9OCTmX2wZMfy/oo2eWz2TZpnEhfJIfCoKOdxd20bIKl2ocyQlD1a2ZAa2wnbfk+HxiErOJPv67
SVPw7VwVrMKEiO6Yp7HHnRPr/x7BgVLwM2S4EbRO6hJoaqDXdG2/KLqvbr+3IWPcKtMS4F+XXCLk
EN4N0w8/ZGPYURMUDUXew0bSj6a3MQmU9wvV5qlO1D9Y5nkTrRt+JPXzjKlTeB8y57Py1/vzcdZz
rzyn4mnmOH0uQr30vpUNq6urO/QLi2aNiaezXnTpOgb16oLxiE5ApgFEuDC6IRMKEgkjm+QK5QHV
h5tRtLtrmoGiQXHcSpwLT2Ote15b+ZqheOOnYmhb8OvGl9rcW9gUtmW6bhfwWuM889WmKefaTxdM
W7bAPWZU/hrFPFhN3urI91Hj3Qbkn+Ekds6mKgO4HNemZd6bpQ0jC/X1TSQPPxCIWspbiP35J0iG
aHC0pFC0hGCCGHuOTst4VK1Rjv+ifohQ8RB9nIUMBRkh43I0hm795vReszXyC9om9bBC19ykweVV
/LCIVA3X/8IdS4BzHHyehhV3nVEbaJ5WpMIw0umzvcJYL7fEVENmlx/JuboNZ9mVKjp5E6t9Z3ib
i/PxlVrW/B4s6s1N5dSmoW8KzEd2htROZvLo8LKeoc8vJA1n9VtcS+7N0PjktX5SL87wIqHNQ0Sr
zKTVgaQ1woZuTJRQesUU2vLvjpbJb6T1rQEnQgTOfb5oFMZ6LaFbeX4+RXmlTZ0rXhN0ORKi6S4U
99A1bbDllwewGdTJZkYE1+F4QLkksNRCBXUWGjt8/IsAlsnVbZeqCzr9fOYMGwWH7MIs/oXC9MFa
9mOvLBrA8xjnMYyiIrBQIItaZfZtco8eL0wzPUr6vjtfo14jaW5LaIJC7Qyr24l2VgVFmxk/5/DA
jSqyScAMtvEzMxNhgz87u18taJ2barWJnHmkTjMbGPnmS4xG9c6o/t9rsPuCj8NDnOQInkua+9RH
hmunHBz1ydXRNy4j8DApbLsVbhrj/C20Sb70ejjiDTPnw82ADitWJE1kONwRYSKOD9WdDUvE9uLE
uX1Ymn50XDHNfUaWfa08kX6hItcfJNhXKyNYMQZMUiaY/glYXxifcPs4+LUUQK/vKx9U9iTUxS21
n1RuhHjHsp05RMgVK0irn+QnfdpZALJe2esmnK/7WGy3Rn7CVNzpNUtUZpD1ishiyrxC1zUa4HoX
X07h9svAZW/MPaEl4BTEhyrMTol+ZgzQvZtOebo4uyGS7tNBtxB0rH2rhlAKkbSu0T7oJxgF1Kd4
FIe91G/X3+Gr3nmVF/HPhbsRxnHucIRbNGtYTdWiZc1IAoE7ew/h6V7w8ceHoyxrdYjORlLSlnKA
nNioh6gqjy97IqIjwxUPbZjQ5ukwDJBotN3TTSBXc6yrSMM3GJXMj0R8+1iF3a2ZE2VQ6MDWDwJv
X75Yac6xlzV2AHdhd5w+01YBRAudqQJJGxWVbggKuXvs6LUh1gHSfz3S3syxpQVxWE0aTPihA+oK
AMYNxD/MpNdK3r27pyIifhjtpVJJgi/Bvj1xyz1yczLxGsh+OO6bRB3Sf4bE/ofXe0wVd4YgxgeW
+hbtv1LUclbF6yE5z3GTBHGmQMe52GHFjWtQ9H4mbjh28rMVOI4t1ItDVeOzh05IK4YkVguNYWXC
2vwTnz3s2A/hYFsvSWO0iShtWj53HuIuQX5liLB1h5KOdaGVtNcTkYhSLWGQoBjenefq9vAzegDG
LuObadiVFAr1z1NOVw+nNf/D5fPYhPQRklJbowWlHqy5mKzxymyzPhkln+ZT+QpZiwBao3E5mjib
Tw+q8ytqxlbp8eQR+mHFOv0rXbCzz6MwlWUC2D+SLTfbIMFiplfuHsRiMpi7aa7OhqO0Kcr9am5j
hwFrO5IsU3k0Zr2UZwnht8aaFx1hzLYcPFH0WJ+7CjeBbPaj1Vw686Pe87yxuIpKXPKpr3paBEyp
5Mgo85jcEGDhK5yC1+A5LP8Ky1sdVErxrzBrOpHFz7gTb3jQwrxpbnrB4xZIkHMbVGBq0/MqPugh
gytoSq9ILhLMgwdSA1vCGkdYumhcnXAPgMGKdGwZ0+b5QUKfIGBlrnHT8jgCj7x7OFqDB8jVjYbk
kYo1o+8mYaVdXJSdtcN/p7rETNCv8PIBZNTAIZugJJODC34WpVjMEqwmS+KGDloGDK6u38YoibD0
u++t+rdUKD3650H9XyL+PbgR1c6EMQJOsp60lIR4r+nhIzPSxNnVziz4CZh5Vpp0tzOEcYMSMHaJ
/MALVehlJu4OSXHYsUgznuV4r9HD2UGhtrZFxmY3sfr4fNwdkbC2nQHvdKyc0cvdZEuo4MfXd0Dk
vjwqSJDUiNkW0yA4qo4TSwHu9btn68hFobglydXefZBpFOy7ykMkkBfF0VEjqdGWOuU0YNRV+aj4
RW/A++jqwYFQyHdgE8hVNoYBw2ngQ8QfJSms7+lOkKmbFnVdk/kM+8+DhsMo+dd+3JLXRyJQKr1a
YJgeJMvzRzqxcaOnhz/Ve76BiInr2c+RHUAt3IkfMeg7RLx+pWAK2V6UUPtkUqdp2/bWfUOBp7lC
bgtHXHutryq198Gu2VS/7gSkdeJXCjAQ2ut8tKSCnKa+fHfm3bZo3wcL8JOa7wiPxuEL5Cxd3BCT
ZQ6FijsbdbCl53EsJyKT9AT+fXJiYN5O1OMYGJmtMK1v7er2oy3DNtCQaWeTM702R0V5YDh496Jw
YOSuoSLOo6wPtM/DZIxpmiTsGJ3b+1XbMJoovsSdk3NBw3TjYKdcWqtnPmA9KABi9ZfgzBwBruhf
Monq5T3GmbtZC3YpqlQBZp/pJPn/KKt6C7lOTrs8Sunx+ekMUsnVbAOWX96WY7ghtb9FWnphlUCZ
15nA+LCONCkqkA6qopn7V6AI2NOXPuNdWaLaS1l1TLXDCZSd2In1GhTOTWE7dEL8BcUncWXIxfq0
3atKuyfWK0v/BQnmUkAV1tg9id3FpaxCVv4yhXJsDHMYeN9I4XB4eOqm9/TEYu+XlSkGv13DqBV3
5JF16GeM1m+mE3kiImDhIHP1hYupvyWbHLJwx0OYFISQiE0q/13BnAl1z76HDswOqokhVqVy4PvP
eVmaUHioyu3x2Tg36/dXclld/mtr5yffHeRc/mhk4ZKYlmZQpJtxOHjWzG68kWhDi26yLuqVyeyS
8ijs5sY4Vqd9cuWCk+8gEoCUckfPqSHOaM4HQs3yTvuL2pZOM7pjZpaDL4yKDKh6mkPECwQgq5/A
88VvLTm0SNX4iUuoBnaO9xxYrILQ6tLKGa79Z+lSHB6o/6vMq+FWyRl2JJVItMp000NEsunG1w09
i47087yAUn+momf69oF5EUQ0tZ5AhoSD0VgKUlAFBAxEb31ee6OQ5MXCos9xs/EfO/YtllZ/NlYi
Un4uQ1vl6sq87yPjNsII85OnougKxLD2m7o+mCnMaGURksIxrY5lfhJG9KiE65g6HU4/qzF4mCMj
4IfJNwORWEJfUfVAFFMWN/wwkjLrtE1TDp5UFWsn1SE0o9UyA65zPMnCi+SGRaIC32VvBVYnOaTv
fJmj3ilNn0ZNiIRIOPKpa5f8ayZSJd5XDm3yixbQye0jOHrE40Rk8yqL9u4oodnbbZRrJXNNifa6
+OSFxgu3u/9ffTeI+OHXuCs5iJkLttHEoe+z+RgMME4rGBvhBDir5ReZeRf8qci2QlR4cQgD0hYC
ze1U8SUM3D/rBfaKKas4hhFKGipMS2IZMLj4MAm5OpRCSSSg5GerMAkAMHjtbrY+0Yr+gaU6w2NC
brVGTegmy90Z/5u0h6cpW8TNu2cv1Cg55rHkRiFryyneCM+y+6QlGHvBMWA8RQeR6wBe/RdBvC8A
4nN0zz9Cibya4Z2ZP4ozsan7x+SvHtPGgNyu+Tfp22Ub+swdA6oPCQ/eai47zh0w8EuDAqKj7nNY
HGsLuxkJiclPO70xhbUKCTHOiM84B2K3+OVaOn/iIOA0OUAbT4h8zEEv5Wd4KLyleagmlIvUpiPl
oFlw8xcj6uWgg0s4oewiZMA4bFZBtzNkDSjpXzrJYt5hvgQ1Z5lHj0X9wPi+V2Z35s3QcEyabAUd
tpnSqkVCYBiDsc9InuJP3pkka7YEp4uImGoU/GiOHfL2rlPMwt9xFW40JJr25eRm4J/0VdjroeM9
XSgZ10RcO45oZuT2Wv01P4VEp9Xi2RAfo/klELnF6hNOGaUgPTi/kTO4yLB9imyijKCaAOZCLMM2
Q0IFmP6O3qntkoKo+Prrn03hV/hjJl0ld8N6thCFHXebeMUb0A7xnemy+i7zRc5jvunhDfxIHIMU
eqTzFgt/ECn8oghAQk8K/HQPDbdk/lNd/4mwnQBUYLMJrXVZwrLdVTuVyCxlB6/S0NbA8KGxP9fd
Gz+ZS26chH2OHbIzAB9qVxJAj+hmtlDS/IWolgxB+KN4ikJUKABHQ7EWVoOX0zjkrh2JjvoBNW26
QyXhXw/ktyq7L79LBDa/WWW2GB1IBKxRdpefXrO6lOZGkLYhCv35I4o9l1cG6dCsG0PBRuC0nUYa
Y2Hzcq53iGeCGRp5ZNGyexK3VY6VN9ra8rACms1sVNgVrPa9Zm9LCEhqx80+p1HFTx5P1wnXXONc
EOEfOomcZCXl152/UodefYGAwR7sLORECqfTUcHiiWevi4vXz35p5nKOnwOa38kTXGTsxOjT90Na
4CIL0S8EspvmWAYhrt95ECd//KnEE9ePcuCb0dCwu5HjDtmHkBLJILbbpxvJzQlKcU4JEXFapAJU
VMcLu0yAkco8sSIa6wwojWbnzU7Cyh1UM/THnVxSRcjQBDyYb8FJ5FDziJEtt0oX9GGAfShv9QfS
lx+2IPtn9/Af2g0dxJ6eRfOLK12ETCs1GygabTloRtb4ZyzjxUOP8UP4YEpVNwP7LSBsvDPUokOo
LD3fE7B3BE3tjhDOsguk6xmd/mbbUWzHPDWsAWB5gzwNyDmDX7S9T7yJWfDqbWGj5TjuDUcr/mCT
5ssuwEe92mHuxFcJYOU04qecQx24h+8PVfj0ZMe0EYx0MC0I222GfsWCBuWACIys/nfyw+/r0hxv
YX0RT3wNjlaEJWm4Av1giXhljccQw0rcZO2umRddHqGmXpur6+oejq0qxToQSe7vmn7KI6u6KuaO
9HVtpflbUmqi0ivymd7ZNUXXTa2rIsQJxrTdVI8rQOg+98S4gb4Sm7Rk/rVmKVVX+hlIguiN6OE5
s3QGE6g7v5Y4mM1JQYEN6gPsyic9HujEv02nB/QPgqChtD3RJumsbhTc7rgAol15i1bPSpO6J2Qu
e+PVCDn8cYLRWT6Orjax6uGlGVjzI8mJLTi7PQW1O2fTbBGFbUzKi+c+TVgvDpcpb6uSCCNBYMpc
GxtKlR7Gk6FFZsPB1mv/QLyTHiIZX5291eZFEj3bMyHXL2K2Ns54ugvfgNS1AATxoLnUL8WYt/Fj
OrLAqoRN1H5hpH/PCrAcn98fVUPLROLmjU7ULSIjQxRbJ8uYb4fshgET7fdzlk3QAAt0WM69d1Zd
Fj9Z0KbK9VL60/qoklJAzS2T75D8rfBUw4FIJwP2ROdNVGax/x26DpWb5qdShgn2uQ3KvBafiFWt
2oiirlS9YF39L40eruTMhKmgeA0GuOdeWamwCqTSlsM/F4JbQXe3UZc4iSzabSwJH84HdEAihKEa
0/9joCv6q9Ul6isvcytJaLrl7bZCelQ9oSmU3TfjGwnr8iCWGFuhT3mk9en98xOqeBIcZo4hex5P
JCWQ6sERGvN4O0K4hoR5IS7tC80RY74X1Rmbl6RzPfJLHnFCisr6Nan7e3KDjNPnXzMan09ahm+n
48ZKmTNOlzSbWx2Kth6bkenQCgrNUdb6JbwyZq9h7sPJsmUbjXT3D9OJ3ziQ4kVF2Oof2PQ1JX3m
gdrN7qe+2RueNZfaWJgFm5mML3zmeXBdEEv97obAKbeJV8TnuBBMlMy9k7vfsUZSb9/cKjVVN1LG
EVMX/DCkAK+pgSVPefFvKc2RYNKnf52CEPO+udulZVwmKOd/I+GvJl7rtnU5wugOxniVn6Fvglxt
hYhm5wvL/ZYVSzienG5dOgzpvBO9FyQShPK2ysslMAV97ITodHcPKYQRdliMX4KtOwMzaJnKLL4L
gN13X//XzwbLBs+cjXMt7z/hzUVfNv4O7l9+frzrbLnDjjJ9A4pHICn1rjQ5DiqUFEI8eDqiR53j
8QLPj+KkfgD63XG8hbRpibTsaOAW1dBVqNG7b0bfFhqk8p2x/LYgPiSpuPUcpqS8ZJt0CBREPRbb
8vzuosL1G9w8xY5yCzRa8V6OKtVmbdIC2L/Lf65d/GQ2q7DOjj2K4etsoN+nm18/PZsZhUt2GZl6
wu4PkavcRiFoY+A2XT6lFgeJRs6MxKAxwzOdbxtA0J3k5/QH2RiJyJVTlx8mbhBBo5nfThc/eh/v
6Wt1SFKGxegEahno3Ggg4x63Zqrfl0Y0Rh5iREL/KgXM1k6O/IYFuvlXVYP5+u1t3uSTuTXzKmb8
NqNww4lUpqE1K1/sUInELzNmxk3m7/R4Pk26TY3E9y7u59p+roKmBbwLxVt/6xk5NmfHGEzuNaVV
WwCFiWghPGJ9SScJHJ9IpH9RjKGfW+FL4wO6TeeG5DThptUfT4e5oeROjxBni5ljPhkiWK6QjwWU
VJ3ytDgLMkQ2XGPBwgi1WhVGFMG0YR703iU6BJw8eBm3JkN2sq9ZJTpzqSpGjB5gO/KwsPTFmtAC
1UTE2fvHNFHfVdxMHoh+IVEcSZDMA+OP5qpqJcr2AbBEH3cYbHwB77pNwk4faNe4rUL8HHVLhYgd
CQ2rwH61AN92vIf9u7jTZ3XV1Sha7jvPFOUj9ViiRjioOMWfrqunhXtRr037GOwKQiEJ4e4wQqbG
4GYa6RX+OSU/Ogq3hwt80K7oMi9CGaLRiU7ISQAqfkbO5cgKohOugbrxwMOdqSF/i42rPclpXhyx
6JNc07cz8EGGFVYtPZ6cDGTUVkN85XT2WMyQjoeSszTzlT2e45TA1GdFzU5ZisuM4pQM7fKjFwIQ
T9KgBueQCLWfEHAeGj5LuDMMu+oxZmwP0pgZYsXDEo4I1trziV/tiP2rkCPw/aWyJT9yjillBof+
jfF3jS45N1Y6GFuaR0pibMMchJRIIQN8TW3ZuC5lVj95bfwnuafgIz3s/IYMG9fRyARFhPTaEEdD
0ZTqNHyZ7m1x/lDFNGfBbh8bRX9LPoVfpJWJyadBGKjKtdKFheN857GrZjs8xMnkZul6UxwEi3DC
aQOvnwqT7f5fOoTLqSYz2JVTuPR2hmlsY03h2YvF7+CGVieFNB7kZJkSEnTk1SEFfgvRWqeNarGC
9Iz9jNy4Ulp55CZP/TWkY63cIhQ1Ud4wdxjXQ7YE1JBkI1mlb9UNlXHU1bX1qAfkXCPaRVWRZZKY
RIuY81W7JW0kdy4Gq1UG1pkV4ZSggOcdLR28f3x+wWcEK/dX4EK8klcx4J7SuU8lU+mq2L71dRXq
OVauABrX7xHq4oPXwlcv5Q2qpzTCcdnjzo2BwpkaLJ16OE74U+PIJ+HsxFYWFmVkop0jZfNM8SMb
A3lL7fwL7RVsl0Jsjn1iDOpsWIsiw/u++tUK0uSo3bxjqNYtuFaHw97luWqSSR7mom3QdUutqH8S
r65T3g5RvRnqb14fVxLzt0odkrQwGXR0vKV/7FTvXG2PIbvnOjNsu7I++IB2FP68Pag4AUPWBmMp
LXbcMqvqqWX0oQNJ68aIOsv+icegPBSe3EFxNR4GwYJE0FZQmpmuKxLdhNbySTphrPWY3FzeymLL
x11xjnF0ppA+AQyRM9tUyi+dinmZu/BZLxzXy0lKHLNse0GC/zw78rqB/tthVdUnx2O2S0CIJmWm
kGSHZ2+0Znhkgp6cCf/zfQxinCrNIUPfSKbiziv0nSXw1bAzpqDWoP6TNeNff8s3Lh0Xo8+bpF1w
kYfgOPqQ8PXOOb/EmEpA2CYIm/vJzmMS4pueyJyCaQPOnmlRR5mn7Uob909g40u7TeoW+mTS0kMP
Ok1SuGQP6lBdzlw61WJbf0e/85BvbpREyK2+a0ZAV3T2BhqyFQlo7c5NyG6kKv3xUjEBq1ioJFDP
AwM/aPj+muFEfSeqfGy3XzXer8zLoo56Ck8TRZKnT0nfdR++P8ibMx1J4hFUhoWlEAxr+PnC55yb
Hx+mgWB/9x2iL4tM1u/rgmGE7C2pRJxmoAaNuobl/n9my9X3sUzn1TmPxHpbllLUJ1stZXKLH3WR
xp8Wvtza+L8LKTh3o5GChjoP1uxjaoKTG4K1KkxUq7ECxJKNDvkbyh6FTfrOkXqzIIsDUKm3/cN5
jOoiYRCKQfkj2E3l7w4usyXlSmwiWxCCVTs6ep97ygiAGNZZsAtTmmdtLvolBg4y+D619fXzub+G
1Cef2+MjnxCDvTS17b9F2wTdOYvqnNY76w4jrz5iDYWHLLkJG6I1nw0xEhEHcIMmnQjmPDS2kPUS
AX9UBY7GfhTQvRQ0l9V4GriFz6WMicpSPDcLk63WfoUiwCNGfLK5NEN/s6Cke/jz+DFtSK44SM5F
OUBh+deoHsdG6+T7+XGjF+3p76iaQZJzn/lbYGgF9GtctNZFnHWfw/0TtfApihsv7SqyX/iFj/9s
6cWQkIodXVyAC1iWqsZrLEc0lpfqmoHrmIBpJ4l3djjw95HRINH/mAHLBGSmdkJod2VpmegZEOWv
WnXYK+Vdrax+iAbpRcXK9jWVlVAT5dOHZiTBLOqVjKYsEBN3z44jsv3rDxzb6OKhNSNdu0lXkFmN
90lZ/p9/jN9qch8WqEvJP51o84hJUqZbj6kdNlmVcf3DLfHEvAZHNDTQp/V2icN1+i2ORZGCDEsf
qQNzdPdcA2esHu0cEHrs3lf3u1F97csbxp/7v1O+Zgr77lj/0JvBTR9goZ0/mrYbtH1HATnvCPPS
IUnacaXP6d5K4Octtx8SPbY2iTNQxVIjcginRB+QI236RbjrJyKzSJ3iv/lMUJ+IB0Muqf2cNWrW
wSZPW5vkODQD6Lb2xChuPPPSpC4slPfpU4cYqc6MVg6S9QE7QBPLyLtf0zR3h+BJ7qGq7SFe9VTo
/QyPwZqEKjrTqpDl2z/KQwwctyV9fnm/uVVYCIF2aR3wW7Uzjw4HjjYMzJPPvWmr39pzXasqoz/d
JYkwRyBHX+wlV+YxHSvyXDCGcx11tjzy3qRvrK7gp9TviJuy0CsLQx6NU14G0EXLG1k76PfaAcVk
E6psoNCK6cX+16Q96v1LZe60KvWwkyitXFn65fPFn7gILIfq1H2hqBbaLg9hwW9O1JDqXharpkV4
dKV53OmBfrhS8buPBHYiwN1WJ0LTt3G387fmkfYhy+EthZP0+KhebJeblcVmt2UbBFZAW05SLX/U
IS3M/kV5tvCrBTn0b8LkK+2JHEX62+ZyiNryEFkfxCeXtPfEydM/5jTz0/TVGqUuQME8qjjY71ty
JESQ7+efEZzqPYueP+F66Yl2tdZBSuL6aFblBdN3PrjUFadRArhZby/dtTZl9VNS+e5V98Hq8/LR
TS5b4JSCIXNFrORAggfdngrKM8dL/0+6I5qDqJAwIGs1/YgwZ8FKljpWcpH1Z886J/XHxc1VKAa0
RsQejcwHMo8IEO1n96kuwxYAx95Jt4531CG59lkWD0oLetWXvlo05ggC7qGBQpsUVureyYXBW4tb
QCLjcbotejzBR5EqHqiQRK4MGKmO9kQLu7oPymRPh3jjivPTZW2cm+6q7Qs/XhKa8r03k9Pe7P5b
1CmXYYq0+wHCNMrjIpTFqq+z7nHGRP/AYdxMfKS08f9mhUg2RtQmlP21nRrSVuQZ/bFfxoAJqWOO
gDuTbYBnEFYHN0z4N8NuunfM9PF5xkTmN+3YY2Acdq2b0PeucthrAb6xto7/r77RBJiUpPavXQzb
fP0N0Psa66lCexljs5QienmDVcbca/GsVRfomto4MLuignSZv2j0frnY/RfPLUQioFqdU/WMxUWt
sps35EcMS7z7CwO4VQYuWTDRdS/sLsRMCx57zH+knV7UZXIhnneG0zWmm9I40D2w3s9nIS2j5WNC
XyHMcu4NFWh41tnI5RArpA5q3a5YgR2QOyYa9IqrAHT5C0nybKNOir/FqEPPXCXLxfiEmfwFFnCB
8qfnf1AQKPOFA+xXv0zPB+p/6evnlvTfaCCN/ysww4rrqz4SDCUSBKQBwnV8IWL78dWTdCYY/4cg
qWa/wMUHxuOjUcXpvwnKF7hxfMwrd6lNbEA7HShwO4aNSor2NpZbFxdNqE9gyqy74agFVparXiKI
NZfdvwsuqs5PceOJyUgTy23CjFjTFH1YCaAkHzegtOSRyVtTD4uXPrB9WqL69CfD08y6wCeGWUip
hsrTGLK+hrMcK5aqFEJRS1ZvTipWNQyoukBktAiX8w8BLi8JjMfi04ZlQCx6mOGRSeipepy/I0fq
8D16MtmLi8tEn53Xy3eL9ms+sm681jcdzPdsl9KfEJpGHtXe7WsTN1KnsLTp1tMovMzoBlRnYF8J
3YdtZKOpVPbQFEMHSmp0oFOakMOXmsHLbp4zUCTRYoHblnvG3nw/2iaiIWWBO8D81iXU3m0WawnS
9JolnV7i/sp8FeqybtJN8vh4cZg+elZu2C41WintlotjrN34jaqqEMflztzCNhBkI+AJ+lnNuElP
Uv3jKqvx0Q9dbl5YPo8stW9f5fmvWANbrNbsXnxu3zXCX9w9BWjaE/RteIbjl6bdpnpczp+7TZxo
HV8uKej+aWCh2+AOSh0JuDvgQiNycoY8Gb49T3YQ8NTHBwdHYZ9wE9/iIW5mwkGyLd0ryaJwBo9V
PtBeMukhIQuXX6YWUEBR7JXBmZS/xsQrWj1lxRLYdtlrCfGh72qeYPynapGF6ECqZ0bqGg46PBcy
EPeAo7VOUD+jUPy44gQTt0tjhMKUgjaABfRIQQb56l0tRbCQIFmMnvILf3UM3MM9AgMJKd4wQNQA
oBZPC96HZAnLIqPC59yZ/hWDcXElejsYeXu6b3tfxXb0u6yQPK9No1fvmoSpliYWGJwzZV/Jbtwj
2YDtKKn6JX7PrQkYj/Lt2FqYnICPCCZfmibdREM5yYUmRIvTgGUcvpmhdjfxd4WNuMwTAffBVhkT
BCO1fq7ANf+WnV0dFf3kxAQ0InscBVPmft7GdXEANn+AGZDUi+d4REvi5Tesu4Qfws6XgjeUVUji
G17Y82n7KaKTKKtxHHg1YYN2g87DKo9CvMgTnkgsqh6Wa7aRtoWMUYL2zAdeOOFPqyqmXS6nyRCR
qZamibf+CzZR56iz79xHlzHaNikKrqYbq0wgsiF9fhRNn5pOFIkxM9qsoRHQM3pdvCUKgL4Gk7zD
TiPgzgPv2/g4VZk/Xogm7WaUDjx6P1T93g4QwAOhzbD1a1mbFHJjhqxSXESXRy8OsNomWrFutnh4
dmtNTN7ed32ZxVyKC882ByaX3GAfNKjkynv3Hc/j1UPXuVYB0Wit4bEP5wwoyRPzftFqt8fWy03a
gjTJTvnY7wYqoE3oD7R38mlL5euPbFODfN0TH4CjD3bfUrqgCbw8pIGch3MK60MhebQ/ZsxQhjjQ
i8zhbx/vqCqbt2TTKZe3vzg5m9eSlO5qO8Hb52KIb9zgsPdXKzEcW9lja1A0n/Bn4QPYWK8V9oIF
CgfPmx6Eq4h1rNR0JSWBz6+kkb7Mm7XM0OPzUNJeP4wfGz/Fowt5NXnLICcUREdkD809A4ttcjRN
65mVLeFtz3/oM/QGWwCBAbSO6CSMW4tOtk5qPQYveuJg4tvibF2rcPPJRk+MIUMEpLzzYMdbVE2K
M8qfxCHqcTZvOc9husLmKFvJgVBuxmkeZRrwAszwOHwfjN8uuyoOJjbPtPgHb0Xkkz7U4Pff9hJU
HcRdtczGM1klFa6nJN+YVKm7SPOoZGzJVUNQjfRlFgCgpKDq7N4n88wJF2NhGXZYPTVtWKrNxuvP
kuoP0wctz4ZPgM2S4S6CJ2XJlirYSWgEGNZwhiMOobozloYrvFocQIX4mC17i6ZfFTiLyuMDz+2x
qAi78l8g6kzUiumvOmhFDK3ZGga/nhnwakRnUAM5++cY9lKUVV+51dtbykRGQAfQRYzgSExw268o
0fEAfZYg5NASd1BquGcbZbzCTmx4n41oULo2RkxBtjunX2Tl2obM7UUObacfYVwc5dMFF1v4mlHX
B4dv3HHiZ8gBQCskAqzxP8RYOS3T1+bOd+0QHVpG0UcFGU+tSyE7D80LHfAF/lRZE8ehxtHTekln
eWhVkkPz99MLl97B5+GG8UdWBJ23OZdn6Xx287eiUDzR0KAW0VL3elNR47zCGzkMNcKMNP+EoQUM
Opx32zhu6SiiVPAY22wL+MOJZn6e44z7LsyFhbv36IF7cJxo2L1n/es/WnMNpYgswnbkr3VnaIKp
BriD8GkCtmrm37poAhz+UN7IJ2KMr7ArUV+X9zD0VqB11IcCReLds22jHRxmCNvzWO8+nCpnmNtJ
Egsa9G+M2NlLb3cpPt+RNmFb8NAfup6ET2z89lNWma1pk8EfXGrrXX+8MgTcvNSpFZUepd51TdjE
twxwEcfX8H3UpCkwi9iHnNnIVf+PhDXl7AE4vQlYEH308ZPVkDEdoxl7wMbaWCtjzwYxLxAQgSbg
+2iHP9bQY5RQvPWLn10wYqu4iieNq7bQR/n6esIusfRHHyAqyI9lAXSbrlV/O8Bnfw+HEdvrqyr7
hwEVdVd/o1WRu0MPKLG62PwZ01/IwczraqRQVriRxV0fhneSOOsYeeHIvmCaKzYRYd/ejwOJHOYj
aCYqESC97YbWOc8bFEA2Pwsi0ETefvbMyhpq4vlAc68lwRi321sAjZd1djftTq3G9Q6169peOsBT
p9gjljeQMJNgovMBikZxpH6y6e8x6lgligZRu6b9T4bJT10xOXx+R0BneV/tARb9T47xIzh4kaR1
zXwRjOgF8q6ufpD9TP5UJPz6ryWZtBaI9O7kL3igZFEwxsMImsD4K+8y9XKKBRCZMC+zRPxDxIQP
OEzE+d1VjYqAqiexIGN01B7AoaCC+cSHA2o4Hx0iu6p9nuE8xIF5Ul2Wq1oSKEPF86ioTmEw4cMS
VOPX6uEYNgikGXExoSo8JReo6qXgSjM2d95sNvuR9WIuyP5B8eAwDlYm/PjAbUg3ILsfbD7DCRKB
LEoSrYWRgpy8VXIYW8bfJaZQz3P3u57srCXnIiDnh1MQsY20Y5pu8DbbioOlZakKedG6GRDyb3GW
/geFj3f8H5NH+w5c9iADdMmF/AxZm8FXeWZR4hvpRuhqgmoQgfarUAqB9SIj+CpHgRzFBOf7oLUQ
i+dJxz70asdoLJnlQLwV7ypTib5liTINeNSUv7oJMOP9Y9wKygrDze9a94e/i5plbXjL+QCgr98L
1Kix8aiUeOYMOrCqoHncZl96hvfx1slUYf1BxMwEP1UaXZTIjlZInrZgMAAwj8czVCudgU50kPrZ
MubQINplucbmaXZT6IzMM2mbki0+H10Rbrn/NO3NWosJTA906ttW7UGihlPCmEcrdS8+0kl7ess0
GjEw9/W6iQUC0FgbKKOq2eYsCKx9QjvWIu28b1u6lfpQcuyt5VY0mElrKFCZsBR30qmjTkxW4OYk
0iQrUEcuoRKegfYa+zpEuGGEw4Rg9iSK52C9q0QxvGqkWDjT8FqdqpuBV7BWa5Qg7FsDEMpwL6sN
P4a+EtBiOD2oHfm7EXQILvWMHINfpE0BvkPcJNHTV8xMY69p4MQQwr7aIZhBU1ND3CneuiR1O8wb
jb3Jg6NJysQACZZiGXlGfmsyOX82X/HIkLyGYVvZ4+OKydm2zQGyPWhUmFpGg9B65b8Ro7bFKw3x
0b1kULU0fOxkuR0sv6+uJD+K/efKdiiZpK48mh7d+P/zIySefonGNZ9hZRN8/UUmcGwTeISuRZP6
EiKW+yX/ShctqXJtbt5rC0KxgwokyAMg7lCRbmeInuFh9GVh/1hBmFP5LN90rAba1iFxj+uu6kR2
NisscquKzqQ8IcGkJ9y0GdHTJLQSd1Xy8D9qm0V9crAWfq8Suwn8brHcMLBXmeabHqqtWbEiJMof
pzIz+hM6ddrS4OIT1QwAWJZts1P64wxA/pqQcj18d+FabeDFHCG/O1kxzVlu1c1EvUsNs6yvq0CN
PyP4vW5ANPwCLkB8jrFoMzBtQlq+vy/4DhD9VE/EAuy+BFHmm2x82W+ZCgK4rtcM292Z8PPFIQDg
vc2FoNF6PgnSQtzrUZZ8TJj64EZfNpDiPf8lk9+QqaqO2kFHEAnadhySeu1JmeChfiWQ/oV9AOYb
jUUzncTlcNCCv2V5hz5WdnGJSIkaKFTAWgwYh9xkyMgJYBQMJmICFm4F2hAJ//TzmJ/geoE/LOkJ
0eSOuVPHJrfM4rIxbK9KYyEg1zszIexljYeVltXlmf/3podLBftv4ygWFsU6jtm4Kd/RdpKBu22n
6VyLOpj6K7OeVJfN0hWIbLQn9h7g0XAEuYa26QYgMm7JQg1o1JS3cILKEr5xT4uZvZi4AfhxitYO
Asz/GuMXXMCOung60/D/25vcwPmBvpniUsrH+y6KioIi/hNdZr9HBiSN4Een8OKhnXA9Vn4W3dNZ
URE4sZw6MjzKnvIQ0bX7Dciwz0CkV/K+udAaueqc4BxcilXkbjd4yGTtMdCbx7A0SOwlCtVB98PL
MrvQwzqtsOPyo/MT8wz6A2ZA4QqYOrexUiAMv0zEzouihBN1Z7g/jq+KMV5VvZLpFPdbx7QP5I4b
bLAzw2wZL0KgMiGK7vi7s+KlHpXQ1mffqjJk98KWZnjTxlrcaXDCTqP+VP8VcaHZ2S0Osw0ebzg5
2QPlr9XVik5TNFB35qYrk8Qa5fRs8B3utl7p10NSICPcJPxfw0sNc3k2Tk5XGJKvTVL6kGS2JRqV
9k8GyqIQontubXDtA3xoGSs14LDlt2sjjH2zcTWlCkBnPVeR4rUGgWJPGqK/tDgMaydqGXviB8hs
dizVw6FfkJqH8jT3v/IVjDd7nWn95JdMyXm8LKVLhYRDcGSgoz/B71CcuG4eZpbX0PhGSh0PL3qq
9AeIplk3/+3JTpKXMe0ObXBGnCv3rwD9tNOqyzJgMU4LsbNqsV0BrW7jOX4KoCg2THfZYRwLbmCc
6RHEGyFuJHmr/pm/RM0uzZXJnGv7aNm7nY4TPSJ/PMLfG1ij5kWz4xiUtKVJ2DHEGkDjljrKSZ2S
HBUIWiojc60b0+oAS8x7uP+/XR6z8Ka3ZbRUaFBpRwE0Qhw4Y/4G7kTbPZVJcadDsgsz4cF8HBwq
h9exQ371D20S+ieOL0NJeRViP9s8Mn+dvV7y1bPWG438jwno53AgLgFxmwC0A5wd1vM2T99ESVA/
l0RPNmQVX/5O/gTp1x38DGVFieC6FYyfl6K1snPzcugo5+t6yu7wvECYC1Hw5zExSQqGA/xz3TqK
M32mDBgmEUf6lbYWK9DHKggl6oprFh61cJMqi0sPMLBmVGM+JAvx78I78Djydu2JVTZkQg8PtJOE
JaSoQaBV07/plmJSzXV2nnkaXtiqLtJ4A3Fg19OENQB4dyzXIoWz1isoBXilWxhIVe1DaC6NGnbU
/Zlo+mFa2u5Yic7FiIL5E0/+TXQLIP+hOciImyFt/q0HfEv/LiWO45HTM2q3yyj02ah5prDtrff9
YwCtmm8imoEvx9ZPY+Um74mw67GC074/DNseR5fCc4+xMJC0Hb7mSbkYsDG5J2qPpSCIt8WMtq+D
SGZXzUSvLWDHwG+aGhjhqXLWi5EPBXQTO6cL9d+lAO9tMxOjK37Nu7ccrx2dUK4pkZVejP/ufsHf
eZcwUfNWYR9t7W4v/MHQ4pVLQyzeP0Oi7hFfEcT/qiCD/wbM/TflxXLC0PmFQCP+APV9YYTzrbsk
0tktPZhl0MKUXZ2TYe0SZwG89Q9oIG1+WeKnX4XtNh9Nn637c6+ClZYFthw91FG0WpcbRQlmIAiI
MPUrQFZE5Shmj7SwLVyjSgGZqOujjfzN2SDC/kxHETNgcaU2k8GApk4F++qLfpXNikvaHzbVcm5o
rgplwaJBo/S+QOQzvcXxxSSdfkAqDrI4DKGo3tstjbPyhboNIPpp9LN2wtZKWQXZihOIH0WfzxPU
wtxJyWPIFxIMTei+2lsKA72gGJcqFK9et8n9mtX5SPXYKEFUqp7TsHqdTKMf/iZ3ZxJTP7AdbYo8
rI5ZLyJtTrsTkPm6gN9FZV3dN0V4I1Vhrxg7lOxJmLmAkLQk7+xDCD0e/VlLV8RDEP5+gNEf70i/
r4kCenfHqysGtoRuFJF/MI/rKehK3dzTYNckqosf/shOLf5JGPD8RK9xIMFRA24/3kOxFAyzZANR
ykYU/Du6xv1qIaBGO0D5W+XmE4iQJXstr0zPqkRIkkoWJJeple3aL90yLW3LP+3d49hsrm1Wmbha
XwbhBu4A58L4SNYj94jz/cP/OIY9POGxCYAnknIdDtwpMcebExabaaZwoz9ibP4sMEgChyZn3K6V
bGQBUD4wnoQ1jrCk3a/zwOVzcm5Zq9fx6jTGlIUTxEBuw0ehuDtHx9z8n+42+G1NRUwbmkvKOk9C
8VjxQDs17k7vcZBYGseQ3vXQqh3Ryo/OO/hANk8SZVYgHtx/K2W3A90iTRvWsDHlrfl15RT0hjCI
hLAjYZHXuHqms/Hy576xQmwbvBs+lDVKbOgLBoJCRHnvZ47UZbQPP1XE3+jsnqRCxdmD2Jw/+O1E
3SAPrf9luWYAmxVM1USL67otrmHQ1sAvYmUDAi6k3ECXHTBN6HQQDyMkgj645Ctfi3gUVLxEdF57
4GxI4wgjNEtz1Qj1nAoBOBYkDapYWTGAnCYw/Ibib3KcoVZUvHscfVKuU5/Q3gYRucigMxr+HSFW
DqI5+Vfiy3BrH3XBmNfGwGFpnLYvvZME60sNkfcarcGCeGdGAAMdwd8KEqHfBh1PyTI9I51Kflja
MSxF9n7AfGAgnZ9pe7WkDsSqQz60x6wipEyw7LaYPnJ0n1p8MW91m4bNrciCGWwIPLGWPU60pqhy
5cAh2or+UfD0WkwLI+DXI3EHetWqE2wVfeNINk5KwkAg/px6BJW7biyXB61eTQ5OLQJByBmPMgIH
A3QTDMmN8zl3hBuByONeKqhOb3NRvUBMBE0E/+LMUiJ8onUH5KaQ6HuDKGq2grQ/gZMzjjZlyASe
xykYNPAvVoePmwqbtoilPmqgZ/i1Wo3v96/4kd5+6lWDslpHSxJ3V7dmcZ+IQhbrlHPnaa+2VsK3
1wF5qU7zWHsF0oXhIwp8CMh0B7IDkPnp0xJ1VhIIc1OWbHGejT3JdSMPlZijCB9UZypPzpssXD3j
FCYnK4/6wtNzdZJDgofjIbCVANUmzmG8DAnP/CL0jdiLurX9nP3ynRUPVQ+z4qKnugOCisY6BAsT
v3mafQo+tCz2gV7aTVVeY7EoaHrFC+imntO1p/FEgD41mGzNOHGj5U42y+JtzopgXZHXlZlB+RtQ
aUmfzp2HDevpbLUTC8TlrFp7YPEQ7a8ilGogFHur1yVdqQre89BN8VR28am3x1Uv2vdJNeObGmkP
0c3RUcB0zGSbl4qc3P4y3xpWQypitMFRsa5UXPeweJwhn+d3hIqYl3ymhARk8x72o8zDXQ/EEFYA
QV+B+sKZAmCvIThD7v7b0p7q32f+koFC75JNXaChmeDnX6Cj3xNGvuWpaVgVOOi5KNLo3VoHBEyF
8W5pXjAniXdlzTCsmL0rHr4cXKDiSZ42wY3MnvntnvXojSpBThMH9tH68Bp1of5xRx4XKgGmIixg
rmy9sAipD5DfDNCQEXmuBYVSHqbk2b7arAtGH4REkJPSJhplgrlZKhgRRdxT3qSbZBuy5RsqxeuX
aCcLivDBH/DD9rn7MUMJ0XE7nEEwxxL2F2ySxwA+1NQRcPVnucrv+MJxBjoIEkz1y/+TNpQ2ACCS
X+39Z1+ZDAZSV3PO4rTfq76xMCM87+e97fJk0jCCsM3p8JDvmAKQgctFF10VUPvJ1FP75Url4+ni
rKXnPYUKs8uqvU2VV9S9C2E/WvEuh66c/hP+Fo1zxzRF/kyXWmevWtJYlWA0t/rUwfxgSohykg3r
RcS2Wne1Ag2TGLYaOF8vVzw6RmSoEnGCwYJWiaSOHDCY6sGSLK0Qw3fu/zXhS/ERuzr1sdwh4cSM
7dPE24GO9w2biHRk/GhtmGnQijYjC03Fylq61M9KjVHZoMgembqbFx08iURJ88ZBQWf8yxXtsJeQ
4hmpEuYhcYNPV0PlN089aGmdtNteQsY6iwNpNwqc3tKa2XfrHLSO32tvYkkkwyT/MHTbvFlp6A/W
3MbdtOWZDbHoAojE1Ynh7fNWT+6HCBtJHuUgUPVfY8rPneYqR+HIDbpErOe9OJmIpTO+MpalhHMT
fg2whSR0u/i+MXHM0LvZD/OAziF02BSpNpfm8cjClsHK3I7lCBjfMZZfi5LxCftfJqzjqFM6MyLW
N6RTnZ4dNuCmjA0MHBfzgZ+y7yvElO0Zun9UZfcYJrL3ZrgjpVoACYue9kU3vGjIqH0wSI322e6U
n5xh1wjVYrYbd/YAXJvD+oP5qnlXc5IOWT3LuiomQ7hTwXkWUBr8SYr8PYdm6oqFxwjfWDzHh1N0
4IhsWGj/gSzMqmJwQYYomMHFR4poQHCBSSr+kNTdvXeq9igt7VlK3JwuTaqfak/xXXz+oRvPFujP
0gtRNFHhcICMozJRM0OP6v82slv3ca7YAB2On6qE2hWOiv46HIyc1AAeOMVQLT2HnR7pv9TGHmTn
zf8GFcTodi7aTlDEXEu9APoK4jEiGrD9bwxw12tusMx2Utd018qjxWuQxjxRyVg0CLXSlxp6/P6l
7K/L0ks/jZEc6lqSkKskh+iR1sJaOFTUV0c7skJCjrT+fWWdhDriVOzg++4Fgqx0akT2mi9z9IRA
CpTeUOK2MTKcktfIi3Me574qTrS382E3MrdrhuZedEfMkN2G9Uh9yTt6mJtPJNe1FgNR9tE6rz9A
s2WxBbLtvKg/HrRCTJCL/6lKb4Z6OtA1O1VBGz8Eq+sxi7txNivVdz2vch6lgSAk0abZ841wCfJN
+eYZrBn3dUyawC1SmWC6Mfeor/WQ2Q7y8Y+VsTn2kXMrSHcjXGxpjw0Y3+G8wRfaHytaSl40GtiV
GIHJqySKQqgQEEuRSeLkq34rwTexjUeRLT8MrJBBUE9BYv8J72ycSRNHY1zecU43aolhLlSYAYM3
PAC6wtoioeQQZj8z7EAxCOzR8sAlC/KSezZkwMDlRHtNPq9SAUmbNX57flrGYYSwZrj6VF6nWepr
Ar6Em36JtwtVl9EDCIE3q4SAzFGGCeWJGoEll2gBNEIs5IvK4fppxobCPSka8VRAPcMjNOz6bcGC
dp2/1XJpA3k0bvEua+ti3pKEYOuJn1UjbGL6J5eUrj011Da32s6iTBTYHo6rZ3YdUzp3hSPy7wT8
7CC0BaBPxn18qe8hL90Op8UvBEoSNj3BwnZ8f6wP9cXtXlw9ZOOHmU0qjRf29E6xNjEZ1TvuMzFy
3FmXYDHV0KEApjpUzK8tHGNkTPeHhCyKPrheWmn5bVNepvYRac5HPZsq91n+mE3mSUwc3nz4PFTY
tjSsRi74t0L2FhEThsL0t+Fd9fYDUg8kQLHMQQxCrK97cPHs7W73JcrwZLNMIqB7Ij7gMXZoGl+4
YPbOkKDGrr7WvOLi2ulfSwTkBJs+cxhKTDr3hPXEov/l0C2xYMnRUMhD0+b1L40U460tVoqYJbBQ
d/dmKlDEaZ3DKwTKGLCt3jwd4vNgm4wfGh11aHRtPhUsAqhC8P/xmKgSCUHnc7QaCXGWBTk2Zrgl
vBucSVP/59ZHww30fu5u2UBBgvqQQvkkgskb3tY+O1Uisxlg9iBWFBtgMhCh4IZdeCb+QTpETPdn
7AHgkpvJzVqxpP8/08UTVQFKkr34q0vy58d13CajdRLLxxvOZxz1IQIqNhHAZHNmGHa0rWoa7fvb
YHR3CgqnQSqylEJZ5vm61rgwi5gKVCBNj3qUsQlHyStdIQ3EHXBExo9ftIoYEs/QslTnnq6+Nitw
A7mngKpH67/TfZCEloSmssACih6ejqbUJh8QyQFfSG7Hvv0mUIUdeE6va8mO2VZ+b5tH7BMBR07Z
BF/zoNZovwEokJuOzNoBD9JDf14xInRbdfaMkhPSms8MUaNu7ig99LxWajXwwzRxrJMOicpGcmoE
99M1Odon7+mUl9c0A4D48EEtUSoBuLSvtY6hEURNr4oVSHKV03Sn7svZzQGGTpVa97gRhNK8KC5s
koSqjEV4wvvQeqPszu6aohLKUy7fRv+KQc/LkChYLK0v6P9cTIHjOVLxzI2g9ypRb4FXNpwZFNS2
K0sSfKti2Wx7MJfeUZMKz7IZC1nGfK0DUKtxA3OmyQRSzCWuXwoDK1T8Uxe319ZokZ3+Pjw7SxjC
v3rMTL95Q87aHFKsW4F+5TA2HRrf27/nK8rSj/A6pCE8CXHBbMHEhgE1mujPhJXoxWeazvd2HLZ3
F6B1GiJP5cx2tD4IGtmx6BC3YNjs4dMT1yf7pH4jgYCBpGkRQqa+hcgfbe02s08Vh7YLZ/dBzsec
n2BpQOfH9Q7LdDGkZxglnK0g5TmaDUPLWJXu24q225/VtbVb0ho1yY02sMIfDmMlm+c71QAqcO7L
OvzJvPle5dtTEQFJmqh3PJ8vQ8ASoVf/82npPpSHarecFqcsU5JI4R7bWTKeY5uAMr5RrYmrZYY1
LsimS5RtwouD48TBhmbo5badcl06vgA3yU41iFx8uKJtxedZ80AK9yXthNt0d7BzNFx+UDSHheLz
PLwjsZX4cBfF1FboWkANXpC8mWR7bj2ANJZzI5pu/xFmItx6vIN3RGEqy/iJd1WPuvqHjTjIE1qV
qdPAzPgdtmmkhkqHo8iVxUyHcMdFsLeoUNy/z2Y1gEnjfRLGF/jxdmjJ5UpxIK56q2bGM10hflHN
2XQhIZ9gykcFeEuZv55NMviUhmpcnQ16AJzVPxj5dcvXkAyh9OPrIAwwLlcWT10KOViIKxIBy30/
2JgDcV1d+O+dYdOhKZqfXFtwU+XO83MK7S9suGzoZBcAeKWamNKNTPARZJiGHyqY62RVRnIjOdjV
/e41iKudUZtDgEDCcBmQUrZYjfkmyfigFgkGbJeLtEVkjKrpy3GIGXKv2OQLlRMMnbEMse2enn0Z
vWAn7nxS+A8dAtfT3edSGM658eAWDu51q3XrYLW8cviXjOyw1+skCReWrLyWdSAJ6iMHK6qKEJ9P
tFbrRjc7Vr1qSDGig1iYLg5sXKLsIEUZsxjfXG1VQyPe+/9/svgZ9G7UfnjVnuPtODfQDsWDVp6c
8wBq9FR6MvINk3GToo/qMijYb/ZsQlXKOUEfk3hi9aKJDCcu4L/R9V1cGb/FmFDEsS/ob2R+pazo
gLuVGPvCwZdcTbOj5xaf6VPhBwM78J7OH1ZNwXDfgthccscWjU3KR1qHMivog8ieuh6Q9wopYUEE
KXIxRQ5uCWdBVp09sfsesVY4Rh9fLNIx6M3sehGLEwL97anHQjIgjPz+DUhz75VjBk7poOJv3h7K
gdFqpKDl2KTdRvUyM1UAnkOeq7DD1yt9HjIKBtlaGS07dRFCS/lQ70BfHeGgaKIMAFxckXcfXx1J
+/E7nq2aO4YcdvczMql00gznpJN5hre6oXgB5H44xkRktgUn7EqIOqSDa3uJpDrErD96/9JHCjKO
3MbbuldBmPbwlPH/ljOQICHAXsDY9Epag0AOHH2iDMn7a88d404aNtig76t++JKEVum76p38E7+N
Kp/gWVSt6iYmxzsLyArnwgmx+xCdTqrP/j6vZOb5jkwlHQx8ocXfpCyZWMyzaTh0S9pm+tadvFL1
rXd25P2Nrhp3k2mmQeQbvGJDg1wzuEgrB3xRkiB8mh+K09IB8UevzKpBkID+q0nNEofKfPF17UIw
O/C+8LI8A3c9A+f0t+fwiSL0rd9s6XnUZ7zlq4Hu5X9xLJ/lnXtq9Mve891o/KSGUYkE8lkABXFu
JwYxQkbdU4P4maRN0xHDLonjujgNwn5e8Kc4C7eTxO1olMQ9/g9WEFlnl2qV9BCulpeZPXPlsu54
rx/qShbEHylUr4rTxTkJ+61CB6GZGy3sT3+pSw45bMvvqtJWoWp0THdHyzvDiZGCppwwapK1imtw
b62AKTNay/NwCRuQEvyhpnHXEWzPklNN757+/putPNitmCZmNs7vyUDTbwcPMFgklJsB5WpvNEgj
BpvMINRt4H2d229K0cZvTDi4P4K8djZ06drozYXk0aSuSuYk8oR2hhl/CxaytyedF5C8pdERAQ25
Yum7LmyxRXAPysv8SKsYTszaMZB7ZOKsCgAM5SRHleKqsSqu3edo8qSQ2/PfO2si/8VG3ibV350H
mG6g7XRDnLEN+nt44R/I7G8DIiInpY8ce8oiI11LJGg/WPv2M1ES81USGodhSwjFNaW9a/j3B1aH
Erjt2IAckGIMEayDApPKVmPOz4EeWNn1Pm7z5Gtq/OjnWOPc7rq1DZlo2aLEel4S+flrl3RSPow3
WVbpL4clqTbniYk9xzLnfZDGwnIfC1D2luxUUT1up4UOc7YNuKdIXfP1v+SEJgOGNmWr4noQbXNP
F/w+6eZtR+2bBf1qPVQvb84tJl1o0gCaRFnK9SlISL+HrwfztDXsSAJF+l0d8+yD2EN9gQhxqsac
TuE7nrKijQOOPiocI7tAsdyUEOglt2xlMXNh1k7i+ViSfb6V6ha95jIudJbxIfv7pHqCVf/LjQsa
hjWMRHKKh1JI2ZaolNW21YAYSsU+SYYlOsyZ1JvLES3VCqvpPzE/tnKnmCnMDdigzJOTVoM5eMRc
ENjrKh08EyVZQxLglbEjlsQN6Wqd02B0twWhUhKf3/Fe5l5u3UuvoLenS+0EXF68iZS+TVIeEJ6O
K/iiRprEgqGM1EfdW0S0dJp2nXchH8PLAvzvN8C2PTKoSesOG+HFT7Pf08JM6/4EJWBfwODl+O7+
/evwHqcWdKsWRMETL4fVXg0Ik2+h8ZczqcmdNSgqw/qqsOLD6/RXWZrwmXvyQ7sapX3pevNnDhXG
vO6ZWsCML2w2MropG3re5IiF7WsQ686OGYUh+8pwyN2Xqv/RCfmR9ZMTdmKpBTocoLGetR0+1lvO
nYEWPB6gu4+Z3sFCI/qSxsZ9xY2juU99XApw0uKHcjb9NU9lvdelg9a3tVo7QnnMN6k+X9PhPym9
KzblzXcxPiEabYfCEDZ8tYJBKOpAfm0yxlCRX1XeRFWYvHZw5Z5HQhgeVpi4OCQGDO795YhbzBef
Ve665QrtfoYWZ+SCwDdCflRaFKjuEiBezHCZ0YnTYTayfS2Aa4XUeXs1Z///o0wVGvM/7NEH3aCF
EyV+A9OzAU5CdDq0A6U5bKe2j5jWk1iSXI6fRt77QxyqkFgZLt0z93q1GTE4ASsicsS8v3JBTwDs
+NNtokXGlcG0DqqpJYL+TnCkoA15mLYC3h8PF7ERc99QsepN7RDGtlVFtD6/Nbcp4TINTE2ZvLdE
kACAAeZEm2zzaylWMXebJL+MVEcwnZSlSUynYCYrEWHf1MIhrT/o8dBr0VSx38ivRGpK+jBrvbzY
ZqLj84n4ZIbj9mOe1J2SNnKZHZ8TQ2Bgd/AhplPUmnE5pRyyc1Au6GYWDttkqN14LPsVBmXGRnWf
2wKqQ/zeys7XtIBn3nQQaVP1DqI5SEeeQbjHye82HVfXKXpA2okRGW1zxLerbuGuzmWVYWZcrVcj
BJsloIZjkjzJrZzJKX8hWLXNYisbujy5ourrCy6Zy8gLk6dV1Kz8/99s01WRijrdWHHZ6Dxr/jFR
3p27ibDkbjvMGiqNjq7UPbcPW7pwr5st6097saEl3MzENPDEXt+CZWGMnqVLUOQW2vtqKPnvu3BB
iyNjXZikSVvwLadjPOYFYcW2a9+RLHbEXY4R0qgOWKml41PRM0n9L8sR+qgjKxIq39KsnPEzSefE
nB9PKYYJUf8ajX1DFy/wcghedrKLYMOIleiWl5yRUwkaPviQHutNAf78t1bEshqK1flIkrhICvuH
vp2RjnhPDs9w/oUdbJtYy/4+Jlm9I9aBZnNy6KsWGQMHHQi8G6yaTKfUwpZMxI57N4itpU6tBjlQ
sjb+3uRfvkgsvbOdcGYqo5kZ7jagXeQf6CU8vWeZuWXqbHJto8redLZfFxld2u4syGc/RIZYUSoY
L3MKXIXYKgAtiT8wCLNXoI/HLeoGBUKvMZ40XCb0k3dUxzhTviJYeux28pa6jhhepzsb8I/zl51w
QGvOYSw1D0ub0jSyIVKajvBMF1VGNiJb6lGa8+ZsZiaWJiygyBt49Z54IKqmR76LIZ36T3JwKqoD
ys0mKIkbsU8OmK+qRL6q7kMlrNrBtCL5PQZD6adK8JIdyOGmUqz9mW3n83TqP62BhXxfmyu4uuXZ
PjHdHWVIEja2EgdaouzHlMiXhAz/qeGfyBbfnz0SbMF/lTVG1XeIJMYk8mH+pD872MdO/b+MPWKE
CHTmHiDtBpjlGBoG5Mb5eaqnMkWYJTRTt2hECZUj/wL9t04lmgjE9+fDSeUbtKXtJnDjZA1Y35Yn
02II3Eipq9YQ8GunRfdHei1F0mRqEJkbqLEusyxGA0ubGbCLkwBBpYr+QdBlQwR6UrDyxhB23o4X
PvjrtEdKPG4xWMOmYwRV2yHSSrmqZ9iYkyW9SQNoyFJb+JY7vVE7llAZOKusn5vVGXUkGAxcw3e2
X58W+wgeME/RktVz9aRM7aomVvEPQPJ2X3DyCxM9j/xB05NIou+hug4hlThbONh0UCFpzuCeHyl/
yql4PhrHlx8spBCPe8CQXCH400Ui/i22bxLE3Zrf4chz1QdQcXM3d4h6EZ0HG5bn0pfVlLrUPPlO
NMvtHcpmXRFoBU06zfXaKdla3Wq+vD/8bvIKIcfIySfN3Z1WEQx+UeQzCJnOo/V9VpcMAJJZ/Cpf
5AJ4bIP0NSGNB475rTIWxVAU3oTeVt0eo2eRK5ozfkSRHoou3t65Yj2Sa75LX6NztJ/E6oV8x/mp
R4T7KNA4Cr8UZdRVG5rmkUbgAccl9hgRg43SGQ8HX9x+q2SfzlYu0DCtRR7DgpdkDbY8R7uTD2i5
pEdCrfQ9ulObtCxKZpqVn6+oCH1DrlkT6cn/Y9Btk8/8F2CZsgnn15GtmoJTy0n5A0kaZAEc48ES
dMRZlrQCTtfEuwnbPO2Z42TlEl/0mLidOq6v2ZVOZU+i5/+DJk/Naltt7k4F+//dhiqR8271AXXV
mEJXf9tTs3aLhqpEm22B2WWMGOrhpAKdestBKifEJmtpUwolSgOGD/Ipjz+/lT29YE7ii5pusRt0
ulZZCbzw0cX0uvEbM4LxLM6j7R73AzBHvUNP2CVgifoaS87QKFuugYsD05kZE3LBFkf1Y+l1J+yC
2axdi3kl2Wb0QHhn4j2MROmG0xhQG88sO4/5wyFjNN84tUUMiOe64nA4xHsRGsT7Pg10bqyhWW3I
lesm0xrf0Yw3ML3CUx2FiWMYqWo/YmlmQsUrJXbz4fD52YpM1i9duf308T5tY6d3/pjBm9WPBLCI
DUySEdk1J4hQplwTdJETTWSI68NKymbM+7y/2sdqwD3TZz3REasX7RbWj7cNyqIRgUgP1a2osonZ
pvvoXMWt1jDy7M3JxOIPfXGJG3/E9ILwbQild9lrNGZy5qlKuNf9v1/LU8vAZPwqTVSY+8YSJDrw
3mMLeZVRJQH29JrZr2ET683rnICMyZBCqwXCEZSmiC5b0z8K8bv1iDcEfBNww0unqQkoR6dExvET
DsoD2Xd+ekXU3Y/Fb4KCCYT4jxbLCNAAhXJnHCMmurZutLN0YlgoV2Ec74iu0nZ+cGVsn/qz570q
Kh5i5gCDI/9g+c4aS2yjn+HI6PkM38cgNuyhHv447NM6N72U8V/jTdroiMmLgb1/ACtho4o0R0Y4
QZ1K31XOjlj2Qq1vae3++/KdLYwy24tOs/nZPmOn3Jj5i4Qw5tjVBT2+ni/m7VgGToOhA/TbNvqI
EaSSmt6Ewo6q5rW280MpJfgRKAeTy4P/k46G1VLoWA35pbdWO09HZf4MwJyM/Hdx7iqfP0SOLNLY
Ach2u/R4osoHOqZmAQb3ibmNLk33RNUrxlrUcNWUGLuCybcfwK/EG+RXkw2wff3cH488DRhBvUl6
5PIJBMj3nDkcjhPiLQW6HG5HM1Rg3gDwaV9rNG01t359x1uW+XsLx1CYqGm1bFdLPXo9jf0JzehG
3GXSH/aisf+cMaLnfkbRn2Ga9Agl8Sm7jpIZB46wQxAo3NIu9/68fWHpeUkLcJThj1Oy0mTbxI/+
qApTCQAkiemeihDICvWYReOx9eXb2gKQ/PyRF7Jzcp0I4Bz7tePS6SLIiIGqTZBN5lDt4ou7xJsK
ijIHH83Ei2Lcxmzig8e9WgqH5UrzhlGHViu/5WZeM7xhGkHijBb37TR7PX04RSS1yAHpKuIAkhyo
UR3oH6krkLyPF/s8hnBkizkcjI0ZqnPxJ2zFlvCCTqbqLuQy68ZOEF5C4Z5VsFniT/gHXaOOjDP7
0m+paFLvCOuttgugeiJYOwzDCH/HDAlrZq/jkbtjtzRWmF96nVMNvfOAhSdL+HpUqINetVBRof3t
YpnBvmnAFwhx97kZSrCdbqxk5I4m4Lt1nt8oc8SwVDOsTtLF4VShoCnX2pPbhxbQpCouybpasSpZ
HN9Pu3ILWAhmyUg7jVXE9Vds93Pu765aKjgtl/xHOKBoqojZH167/UiuKPsWiAFoZn+gL+OUw8RL
tjOGdzUIzQkRqqYOGFAQAZrCZJlkaDV/Z+IDy3UkeXxWIoz9SwLhCuQZEiiNAvf8u57jkE2ipts3
wwal/ebjpoMF2PUWN/NY+UgiWITtQObCnanmwmVXkLVd0FnGAohym3Mtn/u2IILn4reEPjpUOyvp
fVFshGI4tle/FDPRWxGKCNTFLqFOi6SmjJ0B3NljUcUrkJEXJAbYYPap78JBRmSSYeJS2QWOvtSP
9AbSYHQBAg3iAuFXCQ6FxowZla9/SUEZXsW3FWQl3vyfyL/0jRhIlkrpFbxTnpIZzqnFW3nhvu3q
H4zfE+zev/VpfBsoA+t5EGmzYlAwIbsVUhKwuQ6AtTVLvYp8im4gFhec1G4rxsJcU8tgu9a7tsbu
x1S3YZDfONLdagYGCFO5TuW8C7ipBV94wnBF4aE0TXOzvDZKE0585U5uQOdXKmjSW7CqHcf7JwU2
pF2AFdVCTVk9mlA9DMXlcGovuZO9LOmrnj20ObtCARjxTmvkpCNyEtNuUAZvLZfWY6VrI+vikNxm
aX9QHyVKStIx5PlHhII/m0cY1Y7/w3KHN7lMLbyhaJocbmUIkQE/lbsLP3S6EuZICr+tYGfvROhs
jS6zOf+TobVqeu1z391AkGEoKvl7qvHxVwpIZH5ldpR6weROIEer+AlvaDCdPE2RAErlv8RvhTM0
o8XZLDzUSqERKeKkMgqsVM6TJwBCw3+SrTREVJX04dHQBKyoUX3dLNjMzpGnopqZArGsp8hYC38G
mEiYgrD2dotNcwUs+xik6Uwh6nS9Y6J6esTbC5z6p4PKfOaARgFj5Ge32vwQ+8L2Lpf7WA11YXqs
G7eNkcP6YlmTPhXQ8zaTVekZeBhUJI7icIvR7mWRBQjsR1hl1vRtRV2l5RUZ4hfq8ZXc3Twj0bdb
kNnpZ+NvrYwAaBujEF79iRc4YxiTgrD8nYzdvAZrMzxo2v/XhJEJhJr8othWT85M2kXd+zqmcdyN
9dsYauw3X7guqJzP61+BfYOQhhaiXACRVItksTq3wYb0EBC3ubMIVd2AQ9F/OJ5a6JQh3/UJD03G
aNPFl8I7qW4kCl8Fz4W0kLe5Sv2uNLx/ofTS9XAW+T3Jx7BMVJdTRH4vEVynmcNrNm8YQv5cshoE
bOAhDLHpIU3x3UH+xcI5jH/+S90Y2h6Kjpd0TE3xuCXH8llN8TnQySlA2NItsHzTQC52chq6hXjh
noU0PnM2aWnjJFITK9gv0Kb+ZwynL4AMbcc74s8LZDimmUZuF+KApP4bg9I4Vucj1p8OmsgptGXx
q3/DBIlYaiZ5h/OhadyNDZFxYdINZ/zz8Pph94j5mytvPJPJ2iZTcm6btiKB7b7SSC3sWskLMVNM
iv/ns6ctQ+e/JSaWecNqhyU5Qmn4KQ73D11HbAPQC+M2QRx4G0MYlo7kYT0JgEJdo06r+sFs47y6
2n1AC8QlXle2KSVr4ZjClHoVm1ldjLhN5IFLrnz1yzbE1Fy/X9xfP3vDHYBa7hg9w+bsMnz2dEbA
VbYrfmwj9JBFubbpj5A/RnpMm3zom5LZVTYt2R+SJCRfpruf7b21VnQn0omneXhWId1e+bs9hFvv
JNO5++P+a/FgYRTJ9Pf56nTRYr0m8mOm+JBsJPOM6UgVwzmRNfbhi9sv8Aie/NEt90QevhbAMv+n
2O2gjlQOxvbphHCbNQvtKrM8cplxfbL0k+/gaqto4fc1cGUdwaflTpazCTDdUU42tE8Qc9TVe6Ei
B/D9C9bEmi+fnNkexJ0bprGMuU040AwlAxsCw5Q/dOQRSvLzILO1EEqKCRiGCywZpQhkmIUMuPyP
/S79TiuQ5lax8SU7GaRH4GZQwutVI3coEU56roOnR/SNN3xYKWA9WH3IaaY42ivS2502uMtieTaL
ovJ1cBZvIBAonMruV0MtIAz0+mtRXON3e7dQETV2W7at8KXyp1yczoGMJDttL2Q5dtuKisD+JTQc
yR4jeYLEwL4E7lIZOkGuW9+TSK11GaAsy2WEMvk51qWod1VbiqbOQs/4FBUgBd7WtfpcWrlnweTj
nZnncF3mcjT9ylL0ouAFoVCalIcYpB2DnnqTLDcmNPMqJgtGuLlBRkWdgiHROVKSnGewfWBtVg05
W5wZW/FvazJO62+jnihYkqWwoeqM9jlIAZfxf+JfYp264EOa+k6zCXTFikjmL7oBtKcCGT1lCJSe
2ACeFWgRFYZ5iQViQdTjSi/1+B0m8yf4mGevWwADCsTJbGc4tBTo63otZkVZVW4b3t8Zwwh2wE5V
Kah5D3979jAqaCJUkxzNpIsC9RYzrKQaql4ec/c1yjCRcW01IMIfR+vF2fOxSGgSEr2Jss2EQvQ1
k/uyDq5Q+NTPC3yAR1qOQ1A83rdeJMAvbtPPh/cN73/mAGnUNtKMfE6epPkaPmslhEkHzyWobMdw
1+rNbSy/AKkGkQJ7JjIYzXuehVK99YU6Yidb8W5jLBVNqQFFgwVNpPxNbN11tAqsQlakVFn0gG6x
HQGO8IKQQg5smk64lYJ2kfnsWEhMfDsHpFGM/6uhMJjOQkvRYBbvnTk3hW17W3n/h9eJwEqP9A4h
y3JMfN4xiOLZ2M6ymCewRpOSa0wN5ebJGY6wZ/CgjC92gmW5caD+8vIrqB5KIv2Tq/kIicapSE/X
jFp+aA7kDp8BzJoKxi+6p8kiAPcIhJMbX/MzGX56ZwPKlrq26LrFNIVgkUZGH6nyWBuNmZWRu1XT
m7UOJHFojbouoPZgr22g4e/QtilNPdNIeVCN95axLrJlpzgvtCLCwHU3jVjhy3Fc7reTUgP+aZrF
cPBYQ6T/51KkuZFmXzysIOOXUYYlo8KNHaNGLaC7FG69f9LxX210/8BdAgcPur+1hhTPn+p+5PdX
m70IRCun1eNZkIlY2nd3Ph1/fPWkvFHKFUPBUH3UjywtJ0D2LV1hmQgzyFMe1apJ9io+LX8sgflP
qJMtbRa7AVrMdHRPWZevT5outLHffbbcMdY5JrC2bw47lfqsCyoCWIFJk0iBIiV0/gOmfbxMPYdD
9WB5ELDylCOOi8oRVg1mzcYx1mP49cGsXMRFq/oFnzrqt07T9UYSplDY4SJUiyJzuvgmhA0kMu2P
pctnvsyFdpgnCtKCo86I3rnze1C0fQTwblfJKTHsAdRlQQr9+YaXx0uqJU0FywafhIMjuyeGeank
h0O5Aur7xsQ3f6jmkiwt+enrmLPhHZQubRRehhl4/CZU6cBIqb2QG3XJc2d0cEs/V1nteAKUzIkT
YTVpBp6t4exlSMkLI1TDRyIoPFVUYXCR38xuTB6K+2WGrRmKzPTywW0IlrBH7T+ndBRlnuQOX/po
3q5B4Pujc6LeCl/iaOhfy24JDhebacztJ1Dp/cn1eMdjiAZJcktH4GaXbuMRDe+UK6rLxs9G2Ozn
jxoVTKxPGCQjUCrUi1uah9Yjgskmeu+iC76WoJdGkWwejavY9bV8haQCSyQ8EHcNeJuALws/aPrL
isV8IeOOjJUaw3OD1sUMaUl3VnKIeX28fXgqysk5D+HcLK+m6mjuPtfkXrTn60vF7dihCDfm10sv
3t8ApMpW50J0h1a4XtUJqRPtagFAgw6E+pl46z0nuUkc1mK51gJMJiHT+h8oJTK6OIaIClOcePLf
MWPZiiXwzqSXpKY4LyRc8JfahQWGJLQCQT/UxOZfs9/n//8a2UzFQtXV6TrQ3jUqa9IkyI7vDa0e
EEPm14x0Th74BtXUpLguBo+RCUqdDU/Uo+Q7Ks8EnKJ3H0roG3kyjSr+LEtDMag8+o96VCXP10Sp
X7h6nLWnWGpTJjOlWex/D8aSNg1tT4QDA7o1KeU7YHDJXKU9x8okSKbcAhwEfAZzbUm+wMtcfU8j
u8Xn8zL5XUJ3Ln4SrhQu6LL40hrqqXx/huCHuZHzxAZqKNpBL1CdOO+4TzzbTsBLG+PXf71voSoM
QCux0Ogk5ngdSGamCIqQlZMjw9vlCgsLDnfPH8gnw+RujIO7C72PLLdBlV3eWH+qzhoBl8cl9pXU
upkgSInWsWg8Qh9/xjVtWe4bWuagTRhZf0I5olc0hImy/pJbzLNvTC9QiGMXsZimZnCExfg4B2zp
U/vWGa4+DSAurcE1D5nlUOUijPzIgR6K3Zz3i6fkx5ZlfXwAv+Q9066jiowYPY7EPQLmJcllHnmD
+ZV7gbI4gIF3eTzjByL7udakWogGgUkWhutWNRtAKr0kk24feLCCUGkfAsf6Xqu/cdNXGvLL3wsp
u2ORkIBnLpA7324pth7d+JxI4hBYIDA6iIrKTb/UUKTxbPr+Yb3ufmoCNDs5T7eWiBkeMI/q1v//
K9X9rfG33LB0KP1Am5KUnN4x9f/zyJeBPR9J6UkCKRnTAs7OOMBOm3L0tRTt14k2QSpgu0McYcaT
5A+PmEydRKpC332BpGpYGHL2wAcRQVBGztZ3SgL3HJoV6tP2LT83UgxgbtIH6fLPruVx/rbdS8Hp
bTD0aVpIXspmiY6XMWHVbGisGoCXjxH0QYcrTw9s7kmPQXuiBdHP+UF3kqvpJCD+1VAUnOGVz6nu
NOwyxcShooxFr1sWWfInlN5Naed3TlIQoM44o7lUBydvR3Nu/ecWc2TsN5Bqhyi5uBhQ43yeNabH
0fWa+TnrUq+oHWvLP1dP4rwvXlogIq2PhLjcwsPPZf/SzHO3ydDGh1O9OdWnZvRa6gMg6TR0LjX6
TyxUAdo0EUod5QaxyhFYMol/xQPV8yhrST4wa3PMhS+mOrn97GbC7FTv/c9uW6l+Jixv71CdfNEJ
2rnXDtk3PaDhA0PS4ByljmzM+VLzqJPGLZVPjPQTzq/Fqq+JbiilgR8fZl2BDIpMRhchEl2kqiSN
RGeF/OVSPfQ48ejZ1/gZMLXwGSHHpWgSBwq81HoDtUPTJ5l0jv0XRfhPCMCBOVwuGg1AUiHiQggx
RibTbgTMFuQg55PN1CkkSjwx8quLy1aRr43ZdE2inyTr8bqewowS3rm8+4GjWdXtZiLGEW7OHOt7
w6xZItyoT7IqIFxORkzqtLZVnBeaB2U3ENf6JQkWfRAQJMrJErND1JaYCaEzh+qPOBpaiH/s6Bcx
fipsuI+ADoEjur7msAxOl7zDtAm1+8NCujm7ETlnaWpAjwZMntb5z4CSIytaS8h1O/5A4f41w69N
z/E/xIikcE6Ot/Opwf6aOOCtMKtvnsjMj6crXs63sZzosjn8LMUhFk/TJ01JmKqa/hhHTbfLaNwl
rP8Js4J4/n0cbQh3FtmKjHwMXJs34IUeJp+1rmQemrB0mF/L0MrGkbG8VjtSoxo2Pq7OzuVaRVzN
wAUXqgUV4ULjgm28m/N1ornaUGuqz8zggz6QR4gOKvNm+J+29XVfwKHZSbnfebVntxyeHCIIJ4en
9RcPbuc9YMwA57hHtncdO5dibd9tBuhs6PBQcPpcFgR9oSnX+8I03x3fAyFQTcIpfiPRbPw5phqs
XAud4Ni5+PTQVqHgVILEheLDiMb9uEYbLIvjjxIRCS+DxWr2i5oQBveOtIRug1xUDjLDXCVsBYJb
FSmYeumR/lag10dwSMHlGyYK5c4MifnloqjKqWTr+sFJGvw6qnyU8yamj2hWf5zMCNvM+ksOKeGn
DXa9UsH9mBw4IF0WrenemuzjQemfbTG3BJ+jyJRNDkBJb5sP6tqi/DloBou/KqhxwB7GU/MVIGbQ
x1p5+OFfjqilaa9PN+I35wmddUAd2/PEfweZzUdw+GI/OEbVU04inOwr4vGH79QfKhlqHh1gO+mJ
rV9ukd48fMgHuvmQmPCKwTdbX+OC3eYxZ/voGeZ+ldGxFbI7lyDRhJOPW/RKl+EdZ9N3Q6B3XVcu
Fmknt6BWgchUrtoXaO+XsZjdoA4viOVxXRdYqX1dFuhBHDCf/4RjvrELe5f4qctBHOcskJugHxYk
N7iLc9hR/KY7hnHxIirtl68wUyWJ/4U+OIS6I17hPcMDtHVCKpcRsalsDs1AFvBfqxUe3IuEJtD2
t/w8KFCGedeTlQhQU9wDW5fXIlIE10GX4AVzYuBs0Wz8WT5B5NHhKCRkJ/W5F+VnHLKv6KfUsV0+
FvoCfari89bgGgrpYog/A7+Pdg3nK8r9e4PPCPloXe8n7/gYmbhBI0T4/kzsh9gzhVh5hyEvmaHT
cHepDNlXaOXSGOVZWCyiVPA10trvNSR4C/7yXjuwvIXKCFQkpwyDykbozQnZz8UrbhOq8Zi/b0St
Vg2Y9MuGKuX3GF99K0tFRLw1LKIMBtTXn3bo2F1rSLak365IvWhIDYfc8XuEOgN6fnOgwxF0eSB2
RHzpJgR83Wlj1wP1/erAEhzq65JiH9M1dT0iP6zPfpg+KzpHvx5GMsB58ALLjj1R3OJQP8p/cStG
5V5iJN1TJZ0mHyke3lWMAt0zm668sOgUO9AvA7JKcr6OzwDj2i2hxI6nMiYdpXE038GrPzYgP6Fi
3Q1CgrtvADyFh8JjeCVhJCzPNcRovyyAdiMqPbDDXDkxTfzeanr9EIYaeDr4HOBtWdt7zxaQ/xTR
BNAxvr7Yb46uS1Y3WH2B9fpaLMVHalDwYNh0/EcVEIAw/sFD6jUBrrSMA3XAjLNALNmWomt2i0F8
SiY0Ia6uz4uAv4kT7IQMcxyURtK3N0561amtCv5m/xuEVU7NqoJjGFU45v4DtmlagnCPkin+UdrE
6dOzvH0WOBEdzlgtCHn7OHBCBVOpVZPSNMyHFoNRFjXd8HfOOhkGkJUPN+3cizGyTpV9lw/Z9C9r
IDdjqHHsiruk7fI4jPftZE3FSSgFGImjT9vcrnHc5lkroNOY83Tovm+msHe4WcYjffBPbX1SLw0a
khufnZ7aUbSufIDliBYsO93is4QsGy6esUFxodbgtove1wdki9On12jP4RN5pyeYjY595/eiqrD7
yNKalE2OeamdGfUzSzf1DBnA3FywRRTqFGp+eQiBN6fzr0bgNX8mnEDCropHqTSqw1SVZusH7YMU
k4c1REGgn5xoD5f7EawbZwQ6w0xrMoSGh1yiH3PI6eHV/oe4Ei0NQLq6y47z5ZXeQsJJ9jNciB+C
4bbzHuSMV7B1kek7+tYNvMag58eaZZTae+L0l9BznXj6RboSviRd8UikJOHOojIlvoLSQl8f1S1h
CXTVEuzCwQ8u5elWyOh2BkWlML5w6QkI6kakG7WipqdgCKgG5HnP3GOiUBIp1MVse8nZPacRwply
Gm5LJh5Bh8OqvQFPIlM4kofuvRW7sfZSCA3NtUr0rUkqlUeoIIRcZcoSn53HJN7r3/coUdnjWmOO
ysKcDn1vkG6qTVLLeg8xTjwu5Qkh3SDV+1G2aVk7e+gu3aPnJB/VuLhHSEN/z9fFrnbFmTwuRDPo
+ii0DlKXAhW86G4rYx6nwqHK8gH8Q6h/YBD1B4ek7r8nnrrM6ofPT3dumU1l7x79r5cYV6m/yNTB
emisUOegTkMUcFawUjC70IyvzmleVh66Z9Cyx+YvGyU495pUhNWJLkHm1ys4abfgAyD40nP9tyjb
x2vYWcVB4DfUCTpbWfb1Zm+vq6DfFLa5+NAtDkXq+UtmangW3TplU02xGEq2205p5pJkFjTDbVOJ
4Lin4UEMh1OOYmxu1m7gO3+CdzECgd2SQ6XovryNaHO4h1y/sD7zjc4v9hOoNkBkptameMyyeDF0
g0wayhMGkRNgDpgc30N7nq/hm0XfyjZPFT5w+KaK3mqv5JBSTBpk5kF3Nd7y/49eS7UFfJvzQRlC
7+C+nJAUR72vYkDNAOY/mzXeDllvFU/I2Ky+AH5/79oz05enHGzVWKgpYjhnWOB16mWhcKFWDEfh
Vw7LU53g7UXds+DM6mqnPPL+xWuT9L2Nc8dL+al6l/iNmJFkzovabChedpovAUKhTwP0bq9oISOz
uiKoBAQD9O5dPg6ac40iZK6xDAlzcTRjRJxjp9Ab1u1H4myIGcR0HzUXZoDJ7Jqom1l14B2XH0At
Z5JZ8T/+FD8wRaMInpSGoUQtl22U9zEzUt/XggyFyKHEl6OYrPNf17cKbz2O+roy3Zsb1S+is7dR
5+KRSrG04H5ps40tOco50SGuyG1GcDtfbaFD5iAvrgAFEQ5/KwKwRKRcvJq2b1NKGDNcKso4zjxg
vguEEhkwt7REYDgNIPqTjN1ShOY6EDfebBRNJ19giWtq35ejBD9HJz/nSIFv7acv2ayJUcnFUO/f
ustibTv4kab62eidw2NTu6VdTkXfQPTqQxl1wdaQQovSV82HERRw+45rCGpljefOrqokFHFAVIii
/QQlpsW5cn4nfATGgfJT0aaH05+fA9Ty6oUnbOhYT2xNUePp1x1vNACmr5WKSJ7Y6PcWGY7ueRiH
vWUWnm5Oc/t48PDPKvpWw5Hq7rHEQfIIGOoF80fabrkrpJOg637O+o5nT727yi4KlQRzsHPZWmJh
+59WGB8bUtmgFt25rkfmcOUr11GPyZHJV2ojtuK7jSpQEf9q+tpFM3jn7vaSk+ua0Idf8KLS3mn3
cM8twZm6ViBrwaSHtp5MemkH9gWN8OJFiTrW/+yaN8Q4TVm+osLl+tMM+jCGP8kvUlZcS7tDDZb0
w2YkIHS+NVVlnMNgjpKjql8OLgU0cuHqPcTp413LD9LUfh3L/gOunEx/Lq/NCG9WtzTnVTBhk7of
iO/w+fCCPciOpyW/pI0Vh2DBDCeje5s8vIKYhcpNdjwSFxm8m/mbH8qrQ7envB26ZxrrJx61rWdv
eRBqsFSBpy547ehqys6uHsPe2yCvhTcTTD6IilmEGwP9X+Dde8Gu9/bXmYcedw/e+U932ASQweBg
4ED13LCuEBoXRfcy1lHH2SpAhqvDRKMusQyhxlDl2BG2IW0kifXPKyULBrOIpYIF+sMPLdaYk0BH
47iLYcjN9FhyBhcY000gdjz7OyucdirZcUq1Mr7mhqqh9k6C+viPMKvZe8rr6yF1fF6gb++P4UPk
aWuNR3NBdbqFQWFVUtGgNNZHCvWI/mgz/AVzptC6HHdmeFrrJhiDP9QW0YibNqpHEB+ZV23xHKAV
GVTxbTjQVzntd9lZgqFbWG8NFJhc/Jjv9w6XVX4TKKdMIeZ2fyLPgJ9hyqSaNpjiQHJioPM+id/3
3WMHaYjKRIduR0pKgs0U/K8EJzHIClMeslB1VnsznBE8CC8QzQvMZ8FgFH+tVbWgK+EyA+1Kcmkk
+6oZYtEeMM6i/egtPG+DYwR18PR55WY5s1YeU/u+5nPvloCxNda2lthgOl5wY/oC2iPrbKE0nbdf
z8ywbIGlXgpLtuWqE/4ZAOaISSE4nT8qh+d61fdVcZXgx0wRtvvRuwp9SYlq9dEUwAGOU+XrWjA5
7LjLPrrH1dZOaFRbVDbWoqNEumD5z/SZcNSjAYBqhlsb5+WG3tdeujttKhNYnS6QDSQw5SnSJoWI
g/AHyUJBarmAJEYM0Z3P/euWA3hCX9oUk4aBEsa9/GV8aY9+nFNuVNobR6vz2HLQk4saCZUtQtKz
tg97RFK7nrkYwFdZeYgMR4aXDX5sEKRHxEKIcCD+IPd63HkBQgMWhUaU5fruVciwt/aJnXO1EHH8
WGJ1X8CQWlDdhuezqHxyI9vFBQQqFvhhQeZyWEN5WO30WsuXEXIdggUDr1t+J4OmfnRusNLolqJl
xgXb4PIh905A1X384sqFbOOhLN5+hjXaS8Z/7ZYMfN5PNf8UKl/Zr9Trx7ovFq1xH+RlwSaAqcXn
SkKNkX+CtdCb8zYV/gfShECc1o77InZbPhm1dBPjUPeH+JxYuAn/HJmimDgr9gbGU9jBOrkxoHSN
eIvPf4vat4N9jSA5BMdALPTNxUjEwgGY8yWkXMlrkOttm7iseR4C7tn2xyz59Brq/3g0pkuEcqPp
mT/j862s/3JMUXItUi0Xb+r10anvxOxeh9Rr4p7jUmA2CZqy6LfXYZeZ9pKlnblt5479KH9HxY7d
f8cz+xN007rSG0VHl1YxhfCEGN1Y99rSoKQJ8490y7z3eLdYme1Mtlo2GZmF8yj2UyaWzqlkkkFh
s94VAIHIruoOGWIWcpAqNMBoYPCuZV60OY/cCVa+6nqd5+w1FcJB4WsS6RZYdM7YQORWiSK3e0mt
jQGXqwgGqTqQlM60+P1o5LqDfbQeMHIrVQ6+Xh91h87TKeyW2aT87gPrgY88Ft59WrCTWWqjgA+L
yMiEZTKdFX6qomfkfWVepjwpCtWU1I65v0oBDPTyeB3Q8B+AQ4lox72rn/u0UqOAZupNc8+iigqx
XYKVc7g/CGoBghXYWPbezBY72YF9sQc/+KoDsiVc2d72NOQRmBiZb8LUGh1TrLh4i2baoSdZ7gtV
8orS2ExT0YTdTi8HeZu5UmzEWOUbOXB24HSqn2rDtxEHryhF2et2WyRBNNW9VedaIfDdUeFUgJGl
MKZI+Hp/Mwl0Apx10Pt9I7jhCABTa2xqaFFSlyZuo3oYbb62FbBtAAXr/g+wdzAaOhyKpH86ndhR
1YLDnVAGnj7FAEoZ2JrJvPKNCnNcHy6/nSR6/UapQgTTGqlYKjL9n3XqWoiN7mmNOnKvOuAdD3gP
xKHERnLTclEwUgbGuNf1ZpoCjONikzx82/KJR+mK05CemNTaav0kZftycL4PslaJHiD0BaUIOEfT
zm7M54YsbAbMZpKFxtUYpyN8XNHN3DzOLU/0zSngIR2nybyQM/D20FMs6rQzS4CeVAC+1zOHVQXW
ahFgDwtFaqfYDid092zmw8HnysSTDvhRD+jcsNvOcUBgQRHkf64Rbp2v3+Z6EmHPh/fvYVX5ooat
FqoDvSmyZkBAGtkY8tEIt4ge1klevL6V3fuwU0I0IiayaTB/xescesYVm3z0zIoqymy9M771v0Kn
fDKJHlL5oOpZjH2MYFuaMbYuy8N2kdtQdgWcxHhFDZ16bT7UgfixgEhYORqyQPuKpNKfFfDTwULG
Gc1UGKrWMVPplThzsQec7HHdICiSzrMV82BsLZZFXBDItCL0zvwBRFTEDXQFHD9GeOmwdRgy8nrI
4FifMvNIkipQuHc49bu6O+H6F9zOGO6oQqZW0LIJEnqlFsvPIjUWxrwWcFv5VpKxMi8TE6XsmhNS
VyuoAsy4hao61fivoG1LIdFbnxsNaGnNDKjJzffWSjtiCZRfnj1G6OajafQ+QDgL9gDqKP1Cu03v
b6uDIedPT4amhEt3RvqjiYz+fnc51JTRfjt80e//jTuouQeCHelYhLPw+yPsM815tdVsdrS9yXJZ
qtWYcYtz6b6S3+sYh4sUDJRDY65qS03oFhl1XzKBXOfixxiKWE0bF782UCofoWF6Mo8VswiwdZmp
PGzn0jnOsvXCJeyKS+DE0QqOLsHmNz7tPnCqyDWpY8Jo53L3ud0V6q6s1ZDTiK1v0htwtRBAf1np
jGnof8H71xUz/9OJES6UGj1f/sy2QF5++2XT3PGRwL8DMeM8lpbPatNVNVeqNQu32CA3+PuxXU/N
NUdR4diIFQZ5rYwCZ+LmunEHX18TOthyGGvNou7wfsE7ZPomWCLEcSQH/wcLVFDY1lREybCBQplG
0jeHPgKPbQeKbPRAez0MTX4khf/KpMf8oA985uVJ93OkmGU62yuz/hVrDiT3nmNzLHnT86MHI+fV
MFKm7dVECX4zd8bUFEcg+FvCfFNLX7fgqAIOF9TaTrWqOEd0Wx1Z90iT9eKBWuC3nW0E39aMx+ZE
07JxD4ySiM9g0GVbbhamqvAkP2jEB1OucRRA1ex0UsyRpQe/WOXscll5uteuSChFHheOBkw6qtJV
GgksjmAFwgH9mq8QmQgkqnoox6DGJ/MM4XWzE8FrcRv4Kv/bjgImiZpUR9OeQAWRiiDX8eq5iM/W
nRI/kuDHjIquy/BiaWkxKHyQ2gT8cQwQNu1jDFNL44/rIu/cfY8DV+KoExoU1tmbsuWC0q88dzpy
hASj4OzkidxjTZZLLtQaJhf0PgEJVEQoxXC9C0+MnsdQkwF9SU1PgB3yF1paNgbKHiD3eja30TXh
BTwdcDGe40FhjPB8LVw3x53Ztf8E4WNllYZ4B3hcpFCE2lcJdlq3e8UB8mAE4ltjpxnfuf+eTnjU
nM6nRY2Y2NkRMqhHKqOssf5jes31vXYfC8tu/hqSJqcEQD8hUDyw0yb7ujTGCPbzXDxTwoLtbaWv
y/ew1ta+AoWW7zDehH/L0ljb1gq0Q91w2GQP/wnKuIqcMNtcp5n5hNvmcg5CFIq3PB0pl8CHJisR
NlZxUW6+z1YxwAdPirKu0GRNZuEJ+yG68zpYwahSGHW8RkY20HofAEqnxUtuf0Lw9DwzeaJ47gjB
iBm0SKKxCWGe4nWCX+evLo+fDjkGVDf2pxFzJdXO0hlUizy2lP8T1jOSZ6NcIP2fMWUXeMSfPMWS
vOdVtFCLzILTPPsmeMP4dVhFPHfv0va0k8f9dVu1HVP9QSr3peX3aZpHyagDbcYnIsbDxN93iiwi
4ErlIgiJY/XVRb7lmyRM38Fyv/mXZqTsSgPQCVV8YLrhJe7L5WcNhEYXC3lUAMdwT6JpRQAUtRUp
uvgn4mOOAR2zWZmngIfcwogenDEEPHl/JwiRDQ28DpCbxDTPbzFCB3kZw22FBpL8mNLQ6i80numr
OvufFF1sz6Kc5pNRlJG//U4lKBiwrjmZNIBwbF0qkD9XNcg6ywrX+IAchDiyU8HH+RkmLyVYfSlF
vtPeisvNn96VR2ewEl2/4CXEPY5egVw2HpxzFtc+1IeZGj1ptwyHvq/giz2xv1W7Uk5+meuzzCqQ
ySxpbqWna4qyCpBYZ0tgbeAQ83H2Re9zEujFzjmiMM6Xoa7xgjIK/IyRAGU2+ekOsw7HEAjvJ7aC
BnraMDV5GKjtqMZCz7wTeFZWzVIRdobtqttSqJswBfGxmWcpILLuwRjPXcyc9C0Amq+nPwpZz77f
bBSEsrBuM5vm7fHZ97ltHLFLvFcmlmdN46fQqADGYG1TGY7jT3Owu4ERJvIDRAWellquofx69z9e
jNoS29Uk8VGXMqap9ZoC/jXYOMRxWrasL2R8pfmImk7MsUAfjf1mITkdgkzMFi3TZvHuMEb8m7NJ
8iKKCRqS4/HfXK3p1FFBNwxLsKhql3f83GkCSyyyNChIL1f13NWl6UI8iquv4MiJ3zGv0NZ4MLp2
lkPpA46WRrrL+XpWlSACj5MVUslnespGZP5dhUSw7lWIS4j5WkFWIPOxOkL9Hn3uxaqoWIG4isye
rcuS/WAjAmozRFSb6VyXowmmw6aajQpnATHfU5de48YFbRZzwGCXSD/J8jMiHczTDm4gkxU+uJi9
ISbloh/tSnjuVxgbAppUi560Bg7joVuDLQxHuTaDPqo4EjbBaC5CMMWrb4aS604WUFN0RM9sMvVW
7ixDQTrSlMp1yDE28Nfql4s1athrvIOQc668PouheFWPuZSxaCdF19lQxyfuJBtbzp83ICM9pKtW
jzPD+wc3keE4CHfrBzcV307i/9nXeMUah1ow+/H3LHutVOfTaSCb8WYZp5YQmowcryWGzJMMbHXP
ipwrHSrqbX9GVzZGubrQMnwNqaDGMw4Pt0Kh8URBmcCGhhMui4D2RsXCfPtwliaxOXK1qUzXmXMZ
inPeiCZgCYMg/QJe5GCDFyreJkoTZtKY5irga/dhZRiFH7ZHy1EsBFVr2VpvD22C+A0etQCPnYrU
GaUYMbkpL9yx0KVPN/Lcjma5pJ1MW3dknt+S/MTf9rdV07fytFwX9bpSlakQa/n38jq0fibN1lqp
BSd48YErn/iFlqHoL+CnSArQNowLYFJgSB+YSMzop2+YGFjDz89z8hWJnOLyM8Hzt7FMZ10g7TTu
XS8VQEYWOpTI6Xr5zhDCWWIRM7ze090rGDZagfqVIZoQLlaCgjhanrkpYGyVLlnbb/oJ7mny5zgy
EGxYTswADu+wuU0fweljpakTj0ytdu2gsBSKtSDb1KgW8sIpUYUofFpgTt0iF8W50tL6t5Mjaxtp
4OuiyPbc5OhDZr6KCQbRiWfPG3gQagth5yTultnou43gpuG/98LyrMsOuX04Ll2mSxd3U8rBCPhE
DSNoawcF5oolQWA26LmbP/44va+wrirlfYa+LIHLc49Q04Ar6Hw6iwIVNwgqYS/w1T7srVDbS+6A
xtFqQHqIHlw7dKZYRHgLimgt+g+Q74sdtAKT6yUWb90mPxF2HgzyJu/WYng6TwkOGp+G4s60YHnX
sg7ORKcAlWQh8Ib0dOnppQV801sZeZxCpCAANyuzx8dcrSCJCIGp091kxaZgmgQ28lW8S5LhEFHZ
y324L5K3qzvsJDzfxfb/lc4d3U2+1biIWqfpoZ/jQ8wYW5qLBvVFUC5CQtLnJ9uoKzReu8OY/6Fc
1n6y9AL67nGn66YtMEAqZjqbLyXvMTcAplACGKBfHNEx5uTSN6WFJIWhgCaYmJWPIr0ryEvFaNL6
EmkZLHGwhnXqlBZlZYV06m3YI2MJEIZFDw8WUyIm7IAq3vvE3bEa1R7Frz/feuS4QkzFq6Na2d6A
U2y7Z8rVIOKyx4goykeqTzBxyNq86llIZZYUYlnNPAPrskuB5vrgj7M4eLuWP7jTHHdCG7/DuflB
0LlnM0kS5MAmisZBVuCMrlZK3bMM2g6MZsikczYG8XIyZ6BZVaQTqYBgx33X9++3zrzpBhz9hCmq
Ujlki73qJklqLw1c+bXikn2rGY7rEf4kJxG2zHRqVJSxe1dFZ3Uh7zJ9UpBWzg7RfaXxiNBIfpAq
hMAXBIZKu0/4piZJU2Y0MZC8SutOBKs+Czm39i/hKvcyGYv0ls2cusRnCktXHB+OQxEDCxl+ZrSb
Tb208WuA1gM5iBO8dpfwcBcAgkEtpDXkuPrHr/S/G4Aq0Qe/TBnp3He18Y8pQ3FIJVIOnW74zvcQ
tMLlX6injAgAfGdXFk1eCsyvt0oMeFBG1pKqIz52aOLmhDl7YUCKXItAWbZmndzDXnL3RoOWkbce
RvmRSTlt9g377if1qabDFSjdtFYnHaNXz9A2r1gd4Mk3RH+UouS13nRH0LRNEpl6doxwgpzqplAy
ZgCAy1UiEhxjWV0z3W/lQtFdhn4oxiTAn1kWILoegQOB9UVBhTQTt+BCkAYv6GvQd3WYV5aB9GtF
FNAo34mbh1SI3lFGJ8QWzDHBy1f6qItRCCqZmAQ9GV68z1i65ki+u08GBWAoCwgHRN/L3gFTXKGf
KJ7vT9GAxuyAf/HY+rn/kYAv/9DTaX8LKJaesdZZ2uK7mx+wzAuYlKBG2pZs+tYPikSoTxOv44Tw
yHi/IZ0+2Ot5x3cd1twrOxJPjIN/N6MoLYJdFZXW6OqxENKLOmzV1lrSs0C7Z1+gZz8s3tjg9wHa
+aa9a8YW4kWlBsEUQIqLEDGQUH3rNRywFh6TXA187pvXP+pzuRpPJoQgTDDJn26Jt+bvcnj/pHrL
Y6jtRRNB5XzR51pXxHkpumBhpgPSq3Wv41Yo24UUTBxcXFAN8nYh+ai2NvPENbu+h4sFzTaL6KxT
5zo196TryUenly/W8VwwlkrGulf9+YxN70JLbWsrpJX4S6JcDlJrO6FqMVhrFWro0tgBUPEmu2K2
nMEKLweYQIkyWHJZZMzSRkgPXSXYynBU4y9W6mDreIpPdyF3/utmtRHspGt6kAVmSIyzL4DjpzJ8
vQBftxzbpjleSFVi/ms4RMNCTe91PcdFKYKRsOB99v5hUnS8P2zWMfPF3hWhbVuio2+mceFVFIuh
68DmwVpFNTuElsTrr8XgZdnaSKBJGJMnMzhvIEs61uHnlv6h/2VwuGiYURutdEG4MH0gWAFpoGUf
QhrmCFhGbmR2Xv9cg0uw+aZTBHov6S6xJaGC/0mrrmwwydLXafgOI/dlL3co4gsmbyRwjbUbnlPu
iP+pAGugwwfxE3L8afWyNmO3oMi32Ic9Ry/mmpZWSahf+kZhOifFlgrYCEyWxhqBxrZidJAkcwyp
UVaeFxVSwdZzdLvVEW0VXcevzw2MkvnfoVe3ukhT5MjQ+AED0eeQY2LFtq6gdpk+ZFwnE6w6cpUe
2nThAzneo7zxC49ikzJUPUFLShWuoFnadVypuRuEa4Q3yjlfFPUCk3SW7FU2isGaqr5sDyEQvmGK
hN8GT8uLpsu4bcZ8r9hLgT52ip3jobMau4M/gAgzi3X8BU1wGb1XGQVGGTTFmXrJr9q6OwiWqe0l
enW+SbkmJQB0+Lt2Uycw+78odfpXhPyi/DdyT3XFKM+auqxEj1wVfwaYF2rw2+gJAALtC+DMcAMO
HqNNfexasBxNAQl8E72RKbBZ7hu9OD3RSfoyYc8judeSLfnWm5xIqx9fsrRRxVh26Ya8+qnPVC9K
UVxz5suetOONabR0xAaE4nWO6fRUbT7FOmmWJ2CXgJ4gdaRdXPbMVke5gtKLmi/CXcagYMQBVIOl
ygIM/tIrckMKiJ77VQFARi6peZymv4nohDSrqMDtqVbYkL2V5K6NPOip5LWRor/S/+LHDeLo4JcD
CUo/ajNr4jszCImOVTD+nnUlGtdaBx+yEi1Pb8L6d/eU2pr9ZfJOnuhS0qOFLZdRHNrbwrOWf2sp
PPvxivodmhBXozdhcFAcV1weXVBe/hAPHUqVi2gHyDIgy74YXbRk0oadwAZkDtNp8zNGcfuYd+Tm
QBYPFL4rIqxXx6CEvqKwJJVdzyZbng1JbU4kA2F2sqRIlQ7vxejydrcLnUFBeJCZsqDV6W57OZ3J
xjCmMcRx0zEvI7Iu/kavs9VQ5p3+M8b7YdQg6Pxue4lqCLF/681lKuaacESEBy13tByNWJ9QZ+5s
ahsGBvpdOKKRnGokehRpSEQmYQMpnHrS8VPmTyNri8mLxUvcoRKk/cTG95tzOvTiFV2gGDZOFg0N
8sw3Je8y8l9w3KvTRxMgu5NX+g8VI2WRSpLKy040Wy2AMlP0l9d9PdEnnjaOqcZCy0YmjWhQfeNQ
LbIIeJAbOz28EvbDq51CcbBrwy8tT9ca0o0YkUWFND9ChqDORqkOxn46lgaGSlEM7Q9JjQKz2vcA
7LEi6S51wN3azY1qJ79955TPUhYgUpgnzBNuMiXElloDV/XG8AhnY1w0oUaJAl4S8/pbnAVLvyg1
LqMAAPAy1fyrGu0qX8x7x97oxJXsYJrpb3YsI45qYinvptS7LvMRrjhGIq1AWX1NoMQ0fmgTxmaZ
gpZ9AGfgvW1k+V48PILfKVgzb11D+ljgNtk0eyarDA6FQxwygXx+nxEeIXreIoppuHWiT8pqtyjY
4R7DZZCvqDLuOTomOi5zqfBLZWl/tVZbnIgiZOQv5I0LAmunK8VWd135IiHOBMB7vKrL/bEou3EV
cxccc+OcmXug/rtis+H6D9cYi0o7pVDNlECiGiUwmney8mcK7BL8c1wClg/f0KjkvX0ieLykt2IL
5sk6WCO6PyXcrtwiSIdi3vFJv9hY5gt3NjG7MyD9JsaflZmRPPEctpMZkRPhLUnI/l2MJKOWS2K0
fMpeozYEg8khOv4TRzeIvE8exucqy2YanQazyAEv+PJb9NRGWvsYfVNROzfArzjrx1YoFQ36Ecip
6upDZPmUvUD3yXN4SI7UrS0YVYfcpHvlvMOmyfqlO3ATeaDqLMuViWiMiXDheJei8WxysrG+HOi1
qBrF57FrW+f6h+qUq/MLHqKCGLs0dVnU85BoDO00Sj4uj2IvTEou3g2NmDYUJL9UJBZVa8oyZLO+
C9kl5YkLJmiQoMySC5GMgBEGh6y50RAgy6V3InUqCV1rd1twDZEnBdurnbgcF3vja7gY183wkgp0
A6byBUOSgHRKLqmB3LSqEn1XmlxOcMI6dnvAMU99v2PYoZsHllyGoEPYMM8OGbh0TNwPcS7Ouqne
CfJO8hV6yqV36UtO1pcnn5Ejs7RW+zGRJ63m3WLpAQxCXo0v9W051XuYFprfca1B/1ea8IMadYnh
6IVwUVRRBOt3gXsVljkie10BYhlw+F0seidz3X+69rTYGJo6jiz31Cz6O3y/FioTPiI73inGmTi0
JeH0ght3txl4oxaMjUE6G4f3G0vXU+6e/zrgFPGn6Z5ash86tHviNiRpNFBcgwYauAk7M/zllNT1
9wtxgr4+K2h15izFtswRsvP1qVnZKlzP+nSuihGWwXs6Ku40bJgC5yvWs4b00ra36p1a63/Eajoj
5+lDk/UmcB+yj6s0Zpmi5u8njxXWyXRJEwlU5TNKuwe8qkznJebOUE1sqXU6EL78hoYEezBMwm+0
bTwXE1TdzY1J1DsiVCZZ4hZ4X/zWw8s7LpVj+EwF0awvIbWKbC5dwd7ULtPqXWuMQ8uy0ddYmYq9
UiQTyjDc2CgwgKiQbN+Ud06ntE+iQD4UW7vEQciI47Qq32DUy4cBYd/JmN/w4BEbcn6+D50GRWQ6
P3vXj1jxOq5FSooCQM9kuzyGWjudb0DZJeCEj+ZFZAJOICWY8wNQXbS76TjGynPyy1p2kigWL1B9
13ues96PJiOBjNAOyXQLGyDxDrL8kxvNUMY9xSS2HuFZt+e8XUP/OGt3np1pjd48bY71/Ll+ML+u
Gu2dLf49eiDj3x8az1km8lHWs6cwAdr6pRRY01cH2ChmGQUoVCB5gL5IA9UQDrcLtYg5L9TycHaO
3V+zAAXU/opgGkenX3LNWkdBmIfNG4ZbTEXhBiHF6uv6i0SSJ7+Uy5U3o2gVvVmB6B32bM4hdfoS
pIR8/62uceCldwdTudn9qMh+wSOGCdkSkyDCX1qJXdZeCBeu9TVot5FWrn5voYlJ1vVJd/4FZDDS
fUPhWpgHeV2Mdm4fQjxmJns00PLvvqROS0UVvcoAJv8Uw6RKa4T6cMKh87cELu4Bow1xcwwXtqJk
aik8E/3xvi+ZXF5qVuoJE/nBKkd4D91pOTZOzAgoM9FOKBYLRcf1ngAjpWahILzR8GoSPFAzVvhK
H0yKKgcSoBfPDNmW2b0i5Oqr2hgNTpJhfp3tyUJYrffWwqrYs3IXujlM/cVsIC10Vk8PzISaOZKf
fTwj+blChDEiEHidECkgaaR6Kiq2MaSbRnJIqtt/Whw/LRFN/MKdVDJbPMa8UXGQ0nxnhqQ/6e4c
WB/vhDreUQKylmQu7CoKs+L0fC18XLBVBv8ptXAawt2k9UicDgayAfReZsUZ9MuzEOj6tmvKj4P6
OamoBU0prchWm/JN99O964Bm+a6/3tvi8yEnLDAXfPycvXgbeXjbyPtZ9Jml7YnWsP/0N1De//iQ
2KeyzZ/3FjcHx0F79zpudDu4WZFAqle6cwMkQIeQ78OYxo1gAa5KBC+U9z8IOV2w/W+1O/BRcNfI
hALILv9Ryfqpi0CHX+t3AnIwwRpD2AuYnafoYOR4evs+uM3J5ZmsKtXwDHPrBgLKhi3n1JyFgKfE
Hoy1WnP6OkOZjW39yiLw1gvVS9/ZP5cQJ/wjn4QkDvD8RyOr6by6wxDMlqAkij8Usv5fI9Tsx9zH
Q7Th37UUumf4nxPGfVgsjvVpKa0UKtYO7nkFlie0csjPm6WAMARXAmJh+wDJ4H40w7iakgw4gONI
DCB7PmZ8sEBPk9kT9RHeOpRh2O51wKrBIWT+f0TZzjqKiD5MKMTASHZ81aq5av9PJcSGGlJHbCQM
YNrAFRDMWSWyTDppoHM5ezbKAAcTQYSqxg5Ra2SpRQakTvTOnpKCLEp4zlX1k9Lv9C8vCd+tMl3U
qXca5b8bGxnEY6m9DccYLfgB9owQOizkRV4yCkMvS/gmG8St2HBr7JLCNwP8UdW5mnmkgceS9iHD
sOed+bnGQxjSaBAG1FpDlBBLy9FY9cVdb9rRU5GKfPUe47GpG/zPyn68TqzJwmBnnwzn/NLCSh3v
H12SGxMzjzDN9IexO4iKDwYZZ9tGQPfusdukSxJ2PShdksdkPGPuNyIpSMOXH9Tm1qQVvBUXYU9r
TXZrsXHpJsXLVGrnrFTVrKNC9iJPWrQD2ZSOucahIhOsbsVmT2nQRHjsE1vDicgfYgRan9RbpPId
tgXAezuX6YjG3hBj27kTbT2cNt9PhKMgeojwFEvLdayybgE+jY+68ac7nd/bACqcYk/bF0tpDZ91
VrJ++1giEMjKmzT+Qqe+tjNLHRwRzVHRHMU698gFFd7SQBDSad4ErI8us866NLkWPqnl2sDSZ2RI
s75tqDHwumCzRM6BeQPPORZUMrQJ1hnkmLEzr/JMvB0ETrL52kaTwRE/AEXJA17ELPDJHK+gwehn
mPVfVhg32axaUUK+U1AT83knhe1tza7qucBUQKxwEg7a7vKPNGj77H8pvAKq2Cxjf2UojG4G1Z7w
6aCkM8tBWiNMxGgmwezXZUAGL45krfsSPxyEEomJhfFVmakrIYWLWzs+j3x4tusAQN95CMC9Kl+G
ujBmIlVq+Kw/uoo65jwB1btEiIHpC4b0CsCln+AUpCDSc6HszjmJOQdGmMiC3XMz4N496wLiKPRu
XugBM311390gTR1z/xFNqm3E1Rk0bFmSYvgHchE1W3wXdXzdaPsMq3NxThh+wuFmWDI23+M4NWs+
FA4u0QKju7c58kIujbfTyTMVcIf+sxdf4gMu3LmLfnnk9k6Gbfx7Pkuj/M7M8A20hyBknfSTCeNj
oKtmp4TfvVqQoIhEUgd0HN6dMLIuSAx/xJrvxES+l8VBqpsEqkTBAJk6Dg9MPa12nmiiFJ4UyFie
smQnWLq6Qgy0tRCRzkTmfRRCTmDMr+e6sYFbiXFLMdfh7Em5nw9yeYIwuSsJssnQ+rsqgMA4mn0m
d06c23chDwvoUdJkj+NDf42EAA2qGGfEvYzxrEpH0V3uiLtGo+x+69G1JgXVFyF8/vwybhM88H7N
s9FcA6nOvirt61O81ZT5FsmZX/adT5CE1o1/3QS6wHl7VhSD193PVXMe21D2t3BILIX1V3jbzMaL
Fta07a3qLcgMMmNQFXDbr5uvkMt8ekWMfsD5/tINzJNRlrzx+SmC5ay889iut5+K+QfoaYgJCbuM
Ohmzb6A0ZoNN6aLo9JbywPsNBXVWEi3iZpNxTCf/3psf95pcg/vfIj7eqeHg3h11Atj74xx6ozM4
mQ16aVD6n8EvjC+WfHDfHRJ6CZJbLf97wh3S+u5tX7Uz3WY8qPC6ghn29uvgUyd11hRJUlIau2gd
SFeTjbpbWx73kaxZxAE4PNnhaRp/qxEDfwAPDRmtLr7A2DJLqqTmXk99bPC5pM1n6mlhzlEwW2eK
muk5olV7ShP+wudn/b20a32A+a22PT8ciljYpMbs05RlEFoDPIXwgOIFi3kuPCcgfgUFAzzv4L17
twIwqTBzGKU6EXIJ+abZNA26N9uoFSfYDjcUyA6ajlEgjrPM2hHcJoFWnYDJ4BNMKut3UtrZLlyn
71Ycr4Xa+890Vas8xo+dRstEKcL76smEwiUc5ont6Og6pCzgQBYz0GYafsOh/M5FDplnL0/zH2hp
5Z+PAXiHKQKffDaN+FJpUlm3hbRSugIECslD6V9RUyCr1xM7Pd+m+BWktRATh2YnrK2IFT6skGsH
8Xr2vjcYqSbUuTKi86U/mTRRVwB1dVuvRkMSVtcV8bh8tn5KIFuSwwAnieR4q3OnVeCoytsZfelv
6h9k+GQYfYHU5z1pQlsqHhlX8OL08S2MQOmwe04eFbCGq4KwteZVWu0KYUW/iXpX0qDqyun8SIyj
Pw9I/LUHFu23vJq1tZzVyCZMn2w+hUbBEPbD+cqqZgKjZ4NLGnIRiPi6Qha28SKmeR6lPSpTV1Qp
Km4ChjZiTahoKxYrq0WGeJcE7V0VoN4wK0iVDNrQvR1FRPlGzIfPrEIFbb2LOvJTGIQYWEYCHcYd
b/mC5wv6p4GITe+xe4CKBwYS8eo5YWtgcby+uMj9vqp/gI8iS/M9ls6dqgCE99xNE7+0nsSwJAAg
lK47KricplPM77cljkwstoiVxXmxaWygKnVQkvrYg9B0om7PhZTIiOZkCd7tss30khdHbcsSkkgN
a+aQIrR96K9w8pB2RFI4/D7FDxGGs5m40ijCpCiot69prsXKVgu4WxkwtJFE/5BvzInJbn4ffPOE
1RPIDIT+eZU5oNxf00kMkxYXlXUKlb8KhJYm8YJfQazQnF/d+vUSPjk8ApNyB3vB9wdXBG31XWRm
n7oZf8IWGfHtqrz3+kXs7JQyL/nrPFKUBMn7UlI5JuGkC9IhBNHgB8PF6gKRiQehyHLjfrXnbL20
fb5NnDq+21usCAvbtptPsZMc9aQo5MLhbNysJE9gxL7tI4PcqymE6KfrXEWLGlSxqNEaaH28Xplu
zEXQISqUSn2ABlGd5/e3xYKVw+dpRxuAkfuPthubV06btFuUckpVD0Jwt754KH2JptgOhBWaBumR
hWM+17pooLVOJ4UVxzspDvL11Gsh0slPDBHS3XdH/JwvFOpWgFIEDDr2P2gNBQq2/XJw2SAipRLy
kPAnlzOLl50UfOhaaOz1ux2QNonOAwbzuLCCiyJWlMs8TxuMnjiHEoTmTLAe3NNTnpKM9mwYAkxX
WoiShxkdymE8nIlY0wzPZBYjiURmFx3JX21qb4RIMoHb1OfCo3XNBaU945sn1e2yM6bDCERvDc/H
01k8LDSvll7sUPlvuBK3wvfP5cRdjakirCb+4CplQ+yG1CBnaxFtTUHUwXkMwCT2iZ4xAD+6Jk+2
xT5sj8SOvnwMw/H19UGgMEE34k3oZnZz8Gbed4umv0cJm3AOX3Hszd7GnhXIX2WwFOGhst61p+qu
AiXe4hQlSh2ptrcjSz5KoKvcjJeeISkl135mMiuxXzusEAGlxzN4lJr6ANT1y/dLuXk+gomOG337
gNDCeryeWW3xsxWx9Hje2T/kqDxQJ5ZNZqhiGT37GHnukfHiCm8NCozkW524xpxee+N9qTiYu/oj
Zr1hg0Qpc8VykBChKYATqoPqVLoWKTvo7wu19qtuK5QJoP27qxcZVCFVRkSFE9i3vNKfgd6t8yfe
5Ly6BdTblEyfg2EOblWulhEOMRB3KVXTTCl5Zqm4BLW44VnpsHQzwAiaK6SwdB8aVo/jDrzrqG92
HDC9MrscoW8pZKrnA4NTzNCWiaFm/AlZqhbUarBBzaihu0dRaf2TFqX/X5DBrSzoxbKpZaahhEpJ
+4Xhm/jYwsjnBMvKg/+7c+MzBstoGZRS/i3RDci5bL+hQD0Dy+Tfb9exfsp/LDkDRINfqfYkXEbC
464g86yQ2VbJuJqJvJKAs5WYunE8qmCFNSZFzkIoGTU3Xv8kMxIKbPaft9q9NMey/U32n02ir2PA
a+giucJsvcwkAwfMUGAgtr31HOsmzjw+IG5Ey45mdBwsOoPFwTtGYw8q6DAz60RNEibCB5HmSoxw
1+HEoGjLB30lYrE55Bua4JhS3lxP4HyNxItC/70zd7W424IPGD/R7AJsR+IkbhANsuJjkw+IrvZ9
nHIw0A3FfU0PCaPUS8U5s/AXEe3A33qC39jeyBvB4bKoEoas/i6hrwEFe9MIkefSXp+l6TjeNC35
vPyQBxlzLraE1xi26c96j60qQYBxIZJq+2fuiGYqMlpMRA+I/hLYXghFShcuSmnk6EpXhMoj8UQ1
VXjhigDBiFYaWh7d7zLmdYQwull+1HmuYbFEnPmiDrdJJ5O7lA6zINuLugiJDO0yvxU1d3ZRppvf
k4rk8R980M9DHGvGHBbzziD3Gouo84YOp/NkuCSY0DDLSSSQk82qWcGCMzK6GPNj4k232fOu6Dtm
Fl8uhXHCQuYCwbkGly38bFLNLlfBo/EhZvqH0wgyXYeTkQCD67122Id3zdldKeksdd8Q2MWzZntd
VybCxe5pHWDoxx5dROXd0mid7s2HMajve5jYLZ8a3bmoR5eEgurEOmpConVNzvm7RSV3m31BoLZi
RTT0KbS248DqnlovAMLzTuABkX1ZKc8RksuQAnm0RC5BBh2Ki1QJOLDx4WTEV7lGjtF/WnOh0rAu
I7Iux3g5Z+xcwxOXU3qGl7xNgMYYFXJG9J4ihTbcTyBxwJQ2E32tlwP86MRL2gujbBKQIrInKaoD
DSHp3CKJSB+pJAcjePy4nY63oGJH9m4BydZbPXg17DBnP0ItzbUPc+9tBQtXcxxLdqG4uOP9+P64
OpBwWZm/J4ycFNUZ6kg0D9hYi048F0DRX/kPjjCB0msHLDoVOO4vUC9ITmJqp0+2kqGB/siwg3jS
AsHiY+i8C0DpF5uUXYSV/2ZTwIPSx6IoRJX2TvV4zG2TAKqGbqUjK+EcqKrxCuHm9U1fxnK2VmRF
bnolIiWE9scaGTTekyC6jJiQyYY3Pois6jbnBcSq8Yxn8Kt7MkkTUZVSPWM8zWE8hUV7odyxNA1j
yO2+XMuPYEX3VoGDcd393tEEEXTFxAnfzLYmOYO7IwBnjN9e2n9C6NpV8oW2V68nJihEgRQnGGop
lbuYDZeRcgKYGx7LlKlVrYaEJleCz1sP8kTYqivTf8NYCpmJpxKhxwhSVzl0sqPQ/p+djhaWZrbg
2L65QrWeYU0NMoFqBtJf8mY/Hge2e1F1ySVjhYkTZzRHaeDxpUDnY2LpEH2SPrJjw07ioQ+zNJeB
PZZzVIGoCaH8w/o4/LkwzD1vO0KqMPqLA+IRqy134SU5DNrdqwEjmNVuGNkBI9ekq/FMSY8nZBs5
tXbQPZMycJJ3eqOC/akW28v7py/3z9dnRPABc2GJOCLnstwhpNnarqGJRDqBCZsaLjtDoMkyWlnw
C6DTELu+G2fNLP0MwLTPcZRNnvxaJzY0kgihVqCUNAa/jfa25IJv2T0G525KsARgQ8f8shltp0+A
+LHo4wuf3Va8OGFO2Uv/4LR2RfaCwdBvaf9ixKepe/9bxSVDWgnSPQLKlube+eFlqPVpsB85m5V3
DIPMWHdmX2UWizIoCfPgOQe2+iBQjhElKlr8JH7alkKl1WsoejW2tAfzmZcLRxT6s0jqIcTlqu9+
KEjIn9N3FjF3Pc7dQyaItYK4SMB2Z52awUCvbqbKzqXkbVuAsOib6yFfGZwmRwMK8cyR4Gosx4m+
0yVza0BYOYbOefJto0HLB5RoCeQw2Dhi+NbE0gfBUWVUeD23hk1o1WuX5E37FZaSFRBsq7XjMB4n
qSYyUEV4BFf64S74jDc46fj/hmFbRC2jjIuT338SFax8z8S/EqZxAYrCUP7N+gabTB7C9IWtEfuS
9ndmn4gIw0TCKWADudYhldMYfQBnLckS9BmcNTY/PK+1o6wOqAu4t72nz1uCI96pAAiFbMG7SlVY
seeSj1iKHssDeZGWzO2AfgWja957jPBELHNKdt2WinRbWAGUwoeqUhCZ+4xxZ8BCrcQieTkud1Nv
eT6GdYHEaOzYiZXh85ulrva8uEvfqgTBfmXbMqjdjtogX7punrR8S+OHxgRd0DN3cKkuRkUWHb7K
fyMeCK0wZj4Y72WPy8FlLey594fLRBlek25Bgt19IgVbx0/KPgwa4B0qPORzXMmMZ6aAfeE8cKZg
0BPjW0cgnHw5MmlleToN7lGU0wmtkGeA/WAsoYXsySHSCDHjlsqdRUTbpCRDEUxnxjGYVuHNFA3o
7f6nRKEOMv3qBaDETJOp0yfyV4zL5GeYKpPUvS1qxj/7WKzwud2VK7B2DP+Yckd66pKU5hC65uW5
KiLFs6jF4IgQQ9S1BrXaG4C4LpS5gfUk6EgYZjdZ9elDO5oJeluzzTPikCEn86biMQoETY/NWN3g
FbYd3Sc4Aa2UG2E6cq6ZfWGDxm0JBI/zGGJevaN8j42vIj3mR6byJX900uANOc56l2tdy/+1SeCt
S5RzEEsy3Gsy9Zpy7btn7VufVBbDXZHPFE1Xn69x22QulgVEc7XnEQVSeRhRJQpBFT1KzCw3JWoe
/bwNPvrtjH2mIvIes1kQooRQaF6VVAiz6IpswmMAbh7RD7YCy4C3hkxAkxR6yUnsj9A8e1AQFOnR
JQKuWteY5s74gXZL46+EBIxhh4srzX38f3Yx1nrN9gMwWES7vCbHNX2ZaF9DDNKiHykQymzAKr73
bQQeUwactIOgLgpyRliHGcP7aKcdjlEhlD83wFIs6+ozFWOpZ6vSiG2vR30M8G9SggdcryVT+sPy
oK5548u931Tib3G3rCsOYc0ESMr4QUrdkndTDtcRPTzkDILCSYXCIgNMXVxadEdeDECZfmQ7IX28
oIXr4XaP1JIISkbHRFFsgb7gWQZOS1wqmJ8YhxSmx+N9Z2+y313CBC9bVJhTbOwbMfPpMrY/Ll7a
cze0v6N4VzwddaYTzlZPKYRb725bZ1VQB3ZrvUXCNZt4DihheOXIpAZ8dh5cTZealVe9isVuoHf3
+eJ7+lK3Cg424JlQ7wlKa6L4r+EZ8qNLL1iJVGsQLh4xNjczWoob3fTXJzhmL8B+bDakQU2Ml7V1
KItCB8FiGo4zxx+QNzlj78+oB4+4MsO1BTFqTJPM3PPTmYYheAWSO5HnNXW7C8LM0cdduTqLBR64
Zx2i+Am4lXjCrc6NEcgEAi3W2/1FGQ2rWK7kOVuhBp77rfzH5Eis5miyBYBuC2xJccbt+7iiaa3f
TI4+dOba8qGbwddo6Am7jI20ILEMBwRTIescu0Hd74wqXbby7k1eYmXEM548O0if2LE7pN6z7GOt
Y+g+waEGgnHPp6zj9yM0x8dUWpPd//FMY+R+wwFg5oj5xaTG9Xx/zJmPxx/lMBzgDWkqYAZBN2hn
gUFg8A6uwMUfKC9iln7BLEQ8u8EAmW1ixAtd4jY9f4h6ofjFtqCWu7GJ7rK8rvmHwIm6bk3nSSiF
VHK82krhKv+d4iar9iYpnWR5o7lLbKy2+B3OhfRjhypDZgzTIDoUOECO0KIwVeRr2Yk0gx6x2vWQ
7gFycL6/BdXCU/XbD0XEIidRhzh5GMV1Kz4cRrlDB8TaOfDoKPvw98/fwlLb4eQEBUpgJzdCq+Ay
Yfa5Ot8+4RoNTwHX4TGOFtC8G8JDQYqhl6Ovg2tuyKRoS73cur6kj/ejs807U6tLxaTjBPm0oYAV
stSzrkif3keQUKOEx5TtefP8huY8WXW8GQUajD/agb/ahieFclhORH3//6raCmW2th4wTbdUH6Wj
g9DJQH5HFb+URuKzUzRpDfozOB3yj4cv0jplCglS1mDeQijlDT3Drr+ZGJ9fnVBlSSmnrXdfFf/d
+87+3PdW8QIPABgG2ivwUqG6xF/FRht+uesJaXjnaT2F7XX0PJfK5ZlmSwQCy2FFiYLy30MF8Voc
C+m631DUIGJo2B5XTFCaZ8QCnjyhqzoTGMGmxI9aUQw+EcYpw2F0VpfE9bv4VthfOpigcigLy7Dj
nfHL6TtNl7h8/p/PD3vQdYxQ8HXP5nIIJsmY+xWxt3QdFwl0EfmesZVzLsIvs+S/qWClT0t+z1cw
EyQSuuHF3hUsmkK2ua8fESTtn7AAjIu1dZ5e8ieaTQuR+kV14ihmQKFzOkL4ayh/984+HWYwNwcX
rQQsXYjyoxqg4gaMa/PzakdVU6FChXETuk5Jn8lpOWfqHR5ci0YoFCr+lhJGV8vawh9+FUHrCu+R
cjsmaOW8gnVTdYwnnAOjDaARkTQESrkVpN4dePmWJdC8K2HGndBeKPwkcn+gSNcpfABLvTSLBxyb
wV2bd3YyRamkNcUYccBC+GCOT9nfHr+zcYR/cTnhWlp0wZnOtxvweGzOiHondO4fP+23y1CDhqcT
R/LJ4HsOLJPQhUt7gTkfAnNRcKUS1R0wzG8bkMfS53L4tpDLhpWnakUti1hQUcu7Ifi45OvvLMuV
JLI1Fqfsti3Rt9FEotnPymEZW0MDfBWRgCkYDn+r7+oNj+dLAvF/OaSrJjgH9Ooab72yARWBJvHq
TvvijC2XPKXeiB3nCg52rJJU+i1h6/6QQB8V9rCknhyUrmQYIYl5GnZ4cHEfhU7yEP6+wSdsABDV
uwov1gAxno7cGuwm6Lo1EdlN7XvuHxTJ9G8U7llwTsQbFrlpVBGeowTv6EvEgW+mf+xWGdZcMK5X
yCULuMpwUHzeCxriQm7Dn3ATr8A2DdIT4oN5h2EoUz9Tf+ZSO10Pw6wOJgu3buMWMgBiCA5MxZ4b
I3MP1LhNR9Cls5rGOI5Nn8kb3G4/aVyEpzBl+O670TPthGUYVIoUP7e/KOB1gwAxU/O6k56GqYWF
v0Jtuf2yGIWZZGnMv1JgxyJLMQHm5F1OUrA9ndMYoYiyeJPRQoTXkfnEiCJQ4hhXCY1iFuW7dBRg
yhc+ULNZARECvXaax0brR1GN/NbQlO30zh+OzU4I3LfZ7YkD1IGYZfU8tSHQBZqTWv3s8wo20bFX
xz6GaW0aXgPvHzPPGYAM6tPalDB1YRHdfCbX2ezjqSQn7o0101P8gracwbyqmPckaEzlvkJmuhmY
Bj7d80kRDDE9J5hnKtxaW57h2vmge1d+dRo95qluaeVeahDa3ZlWWK3Vk/y1iu6UPAJv7UHbXubr
2xXsILrKYwUvNPNbWz6qAMOo50ynOGgnw47jzgCPr6HzmDTuHPrWJQG7LUvWQTN6O3SKUJ5RFahm
uuKdXKHTdzF9tLSit6xi0qvmNJj30L6EcIGcGQvULtiPgNlYZdYuaHhZR/vx21zq7UTVHlnBtT5C
+Z0lHy2+cJFMC8zY+jbsSgVzBAVyg2GN/KW1Cpne3Iqjm5+0B2OMcbs5iyrihlfJ3g5vQ1VtzH58
UaohyNyq881ETaITf+bFqALmkTVHWf/pFGgm3r9hDIkarZxp9f/HuKAHWTZtqchaPVTxUVK9xsqF
ICCGRleYYuTH0sAqtMyk9EzUjHlHqz/DlrIh4fKF0F+KYzAdA1etz13K8HPHTktk8nUUekmP4SSs
NUKRLiQYeW/da5XwicUJgEuQXNz+tpKr8wbgJbDghVj/dhTjP3OID+8rWk7onznG1Q1kzdsCQ+4G
7F0bSr/hV0ugjlPEGk5FWjPbIEbvZ5BXlholGCpGkPzHnOMMwDtCxy/C/BLMk4k2C/fRBJJ7+cP5
RQyGJhEG6dlvtN3imekmREQH2BDJDVlKxvkl9WXLTXm804+xCFlXs8agXcZR9OGZy781RnO6AsD4
NrEDgwO7y6TBRhaI0mQv33aI5QKOVQJt05INrRygF15CwyPWlcQbB59Kp3jzecOBpAKAbt1rz56Z
7jIXggf5BMYkckKdE7uPYwI1fxQdIeAYt0l1HhAPOEd/MVqj3Gw/PxtO4tGU0YsuiWHS3JA+XWhQ
dEMHFR/SFH9yWqQ5un9Nr330Je5w99k7slh2OMow1AvEY9GpH46hbQooR+sE7GA7oM/gwlWp/hhy
eAQUMCxi0Tp7NAMWixK9Ao+FMuhJXgIz2YBlDAWDVVUBed1vRZ8PW2hlOSF1UdasdCeRFlCZugry
wMco2cymQ2zqSbY3GBSaJIlzFAW7a8b9eoTt0vTcHnD6CK9rtGXFnFK2qU1LcPsBPHDNSx4O/7vB
0PARAYtbtt2+rNst8rpCllAdbCBks0vYpaF0uBpo0Z2s38iOTy6Je/TrBhVu1HTSTepn7AMDKwQu
cHlo8lxgIMfg/hddiUiMdAxsm98GjsOJYvlNcX1033g/q+XyqdfVwH+2dTDPlUpK0R+4TfQAMTuM
zeNLxPK+eYSkRLoXBGuqJLoTpy1Wl+9Cwjoi1xCPS4wsAAOIeyArnSYWOddCqiQUC39BsEP9yP9+
C5hDbJFLNqFMQCXhsRvm8v+RlRiZZy/kmYeN/wxWm8vULBR9aGzIGihts8ThYHERRhvM/Cposn/J
vN32nfff16KELgvxJsFrHqLbo2JcbMU+trG3tJZNbz/H0oOQbZl7yP1tPfXwD8OXUfkpeM+TfvfT
TETtEs64kpZi8kGV57BvfIOZNsDDZ+epxm2S9JwO3CTg2YycVu/k9adMHWwoWw4eb1y+2Z0URYi3
LnTlTGnVXdQveRiM0Q6RMs7qxXawHR4NrVl/cue1PWm0tx/FwLOi7V6jQoFtSha3gA1AoCppTiNv
srOQg3iguP2EWG9E4tXJ9kounInVswp5ZUr2p7KztCNM1IbthB8XO75M86W8uBRPjq2SY++RMQN1
HTe7pHNR/tfH1VS8JXyGICyO9ex15tPqOqyhQSuk7Hx3H2yq1Bx1AavU2w5f7OJbWpwfvTfyToak
+ollRJrE0gIRO+JnmCGMFBUha5J/ViOwkrkkcX1ZqzjizDknsYWKt/7UeyuBV1IQXdm7WxVUj5Uy
/pG6NeeK4I1wFkS9wf601KU6qos/iQGPbvLJmdc0tTzxcIhieIYIDs92Svx1rhZXy8pdRYacD5XM
LPDxE5vD7W/AyS/HXM6p+NUwhuY2kZRjZFBD2NEH0Yvkc66ynHoDdshjCv7ZsPyZxTLR3+M6k66M
rIAZx4syFC6OWwjwBgD2TLuJUee7dNlcEe9HmCwW/nQYCG1wMkcN2T3Rh/NHM1CWm9HU8aAkB3rT
nEI5YXYWpUiIC99cYBbG2sSNYXpoZep5qdye7qwgyJGBfmUd0lCXtIernTo0eOdDULA+avtetSJL
DWTahLKf/yNw3mfkx5u9tdmHaTbLHBZPe46BK79AeWNLbpbfOQ62woB5D2oWYe38s5kJS7BZLPXH
fDyH8BYHU0ovxQpxczUt7IYNHMeaeB6GHt/iCfgTiPM5yCQ+Z3xLJ4ovsQETG2cCGWlZeD8/Z5ds
geWrzbDvrygyKAvA5O4veRwbEv63Vr5GS7/OgbbNYtzC481dGtCOyzK53DZqL9nQ/odHm0EFAw96
lJk2HrYzonWX8RFeTxexRQ261zbmgS4h3C3QOSjPXwV2kPRx5wk7xG0Z5OZU5dBk68DCY5wZy3sR
38ceRkHn/lJm4j2lYm+wZzDag7RqJcN1PeMnvYoWBNm84t0ereNYvEw3SIHIB/eb07UBUBTFBFN7
cLosgzJjXP7mgOTjs04MnoLNH3JWr/nzRNubu0klwFMaMPbCaDPqAIxS9pVgHHqDePAIFDxCQ8hN
YLupUsxYiYAd39xYdPs7ykdkIGeIrR487f4HLg6Ck2CUkLCNf9i2nnq0rTsRVKJF0o+zA2rBEI0C
YWa7w3ppRpnUjQBVvmcvywUSsBO5GEZC2LhVE4hZLkFCIXzTHTVPdMhQIm42RZ52IC69dqR6ZkdI
+aP6qStGIDpHrXuwn+0fzoAyVJRm+8oBUumBzB7J9UCSj7Rb0lbk+kMIATIBhiUxelR5uNPTOs2e
nktjzcK/rlVDx39OWw/v5gm5xwWlJBrh1LYBEoLXdy69Wq+wZxdGLhhzRMXkUNLIs0KMPhswh1Yt
fEVkynWq7pYYkh69QHl9bbn1bTwfUNM/2eEMZhitu83w122tMwCmdsAkhYsVNveawUaYwl/t4g3T
95GMU1WBqTH2gbFmuYsoILDW9FnC1W4tbkzq5i7533gSTg7FQDUuG8KckCkn5RJMPLSyfjdht6wl
3QK30Iu+u8hIcawhl9IcC0XFPp5E33vkXuPTuwmuf9j60eptkVBW0pPQr6WlazLbvRLgB07YlbNI
yAuBWJM6Zt72cqJs3tNugbrnBUxOB/h2lJC1iOhwXY0tMZldz4KaKaHLsP4+3oyO90XlDvxeql9I
NT0BQhWWvJ7IwTU8jEbA9mVTgwIkQnksyKRQthJBWo3Lt3IpovoW/yzl4eNcq6kZa4Tz0Qcq0W/1
6GaI7MRNvMYheB6h0ClMUQqylOEWDlsd0o3xV2kLfAUA9OVlWn679BeXirePJlYq1bC6K5wcKj7e
eme2gZw9XfREvNvnT/3VIMR6omS79ny4QOIZzwnEOYoyLc5issbBPA4S7M2rs17QTHY1qvA4kxCz
8WKINyJ4//juQC/+iIbkQG70wbyQFzTtncTqy+FXlKoOm8WG3cWIryTHz0tWiryU+2YG4JBWwC2I
YV5kLwTlpajWbUB6qYm7pxetJ1JLP0QNeTWF/ujHoJOVHmCpv7+z2f3gYLHxsoJ3zOH7H2IhOjL8
G4C60A6aQ0YoMWNsNUfbgOJUMKsN8TedlhMCHHFAExn2bKQ9SRz9roJZn/5//OTxaNotd+XYKJWX
0CVdF5KwMjU6D7TlGFH3MWgD4LhKJHWoz1MP+UgYZ5V9dkXGWg/doKAiBAG+NegDpRg6FmI6X4bm
nv+JIRpRMtZGGHsl4WoP3sI7ev6qG6DmDDvXh5BEYQy6iDMk8EjnluurK7D49MFGtBSh9EGAPA+E
0wMhVM5nwvp1TZR19cZW+w9HHjPRZWLEds09ZEhRBmEKYhuCYCkiTMr6hOUtBY3Pia/sxRuj72s5
EZnznMYZC9+ixyin5LnNC0mBFPpAQ07FAibMNwEtIO6e5StIwSLsJbtN1tbpDJOszY9msif3q3MA
JE7uNz85hf8HeUAhesVUj5Vyx2clUy8wrqg6hxwPHzVNplEmYp/oBvYCGQJWGY//4KBZVOZe2ljd
MPgUu8/1oSQ+WqdoDb3QJhwB3bdAI9f3gHf/JHPZq2gkW1kUxv+1B7+NQ/SstTXJikyUcRnwvjLa
ZIJtPKkDhFubsu3TQ4ivoqj+CdcBZ27LhcZ1DLfuMIOXlcw+3cbOjFvabiCIKIq+eM85t4GHT2YO
Q2kni8J5b09xo/pmG7+RdnlK/y1CdjSiENQF2BoIjGChh6spbidsiEOaGbvwgwKO6iXasZwYmqHl
55Bu8TzFdNVfLV5qV2S2iOEvrkJ2wiUBcNNkBDMUsRFVyiqxuToSlIjGBs0Jf6VDfFs5AJ+tzAgU
g7QMl2qy6wIBX0QS4/ovt+mtOku14n9dZQqj7j1NBfry+dMxOExIYtQn0QafTPzWHvAFRD8zmKJj
CVi+slb5RyHtrPMQY0WTlfhtxeFCxtXpFIU8JrX5A3Jeu0Cy6Cn+WqHEotY0Fum4vJMaMs2zsy52
jQLqH4ET67plVc8zHltEUBxnHgyyuRo27K8gHDywf6DbYJVsqHXVxyFjyGAPMkMm4OKMN4idnQER
bL352MNvKFn1kE/x+hJEq1fdyOTHXBkFtCtyQKOB44Om2i7udwqyxcdBBvThMTS9UACTP7L6kwf6
MTFp72slfvaNJ6EYfZCjsvcR/tT52vttM8DXRilfHumaBH57glY4GgKlf+oHy0LYG8DTB8wb8KH/
1ionetADVDGnPe0hN4HCG4JRjyWKzvpzEU86Q7r9x5ZtNHuAWFtoKPrZWR10MBHaxlAzICIC2dM2
qdCeanhhu1d3P6KXKgjkVvaTxwiRxhTnmqew3cJKTJWYEwF0Mt9pAdHpbTiLDlBKmTpTMLtxpVGx
24Jrto8fdfDtYyEfd04Nnq8cw3i9FvnwCnln/C+DHA0iJ71T/vE5nzeCX83kR8HJ5mx9AaBmJbGD
jad5GpR2mo4gtJjysgxf91WOsKZTz3glL+d92v/dMWZoQz6cpslp5fOg++GHVPAsGKRDpZVedoUx
vDWgcjIu4ep2Eia/rYiq9tMY7dgawzdLF2QNXi2RU4YpkAVqwyy04AxWzffkpQ4ioYza1JrV3IUy
whBbY8cEvp2szTbJmNZo9W+Z2oKqVDdGvtNHI7qQVchpu6cTR2b9eOiXepOQK5HUk9RAJ/JTtv3z
QAkRGYMCfpBiqTsgL8CXsZda5rHRYd86hniUlSLPB6DE+Ap4T2omw9k2MJ3ye1h9EYE5eDSrO4b6
xAeRrhOFvJWR8q9Lw0UbQDt+S7Rjq0KKn96iXbnD3BDkpq1vHYxX+FuTL4HcjXfAWhQYQ0n5jwbV
h3Uub5osDgKFCuar1JfDDEfxSX1gneDr6v85oMheneFLr2Gm6aUPTmzyr/a8VHy52a4pDnHXbw33
Tki/gKb5Hb2snYVDP9C1Fs4BmkHlrgIDRBHFETU4cDeDCp5PjszfOWW0BPwN7R+U7OTAxQ/wWhsx
fiKXagjgBPxkg7NFWo5qv4clx75l7+HfNRlyx0j0PK6wSDLewqTTfMLoaqdbeCYxi2WMjobGCSs7
mWTB1jc8WEWVB/LnobZtn4hS6DBu4TVXCAv/rgBU4ol7/To3BQue24fgiaN49JmToOKrQNacDx1D
khBV4DlV4PLsA1elgp5jgH/45WLYXxKVgyNWpyE1sfaZw9pwam3ustNtqARexFx2+CLnnVfsypc+
/N678ywmR6IV/4AWWwS3yGxHK+CTva76p4+q4KRQiGANlPR2uiN5SX3VhXglG6CwubXURl/giQwP
/5wPdwQnT9btvC+Te5iHs3W97Kh5pgP0fcEnOWQ+Rcg6uOvNqbyEChjbGvDwc02HLDtEa10dWIb5
pc3PF0+lhM/Ve3z6z0ZSeE6wqlN9AvS12wMeS1SfrojXKnv5EiI99jsg1g9KJr++3mzM1lF/Sx6u
bmLDjMS00GBFoqDOuoCj5WI5juGd8aOe0L8wk2NTy1aB7LTGrP0BIOWg/gWiYbbyFNLtfJKCE63O
01CwxExtujWPEDbcsTDhOGeML+rEnUHdEydOfh8h1SvdaCOQ5IHR1lwnQBLqhHzspdnCf9E2oGD/
/v1+Gnhhv5+UkbCBMLDkFZMDMgLPuL1MCanTZJ3T/e+rWWLfvwBD0YPuYCg9pLU9hfxUFr0tGknw
36e7/qkfYwjOdkQk/sEb48UZ5U7Q/hfjknA6q0HsY0NsAYE1u+X4BX414Q3pAAXcalTu5tzNjS4V
UY2cqYu/w0v20Uu8yHvJir9W5y2MbjH5KIBNBgTB5CIfi+5M5Na1owZIH6xOkFW85Myr6rajjGf9
N/FBUm7hy9bEpXQ2P81REp+8WJvV4OkL2SJFaSTr1PYJdkLCy5S5M8GvwFoQgCBO3TisnQjnTB4O
3hWHLqkt3dmI28YxQOnOVc0JY0A2AnBJqbqDahlPU69ltPpB4s5xLZjs5nH6unIDyvjv7Y5urpI0
5j4ARcZwHa/10k2fQx30xSWo6sxugWs5yKnQ9VN7zCVr23eRwr8qSlCCfPT5myHy1PwDRk45kgVi
xXgL4SVj2BwXs/okZoWz47SpS0pxh9NONhudMLT7cbSaA/JaCUyhgIUWlyIfSFx10aauBDDR/OOC
Ehuh1lvGaTjQcah+Q6SbSvmlj42kL4BKRS0v6Z2G2VdjPJA0/0nmCDqlaMKpbRnmVyVNFgq+Fy0y
KjMXk7mELsT4gUt5FRc6LTNqpvMaOxypwkex/YkCD6XjyjwfezuGDpgl79Z17cCwNiVz0MwnekyB
1rDpaEW6cx/eOhHEhxRS/VobA0s6vN2+oQAaZaYY2l3NDcFKGwuiwe+TXAiPk8ByUrf+YFEflkvU
TAf/eHpPi93hE5BeqAnxiX8+zjfjetC25nwiLaG3fLxB+kGI8UMojIJ0uk04jy9pvAlyFcC+z7DI
1N7soX/SCX9vkst6d2S/DbkkrkJmWsB70QcUhmIYFDoeLdcLuLq9GD1cGVW/FG6g/Ybv+hiXoVqI
PMDZUaq7fh+rTmvFrRQg9EI4OUeUFHf5W/pTHhSCaPkE7dh6JoQYHHWllo2ijHnr9eZpQz+XqK6Y
NBnWvwxp2YmTAQQIOmfnW1VhoOUfCGv8jUeK+hs0yuqdeWFpFU0GqDG5p/WRQ9gg57XtjDpfORoQ
RlaUelYmBp0LfaHa5VlKhohQ7WihokW5XHZY8uTQ8EnZ1LUq1Kcs8jg9lmyZRZXxaUE+bp/ZGYPP
czM133qyMDZrj5hhF4oYTynG/EU62lSLO4lSpr61tdPYFESqmxiKWHw4bW3czSLfFPpfdzsYXoec
ZwU1+fv8E2Qyv90q1RV1oPkS7STNDERf/A04TJT+VuV7RceSk+fUx+LKsspPMablXP6SiZUtVDNy
TJeJpY6d5qO7o3uP2xjYtcymqIcsuXXrn6AQ8MK6T/Y0V0/ylfx2rRBYTWQPTjwco/vQyWDYsJb8
YKbDzLmpN8sf+IfC7pSyPFmaKu4wt4cnzuDzZtOzGCKN3xYqd7n0nEkNqxF3RtBM5j9lDokKyOA8
RaQsP3pSZ0rK3G1reENGE2pEpLJaDecNfJfiFdWF4gOYRnBD8QcedC0CTXI820NUJRGEkRvLSFcu
I2tsSd8n8TtPkIbHV964hYDqGbKQYEzs40mkWVZvMeBQb59URHh7S57PINWHr4lV3jbdohFLw1na
TQWGr6+GW/aZ3OORZMRmrebVMGnKS9n0OxzmPo167EjhcKIOEXd8r+hVhb2dQAX1MxvYF7aiuYtg
sd+S6L5XcmqgDJzRtRuvi4JzAQj2Zp7aTflDLq392XjdH/N7oSH01nblFL2wYHLYUavmNmbZGjev
rRoULgVDS00Auj7VriuXQxWw39oJfmAcb1yUEhDKqk1OUaOsQG8tvmukHUaIeYeFpIAitrokaLGZ
VIhEEQuISV6te4uJjdlF5qaK+DAdxIQVL/2QMAfhnxGu4Xbh2A5xisUkwLkR4H6itMNCvvA4hOQC
/OC9LKqea4kxMgY5U+e2yoO5i7erVhQ+YbJu+1TVEUKnr2h+OQqL0K5LxQL3/9OLcWcxt+QludOk
s1As2Vq4j7Fiz+SBB0n3tx9XNWKM5bymLX24E1s+xp2eI/NjeIAPaf/OGgKuHXVgAzXfJeld2nlg
Hthr3RAal0Cv4BNV4si/bwccSuKxU6ysF0oLCl33Hn2BUYOtEMtZFfpIySVkPFNcv7VpSKcJ2Veq
Ef9NmnxKVPRq4LrxaDpRw6UOITm0xl9gq5NFz08y7qmao9wcOOZZvpoUQfPayqW3QORK2ZNaRZDj
GFtF0EkM7h/xiupjpT8Zdd3C3KbTPoAhY3ISeY33rd2RBYm8xF+PxJ9yEDblw3tzid5Mdm/cFlNE
XNU4IvXyA/31z+oEnJi4MM2wFNora6YWc1tsKnnIgTSbp0bMz6A3ErG9EvZcpj81LK/TTE6Ch31h
U7PdAWFa7ObsMmx1eSQZHQIfKOPsJE0WOrEmGO4dXnK/ooP2fIyZf6/zZ7FWHe9IXFpgU247R5ZT
L9vRozo8hHC0AnyCl6pBZwbkGEVWg9jzDbmElz9VWWguXDzP+ef1/oqr4i0PC63JJgwcG1U4NjFO
4zlUTFSLecu92vrKQXgLoTkRKe1q912Eqstg7WiHcotTlfWM9+jvF861639LPy+nhsVhf1mymRw2
gHat8CccHwR3rJuq6+HK5+DzogYXgOIUPwUBrspt1Sum9oqpHWd5qi4sElXtZt1fdBvb1E97BAmp
fxqTCUWFAD+5+KvNxHL8YLjXHUTAXCn/9AsDeNLh/UV3tIPiFpHsQjBm5i2HVL2+hU/iOGIa3bgE
Wf6t+e7Up4c/elcaMWXBu/Wtmn8oQsOgBgNmb7GD3uctFDVu5a+D19W52TFRbSeXLnb0W6nGxTUe
A3vpWyvJWpf+sT9nxwuXoba7Ib82oghMlauHynhZTWPe0o0ms3YHO7LYEI+/OBerGweKu4fk2XZZ
kc/EJibi8uE3Zjl+GeEU5HDmxlmrWaJ8dBpmUtoXxD6DZ23OKzxyMdPaknPgTTCLae03g5lrtW23
PqdjGKeGa35bksop//kTlpKXG6gNC7/XZIOhT0twAt16d8z3yEsMH/MSi72obDUOI6JSjbARUGsk
01mOHdwJsS37Xp7wgDkdPX9AArXa9hTyinuUdd0AGFF74kVD1UWWcC3LvPWRw7XZLkG6b/eNHOjk
kQN0gUl055hDJPg+P/idyLl6RQ/oJzkO2CXf9MhHi9Pw6iQVDMOnRphONqsPiUpRpi/pnC2wbklo
IA6yBVuBjiQ3Lfrgve4HqRBoqEZtmrlNL3Rs9hrmAunx9n6QS0k64bmM4w+mVVza7QISC3cwJ3Ql
lJy7yYLhJX5e3Mr/3ldD1frYKXuZCheFPr2y1crGAZO2GyHrY6xpeG0q7fygptK0urzptdsk5ISG
T+6e70dspFmYbCfTU4xwo7WdYRAVwcPY0dlOFd7etZOEKXAE5J1cycca+BBOeSpwvzaVGeIg940I
QiVSSxhxri8n0bBf/zSLQKzfw4dxSVgKqCc+yh4xrUCp7aVI5bW6R/DFcoqx9ONGBmSmRHR/J5uv
nYD9ai3496VdE6bbv4wpcKQB1j7DTjnZehj0BUiWaC9ojG8rKqvgL6MTTjLXCX8dbWWzVUBNR8/e
dFt/9wournrrdGrJjI5quPoB+D/MWD5Au3fkXJSSSRDofI5FyfulPQn6lZi9MH2O0JCLHDwiveqB
fWZBsEkjsjolonkCi/gDsQT2hLm7XSmYVCnbJOy290sYxDhziHL6vuwioxft3wuwUfQVZPtpuzLl
M17IxCSilDTr9KCMtQRrPsmnWkAgajeibSK1tx0ynnFtSLzIUGCGiYd4nxJxTC8fU85Dhxav+ZmP
Tyaxnz+LF3Z1njj7cKJnx2qjYgHD3kWK5kb1PUWyw9uh8YYxwGNl9roGfsUZ+fwBSGZH4hgNsj74
m12zmN/Y7cLyDzay3FkYxVbT7VX0LZb6wTD5jFep46w28OlG71UbVT2WTWHYp9cM6UWhACzwEEbC
XH8A84JYeR7VKgbIXtcDUQS/UDDXei/18kQJzay2WMhHKJkPN6mkCSoHQvgiULA/Nny383JRczv7
vdVway59RS9OpkbSOUMgbejnrSCqCQrP8+5bfOGOPmbVEnJEMsypzbg3AK3u8mBNaQxDIddSYrob
o3MV85V7b/KgL2zf0Uis0ZIi3XXL/H8kXHQl/7ljRz+RJRhWu6xsdTt6TEysVraYEHpxDBucv2ib
ayRvH60va4tFCagETyTA1COwHSSiwjyUqN4oPbrL4grZJsC14fK6YNt0k1lzrrM1xwjiqQ96QMcg
ky2ab8dAsuqIKRBJxujHYY/ewy1u2gp7WJALAYpebsfaynSI2uv3u6G8RbVrNpVrEHyajnXK4TKI
GUcIX+++k+aKAOCj7KpK3wzvuY0ltlkpHDrI0DfLvdBAlXCHso2YAXFyR7fmnjfUuyAr6vCQWwwP
FWI0PVZEZkJI+jCQG24APd7OwwWD9ujmSp3vxRIp35Tg1XYxZfxef2UcrhxXGnhKrNXkG2Q3kxAs
I6Idb/kpy4WCGuiTV90o9jDFLIteXvmUQWgQvEgeneL3avlMBNAiVJa1UF/PqCyivAGDGP6EW98v
OS+llVEg3Z2+G4gWXNorHrnZhJxUpuAFAWxFd6jiWAJYefKHVJuB4UjQAHmmn4eItTAF5GVMvGFL
YMbxH5/8XyxQqc5SrCQ9vyoqRXXv6+5D+G+Rpxag5K/re7j0VtZjH1G8scR6r+WnR52pfxtdwt3f
QBFSjTfFgDNGcK9I3DA64suXLHbFS5modonQ7q/T1r9JxzDp0gRiFmKSE6hjH9C69cQLQyQnSPPy
3Hs8eRZU9rDX47nt23ZLa93q5jQAaUeyvkmt5zmVeWkm3e62GeFl3DrtKi+F2I1gfeumHpurjcyI
fuwM5SZIcPmquM9MTZd1rVWIegM5V+nB2SO9Qlc3dCXuLhLV1hAgxZRiQLujXl2izjMJdM/51stD
HQvIUktdhDSSBljay83QA9QKJjLSeeio6cnmtlHhywheqe3w/JVFfRWvM8KmKI1GZ8txw2wMeFbz
ZDt6bEc5MOFjJRIN1NxtXMyqJNBEsiqOK7ekn5pda6t9S9MjlAJA6IsiUoDAbN0BVQK3/YSCaxhc
RympF7xc+ryc4201k7vyvZVeswgFWS0scJMngSXx53hR5aK/atIKg8c5xH9xiV/x1jD/GluIVobh
VLHE+FjM70vu8n74zEq5+wytw2cnrXfEGOiUBPLoJ/o2NMmPtGpIS2GT0ID0/Ws2XkmyBdkd7bSH
uH/0rNBpoH/KZCywGXDqSaiGsIeQ3DFgnMaKZkewcNNStaF7Koxpin7AWnd5ob5fxemhLMGQhQlQ
BIu1T91+m1tLgtemNVYw/S319NCftC9xtPLQQT1dLH0GOxjUvx/41tYSh39Bm5WUNBU3mb8N1zrd
u+2U6lphd16LznqSiA2FL5yTBHTHSid/44IsSs6hzFPk9Zjlh29eHl5/vbs0DeDxRhMJICjlJl8r
qnl5GyleSmJq4IiLrTq5T+4W5IuTtUnbQaNII3+L+tAHL4ZJWK5g0abaQACifCpsBTLj6bnHqMkW
KGDfP09elNx0lzHB+jupL2f5/rJYKkAG26XYetIb3o0fM+KEDQ+Z7b6/hT8Kbwj6MYWdhsT6H+md
8iClIHNI7ujZrU6/XVNd6YgtN5UWUG+8Zp/SVvap4HiK1t4kRBknpq2o3kh70Rn9YtEE27aCoEWK
X6yXJzEBUY7dAq8hjNYuPRUv7D1DwUDt9c7v8Jto0k1KIQTnA+Nhgc9xwSxbvK4UvbkGTysmbwmR
RsHag0uuRtGH5Apk3MVokWAt3rPGCf9Eh8FQErhP9rVfLtxocUggEMkneqPmnnp8QRn6SAek1R3e
xZFtWCZsBR+Q2K8ZssyVM2+XnSQ2w5QRLHs7Tt5lO9EDAF3obSbu5Vbd1tWnjjQD9oYUatj12DS8
mMGpLlWmDFdX2UHVLqbyXRD1flSkzC0ghBh5f9hOD/N671mWdqs/JhKEtt1GF4UL48waEdkSQCo5
cA5s9foTlhq7mUiAhB7cBUVWVejeGSpE+odAJTnwdnTEtVi+xyNk/TYoCYtjlgcqBhdkDTiRxTbF
gt8EtHMottp8+pwugXru0V3VlK9R4E12XbmYnHZk+fKsH5JyZmyFxXA1OPlLQLSMwtS2R7EU9mCN
lEN4xGJ9M79n9w6NVhTye61jFTZ1cqeHxhhzsK7xX1clmH6H1ZowunbFCoaJawUtyrv+NAbNEWbW
FTaMlGCkC5qkk8tZHgEo80Jv4p5Dz86wH6+qVkLludrApx7Q770xcG3QFfYPs1ggohJs5Vfnf3Ji
i4D/OHn70tjqGW/KE7GrPpc8bwGBr1KgF18mEiWj1XP2ZTYxiscYOnUKV7dtTYVmiyfjFOsFi2TM
P9koCd0AYSUZKWDV6r+wAybLj5+dF/TTPOvmsQy2F/puuU9NyhClMEtFfx68Th/tEZIHXDOk+nVC
1TsbtjvOKa/MD0fkAFAgBgtSKksqhnwxcX6PAG0VJ1xK23G95SmybXQubnfNgb56uom/uf7iyKRC
aaMUxegzJlbWMSUjPDtl85LtV8CJv+P6CDJRTcJMBBiyPA5/jMZi/B1OTBeS7ESZ1ymQtkCmkJ6g
OiLsxFuf499vtJJsizbKJpvIRYMbJoOfVz0WB2qInuRGaor3KkSn3W4qL5F6G3Nb7ENAJ2TXVmUB
DHSMsAxOPsKjVzn2fA7xpV9zKyJ7V33trXLzd8I3u/8+1T2twsgbm3VY2PQul1alMH868uGJ/7MB
zR1vqzrtKBh+tjc2U+txsI0AKe2iti+gG6CT/mMKjpbd1ESx8XFF5It8SOX482p67TNiGzBwPN+o
6kKbD3/IxmuydShUztrf/zJgjYnzbWPa7XJSjC48LrzRYGpy+jMnTiwduEyTQiF/noMqLBiRYZ2U
SOao8Or1lIQOmb79Um+dsGRUdPwCKkTgpNklxW7uYWV73YN7pa8XS7/TAytspYuUEQbFJcTxuRsy
iFQHjmS/H9dM/dfZd/C4ytVeqxTwktNEwhzCtaT95bzFLtrnp73O/63catkzOIJSwHCUUjEkWF1f
8EiKO6CFdHQ2Wj4GFEXVZIpTRG4Bkre2l+rEkuPwX21J3q0xcoeKRZuBE+FtmCB+DYwo6bDidNSk
pDmlt9vY/Z33X47aDyQS/hHN+TfiHvKbwyUu/YOCB4oI1U0YyiiEiNBuXwRXfi0aL1vIDVizgRjJ
qGulHj7G42DmPzhphTeH9f1PwyaQvx37Qi4DUdrWSKVJ1q4XA0T7+t28EIXrwd2B4X9Doeqw7v+j
WC7x12TPLLh1l2Qmw8cC5Dm0NDCvYBeakqvrDptisBFnYffbE5kMvkoUTTr/pfut8YjZsXmgD+f2
aw9ro8BUw31hOdne2i2D1yl67qqA4LEEmHGNzA6zyyoFymqHw/is+LqmbXCVLyVUPPUF8N9+j+Kr
VFZTLiVVRaCPU3yM+nsPkGFM37xqUjgamAhyIZ94AWNgmZzaNBzBq32IWl2PQe2QaTA6kf5CUvuw
oUaFqsz+n2zQgbFqaHaJ/a0zHWM0ZRaUfuTQyKk/muCy3qG+4ifBYf6hqCSoRo7eVG0YcQ9kpBE8
DlTThpTGunsFMB1ySDDchcfIFH9jLMOLPbUeRIZexdLq/T0xgiuHWqa1TjUjy1nBD44s/B6oWraJ
FxP5JFPnU81Po7XY9ykupTfHHehVoUvJfsZLKt+61F7FY7IlFTH2g95a5+J0bWFYzdrSicUwAREA
GXnBGzrDPHZ9gvCuNSZhAJWSL8+NjDsxsj7BgfB8IVF44n1ktkVfVFADK3MU8YB/1175xI2hLHsr
nrJZdVdQXmIPUzy+yztFheQS0v6M++qva0ZzFiZbn1x16dhthWFZjLQ0lNWJHCrabWcy7qW9+9Cw
Q/LDJWfud1btK6O3ojgPsl2bXRbeX0FtNWJQlApp2lcMuHIStlpCyeC9exxL16AEAuQwyn46/S5W
ANHKzCSpnW2L4rIONUqLTpod5DUqQ8kESDit7dIMwgbKGtytn1AZoma+7bpGQLuvryxxNflgDFM4
W75Ba49sNj2wDhOnjnEO6v5WThkkFzBjhpsv5n725XIVg/G8ZGMxSeRr938WBm8Lvg06TiuoMfcg
uYyZ8wu3J+QTHUh/k5X9/zdW0ypFcKV9BURA3EtdTxB9cBEqdvO5Dll72UXjanwqUEgtdso6saof
sJmJ4EuoDQzikfY2Nk4DwadvfU+bt/wsd6N1dTKy+mPEZ5DvnobQqTkmAsy/gpdJkMOoDV29PMsp
eyLKFtA2JEI8XLTpeYFdE6RkRh5tXGKdYVRtm2wV8X8Azr0lW31TeNq0iW/oATm6MPVG9FND8biD
ytWeU080UE72os5rqA67fMRnPOZxP5RkaFpdvuUVcVnNk4JhF6B1038PS9/BG6kWVdLI9oBOMc+N
Q83pQTcxdokxU5RO0FJGuT/fZGE4Whoyz1g/ExehHPTlFtr63Zj/pAL2LsZgk5OjxBz/f/hpXB4w
en1Nn3mWFGTot/P2ZvPAS679pedHXJzcCPNDwTQfflz6reIlRj0mA9WJJ4EaOYq8Zv9hLto+CnOz
yJr3PXnfz7cHmXx+MjQ2L/hq0jLbkKHgZwLWA5RXcinX9XU47jmgLj8n7ADNo25isPJd0LzbfXPp
1sM6/ZOiIbEfY+QTW2DFTKxCEwyHxLgsrQsRGV9vjlD6NNRg5dd2cuMiyfZWuwgm5GeVfpohQp+B
jfJ5+diL9ZsDr7AACqeu0JHofZK7r9Ry0TQRe9MnraCfcgxZjOSixDznpcIl1mmfrJ/gDXSkUEvl
LaF79uMwLRG9ZQxsSE05kNqdkqgp1y34apPuLG/S1Kop4fwpmEx2NsUFrrgTy0rlX1BMA4ex6yM5
qGI4jVmebbLFF/4Q0sM1whmNStMzXxwbC5oJ4NjRMFhWdaXabvqhZrkYrBlzISWfv5auPPD+tI9V
y2XIi6tiMJipcusf6iN86u4ENblgoCMscDQptCc/GP/XDQnSt4+jc86GL4wZIKwUsxIeD/aIPSqD
CwiFmwiVcpe/7y+xCORLcwFtO6w9WUPcUhfKP0FD/ZUhqBSM81UIbZpR78f43uwilJeC55dTmJ2S
6+bzNZu+nXH8xzRKVz4V/OnApyO1iCdbN11EWGD4UJCV3rkDzE+P9iflXAKKS/vIZ/ZWnUTfjOuz
vNLvRH6ZAI9JaOFEWERxfFoZ27RRYY/qoGycB25FwUhVShjtd7JXav68xOxq6ljMkeYnYi3qa94f
pr8zqFy5w2e9/VL5s82yaZPADIisqhnIvfMACVxEQ/Q9IjmBqtX3+yAgvgIAEOXqGMkgv5PF6dMc
p0LKDKdidk5urNSmMqiBOPYHUPQdwXid+sQXbF5a9W6F1lalePIr9/JtqEwwFjZyPDvSBfFTZafs
mbclWoqb9R0nMfTXfYtPVQQGpF2OwRz07eZduUSNpvCAha2/2+buCkeZgVY2RKL76b92e5OqW04w
F7rQZxB7HXVaYD+lSOPZYT7/T7wk0sVTkffrFvkEpuhUkoUInGr/GpQLrfMTEGic7eWO+vFjepiT
aiLvJyqBxQP5EmKz8eS97g76+u62XiRpVQiF/nMiBE3C+SeQPdSy5PIXkqTg8YfRWXqD4I+BCGtK
CMuXennBk0ovU1sBO9xZbd3ISVhIyVJyuMeKjS7KI6UH+kvXbjnx/JcKvU+9kz7NxYNlfbx96BSO
5xh1Vpqh1Snla/N6dHzG1Zfy5IjiNiTAvxB1HUkEVPq1nPn6i6YMyReMME7xoFDFvaRoYjd8i/wt
xmxtsQd2IwvOsiPl4ub1YumT6MrxyUlhiMWqvCygDwbHSMXb4tODorossuo+FLJGAwrv4mAPN2Wt
n1YG185zb28Qg+fcEMmHdPJGobvgQx8JlfJ/67eN7H39GBx/H1riYSf2PbVuF2+uc1/IDa3hjO9m
wQQFsy7Zoyr4W7ae4fLycmDL39KhDzOaC/8l3tEEuN8Eu1YjeiVD5doAjDu/sPC28X2gZIzdqHvV
DbanLckhC9i6kKKGj0lsRi0wE3MbkWzmIO7Ph6Um8PXDYqJ/2njFneSwSc/qfWUPteEDBnpbtchh
M9e+smHZFsls0ioxo7d3pp1raGtcUClNnaJiPtM6CW2FouGjrejiAe4BstlbgsGUscHi+IzxK7nS
DrhGJiqCDQS2+aaxbjU7tQJpJS9Tal4vk/cMXU/vnwV/+5jTHBXEcNAIX2VYR5kGeusj+HR4Ffin
QEd6ApRDsb9aPgtbeCGM9IECstddtKHixweoKFXU0w7bE5jQK/bnFAuN77mhsgBpl2Y6eT9+47U5
901i9Ism1KcqCNxw+Jy1UE4CmFcmLYeS1UYleSkAQR0l7kUO6qJWEGG7l8OCygfF782YI3pA3D2P
IsDKFKAh3USNJy8WZYnaSYfI4mZLO33EFsFgLDPGwR3x4mvQ7lpYWBGcGw0++xpCfBHV6etqpa97
F7Xv3es0NKFRnTQW0HOEpUUatK306wQnC9apLpVLJwZeeobPdRtZMIodcp7mtdSjz87bb6HmxjfE
WxCUBNgMxiGjGkMyh9IUY1LrfXv2rmLuRzgeT3ce3Rq584P2ECNBNEOTY0d8VOOSD0zkLaUCI1T4
up1C6oD0GqIRx9TitaxxyJ+RGSsJguyeplx1rRTy69rfvY2rJqP+MmthP8ia+danOf2oXADQXzs7
yUQ32+DS1xo3j5OS0gjfOUJFYAbPOmcV91K3FJSZcdwMaoP336kX55Ase16xK6mcAYFRhkkJJCOB
WliwklCswJ1nXOTzR2E6gQJuYRdJpTnTXs7ol1BA/MYH/2GV+enelXM6Q6SStwwqhpOApA7fz/y5
8LMkWMBy7iF/yFRe55FhIyUDLuC+Rty6H5m1iri3Mhflw3ZwiX1SpxBozmoFrKtUE5dI7CgXqiyS
t9mwgT0rxApRSpMxiiu/A1q1uFpoQOWoSwKlV3Rt606NaRCkwDasJZJJe4wSz+h2H4tOW2jiQzx8
75/O+3JFnE1HQriwarnRJRMBNHkxVDvWsDPPbGF97yW2GctutYiGCaDd5qq3csGa0YhlobCLbct4
a8Jg4sNb4yoHab5dh1f/CuAw9stFT5+kGsNOLTdiQT7Ipp0E0TvruvGuY4dPUwomW5/RRUdjg2K2
T2edyCx/tFkE6jW4H0vE4g6orsZDDI++zhu5FvAbfnbR8ioPNrkJPSwkSa4ifYJxIx0L1IXqe4oG
5Z/NA2C0bD/7uenEpHjPjqetwZJwh34LQY6zaJ5CdCZPVdJCGxcZYSJQzyc3e3AwEkFpfxPROgIG
okz22xBbAdRwFRbinRJMPE/nDT+40iowodWyDo6Pu/g0sgbU9AciXPdvrbAmXCDBad8IdCcsN4lG
oVgYLhlzRMiJ4D0WO8izEsiZJvBq5FpP8y1M4kADAf6qWMlWLI5SQLvDpdSV5V+uaGd/PLyYYHWn
G1svxsV4g8s6DUuZm4axNy+2eq2sReXI/ixwUCPJIVVFlzeXtSoj9shzgoFa8BSo3XLooPPbswVg
YK3x6UhFdNuQnvSq/fn8QKSqGgMPgTg5H/+hjMPEYE+O0Pg1LCzpxjI7N9g47R0JLSLcHsuKSC9P
XcvX6j8kizH5z+nGggesI9owUc5ZKe0lfM/ExwdGMC8o3SBUlFhCBg8iAqX7BJqC0S5l1XnvChNA
ML+cEQwV1SB7AKRhNhXZFh187BXJWeHENz59YtaQu6O8+QAAvK9ynCEJE9s/oeSe43PrrUa0Q595
QbzOQI1w7xR/f+xCO2J1szmEnWPIjhq+PSV7KuWxDYTYS34hMzg8V7LRUKj+WihMUugDpheizTpA
PQcSGWYsmco6aRz5ECswBAB9Cq2y0fXbttHD8GIHRaE/yF8ScBnHpSfYzW/tevqW59+SVoCwNnlJ
9AIQheEuFiy2/5B7O9Kdn2v4wGF7HQyBYXlODz4lxCwDk+T+pfAZV0jfPwmTu0O4WbeJUadNmzcn
n1AYj28MndUpubczQn024udSYHiGsL1weY3Sg8dlT1ub8ScAJMIZwBJ6okKMYd8KaoeZRbQO1/CN
v+6kyWDZ3Ei/ct69BmekE9eioozacBizg68YSqatAK5F5nH0HExhZpgmgmAAQ3/lOug5QwHFLPMD
ZO72GDVyLGw5Wf2uB++Em7QVf2GAiFlYpW6bgR6TLlW6rrRQ+jbM0YDG8BEc7Qx161XiOrsqABhp
R+mrXxeOYNYX4RX/tbN/uTiFr9wtnvZ/1OiIBRxhIBZ2q+G3VvAUQWibqNr07nDAPSMb6ZCkTIPo
OXCoop4BAzvHK2wRhbh9fXPgMJetk881Gl6I6+SgTl1yXCsE6SG21UEiu06VdXoJkheiyDF3cVTJ
BN+zq7TFhQnPgva7/E+ss0wtJp2d9rhVeupsHTMp4XiL34BfY/9GwFd2z1bsTSs7MFcJ9THZFMBL
DyaFY8BF0eSRqENkf+HC2P6CrN7Tnb9MgO3SDdVpbKLaIfJMsSz0UgCa/zNCMu5OxqwQqHsiQQrs
krlzTRt7I3/jwWxqW5r7lj5x7uj8S146D+zME4GSvBLXjl+H4XA9PeOKTh3SSVhtwqbn6zljgSG3
9XMb0PHuxehXw9yb3lXCshD3xPKxFNdObV3fNgwrxRVmuWoSmT22cYa9wi2UmDn8Fhzs3seA+rtQ
a9kq+niLz6fLRXSI9y7JLIUxuDkdZq0JbbNLXE8X1qwJmwhsZsubj9PxJn0gjyodBAU/SFyCerL+
ZM3YaO92YkJLvNHJk4+MEa+KvXuxOtENRRqGt2hJIxqPLWd4EvKTBBCUp+36YpaZOIn6o14Rt9IV
K/+aja6s++lUFAxCqv2BnCBLxZnIAdc2wvW/1MgN5ICSMi9+GEn3gib3ds7p0R/nM7AVfaQQWn0R
GCoKtM7j+xJSUlx7TF80FnTt5xINVkArgc9GfuGdQzinPurkCWP06hQETxSX2DS+sxV58HiyyzRt
FFAJ/SZpsGKUdrsEDhXBVlsPMwMV0EJUi65/hD6a2WPs7C5s0rYhnR3dD7TwbWJUEmgnpQkyAdU6
k+twKp2y/KIRScPa1vtv3uV6+ASAA8zvnfMAYaok9Jm7TuXQ9gJiN7VKWIbgHA0bOcCYaPDtP6Fl
pDuaMiQzTYVMz+jbx/VK3SMjWDrUclBr2ed/U1+BTnRO0vxMrczSF3PIJ0Pu5tlghY51010Q0HUS
IwxZtHzpQ7sbiSS2jQ/tNnXaoNM7d5DxLPsAmRZ3Frfmbcb89KdRmMGygJCdFPx9n5/pPg5C+pdj
w4qGwqFtLLjIMjnc5bJoV+GluTsxIjhthH5eyxy11B1KOJcF5e+h0e756O8KvExpU+2tBaDq6OOt
wZ3WqPP/s+A9FKZyhm3pXdXp3XmmcbSSNY9VDA82rWpimK+hEfGkx63Jyoz9asCvunyAZ7KBleDn
079KYhcTLt7awQYJDcd1rfpFHw0d01IQI2/LC1T87lFkE/I8Bqo3h3LPosTyvoPiO0NG1SGPhCmh
kvz0x58TTltQGYhUevv6YRERhLiRfxae25Kg7Eo4Wae5ITMxTG8vW6Qw9/YXAmjxaNaMQsbudp8E
Qx/jy8LQjdcXot07B98Ya9qdRmGf4Wn4LZPt0U8he8IuKqBnwwZ25Kc03nO+0TYHyxMiqkbtBFhs
+JcR7OVGsH1l4hL7HdmuYwkfp4T30O5qLpmo7Zyow+HAVCtTYwuy3BrBJhaD2cZ9NdGkMoSFiz5N
bPGBXIeuYw0tLIei5fu8Vnc7Xe9LLucrGF8FokG4Urg7Dz7EJiq2Ln7cc/8jG1dK8ummCfjf5BR1
+yzmbog2uEz7B9s7y7nMqzIbtJdmxO3KmIPU1ShxvqjflKty675SzN6QEQZsr7chlPaBJ8py1TlO
ote1ffAK0UFldIHSOgMrBuLzWihIDXpCwxmycfuND1o08be0AZmsD2caaDGP7uzpu8KPXQIaE18a
3Q/uVWI74wThrDzZxewpbdMycrFTEhwtF6X2CP3Hj1ssc0jHKsndynLrB2nwvyH32Hd5MgbGoRY2
6RLtSPT+dIpGhsFvkT7lJKSNG1JE8PIhGx3Ie+qKl4SdvlVoasMBwlTHP/SKl8UKXKTZa7Si3mWh
3ZB1vjtp/NoLvMqSbF4iokpvso9AwP3c4+U/kUr0gg0dVlrVhh2ym40VKKSWPcagClpX/mdxMpMN
HXC9QrhyfDVg0UIId+zxKB1QM5R5/k941BEn1lFLU5W+y/yGwpqRk6LqKF/O5Un2/H205wIz5b3Z
RYHxY77i7xkCJi13Eabdy4B6/8clpWdEpghNpeC3lxLlZebr9WmNwFodfs3tsNDQLpYrFcqaWdbu
SVF84ugxe/apj91PYhAF1PtO8Cs/xaAV6HTSBAFosYw4jScEkaVtl/hvuymY0WyOJ4u+r0rNa8nd
H6khXGTG32+/zVFA8i0KdC4yNeWN228JeleTEVWYU70G7aom+hZp4G4h72Lxlgvm4yO1aI5XtwG6
cgAOTUlZO+aKqtab5j8blwvivBfPKoDlEli/sw9AZYPmelGbrE9u2SVPuTlh/TJTftg/lCz2eyag
FwovThGUl0JaFb4BWLD4loUA3yeZfIsI/EACvcOhlpbjReBiMkzf/RWGwiuXAmMik7tf32gvrdGo
Urtuco75zGNvxoowu69Gjkm9Eal3zKbCNvPa4BdAsJj0so9BYgimp2JG6dxYhmsc5MSAGuqnRCc/
AZR1QqiqeG/uro0ulCgM+ILAfnQsG4e0XEpt47lOQ0P5GHtlvpws66iw2N0Ul1JmffHgQOtTdxMq
BIHIoRYGwIwEaA/YbejJ03blfaCjPgcCAo1PtI1485/haKTP0Gi+3qNCgrhDSYe/Prcm/iXUeSHO
fUjgHP+0pFnWScC1aY8xmflAHEvrCFUPjWZ0vqpFPgk8AvyubpurfQA4OOWxVyc+Nkvf6ItpJwnt
qyMUEfbSFZ9+DVoAJv1T9jMqI8TBH5BdzOiJ59dROMPSVVTs6oLDWwM1dFt3d2UyaQj3rKpARiDR
xmA3rYp4GIcAglPuX2MlaGlFNFwArJJtM0CsC6TCkun+W53dd5ro2MIobIlAl/VkKalHLjHdv6cG
88qDiEOX12OCyIKtDLUJo2MKY7vFHg2DhsNJQuT97z2CHpRLiJ47xjWUqTxPvA+X8kELH+BIxZ6F
XnIpZDKwe4lA3rvqgbyKPY0cIQtTkj+zfaQaR1e+9AJy49bKbGy2sLmmb3So+lr/lW2JZ1+6toLr
5C+slkDjMpZNK1v7men0Yj7CqWDGm3zMNYCKZo0tKYBhP29/5Kn8G1olfejeMSSRJtPQajAuobjG
MJy6T/eoDfZYDHnEaAwyZQKmod+PWblTHe+FKXJ31kFk4ZfN6vKDD6WrmwA0qgSjC/evUjIlMRxY
QB/yVA/z5cvsW4gkon7vafRhFK63IFABRL/JT9ZixOm9prOSomtohMOEdi2oiyUcvptjxBtuHIHK
BVQ84cUROQK4LULQ0qurefHbTlMoAmL7OtcIMfQuIexd76uAh7q/BR86kuLItnvNQScgMJDuZ982
4IdHGLLgpVdR9jwO1PooKNwVAxBbBctduFjylqvqvE++f54UvfDeUVFgi8kDo9xghgFWXxhrRkhx
rDx2VNr7U66PySXlKne+3z3k0S2KYnoFy/WsdjuTibaXYaItLdbFKaCZH1mnmqSUXRmExf95bHnr
6V0rQhgUZGFp6SKZHoLjMiE18ZkVTn5+zLN5S36Dc8h2mSz8sxo2gy7PNNr9h/e12rs23Uyv004y
cHXrGtYJ2O9tkXFQd2Ea9NdKKYsd1nSgBQJkXuEYxII6H0y7CTJDikWxtadPmNdvctL1me8pZ5M6
OvkAKEsS4c3qkcCDqLVRftXErRC57NSqQbdHEYXYYJDBVZwzM2aoCzApzJ3m/UMJPegiDTA1gm8H
Sf0dHOvT61T2KY6afe2Bj097An1ja96MDKxG3j73rICJsxnddLaTMJHZYIikMCuXCcuMRqJgObAm
wJKt3SsY3UOMxkqUJw1enw4qUUYRToLu7j5pLRAABNSMfDymJO/JfEEUKhWNqNkLQ3BI1hxDlV3w
JmngoicQu9cw7gSB8rcf+KOb+Y0AM5cxEHs4qtMGiCfjFYqPKn38E9stn5y9Cc9h6Btp+usu3ojO
6uESEWNm5thaYrsckMa63IJD0j76ptiewmelFBvMGjTx1vh891Y/fMazTKVNZlJssbs6CPoU4Fpl
xsxHKUKtMmHPtbZr77RW1sr8LnACwAd8SCVisQVdDwJh7LMKsLhqoBCwMblRpTwVVbJWVjM4Yez0
KkyuUwcoRvOSEN8yufVaJ6J0Jvnkg56f69Fur6k0bygw+g+mn8Dduogsp/Cj9cMz2BdYeHWj6SGe
E4KUqW9f3Wcd/SQEqgyWwoN2EaR27l3Rxk4VF5HP5+JC9xFyQWU3KqP/aOnzYr2fN0kzXoM+dttx
UZgcL20/HT1tzx+ZyBlhWU2l0n3/AI81dWedkyF5KR6Yx59HYa9m976v1GhH4SzDhS/nKw9LsIHr
clFPKgVocbq03mKvcwb/dpD4cQgmD9S9JSorS12nIsJHdMkUeNoLsdBDSA+hjHwJXH541kf5yTc4
ChxIOSu78YbpW0RHXkNI3ymXfhKve8CbPm9Y5GrNx9QPvtxhSjrbeIEw/ry8DpQ0BZmrCnex8lph
6sJ9zWXa14I2qEjVWdwzRPA5wXRBl64MpsXyj8ChMuwV7XZznXOjKuuvpNdUG92e1YRmoNOI4ip3
Xni8OuzLKd4kzAtcwgvlO0u6omPqPy29Lut02FfOe3gOQ2IaATxR+BSX9BeyNNMZnqsZha1JyTYF
Hyl5Nxd4nsMBKvHM+ICshyCLGjsejpI1o559CuYYm2oCbKbqwtXZwwh/503cX1O8CJJfWHmLX6Ou
UCfLclu3fN7JlDAFeyfUVPUZxOVYYCE+ay7ML4//S7waFKtz2/SyfyRsEOqWGdikvRXnJ0CoqAxR
/EEqZLCh+442ypOzgqpak4xsugUl5nr1v+sDwjnIDf8LEYQ5/zp8YenH5spVBIL0n8gRS5hhhjL5
5r+pHvj6KRBsgJFMQoZ9/Igln4Hxgq1iE0vLQzj9e5gOfnPUrNCIjtK36ihhTR+HPRqvT3Q+DehZ
sjiTbbmp/FFZ9arzB+37rt64bcvT+HAusEqjBdel3w5FQ0UUFNoyISx7Ms102KYU9RnurLnn1uoF
+Jq6WF3RhTvRAFHey3jdLkbfZkY/iNhHCse2GabWTaOO1rDYEee4iahPKXZQl3+Kg8J2b1Tc+yVC
tiCWZHcNT8uQkQ0n2CnYYe+pKpCbFaLJEj2aZ8fbk36NBBbzBuWuBFoyJ7A3jKA9R8mA8Qt++tWt
sROu20bVM4D0fq2I4koceRHyv/UsLuN9ZGe7hjENSCisYd4oCHEZdj6dRgrkpt9xzbokP9XsLzQ6
VOZqvuW7Yzn94K4qDsY/KwJckKplv0QSGc4yvGiXRX5IOKS7jOKrDYNeyO6ZmzkNZh+LvC0TVv73
JaC6NqcselWJ50pD5l8ulB58dy1Jccek4X8uE1hThuqb6MBn+wq/yyLmyU+S0FJaKb0sMzuG7fCO
HyIr61QjRS/t4Df6TQnvu7Z/w/WaQGijhEjnxfnzRPY6vVFqOFR/72l/pauk93U+YUCidOT5OnAH
3dMd73ZjkLPjeMErJAKlugdXQh8ck8Z8+oYfLiKglUY5fhogAIehi+GYz8cBpXr4jfJVvpid4s3G
JNJHt2C3HdRtLqLMZBOZ+tlcWNrWTeg9R5wDEnXY9RxDIySPVJ3wJeEgrfJPxfvcr+8AWZUybIJk
LeynWc7zFEcKTyDyuxCfwOcYx+V0yLRv3j4ekJIEE0FK1cEC+gFzwqVIIJ6WFaZFvtwL957Rv0k9
6SOwowl9F5TeZKT9su/4TqbnG5AsSzJlImcPOSrHyuFK0V9MdWBnNs3LdKHCouZnLU5azu7Hbq75
g4F9YBnetN4oQTNFPa5PSey19tEGTGdZyOD6eNvM0WVn7eYxYkZh1l0nZRKW4AJCv+eTb06nzTMT
aQVsLhKa6g8hP0TpLd/a3k6hTmF4n6BBv5ZvGTnjFyT1oE0EOMEDMmuPo8zFWYSqBS1Qc3q6UZcn
2hJIyjcWaDGf6vHbZcOqNpzTdWZkFfBAZEBh5xKheKSE8A+aZ2DsD2a4w8++U+U1IBxgIHeyadBM
5UiPOUpidI3vOy7D9vEmLUsf8LUqMlwm/pYEVkkGQsOhjdBPw3NO2tWZC4YDNP1lW6UcC+k9g+5L
2umUSlNGAz7jlunlngpf729k2QxwmAIrkyVzaAgS66N7D4dL8ZNBlYFIjs79Kaz9sA8a0JeLf7hZ
yzfUIajb9IMPuGivsR8i/oMA3SHJAz0aI+FaLb8tHN8RI6YehDsKsERKgDNJCCXrQE6ZrWP6W883
spt9uoiD0fDSvreAQrpzrsfgD3sZq4BePcM4wPTJ3tdKIimwvZ/k9Wx4ukGbfOApBKGBbZNllYMO
L1iM50AZPrDZNfZrqqPEbN6Wu9cyGpDs+mEeL66kckH0vqoIglZdevl1RHgTL8ZY+NAnSxn9TGhj
T9kVj31HSw/hszdylj3FBBDz7TDJWidUrCbf/3ixP9hbBX/3cMPUU5gs8es6FUSgmw6yowndz8TU
gCbYB0KkJBuGGPmFGEceycp2hQ3/0QbD5IBgTvp4E282686ylxWZfUmEIywsnHg+80IYSlS8wSQc
mGXGoKrkkoNOUM4fl7Ak5wcekfwrbZbVHRb0ikv/M5pbRbvSNsxIg+A2jnTc564DvabHoRTdTAnZ
4iZRMXy8hq+XslhX+sxHuJsxLxLyHZwVY0SUTzMESHcf7Cs6e+2baH4FC1G/FEP9GJzuHGg1Wobq
hYXT0NUmc9ET4B3mKE3moig6iRNrad5fBO0tVX6+mdaCe3fBMDf7PAZNdChjRsKKhZexvMtGwLZE
LJggtf7pPUFM+wH+LDoHwq4iv3/RKmFO5FHF2hlEqEIq/sX9pW+rwWn1Wt7ZDnDVPf9UkFMKaCMh
0squl0nOidiQWoxHkt/9ZLOtQUa1tNS0rPBNMkrqKEKr4D1f4k32H0lpeZEQpoDFhFBewfX/vjK+
1agaHqpAtFA5N2WdQkKzYmPAVluG7iJsy69o56I6R0/bhpYCIZoZjaya6MnAEL3k5XRYXvWG/Uib
VyfXWUW/oEi+Hc5n2gwx2OGCMgvAynKy6s12tkvZSH2jQOx2OAHbmejVASljB4VOwlI84MsxTm+p
gacDS9UYwRyomtsEJ0q9Sxs4+0CvImrgg6e4/3RmOsLRbAL8qKeFNzdOE1Qg/Z1b1t48Q6Q0Qn+K
lHnIwP6qN2kChfIwROIN2L36T5es3pAM9h9Fv8v2GFZzsmmyUvZ37VfjagxajaWkTwJKuA6Erk3z
vzO3tDdRDx+s0OoDIkjlt7Z3oVAU2YVY9jM7JjvovnfxwjevC75U/Y/nrqeQOZmmXZuz/ZC1UOmm
vo7rl/nWdezRdiXWoaqXjl3bDS8zNXf3hScopQoS/q2uZ5m0Ay+l7FWU1aBqJddzOIJZkXAqE/gZ
9v+YbDtGSLrZzj3Te/3XmoO6PB5NgAyVPcGQOCrz4RieA/oe+thIy3eoDQnjvSyPmTWlIHdlv8jC
LZ5RZE0GvGY/GTAC5ToB4deh0jLY4RxpMTlSxjCyNR4x56tIT12pm0RQyZUUf8PjO6rJlcVDbxWq
9+vNR19uTcP+IfWJIwuMOpeQvPrNiuhctKIX8zu9OHpbafPmS/2tX2zXG5nPpVk5jsHFKVgU4Grl
JHOmcDgwutFjT3/xRb6ahvCM5o1HkySq4XLN3Tvm2wc1Smy8qbWVnDZTH9iQmqzXiOuNpXvyakVq
It3aO2P69i1rhHIeJqkj2l+j5XilHrnVV63D8+jX4wtZYxuzj7fpiCaVzM4vcE/vqpXN0E+vP0lq
oc/238j4JzOAoR4uGhPdbyyvJ9l6CwHkSjQDunBP80CVCyFzTcPq9MDT/J4vbmqCXSgJ0oRMPpED
1Q+TchBZjdiDvLztX6sRislerv83IA9NI+6ZgJtPSQmL1ZlS1fEtbjFV1clmPt0BUjw3DjeNrdy8
bk7sAxGnHPfiZo8WG7mZTaYMEpylUgzpyNXenD+UImabQ7Q0dUmf47QwtGzD1xXnvqcrlDynxN7c
wBWvpobcPiiU5XheB/Sf2ZxXb3QmTpY7PIrjRdlBglcZzZRpkeeP8bkuzVZreo7m9M0PtreLRW1d
9MR3CqX1yT5eT9tW2b+eJ50tpaR+MPSJVRSe2MInpRCL0Kjj6SFanfZ8IpkS0EKtILPKikoXvkBO
NEtnlRviPR9tZmljXhtVMW3QLuRK7MERCmfdrYAwaDcYB0nPCTEj5jnobCoETbWrwkU6u6JRvkkd
1aaEZemy2wr8jwrmbh8V3eKG1TvjU/d7+xDrvSoFy75ZeSMufE8Q3hwD1GITAUQc/lhnwf4Ievho
z6laQWOnN7x6FNF9Z5KtiFoDYLrTekTUwTF7qpCiOxpaqSgVZcP/aG1xN9pRjlmWOajIqPI7NI59
PXrRQjA3cltRl8UFbjnsdxG5YcAFvgHwaj8o0fYtiKYiUfRENDL63WVrZdUlxIItKku2nfdlgxDQ
dQZZWd+Wg42j8pub8KIIPuP3NCqEWCZKLaHw9+fMudpjE82YUY8Frv7qpXYuaQSEN3dJxGzGPpq/
seCRwULT4r+QyOeiwLHeBV9El0XB4kn94vf3uNeAK3IOn2Q4qarJEhcYRQtME/dvjsAIaVcGOevM
UD50K4XjmA68dsqWQusGEWhQ3A935iD3ZH1lcA/3B5rH/i4O7G5iRegcFP+dXyuDBcivYvY+iGX4
OZtilAi2zp5uYnu5abnpl6cI/eEdZFIhJvdw7Z+bf7Ix4ccgLEUxeB6da8Unw5mrIOrRA+f7BsYA
bjEp2C5z4yYzOFtEXApxGzy/cp0bKJhBPFLJ3NiSlGd+SAmo8wzFVUolRZW/tFgftFk7BInGe6xm
DieYUGaJAFXLRl7tRjTyL6WU21yjK/Cn0VG1ubHbyYT+H21+tbp3YyJIASOUE/09XIE7mwre+uGC
6JsJbzi6SmEDmdgRrSqdc/lFufZvciYw2WGodALZzQJgvQx7EWZmZsgt0OGiHSmw6/emlgp5xj7d
ub4flE87kVg52+rhm1tE4bTz9HrApM9WLcqIf6PbnUlLCo89UtroPgsxzxqT9a+Hp2YtMumBMESi
HK5sMW9RjwH2FrROn1jJJf/NZNTF1wNVPvlUFFOqlxXIStuCC19bc+1wWxGxas/AgC9gNHzqrya8
1BRlDOXy975hEpyJ9PiK815W643nkgbVmIxkTw1+LbkqlDQX4uRvOQNBoinca+ltUSmPBYHokOXI
GBr2VAzo+qLIA0KCv99UkZ+M+PSR+xaISdBurQxcZbZo5qd8MQt+j8kTd6pQUwPXX7FpkQxFenVc
PfZi+gc/nbKzYvt+IfKYokDaohLNv1SEVEPBqOOFoGiiS4NdsjdVkIWiJZwmIuuJABYOVLh7/q4f
zBuX11NpMPZ78IORnhg49uE7siDi3WseDVZKN2C56kcPqPDpZyqTz4x+Brn8r8Ya86ZBefIjUDXl
Mnf9cVX0SARnTFLQ7FQK6pOo6rKr5ipxnBQrHYcta+AZzEVYWvxoXNoIfLfwal8jGpfmRXY/nAOu
EBXt5V3sVBFo597hOmcELDLfMZ7LuYxtagTLBuFo58pJtbmcL4/YnqiIIgwdOvpsiSqoUG5t/5Nz
7aahQfS22S6gbRXesHoI2xGk93MftbHWP5/b03yFilFgfiKNQRiwHjDqOq2S930F+LuutSpQF5YX
j0Izklcp7bqUPT9jMo2CoYgRyUTF25vdqXV0qF509miXjn4K+7FhhpENdSdqzenTdbT4zM0EspZZ
uB92xlbHIOotNOg6fN7pf0ncXKL4XArj3YMwyydTcCdENGe1ZuVSZM52k1r3h7/06v2WwYId9wbU
hWyzGT8WwiZ4Nw6cpRAkX5towlAnZdQ9Db7OoVFr0WpUU36hdyJb1e54T8T1Pk/5Pn63zI2awMLF
pZVUZ9WIzMUntePpMk2oKpffZMw8nSg0i1+uEFwPbXzf3elWmq4Ron5TTOEruJa32IGsY01gtZq7
W+bFEXxvogbNY1uCXOohq2rka8MHdnngJmaGKqI9TxB4nkA95VXPmqgaJSZ1U/DNYrI305armmyn
EZdfh052lB2aY0uVMwT76LYAmW8LoS11ZbPUpkKcMTjGw1VK90m7GWsgM4Iyu4wuvRyWZGbxMU5v
BXfYDtE9RaMskQzo3H7P1uE68nC2NWjG0XG6TqxXGMAwTibZRhrJKtVQ4KJ3vF3F9b5r1OK5AvCm
2Z73bo1tBjMBI/B4Hpckj3Os7fDKsrI+hiEglH/c4K6Cs6jAlc40xm01uzpPYa51F+cJQmtzkT1N
Sm7yPDdWXmIpUG52ixjPWtCDID1SOXeKP/0e+lzOVlbtWA7X8ZXp9U3jeKRLWO/5zcJWQDPwUIxQ
zOmM6pirTVnInkQ+dnSSMaYVwq4h41N8Zu9FpGR65mMLrS+xW47g4CIcHgJzuEUgwzG2jOJauA8x
jh8W3eutdGiQt/hAqa55usyCzjkFg4SbHHLpmFkOEHcx6DfXGEzhh3x4JAAvq0XIkdYSGXlauDUf
YhHwoPtNJDJ9/Os7VBRlD6Vu2u8liYhIwGURRnRofaRkN3CvIR/gbjPyH2xm8xB/EVsPfl5pCrrE
hnu1f8n846wu95lh2GnI+bHy2xd4u212AuKl6I/QAR7eORkfGXXdUPclBrc/k6ifPEXoIYkaWLfM
JuEUwvc5UrT8zEMEV6vJvHfxWvWwqeUQWQCh4sqLIpAghdxwdFhz8Ltv2pOCWKHCDA3GKt3jwmZ/
Kbrz37ZEpbvErjEIuMZXdOlYnSjY87X6n+/6urPgNdPvnyUdMDW5iN2oY4D8GyZcZHTJ2H4/4Llw
ryVSYsgJo53Ed0VtmDpawjmrPvfXANvO74aNrdSSiARL/KncJySLG0NGNaeV0Q5Rr8FblsfVw6a4
uD7Zt/L/f+ClyqYoJemDEiYUlE7rwNQ4aFBI8v2vu8ReNhUiTMlPpE0sfjvgpOCeJyz9FbKUJsOs
jMwZaLx6Ztw0njU+AJgq4uDQ50pjppw0swpWQZYoYgaeE+IVEq1Wycu/4ikjIhUgGfmQD+wRuvKG
UBs/FwGhEcxMPNdqKwX0KXqGbf3lU0/vqrUMaLpdfFfQhhOpru6IUFZ5BXFaaIcZ8cIuJ9+fnYsR
6RGn3Os23Dt5SKS8upHm3e8Q/qca5D+MOoT6dCW0WGroh+b6ZgmhyfPzGWz5BDE9/wxtGPaIOsGi
MT5zs++1a4wB42WaoKceO3yjK32khh+NVz7UtBqyE9J0YwTBaJM3spHl5So41PgoFMxWxvqFDGJs
5MstiYO6DGb30ibjTVugCXxHfjsXrmgfWukMTLrcMKikj5Cxmvsq14alfW39r//jL/atJxSzZe50
ZkuvK5C4l7ANEY++bLYCxNrQ0Kq1SdIyFblxvlEHqtIUlQZ8OLClFccDrC0iEF8OgBsJyuqp3ec3
dLVpWmeQDo/yeOzMtlUiLBiLmGQCjOCxt5A8U5Oab+sUMQ/UOaHYhaweSc9Vc2U+Q4Jfd+Eloez9
o1JWfksDRN6hgsegg776pyENsw+pdQeapqix1mw12u16odr6rEN9XuwS/9uNVacMOGAJ5ERJ8whC
1nXXtX1U9LZI0+JitD2xbS+UPQcGuaIWnE1nU1/y90GVY4KZB9dzJUJk57/wkqmXX86r47uY5gVx
beq3LN4AkMSNqF0lYouaSXewijZ07q1SKeISybMman0/mnfYNA9Zu2I4uqWCF3o7OetYEIuFV64E
d3H2F9OCJgc1w1osV8AZDGHdc+tyaJ7TZDtOnVvdzrqKgJdanz6q6YRFThsliks9WjnSK3W7QGpI
Sn5e7iAc7ilRUSIUBEZMq5eJ97KyOZ4xKmz5LJgHmIE18r3JyBbTlKR029jtjbs2lzcRLsqtl81H
Twjf13FpCPcnn/+5y9inP4cX8musTHGeHCrFodRcP5/O1xaoebwIzyntNWqESJtptwZQrU1lGd6N
aOPJxZBR72iGdiU3ry233CgMIMhTo/JtexkAC+OdKshT7RZSUKJUvb9+4Z6wwV1SPDbsg5ZLVTLq
jxWG4NnSxZAL7wTUB6tRiumvJxvdbYZ1MaciCcbb31/v2RsVzU3ngo5MXqWuYl8vb91CDlnweGvp
Ot8TYyD+t2wBGCbrs1yzZFhDaXGusc/RaUo8o02WBd6ksPXFkuruszFhnPmCCsqmGx0jhtRplqMt
KHXIY6yqCGBuFsCOIIt63lOUr5cGwo0F2FnH5o6/8X1ahhaZIie7Krpyd6AscKPSk2aLwyWoUpHo
Y+7tcsKZABYtFOk+8BUhdX8s0AEmOL2y26RUP6W1OKtjAmMRPBfyeTuOWy1xP8z+Zsc1A0URKY2D
90LiVXF/WOPKa3P13Pdg/3MUSpuzXccp4Xvme8KpdTW5ugu0MsBYKKzXbOhUwEcEBmybe1th7w11
erxuyfrkw4+UM5blS0dTSxoBKtalJ34PYo1ZHeHYPyV2VDoMFcGmpzoiMYexDFobV3XGL8cljAT2
NTUizK0U1amv5rPdyOWqFBgn5A9/7z7+wQ2dOPlFVGV9QsTl1S924Mw4YIaYypjXDJObwz/cv6Dy
bkTXShUOSNgwhea46PLKF4qShDiXR/13WuDRmHbBBWmD2ofWoaLfkbps45KX5mnb6DEjosgvzUwJ
UQu5Z/tlVUY4NKqGntfds4+y3abGcIC+9T1URocNBgEuC7PF4RszwGelvbOx8o9A8hkgMX0mhLi6
nxtOzeYOYiR9aoINyUuJaH7/M1pH+ENUT6VN1cEbxaIoZWZY9bNykPJJvxehnBPePrcrimSbBdeS
CjfJ56C4hKEtx266ris9z/Gc15gCUMUI9cd4AFwAa69Virc6GBx2JdbRhoJ+DkHNBJOC4F1DlUyR
od0vVRaLvYLp6aspXsXBWA6dSTz2lj5viS/Nwkyr7Smn8e8fKFwBVUWv4tvs34ndANj00vFzb28G
YNxBiLvUfofG02NWB1GRt78jTimRFLkMyCBU6/ROnZsF01O+/57880vGlajpddiwIhL3QwxaGrMN
kN4FYnoxJg9Fg0TqWMSeJEQmnlL2uDgqNGqRyUPrTJip1JKxEReioUMqDLVoGNr8ak7KsukNk8IE
AGJT1Qy1k5nEH8UTtLADj1K+RoMrVaiQg7kjtLA6f5DZIS1G3DAPw8EJWUunl0UfjiOfQ+YP/XqH
/Tq3G+pVs01Rg7ff9y9aemyC9Mmqmxz0zJG9dEAUlJqZfQ1z94xc/QwStwwnaCD6nooBmY8IPWK/
29IHKb30YWc+Bs4vMp6d3HBxozUZ/WUcPePtxZhGdnLO5qfLwyzsCKs4w+qjaTmlCVUYDAwJiJ+6
w4S2KUbjsidRR3MecLVzdxeYqTZWOzdoyctlnAlHerEHmucQ47sD+wfz5GHy+E151oE+9xLp7gaH
MiGF+izpK/7OsOu1DU4oBMB7tP+EQtibHF9PYk9SC34Nv0NsbWXOZRed/prdjodJexkdYAvcftv+
dJKOongdQnoSAlYQonuPyU7hcb7flW3mrySOczVHUS2swhk6jOiq7AkliqStNJeWWGnyG6b8ycZC
npKGY1Di9jPBAIO41U+Vx0jgvv16QpevjbQpv5W2rxGz+vy6NSJK/CHUYXRcjWuSWVWCx/v+sXxl
mw077METforqKOavc2DTNby53EMOoCtwmCuaRiovTkAjcJMBNdF8xR1Gpi1RJe2uA9uJwOMhjpyq
eWSbOSqQGrOQ+LnxPni+N7N9tgWUucIateaWKAa6MlCNbjr6ic0MKhh3MbKlezgTip/AnvBPiZo3
s3GYqKQHvOeOv24nZwni5XnhBXhRrryrQaHsz9MLNfQDG5h++w22tbdg5xEDWu+Fs73272xcBOln
EmxcKVtqXEp9HshwFvjtmdJP3P/Hq6EsbJ0nKRPORK4lKg5Qs+jaGMXtvYf3OJug7oV906+lBHkN
PoAjrkZtT7QSWPyKX44NwzOb/061iXzEPWlfcgWjL79wAylg8s5kwrrGXANPQksOXtCvmHYtuai6
4eJtWyt0V7nzo2chBvorW3V+tCNd3bT2J2QuQM0mXMtjzZqooi5Q5VuXP+MWc3ayQhJsOutWxsGM
+ih2zN3wUgdOPyYpQF6lTYR1BvypVVcKn8dYSrDhftY2IxyE5y7WPA8SicUhUZ9L+uPUqpOtwc8C
e0UJRCgHTsgI+qGCWIuZEfkOPQP1hCPRYPZ7KzZAKInhJ1QQAXOqAOXFwlVTY4JcTQQuE6YiS13G
mOSnnjF90CR7C528/TBKd9jh5yia60M7ye+T5yI98H2Ca7J3rD3cRTgNtcWJvUjM0fGFy3iPRxYm
lMFoc+wv3smSynfYdOTIvP9m2ToaAJCHRmwY/T4irn1IyBsGan2nSRGtPKbUOT4y3pjrUG1Nm3Oc
9uDox6DGvfMzlgqv0q5B+SbhtKVWtSEYAPJbtPCRukDH2mmAaD67d7W05cxEU9ECGuhJMuYSiHSN
pEXHpkjkB8cXuBa3losM6u/WNuWingbhlbM/kw093pYyGGt76igpeMR1SCdkSDu3dK8PkCPnNSlg
RZidjLy0ECQ1wySLslnrcMNkkqdl5GVj9zeOjSNV/xaAU3Ty23heIrtjstvu6dJDj+C1WbqaVQ15
xJjOY4pi8/rFQCWEsxFTmjyn8ysdNVlPj6vtEZuJWGmUbWE1ZKgvBrXZF/5AVQN7RLlAykz/27Ej
YdIbsQ6U1QoW3NbreSYAwAfhObatVFDR5o3BXg3Cb8Oldxe398VESmC7LBIIh96E5d5rSruTg0nO
Ni7VUyA4LupoIDhdbXlOMmbDoAU8HcddDLKie65aMdEjkw3ZFIXzX/q1t46YJfuYtcCifcD8G8DA
rl7PZZq1S+/6t4h751rsrcjYwTLwZ2w+w1kq8tt+KLvKromFYQ2by5osoiLQ05ifwJ+kn/g9VgMe
dvZvXxTVP4S1B8yd+UsPZLd3MsNsNKZlDl/PFCm8NkJaw/arFcWT9GPcDk0Eh6HP12tf6dLEMGVW
EiFZAp+7SaRm5/qLgWu0y6MjaFB0n824DW9boceFfqjn4M+dG/zsNFTCN9KBc044IHhOalo2/6qH
ZRWqSUvxYc0JC/m3P8NeXn4ifsAqyw9iohDGlXkkVoDHKTKwIHumG39F+Kcd1JoHSz5DtvxdcTn9
sqZxrx67EO0lELzzU4U5g6AOuZTVv8RgIc2Uo0ToY79+pUI4kl8U7I7artq5NIKEzMYgudqthxhT
9JxP1Qf0vMPNiMPPNzb7cRHwyEW7mBcrPAzW8661WdCuwCQtA2sELbKA69BPPsAwpsoxBVjzSI8c
5cuJm7Z/UjanQM46v0vw+ovTXslwNBxDsoQpXbr/8ceVnJbRVkmomOJhNh6c7OQVEB8NHCfSZr0J
dS5Ot0d41OrbAlNv3VSo6efMLe2REBqRfvAGvjO0xOJfdOXsRfiZPIyjXT4bX3vscsI/08N1wIG9
Z+TmtmT7Hh1DTOwQ9wD5RZZCVAuDzPP1HG8VMP03k5tEnxfycaMp5VDfxXtcvq74BeHflDwI/Gar
JTZBKW1AMMl1bYXcFtZQ3q3wg1ghhw6V90DCFOSnQnNIorJYqo3MbJWzoqNksVN7KmPwxqI75Vy0
zSJ0w4D3C2ER0H/tU9jIV/ks7HsPmwe/xTAOt6EFgXlNkPrnnR1Qe2yu1O0wybclo0/ELml3LrXX
o01En/0BJFc0jU/ENt8hO8iL8b/gLjYwAqD6w19FF1cg8ZvAtxmcTcLDJUVEhgBxRSja/mTabRcN
fX2Lt50SHNbO8voCvOywLxc7FXL7zzsJ6II3+NR7zoXWbojMc1T+DrHlE5gbDtqzpI3eOrTGTVRX
Q9nudpFrVlESRAf0ZW/NRX985NLwJ9BlGoopATOLpWxWVnaXAz1W8q+LB1UJ1ieB43XuxXFbFabk
4vk5TC8/TnXkk1er6hRSfbaXPTy8JZ2lmad8+r2tNmKgLudfdOYj43rKxActhV1CVed49uQDc9bK
xKpv7f/FZQQgrwmHhfGCz8M2sQNaPWl6cp7BDLI+tfAbV22tcpWJKU+zhdIYWi2pjoewvKPvp3On
FOpRRuNIDVtQhjxcnHfIEx/DXGzSrr/wce7ep9S60aRY4UXnwkySodyAotFx6k8rWCHTdAbm8VtK
KcZrbrmU2LuK89ydy1U6pdR2uyHGWmR2D3GFyRA19wgraU+LiZwfGVu7xZbuXJNuW7/dQLCHkO+Z
CnSORMMScHX0fZr0b/1PXF79lVLNs80zALOAjN4wHvh9V2pOVC48BNV1stMEcIsEChvVnVhuGXPu
M9US9+ZvWYtX9MAqnDchptPxuU52iA0XI//V3pdK8Z36/XzGa1tOX+bFieBm5BxCBPY9Wgm3+aK6
0naDMi6iAiV9MY4UgbHwYoOArFaegLAgYG0/BaIbfP1oLGFwk8O2Om0zmsYS/wd5hWtal3jQnr3m
EM+Nj9Q8fStkZ+yef42Y605Dj3FXxNTiMPLJv6uEKwGeohGHJGEZSIJC/EWLJZKNes9J4G86NzOu
/3t0K4BAEEfeqbQeIklYq0ftADRouhivyB9p2/yumPWErCIx2PHs8mNiEAcvi/ShSWETcJXkSV1w
DkIpw4zZWNqt1TURs8j9o7GP9rPeuRdCYbmco/siloF+OPX4Ns4ijCwaFVnVP7gl9+v3WyoYI1Kx
uC85sAjleqy/2vtdV0e6Pf3DQJAZbemuqxVmTxZ7b8cco4zWskrnjK93LA0cdy0OYONJ1zKxgqL2
Q6sJCHCQ5c9/bFZ3YXc+i8TKyvViy/k6v/arirQhdstesMbMyYzktHiiblbzNFUcLn8hKz4ObqDz
cKGSZHLXOkCbXxT/GBIDTcY9Dqf+9tiV/PW4PvSKxHh5z8zFMh1F+Km8lnFpwh43dmRPw9pNbQ6m
t3FjovNfWmt/0w256vdgesqQP2vowzXEEyD8WVllYvjsECBsKjOC3Knft69IiJjkmheZMfS6aqcs
DFrAwZYnAZFcE8r5MpVcrY8PrTzk+JcziiDUQRHAd3TTURKY1Q//7oyDIBhg+PbrMJ2njRuHSHZA
/G+eSo8Fvph2aqHyBQCXJ7zq+nvfuwnmObFcsq4Tc4eP38hCofktTcX2MY2jLWu0MxBPwVZ+3IBq
d6UepM7BlBSKWzBy8E8ce6tsA6t6Zf6/41TxTSUKVLJNN1HpSLe0i8T5H0VpwFZ8dhRG3ArnWb8l
CeEB0mGbn81PTSZG/mVjFQzZJXwODg6zu7w6zoJ2NzRNj8F4vIG5hBONgoU2LcHrolq010biNAWe
16qtFC8oDE37Avlug+KQS+iCS5oahWpCaXqus0SDrqlxO2Rg5KKjso1nUKsc0PjjTNsDqtnyjlbb
Vjpas2Ct33vgCjJ60Z1XfTBunuuMM9TTtbKbcNU41NQ26AnzNKWQpTBntumPmLZjSwMZ/XEhjeCS
KEShtcF0H8imsf5cV3MiZUASKZP0sUnoTGFEzOgPGUl+6IL/AQaiRFZTBFI6OGOh62sq32a5VUMO
Ufhj7xI15VifPhDw5h5wbPg5nWvEL/q4l9F9MfK/4LMmLv1z/c24+jIhg+/3K0qQm1amok587C7C
rTbEwbnr4bVLOexU94esSZ7JwjmBwA8moM05dXuT0D4cf3mS+Ey4vIe+ivZiTKUBjXlAwrxhm/Bv
5kcAP59yVyArCPZrqsZaqoFlOWlOCff7IS5/WM/7k4x1aHJ+yqmxPnTseMOef+uRP02/XmQnp09k
SZcuCZGL+KUJeEtSF97GEFsmOQVf5dzLt3B8aJsTKTy+cDLxnOjiqP14Tafb3fArUIjz3KcsBZ8B
lfvDe/oxhqu+zQmwTLI28mqxE6KuduWPnMawYIByYd//O4gSpDwkrQrZxhAtzTQgq9DeybYoba4S
17/yvmR5fADoecqt99UL026lYK6ULp+N0swwJ/GcKWMNklpiWn0qr8QkcCP14dvn3gRuOhtdbgBJ
HwGuCBQNJQ5dnNL+GH1VaObmqJSnIcjQTwYPoLN7qo3ROHYcQztT9t+I/WupHvEA40DId4cQ86wW
RlympxPok1WGXykaTcP0eveNXyFv7mL/obhwyLLhqYM+PLRPEdr0Jg/MsXrmMo4SXuX0UdKyWDf3
a5QUfqGZ3n5H1mVeDci1RkQ6PibYtXadRRG7ZZSdaE97cA0nAFkyJMM1StGEPNUahKH8ZOKASckJ
95uBLxvbh3d/RjsYnTgpGH2+Il23Af28gUua4NlSGz5KRmXXUvIeHdM61pZjvwIOshmAfh/JVgPV
62NU/2p5UsaPS4dk6X8TEmzLJRUkQyhJSmeJEqfNXaGTfEXSQeLo+vge6fP+Jg44pnOVqpiL6BEX
2qFSGuDfpA/sKSztEmcajM6ziECScQOPRYN/uq0SKv3nYv/nRE3Z8mkoyBOrrt49CSOH+AJ7MJgs
Y4WWfT9GHKA45mRv0D7wpR6GiMaFnUjbszn3p1Mm1XNNhQBrRe9CXYjttbLqoKPOWW79SdvIXSBZ
l7UdxfgpBNB0vQusVkMGyEogbohCb8U41lbRmridBqwg9ewLMQNhEf9gWSPfUVDU06yhZ3t2FHv8
HVZ8pCEzcZ7X26pAhz+ra5SxCiZuOYAhPGbocLDDJevb1p4IGPJ31HKtZCVmKp7Usk3KnuVHyX0F
E91uIDi/ZFXeDHoaIe/pKLJoaTptoGMQkyiHzd143k/7iKUI3lQHe0q5l2MXsTUpVnO4tmoX0nK+
YAwgxlIMDqMvWfuTeY4hKk+3eMnhU0BqeziAGp7ageZTfwcUn9JhRvCc96MbHc6GaUPju0xu2DUc
ALQ2l8wuDacIfaP9mdxu6RoENfiXVHBU8rDX7wKa6RJaHS4Z2iR+Prv7cBGZzMX99c+FTkKLRw4J
tmHcS0XszklU8RcC0tWDE8XdQgNnOE8/+vZxm43vshGk5I3freYX2aYLW8j0XGIJgqhXJlbdnxkp
7uXzYvlZ4skXXEgv3ls3arhk0qg6l2n2Mi0UJp4p+2Ksqp1AI1yMntsNNyx+h+90P06T3FJZOS4q
QsUSGRBYAAV7VJkdioFwG7PqK0TZmgU1V6N3dq5eRQJKPONYg9TY5+WR3y183hi36yeknhnE95Vf
g2R2mpfUbJNElEPei5TMhSZ5ram/XNawzW6NvXppI270ilSq0Cwa94QRIlk9jikXl3PqU/msJvyN
zgxcw3Vbqa72mv5WNujS7Vi4hpuKhaYS1F6heha5pdW0M4KsrPDmBWkUITwYZTmiDNXDlNNoEMrC
3xAQ/dy08Jw1DsHUUlhCpc0fyObogLJKkRP1iuQ8rd+CIsxlrAqlkhHsNJ7CccbhDE0MkYnXsnm3
kwy6jQbpzIrT24tTwJhBb5KsWAR9UaLT4RtbwfpyMaXDBGy968J2HVdtGJ+yBPEKVVRTyyHW90k2
rHg4JjWKF/oLdSYmvOtahfVmrgCy/ms78eSgOw4BVaCK0KJnrgLzAr/iQ7B0u/kK01MS904iu7N7
m//pBlGgHMxNNC8SDUBiVLfJwyAAxsHKVhwW6hv1RntAhg500DHUAXDPI4Sm6HZTGUDsGR5Jiyin
NnHEBWBvssjgGExaJOBHdmOFrRN27IGIszsR/84AzRdH9lL0rR7KXPHgjG58oytbBlm+iTGXKZvZ
3ga/JHkXK573zXGFH55Ak3PHfM9zZQYbmdZARRl6KVpCX5L3x2y8kN53yW+CaIwci1TDsPDh6t/p
vnN8toBOdOcH7MKJCblK3LZA/lbxBO+PMQpr2xVNqzhyuY/rIgVJEu0p28/aswN8lkNb8GYNBz2y
MzxZxOkY0wVQg7iq3q/1gqK500ufGIj85p7pTY6CIvwMdorYMH3J7JnlPDtNggIKIBKBHvlrBzQ8
94gbGHKGX9+Vb5UgMEWprnkwUAG0NcU9XOaT7noFUoCPZMFuFaig3Y+sOVRzl/hiVzfp7aB+MrKh
MOmOxzEGS0kafIdTru9OBY5EEg0w9InPRfAf+Ba5cwJtittJMDpFVlwLvo6DVFYAQx7ql15mlsW5
OmiakrhP3mt1T5Fl8H6yB8wtI9xsI9QC2o30kZ6ei92+r5nydBI/LocxtsiH5TC9ePJO1yydOmOD
V6DVZyJktu0P88jWhbYYo4GlgOA/mYsUd/yFGEVj3c38xlTCUNMeLekH0HsSVSpu8mYioOTOw8K4
iA8BjQjKQBM0CSdc2ZHghiPI5fyf7KucszOnXKrhAf6L+KQl7/l2RNJ+uKOX2pUryCC/EmMWeVHQ
9uossz8HtvdcPWB8pHJhIbkrb7SMpMmcqpfIJuKS2DkEKYVSS8WZEvt9Ar8HFxC5mjxr6Wpr/+KK
fL2ypSnFpByeFNhhIuQvaZxnnaZ1FoTTGU8ZIaZJYYhC2XSxQnMSyWWFMY4ra+unwrH1bqWp2Taa
gh3xWq36Bdgv0fqF0Bi3umXP/Q8dkRbm5TVKprwtuno0wtEs2MSb0Hk7k39YuG4mt5OUJXtVAH4g
psLyDajgkMNKZMTFvN7HtmTp0tz6tAAXgvCR1wRohpk72XJGk3G2zWU/k3cp+/59DnejEHOdN4qo
3h7Q0UoIOijbw+giCVsnGyf/us5HRdyZZhYQiIOcLOZ2R4vQAAA+cjCR1ay7/mj9fn0tt9s+UDKY
aos9cJVWn5riiEjhZE/8GhpWR2YSa3N80KlnEIFjxTfi+olrxvZ8kroDll2+OMXb8TUnpknxIt/P
xtWVHynlmED4YvrBM1tFj/mb3JJPddsKVl8/Kub05oM3eJ+tF82DPGvwtgLPX/hxP9+txgIz52i9
9W++jWWkXmOUARi8+OGQmOobPqT0WUe+H41vhexsFURT4g56JT2kRb+aFFmjInUYUtjMjI+kflGH
1tNVKkjwiSr2OgWdR13pYxqkQyNSs+YzwNumQIwKh33SL6aN/kgHObrv8eyttAt/nOC+Y1pPUX+g
D7uPs1giJU+FN6+vHRa6UrweMFpbE71mZm6DE7pVnQXecOv2YtSjNhu2BGdfdmslZSmzy6MDIR1h
HPtPSkhvQYSlqKLjod4fs9dJnhAvm46c9tnny2rpcbbhmtGkhck2lgqb7gxMLjfMkGjolrf0VawW
pEE3rm48EtHDUx/OKuNWymRLIvRrUZDHQtxvRpJbwBEM4GUFB+K/+xPyQOloDLlyYW8WVrHBfR5n
0hiu5orpEoqui7+umQRxbM3JTXkbN7c42vJxCM3o+qAlqBNmrCZ8L0mlE/H/5hzDj9eDJ48E2pWW
csQlrlZ5lVydacSvsDp/GoEW/eLHk1QU3dTId68qCal0QMlbdyWZ70GOfUT/ss7LxVqs9L/1u/9p
YrpzYsmyq7ijAEgKAFH2y5Kys9/8cSmJJE/XEI5JwNYK54q5Uoa6j+DJSt892/SN+RDjpt6cHEeh
+GGfFvoY8ESrg78BawBnIvDdH7OPY0tVqwDLU39KxKEl1Al8nJ4/r96ZfypUtvM64uU9qozoq5P/
I0Kl5kHp/Bb/qJYFxRnm4hRjD064pB0G9cBRL17+HxpqJ+ijJbsTyVms0AtSPZEDKTDyLNd/mEuu
Crgj18OwyS/fM+o4e5zO/25rAU9Y36q38xZVRYwY6XooJZnbTwoLQ6MXhj2X2TakAH/kJ1+/KsCu
d9ihtT3U5aGbZr4du1/tE8Dt3ro+zO4gRHESNvLLIahTIEm2AaCuRSWhMDqj+TJG8NwGyPQTp/Ap
Kx0VDf9uEUcdL4abk8UYy7OxrfrcnZwMd+sS5f1aUUmMseo8g/nn+VE6P/vcTHQLFupYDKZ+SNRK
nGx0OweMW6DubXyCHf7Ou0l01j6wVG3svEXpYdWNanKfBeXdxnICV9HO0TlXCLXaEqznreWcJJb8
INKfyDMpAoB+1cp6U/cvIPLW50G8ozjMYxGNpFw7Ql420kbFNK1i7UvgeiQOnB5rV52EhkA1SzuJ
Z7Gd7qY+KHaHpKTP3xaAbo9eRJw3R5cl85axx/lANm8SEZJFe4jltlOuDiNqk5L6CpPnea5MEqOr
soIiJwQ0HcxDNJjRWqkzeF1u9uruX2ytBflPJA+uPQxnpwEYSM22GkWU2QNhbQiYYjB29UMnA4bJ
/6ozbUYwRRjns2fU7d/Uiyd8tfyRLDfafFCewtPTroD9AekvXxEpZMEqgWBFN90g5LwLaAwoUe5G
QlpazVckU5Xp3EqyJSengW9ddDLUWgPsIn+jfjQd+y/uDE1IQwxZKWnqjhNjvTBRRxEpuXAlZYHo
LXYXVYT/7N4VHwGMKu/Ck8ABpcRxQfJyJYK9qjRO/ogl3DzYZ5FBm0WaXJUQ7m5qaEeK3UbKAt0O
7LgSZuIZi2IxC3az7N84z2o3yLVCVmdp5ievuNSiZnIFZs+AG5I9ZaPHo5UhRnJfXdY+nrUcLFzM
z4+IhIfDqawuCVgJSA5n/iI2gOEPjMCedToaYuLhPboWhsGdtouaVN2Aibi7RpgF2kQR6oOSmoeT
pAoZP+LSsXLKbb+oARI3awF5dCq56k3u8Ttgcg+gXdcxZwnj0bXqIiW7ip4JDEMiWpop6Tfm+AC9
mtdYJRwGqRZBJQku1rtRcSVd2c3RVMHN0eSNEwWfLDrXcGqZZ3Jh963yKtqJviZcueDvsrlV54qG
tTDvbwPMXkenrbQWqqIMHufmnbM6lOFJ8jBq9V9BOFypAAt+RFfLST7X4AqsFjcrr1uAZwo9nC47
qfZbBdyaF9DIg/dbo5LwnCW0BCD8+j/ELT4pCbsuG7DgWAvn3pg6IZSIOVJU6fSFwN/Ff8w6o8TY
mCLJ9Pqc+3ypIZwo+7olMBxrYJ3YQapy6Phs6RpOI1AFCfto9l5eDRXfUCjWX2CQ9LDsg1CnGaEG
SWsGcW4uVndazAYcD1N5VdHpz+0EPVF8cNxf4pr+uYXSLhQ4ohPlC6rBxrP2MMvwda8O7/V/mYwU
Gcl18jUp8BE7ckqeT/CpUnhSyV/6saExMxhBs5/g6Z4IS29s8i+iS2SApF5TcvgHqP2lTwju6+sY
E/Ydb1oMmMbFZW2BpWr4RRDPLYtmMD6Q6hPvruPg+ttTgPrS+BW2F3hPzHXvt185vt+WC52yGtkK
nVG4+ypjmjFQklRqb3saLjJu+qRt8ywXOVN3p7JrrRKJebaxXyDJZQTNyxVCVDbee3F+5lDFLALz
UHLWqwjAgMC7qc7uEORvH18AH0i9TikjvRWpBJbK9Hj2yBAMwhywbRnFcTuH0oSqPHJcyTYckF85
uUKaFfq9SOSWq8mofFwfcIWbkf6V/aZlV47lPpWldrp13jIv/Jt9iXzSKEfLZAq5O0VbOzhYi067
UrslkMAkBzEYSj3sPegoxuBT00G4mmVOD0yI7G831ToOB+T81UsidWYsuEdkvjnz2+tbZHp9cByS
dMRnj9R6iPSJv5dfQZyseG9fVwMeF+poQYJ3IczUcLvKn0ucfgKY7pf2hBpht3AwDAmGQ1aAP/Zn
gB7BlXZaie1M9sOmABqsP2GaTWE4fdCDwflvc89Yanx9rt/kMlSDxf8uCnb50xxzjPICIsaGXKuh
6gJw32iyXFOjT8ZcjmlpVondYRSe3G4jh/9gxQfdZPHR5KI9BIGlqkkidcZFcTCBpadq8pNhkmYg
rsfcYyjX755r+4uO5Nopn2SecuMUp92zvy8sPUb6nsHofF3cOh3/ll2I0PRXdHZ0vpHtfxE8iRWz
WxDo83HB1782moCJcMMpY0hK/uMzBIFgZwYCHtom2nxmYZYq26tgfeRF63s3G5BDg+/sPYpSKF8E
mnpw29WsBPiW3S0g2IC2y68AK2dGDmN/tBWYjXq7KvvH4ZHT/R6OfEe4gQd3F1PRi1Kk6EvLYEBR
DBE/PTtJ4lK7Uo4ZkpkQXlhjedmfSx0RSUlrRNZs2tW0q9ODtNovezwdO1kdi4OsbSVme6arYsaD
UECf4p5gExYyM4zZvONt0+Gv7BmPKqFfHb/cxV+Geh0BAWL2RBXp1Bn8yjiY7rBG999ly97syd3M
hvoRQSJ3OyhSUwk4wqf+TrnYkMzk4IzI0Csoj/mQYeiZdWZIbSp5LcV0M8dMXo/6kRiaPXUpHBT+
pzfUahTxQExkGjP6nI5uUh4MY8GkMBEsm449NzCW3gBquKiHJ7uYicY01nbMKfiiGIaOwjB8Udhs
kRwz9J7vYht34KejAlQx9dvIh6TjTZPrjlq7pGUdAWR2SHo8qv0F/lXknTFPzjRgD1CpKxDOLR3o
/J+UlKr4iZloy8tTS+M+GNk0/jTY9dYi6CTmC2ptQB0XQwNSQfxL8Ek0IQIDu26Gxp4JLJc64hhM
w1rUdtG4u5fIa93J/oREDbvaK32W9KVwVp8XtkpcQjFRWmow9pS4D8Xgt/FEBbPkMOtImzw/N+Tc
6D9g5uaDcBdwWtBnfRWqYtkHlnWUqbsCAUXBHA1BJ8fR1Jx/Fz2I9mP5XEiT4KTd5O0dktpRz27i
MpBZCyaL4qyr8V749sFMZm3PmL5VOhY3BGc44ZwGppobTC1EqRltyTz0LODJNH0n0FWbFyzwIwzJ
HAJ50T4VTxZkRaHzZ7uUKJYMGiE5mb66jMlbpse1YiokUV9XyNZc8XaOBLy4jmA+Ra1EJTx0p1oJ
zR/hBguON/FY0BWKr1WkZGNbu//IvHaoohsw6mGcmc+n6VdgehCXn6664Ed0RtyVnhk3xVbhCdx6
YFk3CtocR74OeM6nm5495VXqZJoC2BsF9Pn0rXi82TJEHpycfyha32rjT6wpjwAN6XaQ6QYU6b0z
Ackrv581LiPjaxu9j3K9njdtTofRBENN3mSENME1OLUmeCpb7RZq8IaqswQLBKqYFj2HsL7doSXV
fLm8B6MN4SPxNB3VYKwFirF0TDkVmIpD8/vB8Y+q6gnbaf7R8XizOQi8/ZdYHV2wjKkdoRBOIB/a
t9R71H24ZzVKQiGdrWcjqoaWFVajQJk/EtxR7kPZ7unvCg6gPHJypSfIrGzp/0PjhuHJGvJC0uSJ
ICkJUIvYVyjEhC52COpIa6AWdPkM77gun+j0+nr46NH8/uK3cEheYyAlaxgJINcudis7/RE5WG3p
l5QxTCzmK1VzgRKvqSGl400QZRPBG7rJRy4JWu/vKTbNZtLT2J5sRoL7sMzfF+n6vVvLyqrLsyWt
g2lK16g5+i2E8P6PulifLfGTIKQRL268XbZf8dXMeGGoyv6n4NOWodehgUGxZ2Ye3+ub2clOyBHk
eeFQs58C1qCmpIO6h9WvsoIHnY3KeANsfJgZFovTVC7EYUudWXPz1lh0e5YSoIIPtHeAJUGsUi7V
hir6BBLvsdTc2sqWxRBYmslFiXJBZ1PIFXjwAA/2Og6YQ43QkhK5NH7ZY0J6Gsf9ci8+p9cPD9pw
K8NOa4IdLwGf1aj79GHoxWYC1i20Qz4OkZj6q04NRkk6CDBG5CS7AIlOZ/TFfkMV2hRQa+lhewqM
hQXuCCL8TqrGZGS0D4iW6r0oFpvwLt+l50sfdq7ZGSxNCpiSGwgVyN7T2H9OlClO4/rgpwmPi+1Z
GeWCeHGBcT7Cz4MFebSiSFfH7GocXeHvpORzsESZZCxA3ss1532w4Qcngc0ZQaPP46kIgvAOQofX
g3qpHbiQPvmr9JCKPhWopvDDK3RXJw98mJzeMhv+LRi59v3U3Tx1UNswUz2vbDUr2MwD5HkRoW8C
svcmTQl0wSLPgNtrD83/HK2VmfFLnLrD5DSBmCZpHJMSiDu9SqQSbFpqs/hspZZqTkDFV1lFFlwG
kmAUu8mk77ebKjPUI7BG0AcaJ+gJZJ00+KJN6FRtcyOn2prwFyVN2HMgmARFD6KwzXVZ2+nerHgw
YNgc8QJwgApSm45+KqWKBE4DB0LcUIIldIbx7EciVjiWOomixkOcF80UrjcjVkfW3tceUjf0CBvY
MDz+WBSWViPs7S4cyHjCkeBI8DeihpYbcx7MTjFftujxWl6N5Cug/1Kh16UKa5Q3JkQFoYEgOfT0
nA4bBOG71C+3CYPuMXR4XUUAoHhmUL9HID0OdRyCl51ySbBR7tidkOXThtYobm9S/0nHspcaQRfR
ZfVrUxlp7qxD7CP3SyKuP/R6egbEFKGEaDoOeUSMkpgJzRkEKg2KBU9RZ58f3WiUdETT7VfAXFuL
mNAta5OUOMJBekKhQClmNotdcv3vjd4RHTwhVPCoD/8hmgRgLK9l/caE7oS0BzeKi06S+l87Hol9
njmNGJVvTez9WSQeLYt3Tx3QtfbMCmrD8RcqrB5gJacC/U147lZIuYKLm8ZpkjYUhIbkF2Kq+n5D
RMtcG5zYpj9rwWqtTwO5yBDB8tECOjCF/1Eycu3hP09G9OrOJFUodUYB4uQWg0ZOWxBtHGaGmyrI
6/FNVSHrYdIDopThDdKkq7+f/4wn2X3Y3q146FYSHt2T59X/D7JQhXCBJnw+8qqn3ToDdy1mX5G9
bKMAgiQpERzQ8rbTswywh3P1v9ABqPkLl13RnkEPlA1l+PFOQT8zrtiRRqcNtluHZWttxtLgLHSS
32QQW5BuYZBrimnaaB9QmgRiIx5MiU2QvV0yXP3DTOddIIcqERDmsqJAGJTA4qWhjBghuORlcl5c
om09rUjME5yxccaY+gmuFUl7lpw4lVIXWN+TExqBJ451ukuiR5xeyq/fZkajy4SHnUzsiEs9WcZu
7oTqLLJobD5j12NOn4A9gMRF2UhOOLqZ0wYdUxFWpG13hyhCOKrPmKAl+SNRSNM+8EyDTESro/q0
BhuieXu+filWTP+4PLij3TVr/S0izY1j5C4QQQrPnC64gQssQ6HEjVE8bIepzC/B1a4Bp9N2+dwS
hAhKgOy/B2vT+PaW92yZ7AjmSJJQqff5vrIT6PkMuuVcPc/hSFc2omJ5BKY5cguQYacBrJrd4kIH
rUZ4TDgdf1ykWVWTAOOu9K2FOT7ewecjF3QoD1dQwiuWIGLWQlfRrE98a3HDYZgzC13y32/yo5Kf
oF7v8nWkDHx3FdFqD0mGHNzSfUMIE/Bg8pY28TlX10jI1pbaSo8Dg9pEs3mZUcEAvMHoStAZ0fr/
H1wnr5QwxY9gLiJHMAKYELkYEPH/qeOnmqD1ny/qqeOnHdkpT9eZVxrfXMA019VZ/EKKL2CSF+yz
Xj/luiKmq3Tp7uY3Axua+0S9QpxvNLo5ULjY0L4l9KdNWLmIEL9uvmHSqSL7FZ9ZlKJLa0QI8RVL
6tScs/wSo5IUFZXda1ygeNplZQrr3PjNFyZ09IteIrRpvarCeY5ZFUlDwEKkbrXfNRD35/cpSbHT
8hZ4DiGpq/LSMRP1HHgl6ApWVbJjYQa/V1xv5PeteOmiCjyxEx+jlQW3xuuR/Zlnz38OeNBZWSYg
6qwm+iBBPtr6GeYn/mh4o7m1v0hzbhMs5wiDZyYtaD2SapRYslVIQEeh+ok/49YGeHkBbaTeYV7z
sOr7hKcDtmssbFtheEQpiKncQoflEtTxBqLIYZKhTbxN215Mp4fcMdOHANwyLmjcYdx9qSJTUaTE
FuUvH9yVlQoayfouO6ABilkCBHkb6cMS/3ZIoNgsaZi3cKOBVit8HrbWtjSwVZRWXpgMQYQXJR4d
NS1RF+i7Tkflz2fIEgMjzXeF0/iJJh6A58hzpt05VuKDlER8Z55MSydTsJKjwqDh7Nn09XVvNAjJ
gFt0fbZDdrS1Zs+4HaxAMAeef2esuwNA6hWUICck6Ffb9/2kkCkrdG9ETkZi4Hl8mqB28jyC4pGp
bXOqr+pX2NIcn9GUoBu29D6fH5e7v0mvy1S5SevtbxhiC1gG64kqUXbvKEsxtYVmwWkgid6+ETTe
2Og8PhpE6DXpCrM3NdhrOpWrlQJQNxrO0LEiCm8EhNeBQzkJBx4fmLmEeA4hau1705mtrkwhUOaJ
pwCFNzfShZ+aqy0bF0auNU0kWP+dlFo3vOyiVcjojKB5cpFjUMj2xvZBlo3aCLfuUdXjfGybuqDr
HODKmnCFyTZ7sb94eloID1u8pU99g5cLvMKhMMEG+sb9qbQYoMahJRb9DSHBrFReSJkPpcl8wO5j
HRAa+1j8VKFjB2IWcmJUCmBD1R6Dk0+lxfeCMX4KTfCnqhlCCzSsfiBCizGFyK5IYZNlKkXYMD4I
jOAzwZm1SLe/luA+oLuoXyzs75P308tX8L3YEVhEScJh0Zfp53r+V6KDy9GT9oZ6AVbOyliZU2Jk
UjwkzGA9dZt81kCCeJAnikqMsEmNO+FUotT0AV5XvqROV+EsVeXq2LrNDfPkADPNiiRqCSO2/dG7
tQRdHsF4XTDNU4uXh8jPTdd08hrx86FgiwQtNo/9MS+1RrXcCK89zHmqhsZoDvaP1rT2dinBxOoG
eeomMxf0QfFO7czVgK8HcE2QtwM9OBhHIypJIlK7XOdSL6wzbBoZHO5sz/eeMrjqE8qL1+nV1HDH
uci3+hSMwMYAWKWyKhDVUsJw8YiUf6pav/HV+dLz7ftdbrX2TdXxsJ/8fSZPQXgqOO45BIjYUnem
qZv64IY2fZgLuQNxmFqN8ON4crHLv1dj/h9wL53w1/s2Ld1kqGUN7RssyFZvuX7E4TIM3A0Z/muV
TyHpbx10X0KZekoTzkWRYNHfBe4Nlhoxf+w0fqsvK1Oy9YOuxgbN11h8C5UFDuWiePLlKJjwpROO
xSVh6cCaprFp3dejVjTZAYraxklaVwzX8fz8JWOqz6l6+YvtL18X/U65TlDv/B8TS3T8GOWGA+SA
TFs2IBJ6ZqzmBteZNPcQZ0GLSMIqEEdBalzaervv7h6eLEaqZ9rQ7xhRvuPSmg42c3KjRqj7uZGt
T682Jy5zQxavEmHOpWkukDCCyMUSNB23gqdVko5OF7GKPWqhenb7JwfL/V0pFcHv5CoKT4mfBb8N
Bcs1oYThzBv5/8Ltly3+STum39vtsMe66HGcCUcVDRJh9aw6R1nuEKxWiVSVsD9+3kf0QvgrvOMR
Bx3907M2wwXKgk3xMQ6I0LQbP/O3V/+mJmoXSwvWfFjSNmU9N/zU6Ww9LbD/3gdRC10i2skZVoK8
kNqOveyw9Ynf7MYH253CRvYMoFFX0vEMkB2okp8bVxHzMOcQaYivSQUlmI8dzOk8+Rvx/4/dvcfS
kJjQ6iwcDpTym1m3nr3AuzutAowrozqo7EjIS+O6/I7SULfNoNWxGyjrirdf+EHsE4krgg5Adodw
JB9OfV4Jd13MU6uR77HRHFwA5BZVApLajDUdeoCEAJO4ZM5Th5RgWNWakEmvYLNlZoCSfJ8anB67
T/2muUs7tDusC3g5Q4VyJ6Z688VJtGZ0TTq1+BUZMWHWd8TdmCnHe0SaRR4ffz5MK2z/2YgkYswl
eQj4SbpgP1sYhNTpJlE4yBrw3Tk2RKAeus0vuJnA6ayTSnwwWhs02TIIBLDli3qnfswFVjsbC55c
IWkwE+aiujqmDin4DhwYuc5BeNHOwfzEgkbUQ7C9+fu8h22pC74JX3ahAxNtGM6eC6ciTrIo8aNe
iBa1M5PBFllI9rRT2uGawri6jcGeSnJozjJ+4eGMcbQRUjHtF11xi36g6dhAmRWF64ELn81evPoN
DzaqSZidrVEC9klXw8dl2o3FS+WpFlj6pGd6fP4WgQ7zZMvCKYQCG6R7tafT+tFo2vQ3gZhFFAK9
SK7ODwLbkrCvpwwpQT9Q8AX0BAPchsv7NtTXconT12hTOTsrhd6QxspKCJ1nhlEhmHxDLvmjzT4b
HR7nfcqsRxRoHb6Ydvrx2qfJ6tlgDITpSVLpoU6JpaSo/HmoCeFjoMI+sT0PaNiVgjRtIyuq6cu+
/WBM9gnHYFrtWD3WISsni34Oz2Jv3vDqGTkPMXCWrih+q80GAjcuQvVbfq4CdVrL6+JIt0NoGLhz
I7TVreB+O6ldZ/0MHKBiulAV71F6JVcmSaIloHZFVj7Toy+Otwm+4ezjQZoNkZyZLpKNDT/6k35c
kuElTtAPABraCmgPDG4V91MXrD3XMNwOPxMQO+gVcG2PphtmUctWlOYcf93TbDTsPo4OVaBMYuIH
urqtKMPBAougPmYnRVdwgrDxAgwqJu/OG2YY8R3Qs4hbo4sETM5weKcM4nVnt/N4hS2jgRBWBC79
wTfO31kT7wJkGIR6zaqr5tvJhJHRuxcNW0TJkVhPOGBbv8tWTz6zYy7XrYdaVxAb2tBoDYsrmBmW
p0d/IUI13ZEXVNjv05VRAUinEBBOfGTFycwLy7Vlf3sYrFYmD0lQ3zcTRKxlo+rDFLmhnw7CbVe/
Rl7/TvSkQFIISb224/5yJ7dV+doH3zzv54WV64V0wxRmJfiF6n3dyLfpAis5prGptka4IGp8Y0ac
JY307b9fQ/ld/ogC0VPKQ+9J8/owJpqZ6CJCr3WtJzDT0Lmtecy74oXwls4+dV7A+8w7Xa/3orDr
zuQwk5wBVqlQtztnHt+s2cMzooWOwraHaE74CQWM1Xh8usw2mA1L8rjfJV2d4vnzhB1y2hlHBjFq
H/fZelc2NkXcdClVNZlKm+YrcAuPvnPI3CFGjuUNVd/ZWqrFLmIxvSHsYsVhI+j5df4Coh4ywq1u
WgDfPsGY82VZf+CRDfRC3jcW2wgagO8HDAUXLnSetYmIAXnKDMrpMhQu2FREmixXTtHonAH8Ld6f
zWK2GofTFhYWmCMUePxB9cvQVh4Zo6m+GcOWp7x3zKCcHxzzF0aFHZrlgEqRw/qeMIXOlBdcDaix
C3BOELEXiYhmKYGyrcaE3v2dehUkVnBKy7ojCTXEbcidAv5ixrOb25PJxPOyK32qBMsJHW2XRi8k
ZksvfRW9rx6JcuNCPzzN0fCA1pEHQH0P5yJjCItBwFTDNxKWsOK+4V5ZaRSUSzuSM+Jvz5aqXKA9
o46J+Er9YxjqUpEy9trZCZYoYXRKSpjevASgIiJFEUvrYKKvdM9WNOFblR/mDMAZmgonJXFxGmOL
RrlderIiD8kec9zIT0Cg73ig2QyqztJO+aec7lpT7xRIjHhye5yePwh0azf9a0EhKMFxRbKYwTzH
a8JXTdfHKBcB2WnX+AGSCp3gAGPlOs5fDnKsHVPA3c3iaIihnps2BXig2CmIze+T2XkaR1E/H882
rf5tgOdlHnRQCRoKOKe8jVZq7MGfPdY5GHQKlBkOPrjngpNIJLVHaeQjJ7bn3N6Mi3b70+PEnMIR
eocK+xwPv2KRBExqEot14HxNKwMVzDeuO1r7Wr3DmF3R1eUGRY6yOt0B6yI/j7fejZKQuZQ4wx7C
QKNu1w2KJiAWq1nrcUqnOTjHmtYjLjaG8Z26NuUpVUrgbt71OxBB8rcA/i4+3cwH5KBjyO/Xdpxg
k2q61lVA+b1ZNj4d8PtZdyg0C+2NJ/a7uiPeBH5LGHTEnvs8/3i2zW5C+5CduNt5rEBH/JwP9UDc
HeLMHmwPF5gSyu8C++Wm1zUolJsPGz4kA8XNEdz7TI3Y3Y9E/toIa9KK+v3Jo6u7kmUzVobbbDkk
I6KJItZZS311pAF/otcxhf6fUxfN55M7bQeOXEuZWIL9KXd5nQ7zlhUt10WJcX3ZAUdH0B0ePAnt
BJm9w8/fMDr3oQxkH8li1k16NshGr3j3gfjikPzwzasfASA9z3DYYnh2wgapNbXpKDqSRTpOu6A3
w7AHfKBj3PcRh1c06wD9L6nNhvFwKLR/yec4OWX+OyGoCXc1PV3Jk3c2nsQCsInL1VshsHXrJPli
d3U+Hvo/DvQHB0kFjgXwrnCy2V2uMk46HRFNo1Cr6r227iDTfi6Y5mYBgd5TGhVKn7aIg7y6S87U
9kD7fVdF5yrcEmKxM9/my0SrKq75ZS+3Ir4OmnSCpzzKQRpC/KMN8xSiuErFImpWDrWEOwaUBOjK
oc0aZBM0SZktQW11h8t6ZK5y+8M8y019Oet5ZSRrhJMpffHah1O/LTmGIfbVh5Hmy6bQQUNEOkNd
jYRcHlDWR++B3dKL1Qp5cbzbydW6vRaBUCEZYdOWJTv9cWQdgBNNEXQ4HrayWTkDlMmA10SkRCKw
FS6FBHymPSXjhnJ0if2x21LBpSL2YU/yWglmRijLbYhyPvcMAQzdjPXQgWJ8kmk1MJhayZqpniHj
GGZ4tYMEBxS9QULky/xVF/SVcbdChWNrnmZIWThgtA3Sxnf4s6ySsJm2cJxPtQw5b6NpJT7/arnx
sddJMt/I7/xEHYRkXWpoLjTVz8tRft1+ozZkUkzOWDPPtyXXXsQJrlBV+c7lMRDZjZoHuAYBQTlN
8lVHEMLL5ROUZVA4u2uVNKorjiUFGEx9xi9lNcNgJGPZlSBmdZG2soL1mOhDy1Iq2rOwT06h7fAZ
WeRUg/v9DGhFP0UIA90oKVP6IEkEShpA4hD2zFXiUsHueHsv2sxRB3t54fxnzTnHCnh2Ksh0886M
UWYDbbJieaX0otjHImUTSKy3iwtU7dOR52k7jItDTONRrTPL28XwkHCepxCYAgiO2D66/smxNHlS
Nbv+PIIIQ2Zcww/PetG1YucMXByyaxpHgOSotmaxwUI64chcelYPT+VhVcphjbl0VpNaEAOuiChE
ZTPpWudnHF5g2N4sIRgubroG5aSYuXJaMZrl0kqoxXksNiuidGLRL9SAeRGo9znFP4NR4SbHe1os
d7rigRqjlaejdqG7ym3+fQqSbYxdg50lAyvAsqGLSvUvHhXyA9ANs0TSE7AOUjJdusiEON7Jn7Pz
SaRur2xcxGKNfLRsRs/12MKCVQs6feklfHEHTQdrY3siTPLvcQMFXyiRxJyAhNsRkUSyt4hptir+
WB43ltp1EfezVJxdwJvIbfd7FvznDh+Vbt8tCsDI/sZnEUJiOEteX39zmzGtSEEXBxV0Y4UAjRoA
CAU/pO+Exb394LwIDBKgeY/7UapAH5XKn7xtzEW+XATlLHBPEVW2+GFusFJ+ZiR0UKlBz/1KCsER
fQIqFXBHHZnP2XZsNaUnpA+21jFSvTq3uR11Xy6cj3fLWLj8ut4o1M2o3n/qLXT1WqYEgdSCW6P/
BL/iQTFVHZaAfhFcR0F7hdaFaaJzPzZS5ZJaVJIzQ+Y6XO1GtkbFEm9knU4GpbYc62OniAN7gDsu
4o6mW3m0UrxW3R3Ba72MIPPGJAuA2B9UOe+eDCAkZ3WNX+VsMx1pGCwOVIr/be96irSJfOObARN7
0dNPLvCSqp10jXLz5ygUXE0sVkblZV9CLgGOXGjJo2Pdg/fXeRaYgACUuHvGTDPnrMJv9kJ90mmB
7L4fJ/CFfZ/bWfN/XldVvYOIf6XxyTmW+Q8+KDaUo85GRYY7YBM6HalbY0DU6T4K0NKNBX49NWLx
q3mU3JjOErjYuiVClUgWQRsZPeALCZj97fA6aAwtMp/ikO6fP0ismZEML9nKSGJWRfJ+lalYTMeC
yhHmuD3b8zitqMk/QCQrKiJZTVC+5Y/SAncZ2mAx+gID5bypD0lb70GovlkU3T+o4jdWpY4iwMVr
NVc1a7lCPs3nRSDlQRjLPVyDwLYD4yzgYmBPLrQvuEHs333lBWVd7+t0k0IKA2LEQmuAAJDgPtiI
xnr6tp5HFdDeFEfYJpYTXGfVKUbG0BMA7YWt/SN4w0FJx5sn2NP/HE4sPqAtgsz+LcuFcN8BEGhH
ljhQx37ATP8ELb310p2XzbxxnqTVvCNzJOfn+YJh2QBQi0XPkdYqB2BpXYAnK+8JBOOzPdLFvdka
4tIhxpWPd+1IsS0Qqk1IxG+L8W25q5KKTMbtqlZRH/mDzp80QfcFiMHNgdaQAwEWY2FJnh4DKcj+
TYrC/c5dFj3sLeEp5q3ZQ/YZUKm/tOYIX/22tYQTvg1RktjBR6WHEdT6plTQTcOn+cvOH/T/SQln
51iY9Y8cZDgWGwh2YU/33SP/DdBUGYbPWEC6YkYiTvtHKa9ogdUdxGQpSuczAJK7Z1Uck0aB3sk8
2x31G1rteAwj731tERHhkBFy/cUYOELJKDcaDjD5CuHeKcuoEAl25QfXg0fXteQ3dxjO6V/nYdMo
ueK7qFEv7ETmJgccNQ7DqMMPZEWZWwM4RlJw14X8wvE4aB2MnXhKKjxhfGdYeyyTiFgtsQZ6kt8m
i7uWtOj+rMKIV76jBmLhdV6p2rQPNBpd/nrAii/mGmN/ocGeuJcbcXHb4jOd+x5uHr+Lk800ctrf
Lei9ukubBBne0WjSagX95UHEaUH6EEd/QM64QeJkQrW2jLvF/3iOXabsln6SrSifEr7LkXGsYp/i
wZ12TwsCSpfm8v8GKs4yrvKhNeswZ00YmL1fHfNFM2D0qYeu1kusggM9SXsUNl/rIe9iO5suzrJV
/zuv/Gn6Kj+hLkr1OjyO4TgfRFVPBuOBfscp4n6oTzMztiQVK8zR+tsg3ASwFrI7c8qDLdZ8jPcU
efMv6W9PMw6PVpxr7pHYaY6oHxUL0txRZsdXDCW8YJQi0iASoGICx/OQ0A6v09mt1KalXdIDl9K6
u89Ug3hwJPQaC8maw3c8euUCanIoF40rFUoPWy2xNrUIyW5QoCC1xor9Q2tOzya3eAlqrDXxBJdw
n9SF81ffKpqViz4QBDQUmw48rRz0hbqFRtRfL010cf9FPNzQu5APiy/XVrp9Y/ulBhIHV4QZqitv
p0ToAiTkQQgKc5bT9lVeaeg4zHmqr7lPP6gZWn92/2QMcO+XYKFjAyxecNhOq/3N98jLNam44DRo
WwFiD0BI+Z784qb/sPmZHbHxnLJVS5uyyKb7OLEoQeTqudwSSCzJ+g7HSCkchBmRc1m/Su/RMTcU
hKw9cAk9f4/ptHc7vYbvHb0BaHmjM1h8dgpyGo0tgTF3go0ZveaAHHO04Wa6zA3Rlm7kRyLtigzp
KX08hKBeyiqDS85Gj6kZp0MYFvXrmc12sPQCF9AEiLNmvORnaz2TlHmp+kl3/frkvYWl5UcDaiRa
0l3N5qC0Fu1q/BI9kqA9D6WY/UJrR7j8ZFD5eM+VaTxxIptqHe0UDqr6rw5uEWFRyFS3vgcSH0oy
54VWOhfZVqsNMmEE1WnadsAKsC2LLEa+NbZdqtiXjwQvosdJ/LvJq0qlHBlWDZSNkkQNg5qSeMV4
sKNPKuQJ4aoArXMTcPKNvwaJoM09Tni0xcrlhlKIYtmT2xuLvH3huVdNu/eCmYONp/pQzbllLoOO
Ld5JmmhE4vMzhocOxdtU3ixKrptVBpgyTHigV++t9RvEkfsiUmao+4ET1SukkfOg39EHq0o+ran8
M0YttIK6BliH207lpcwBBZEMYNZ4IqjJi6SVfh3XtY1mtXFvcBd6FlB6rl6NShz5qg7RXTWrzr2s
yJjcBSK9DT00Iq79gar82fOdFrfsAIKgfVC9ej+1y7HW/Rvy+e9S9qyeY40CL9n8uH88wnzdYEdQ
fPEf+hKnefYkx2rL4EqxGznB4LSInDRkFT1kDlr3Q19MIv694fAkAkhUKgh1uWf1ntZW3AZ3gmF0
NtAX5CzZLUtPgN0MZ/X8uTexVaAcu2lgDRRIs4rQqZcnmr1QEni76Ssk0KnRAvWwFIPm0Zs3+9M/
6cScvisqX+6nOEI1fIB5Ha4xVTjJ832GkhU+evHL81PQnWupjzq1chilj10RUycZb+LOB+BrSLmd
HjzNcTeRJoJDAfnBGtckUaMf0dphX5i7LUoQIV/VXQIckQyFOtegEJEDWteWtnTiM/fEJ8GaxSIR
chneL94cQ0I9tadHdbyVT8Kw65DEeUxGxMJdkVEUduzjUfkSMTYDeyCpCWFKl8c4mkqaKX53dKpP
2F0eQYPh40MZuyIYv0CL9t2ZLpr3oQ4vWevkgX24XR0W7sI3NzIbnw9tqUooE6RexzIotq+u7inL
RBRLwjaFh9N1DITKBbEkSALx2ACr96zl5zvI5d+9lQSnofB/nmJ2OFj1LqZTrtHXnquSVuQxYILH
UeuEW3tJtbnbtYR+gx61rLFWznuampzthOkjZgjfENkTlpRJsI+3Wau7uc1rvlAtY8++sqv61Cbk
C6buaBsS8tGbEAmst9Br4bzDEVCpwd8HKqNh1zK64NxVlxlb7vcxkrXUdYIEeyRolLeRbpj8/9FV
0LwENxOZRSQ7AMoiMweMZ9lh9O8RD9Yrq/YUyuDOhEhUAancq5MA86/lLf7C9k5fj1H+UG7vgYKv
HvJWJSZv/DKTqSzgs2r13PBsyWSJM1dr41qtwRAKXQEOBJ7K8HkbUEwyTXycAwep8gwMUE3k02D6
Qzb1/juPc/+S4k1+Q5G3uSyV9YSZsGuq6VtDNDN0m6oMVP9QNC7s5Pk6uVyAtO9N4QfzUSG1NPCT
nUiMaTAkQ/WOVqfkwHxteEE6HUWyG71cAD8/nCu0N3pPSIh2gGeO2FUWkJA023cnFPpqaIgyiu81
okytWJO02OmVfYIFEk05LKPruW4Aca8dhFNaZ2dQ6IrVMe29H6l/JknlIaDKxmzm1QJUr1a5OCpu
WjpFmmOSLpKxYIa6vf37I+DUnRAFqlZeEfYruTFtNzMwOFTF11WeiuBlAIM5ROAznb+TNmWRJyj4
n820yFoqHblEae0+cVtT7DBfZwZFfOANo/9AKF2+GyCuPv9J4DFpEkaEpQj0RLTmc7H2G8KeIh+t
vwHkOoG4dL5G/QcrRmhnleOFaSWUeqj2FyR99mIB6e7B5/gAYkTYBviA3NMFp3xxi13B9DDC5mcz
iwMcv+67QNOKDyTZ6/tvVQwgra1lnDEUk45K5+4KZapvrytnucgHURFvbTboSrChhVlns7nCYaI1
0VSBUZV22n8SOok8BMV2CSn10yaBGy9HZb0mR66Lr9HQRjcmDLvvUjEXiPuuy8CgTogTkSGH5uDd
O1ZOiovE5KqbxFdj72JsjpGRMNDfYggZNAvW78UUvGqHwNCULTnO6Vemxg1cjtvI12Ps91uh+YbY
2W2cvZDdA+dD4u9czmtR1nGBXyUjpoOUDmxhYuDiXRP3DACSIUU7erYV5hScLW1bc67m8UzTmV4c
9CxQ39naNRcm0FSLiBsE5J1pXZ8RzNyDqpi3jj8riiwVleXE4BYMJup537GCHtPFY1jSgEJLpo4t
TXsC1gJJauHQ3AlWonVk/GXJmGpYQNqN+8w3v6EwHsG/wQ/+RdiC6XVF4uoz8g/oQOb4QHQ/XTZ+
o/rtjpM4LUpvO76m6t/aur7ImuiAD3UxCeGL5IyjNNIo5OV17XU5CiDOLuBPLO5R/trnjhfFjyN0
UzLoKicLEAe5Jpz2a5/A7HkkKL6gT70k5f5uZgu3btkEfVDqK6Ymr8L3lyOrGIFX/eU/T3xX/BEU
70YfKod27tjRevt1eNvFfEnvJxZWjwHABDUlK7Zepk67fqMIjxNm2izLyY/H5V0wynMONYVBG1Ob
nUqDLe8sGN0Oi39XGlgDROeOjOVD8ZozQy45aiwat6HzpnixJVBH1MvfPMcHdg/lBN6npvn1L+wm
hmIHz5p43sOwl9y/j73REDzm2KKkkelL6gQvrYIi9Jz9pZsB5nmHTSb6i77gJ7xZGw8FBz1ar3hm
5SgQlSVSoh7aZh8RlWw/cwhTUbzCUJ7ttcY1uqyD8M2GL4GABtjtdbjEXP8oeNdKHq+xgY+yvz4x
xyDIOrqlqs0mdU7rVJ5y0zFdCaPcSLID7kZqtWmYFKvQJClevtFdQz2ouVKSRD5alib5h2mLaV96
UyEx9c0LRcPrJe71eShLfRK5ViiGZxXZyCKM2rlzgmi0aqlKIwUPsBjYh2j88TpPnG7yRzooItcM
xhj4HGnc7T5GpjOILnqVRi/L7gQ0fy59FegM3CSI6Yk2R7Yxw4YFUS+7wQ4bhvBaz+7BG8LNhE1C
4kZAc6z5kesIsiN7u1qqpBtX8mMVxpiqV7/pPO1SDWD0gweuH1tqnwfTM3j4bthfghN0eKSQrYih
lrEe8Wstpc1T7j7KPNm78JtJgx0YoV1Ny8WjAOIo0VFFxD+7itzYEFL88iGgfgzf8OFP2TFsaeZw
6Ddnip78Os6qw970o0Ue8CainHL8WEbWhCLHY1CXAa8B1kYbKsvB2JHtxpnCo/ylv70jw+dIDMuk
QTsnOQWpazUZcB0NCKu6+42Z9KINoN5k+o9/0T8MrhQe/GSnBXRVoFB1Pf3eA0Kkj1AmzetEFjWI
eOaimtuwJWJu5cdCTDZU01jIQthX9QbDjdbyOXGXRQpE3EqFVi5uMlYgHEeO94Ve+H20KeUvs2hz
ByS0wzjLIXozND7Swyo3Ap2si+mmSdZXOdvZiTgokM5OyneQVZI8ywDNFs+cS3U1xwwMkVHoV7ve
RJcYxZzr+oKugCbjxYbNPH5P0MtnbwFBvTDEItjNy0ymuHpnmN3AFzKJ51yrxtflPUk4WnEUJHMn
vtfgnubNpnnK5bcwnWHik9ovmrr9ZsgRb/H5jQbKXjfN0WbVvDjhZXDBHmI6nee4D2Zbhw+F69Dq
M6GjcR1gDOORUjGXvH2xYRZWLoaf1eSAe0D0CNqouXrFUaLwHUMy3XXhqYwtgRhKSQIseNE9GJPg
Ptax2D8xpMJ6pEC8qeM08ykxYifp5l7kFsEZwZRn9fU8xGkoVQPgiqS6SZzGbQP1wPwJ4IZvtJ1B
3q2VVzHfFesy7/w4gBYNy9OK4JmqLcxfVssyJ4CS5IcKbAsio8TWEW/gemU67LnSaj79/1fJNd42
jVY8fjM8b2KJjZLDfIxTlVxbCpUXejS1bMCwNfGpk8YeDxEjXjTEzFCX28ZLgVaGbtvoVRO5ayZT
8JcluCAjIstFAOmFwuebVZc3ykdCMfipO9fXtl7/bi3snaEHx5q3fdyQL/DeMGaPJ3EHbAruXt9X
as/eS8AS7KnruRvHUAHmYj9eITr9yt16A/7FXb6IxDQUKCywsrxH0sY5jgFW5D2PiPgefwG6Q8zI
TP4e6DxYtkDXdUHimumPLk+MXzaDHkN+9Z+OPF3O7OIoEVPX5snKEZMAOQpMu6WHuggmsWCqxMJE
QmuK5FcA3XTwbtst0D1JMXzaWQTEun1Cld2kLO/+YUGkgG1JJ8lHTKKj8LBXw4kXQ2XLEnFV1UH0
fd/zssclx/xqv7SDWPVwfD2q5AKwOTAObZICPpmqk52ftEKIPUes1bGKq/dCfVk1HrLqiKgG8Y8g
Hdi77Gge1FMrvIWQxDOJ13IBuQJ3nvszvSzU7vR8uwQSQcEochwiQ3yZtXi5KhtZc7ODBezE51cL
K1SNkB12O21jut+66iyDUcQQDLzHdSUbS8ye+VguGT1f/1bEXD2olmLAChau+z2WK6Nd7IFm0OrT
pP8XENJhmwrv7kBVZt6TV7Fap2LyjOu3PaTszxcwbgh/xNCT6147l60uAC0Ym8rio1AmgIfREM/e
RtKRQsIhGAK4j581DrpqiqgHXYmKuGp79ki00cbClnqeVJ6dl3/lhPoQnulCmUx/8nnNQNhDbsPa
RPwYSZMQ0ZyBONo78YFJpE/BFyl5LEtbX1hkkvUgj+hOLYudfHvpu3VTjTTWI8Kt3ij16BOkne8n
/t5HQvP0mWP6KhPjyMqumuM/u+8/4XqjAqRprffzSTd37YhGXUkH9Zxkiwxg0jRyk8ov6mfzWSfR
9pq57I/f7HLFdf6gq0HUxCuxc9BwlDw1q9R98jImPx6QsfuYK0oBA2bLedCoN9y3iDydPK02WPki
gcUZcJH5qeqtNF2ZwIXb42Spzh4AmNYatQtcZFHVO3+nbIu+IYJDLRMxa+KtMT8LY/0DKtNlLirO
D4xPgqiQ59H8ses/ozk7H6g+BGOMuTM+77HYSaei8o+PbhcfqB6pi0P0bXEZRvJO7KWqInXpyMOY
MVID9PON4fJGOG1Y/hOj9wp+XE+lWKYfArUXCOow9VqWOROw7ODAklnE1O5mDqcoSOE17lmTi55C
kRwhB7LLYFdu5+NVsXU4nGUhDaPcnXCbZMAdBLHnwL0S7ktNlVkQnEpyBtvdAiWQwAk3CwHVpTze
j+TZlCZxROK1G4XcU3w8iUUx8RQyhZ0Dq0DiCdfBe+54QWjAWH3T9rRgvvRii2mSjdPsRYJws4NH
TxLuCFoWRDJMJNN1kJtbu9SFK/UJaEqpYoO8Ia09OH7bYKFL4xyyTd7SaOJOh6SoK/l9At74toPZ
ePmvd8EFYAJh9Qk/vWmgB0K8zSAVGDCboKOnJrQqnGKpMgI+XQ0aYTpzc3TJyoQx85GB7Iw93tdk
XBrLY6DOWqsYvvzqOw4xeHAjgZx687DKCOu0zD06mXfyq4x1x9c2Bxnfkeq5x1e+ov1UmHohFNCD
+JoLhfHeci35N+kS4tEjars4eexWhedZKvFMgyYy5YIKi7t2DKMcyeNmFFemkO+jSEJg5XOb+0sM
lYB2A1kfeM9gVMy4Ewnl/Ig5PDoDKBZIQuZ4UrZ5TALyehsZETtsg8TXbIw0cjR6jp/f5fVx/scB
Y2upGgQ9njyMnRAQBvHorQhNBDmmm5cqGyaqeIkZZfZLEIRV8WqGEHT0I7Pm0MZgEqbc4oDw/MV9
jeHhij29Zfq5RUiNGaDzUO0k/gyEeplBwXKm43HcDTiyKqwl+AkBa8+ghdfcVgHrT4USjf5JEDab
wttcx9Ht1o8Bp16UMxsYhJBz+EFVRwMhdmPZtxd6ppYyLXyWGXGc2wX+7Jya9BM28XKBG85wBxwU
Bh6ImaNrxxVv6rgsLEi7gB9bttu3InRTa2jnOFdgAXkmrB83RSnBr0e75ezxLoip3xvAiUulnSkR
vJkgydM0aq6FTZ1HmNFojQMm7Qh19QLrdKwodUwF9i6KIv3T50v+dthnH+m+5Y4twQYixaWetVvO
J+4vZW4ek6UOu2lXwkGiJoqasMCcgseBxrSMpsnUUlMkWSGMOnjbcvtgdBoxB+URSoU3CSEezJGu
lqvy1vNmdE8iwiRnzfR0iZi9ZylrCxIWNjLHLGlzpyLs+hj/zCDqwjeKNyEOvbO9//iJgjl3gX3M
1vz0fGAWQ84mdDVdTD4vpND3w/fbUB8N3t5nSy6H19PAkEL8mSFjyOoMIgOs3427MA4npGXlHcKh
R6yO+INg1u1cFaxrXUAPbZw97b3ph+1UNNutoVxpUJCZMtvnoZozHd6eRd6QQ3dLNdl+sOFJE06u
wSG+7EwH00GiVELtT91eXCpWQw5N+bYHxReYKc+n0JRw2TNMEOuiO2Ah7hrrlLeTK89evSDP/G5g
y2UskAwlFy7b+xb2iE28uF5s9HrYq68qr5KoqHE88ALxT7drHcLBvogqxTYuS13nLVuhCBWjl+Ba
8nSchDoAG0DKVfuhooRAYNxE0Po/CqFCBc7WTO376FDNw2QqsT6LHI1gnEQM9gZ7ir8C4mMG95qu
3SUp1GY+yUOdVESCZ87p1jzvHyVXlQHz3Px9E4Ap86pPItgi1qVxfyuR4Gj/Eb6J9Dca+ZYgxiHr
b2HEsvFWn70jQexiA6qmPaKybeJvzD07dmPD3zGF6l41iWlERoLOlIQz/GjBBF95i+YwrlKP4Ilw
EjfYQKF5h67w8TxdnJa7+hiuDtSe1zwYDR/YvW/+yfPV7MQ//QTzmjv18i1b9cgmvf3HTfgZml2P
K0G9zv1meEqddPlHod+mRQfyAyWjqpiXEenSPNgNvIybnFfxI2Vf+tFckA8w5RkZZDqf1ZdKVRlQ
C47QeKBfNm6tKogzCuvhFX+4gttendssjrfyMoSVp/eYkTqgVqqv2opOy0QJTz/RD7RjXCzck77K
Jt8DBE4jdA7m+padbJr9lnEZy9QgIi9oDqYVRhWEVWYMWIj3+RddafjtpFz/mPyVNb1F68O+7TSz
t2Hp6+AIptGUvjHoLZq3JrPvkEWmO3Oq82ReBrMhZ+kjNheRxAJU0dKUPVQgIXOASLMZkcfQvnum
3MdmURX8UyFuO4quwQpTnpYvg56MCQaquk1IPeD8238QbJC6Tzhncx++Ec0kgvbMQpR27+QGfyq3
gR5qLKaRVtOKHYOXgQMQRjI3LOHQffxOB0J0ysyWHi1GMY3qjo/y3XCksGpugiEFsbkSGg4Km4dL
kWcOhxfN2L6d1R6JA3iP7wvNTB8yyTDKh0oLfLtcjfExJUww3NECGgdkGB4f+6WXbxC1dBBrJy5h
TNf4QFhXd7iG5qf2VF1xEvqF3vIoU2x7vZvY+sdm/CnOgHucB8XCvLmwo0ALLpuHJVx0iMkj2lm6
1Jd3nDsU5p1biF3KJ4kMJ7Ha+4gxNN4bqYo8qhbTrjK1ub+CH6u5HGNQhYfZndy0pj3B9NPTKVcv
9n2ukkW941ApnpfZ8FGJ0Zvi+8W5g2S2vf7FC8H/QpypaMidiVMvArKoPwW/u9K1nWffD3PzVGCC
fOKd0KDAJQYJ4ERqLz/LO8G7Hkip8yo416ob2aD+aapDW36Ntq6B4OgkRX6ANr+mO5511IlsMzcx
XhDGduB9znZ0TNH7bYthWMIpJBYSQ9w9m4rH9ePBlfapry32B96B6udCpENkRpmreK1vZykEPAkT
aLqGtlo6Oigbk7Sy9JrQy4wN2UgE0ndHwYPYUMkboEh9dUPVYYboJc2A1mU0mAwe/6BqhAUwAmu8
4TJbV/wjtKH+hUvljFC58IRAf9EeGhnMmN8uzfE8Ds4vQKuyUSP3EgRNTEUhpouWEiF8bc22GRVF
qn9taT6DXwAe39/HlJ8GLh5lC6rAfJXWjq0/RS4nYmKuwe+Oz3bZseXLtd/jETKidDILxUY0fbJV
MarHxMaTdDpFLkOtZo4nb4h8mN9rHK/MNL2KhLAZvoRUWKNkoO6EM+XmnhcSCzx6SFlN3Z/KUvqG
GK87cik64P5ipEgM5YMaEEnaC9xzqYhnmmN+mmhB/V0ojy8kgGY11xNLAkX+NCdzKYPsdyrT9cHb
RO+Xa9x/VXfmIo089g8inMfpehkKA1+U3r7CDapU6xenekq1FUwfKlDJ7PpxwKO8pQAJu7npm6zm
emjSed9cX9217JMYb0gdeYKYzBJesp988l+S/4qlgvl6jGTWSnFkbbA0DG17bQ6tHzFVC1U/R7Nk
UDyuxBzVLSw0dFBLjB9e1VcNPR7uF/xHemPKd2MfdJpzKgjZCbpuEllNdaFt0DmEuQXMm+KghwfG
9eyfUfCxNmZwImQapqYZKbF827sW5IbsWIyvCvCE+DfKdc4sN3nTfBQIsXPaIJr0o980NqIyZofS
ncElKef0B3TU6XCH9aL0RCwLI6r+05OA32vHVS/bVHaN+RRULY09zmNUxYwXhLJ4oYxPTZ1CVy+J
047yfz9ZMNT6N0j5u7TDdvcOFv6aW/dvdP1uCS9JsYZCcJsN4ZeztkWJ62JisMAuZof/K0accncA
pHH4xO6PqdusHNqvtYW/fU0MVl18X0/6rL+3m7mFTsGlaY5h6lPonhTmhROvLlk/nHI969qTf5pP
AcdD8qFG7L/jyK2aTvjnujNCcHSPRTM0y71EYOu4LhiAZ+feLA217kiT5Jx7+fS4sAidLPtzi9VT
0LSmgni4CRE7sYCoecM81DrhplnXPHqeYYE5KoQRPVyw3fBANo43F34FAWbI+5pAs2h5HwAnGtO0
Xf5OvECCL/t0WS5NbN8N7X9cLVTU7BAMkHJmFBXmCSsejFvftY2iFd3EPXkY+jcMoXqzWJpjxgO1
gGDOU4tyqdUyh9ZcmZIcRKd9UDO4NddACkXEWkhuNX0wFbs+itObMssF7N96k2z+hApnaqMZjXdP
LQLZai6AeBV9UnZOhcA1k8RsylrIeA2vNiPfP6MUUuZ00gYkIpqyf7UCZCoJMHOJwJ8VTIl+SXik
Vz40gFUVhmdT760hcR8mXfW7lI+hyhUvq1DdUF+rBIhc450tlg/MhkabqmskidmQWkEaJdllbSeg
kIp/FMvCuDKXpOhnsR4yHLKW4heycVUMsoY8j0K3gvZrHQiJte46U9CZXO1QpUR7tJOy4teAeg1S
P/Jnn89jnPMmuKvJ8D0IiZXFoIZ9h/V4x/EH2iUZLkdCmgvAg3cPYRFpDzRVxiS8fwbCaP0HA16u
ChwYjyRxstnjUiaMjfVn/uNoTnFoFqojSkqvQ5rCrKEGNZE9lluKnZsag1xu6/mm1jHcMHUNOkSL
AMMLYpeVP+mHJ7gQGhAoThJbhfb7vaGRx0mSHEtL5qC6LNCdOZ0cATBF+IhL3eCjIHtkzqd7wQor
7ZNsTHlNLWoNMuA23wqt51nHJMYTiFlyUBXA77mkSOqTGCkyQXTWDAvVWoB5h2GPfsj8MyQ1aQ66
wXZhbkHAtHt7MsVnT0+TMkSK2+dQVrbUK/R8fkTlU6yITcwEyeotpQD3xQiMnqpPXIb3i/X3KVH6
/1OqSChqFWr2gpAYO2XyNS1yGL5vBZ/kBv+9ypj8Z++3UVzv2IUF+IcrthY2muJ04rEicEtxtVsT
57JigsN/Y95DTuj1Ev7YCD4sxUts+vjCiIPl9HfYIS0GfNv+QnkMywgnm1/P60KkMKrtgsqS8mjN
YqBmD7suqHsuUxQ6X5qw4jeA4RzlmoBU6aqoXNN5LnfCdCQssSWuoEvrdIJUR/d9Plh2Dxr9hMm4
MTKkqigLWmRd5XDm7diBb55ERKQUPX5dmDziJ2YPGCSSx8F4F+QMNJNmqUbWhChnFTSC5xdG2Jsc
3BifQ886UYv1Q4/dP4evrUhxHeCsIfq0g40gIh/ASHx3IDMsS/PgK1pWurcHdvMgZRIFmK0aHKmo
ZkxhJG+U+SNCPnk4GV4R1EGr+E2gek372udAmE+XyhrZuttHjU4Gbn3goQ9FzRqBuFB+jrqpwkxo
ZZQOhQT5qwZfiF6GTRcVlncWGPXRVNoNfYBr7tj4+n6Xr1XTm79Ug3RDYpmxBuIcgB2adXzQmBZq
2jT7eMHpLt0y7rOdPpfk+fC17cegKQ5dFn21Zci+z/T9N+KOvpyV6lMxAukCbdzIkIk3iyRfLUhZ
N6EQRC8nBHpXLcb9te7Cp4p2aBZAoM7LqVlw27KeGy0icGoSxjkXOkRZQoq4X/qGmLwFMGBisDCv
VGhzehFragOlOL/yy4QjuzEeB3mxIEVOexhtu4QfDqDbUQZBsv15hACkSPXW1MDLM7phFE7n3ifG
tsyxlpTtJ8DhLry1BtGdHZ7BQFVrjL/qeQriQHL6k3PMPVMpU8Pt7/n1Mq1ssU6zA9mRWmH/6aM/
0AiO4YnpGpSHQA0tH6TsJmsed9T48s6GtD2sVQDEA317uUZqES8QhioGPvi7mtoDJEW4ez/pa0q2
GQrV9UFx7QFqt4GcJzql3G54DIELk3hJLltpYH+x8oiKGdSWqcBaUvKTIqHM7nNZQuOcdXOorwbM
46DMjN525OirbhmosjsZgFoh55WyzVZhLX1oytIg9Lw9dSdhTsXIqFF3GO5L0Nb+54xUsHTnKSOF
6/UnzUu/xG6BTCDZIxdt5Q3kCRZvv/7EWGnCFpO810k85pB+TzbPJeR3H9ur1ClALRKDp+tJ6qru
0CozNtIqY5vYJtEM56vUI4STONMdYJAh8BrkZ2szvfJHDWq7++7TW21XmQWYQ/MgZCcCJcMvFaK4
yH/wcGy650qPQ5+h3gEOpkObuRNowYId9g+pJbbi/vIqic/yf8e8YEDyJhEUx+8Bomko7DjtBzaV
F6aSOX7LfXbK0sPZC8zEp9Xob3dwZgHM5PD8QggrKwEWoxEuKXZmZMgajfLEKoCXJpwiw1bPGyS5
nEGS6xSPZtqe2xZ467nddIy801mMBhR4PzQk92h8dERfgXWyDA5Gg/9wkCQjCKSkJCy44QVjw+6N
wvkGrwbRESZumeAI7cF37J4BKKWXl0zqcVhBkCNgoKCBIXZttxQXJUaK5iac1AbPjJtG1u0fo3hV
BzGPa2Z6REbV6DQlw+VzQZXj85fIkDjGFVzyRqsZB88CaqMrrPmhiIaB0ihqLCnV+FPccDaWzAzw
hYtr/Wajv7GcTs47lL9SCMLntaANFq2vDNHK3G3o90wYgYzIgkpBQpIMgMr7GEaprf+66H24FO/b
X8yutcfQoZn9sHOniK/HW5W7ZiNTYfr0k39bAIx9XSRneMDHmJOa6NW5CA5fHweDMDNy1a+psGaW
DMmXN03Owd4j+yAKi6xzzm8PFgqblE3EjQ3p/gXF3RbuFiYXt0uYL/oOYxhNhc/HKVKgqVsXU0S0
w35PfsZilF8cgYuGwGvqJrWtVvRiLq6j/crv4FHEg9Wzh92ViHbp3HTuFMPF+WL1qygNan/u7Osz
yvxUry1zHWBvgTslGiboGuo99Q5vTa4ZsR65kvA9DSEq2A4Cl6TFy5AobujqgQIic3sSWuQj4b8K
8O9VHziNY93O4hZnhbkBX0nEZIy14yc2vJ16K1pgVFDDl7TBa6iNSP3Fs+esGgGOb605Tv1GleNw
U/TRce5CxAV+WyUNLRs8KxfM/H1CD1kOO5E9tHTlzeS+GoDMeMQJk6lNsnGwVhqpgAS5G/ijVidf
zEQ3kfXXC98rpsr+XEB4tMyCvJSPoW5j1wVdP2uYcgGoWJjyke0K7ib/hTQXFe8q9IWLAqrRglE6
IzilXmop7QoZwboqpvMltTHMEy3QV28bnDxy+8PVMlUACiaYIHij8Bn5bf0/gnoDFhGMKUpQZiau
Vybcp3LLZheb/ZN/BgvL7ZmZOO2BPn4wOvQyHYSfTdhswStMwsyXA7xdpQ5mDfL+/47PpvO+MOI1
rJ2UA4+QppW6DBuQI6+jHyqreBYXQUO+Lylv7TX3cDsWrX4m2lsbxZQ0FxTpKpU3vdpUlCuX5Fk+
NR+ETvNVNYhJbSmSOWModbXk55zAYfgqZ2YezSmb9K0nhvkLXy9An4RuFSr+BdED68aFFwxRDmcw
N3+yG7IkM7CIOTZS9AS1enBlOrqSNn212uASdU3ki0e/wFmyV374GQgZiqd9ZWcL4qLNW5Mxcady
s/AUEhb/E65hu7fg/YZVRK0R8FbOezbKldWeM7MIAKjgAWmpQ7+2dFshcA1I3yDJagiv+wn1o+o3
avz7DLCDhYthYpXM7JcVPATPp01Ve1ti1U0N0L3Lw0w45T01M3JvcXsfYdNK9YOgEbkscosB1tYR
Nr2E1FmwSmxLNunNIP+MrbUxt0EkQOK7epkdQi2X3E9fJZ8daIiA5GqiFhWrv9oI8cG6WqhmPkNl
8qWnDDePUH8GidvI/mP8sbAkeTR285In9LsNaVoQ4UEfjsfTP6OPPZhcxYryLEL9tlT+UPfFqUhP
BYSfFXO3b/ef2c8uLvC41oIKqKHP/h/kiF3/qgCsJ8Wh0ixVLXyFDhnA/CrPZ4DTFIde4ua9IE+z
anxscOaPmYnlIJHXcKiBgiRoqKqoHU7MrxGRZeqIHGLeZ7IM2Yv1poQ5d3zOlw6dRr7U+FjzpAJU
O+m/hr6rhZqsSDAyBZFfMuy5dRvtTdlX+wixcXLtbEkDN7puBCJAzjiRjvye7Tk6bd5HSlTW15Xy
6cmB/5CKtAn+pXK13B/mQEsznSdE29fAcK4d0JzMAcoWe6fBO0EfDH+Zbd/Zlk254fZV1P86QBLI
kmEOIm3h52fnWAddVZpBdCkBxU3kd33kCkMvreT9LFlko78/L4PBZ5KXFU6kyWVOCCrSJjOJCxFs
aMNQV5dw+PFJo+APxvHhy1v2Wfb0m/NPgkkFuRRgxndX430r109o/iVa5L4Q/6k62hLsXKaeGxvS
6Dg/Oo4DW/2KrXGiGZyXpgIKIDHdgEW9wdjoJxKpV3yzDFaovv7TpEpMyj9b5hVxrO8T75rGnwsD
PFuqT1PCUqc446bnZ6OB5Pde+zb+Kdy2NX6xTe5fWk5cWiFXKChORmkUNKzgJjhxn3tW5F3taq26
T0qPGnf+/NKVCaIktmPdHRMXwoTdV+5pSB5+EH3qmeJweKdScen48ezXJlCRcUGBmx3e6pzLNJFU
18F3QQvLA0hPg4ZEfX7GrNDGO8M+DS2WBNGTtpcS/CmOmxdw5rSsIxrKwFYkV8Wr48QKVFVXhTFn
3GgqkjxKJsU5m7+IX0mdzSeUSw8xDmOdQg/iFg+b76xwTcEWv+3tjLtgaNaXuAUxHbAXe+b1W9D/
oE375aqgKHTduU+T98JZOQJeYnBNE04gUIv9X2l1Lwe7n6DlsjRNXRZx8zmTFj1e9i3g+nbfH5D+
/N+8lN7HiupoCL6agC6E3ZzVIHJoaEgR6eljq+1LN8nsXU8lYO3GRAl6RI6Nijc6xposWesr3Tz3
yv8UxMXlwuxjTS0dqd+e8X3OiT2hNWDSQ/kvLCGETqT1wxhEGsO9jAZfOmELeGLoFNoOWY7TsnzD
68tg4ExJ5AXDXY3U4ggy2RNYQi4MYGDmaZQ18Z+JbXGBbJv0L4VyyozPy95CZg00UANj/C8AI0a4
B3/aj0kuwIaMf7dHUtS3g6+pvc6ym4dfXn7HHtGHZK1j2S3Sf3Ji8Cg506lfBunUObc5SFpsNBy+
ScY7+BRDSRHfbLZ8Gh0p8zM96nhc0Rawo2v4a9HUH1RIVU9TOsd1v1lhmQXbKQqSgglfJA2vevCD
RrlhxkwagkAiGnGWnm5IWdLLfxXjFfPySdCPgopUxRwcmL8p2WpLCy6UWDSRNA6FebbcAKQqHYQW
ABA2Hj08NajMOl4170L0ZqERIMt9+BU8K8HvAbjcrgmYDsJ7w9b/heiqWCYj4WZGt2foi/XuZLlq
ZOy23ifNI5Qs2n8pocv3q5lMvkASjNsvEnrgkPTj4ShKTXhM1bLK8on43L96cKaHccBLOK3jx7Jb
ZkKlCJUTEnJ80w3dXXOggmzQI6wkSC1pBAR/jpzO04sasjDtJYgY5xKimurcUAMiT4soZIs2t0jc
SIo8KLrpn2AJutjjINoZVQUfUgNgGZgtOZ9OjhmnIbtI1T9UlFkcDSZVQ2+GOkSWzZu2i1FZMYGe
yP7ea+vqVbAxLycRNmY2rH0Gh37MCbxzZu099hFvDNf4X3+wwR2sXyxVjlPlM2eq1w9EzmSroJ5J
o6vr0HQbQ3s02vXDNbAWjhSu5v3HEAMl+WBuDEZWeFXucIJKF9B5dLs1FUdQu62AFPN+t+4mAsE/
XwRqLHTmih7cSGaEdqsZ2tLbUA3+I9ezPGd9FaCqG0Ol/BNU0imAbpzytaZE+I1GFbJnnuzPYr6J
ShSmqJrd9/DU9hcYMqgCWuxxTeh39kjV2MwvaxUa9Ba88C074kXXhD+4bMGVyrMtN0UDORuKCiO2
6fv8sXVNBC9wfsZI3vdVi0IJDq7FTL3l3rtNZhv/HQAovqeuC3+uWXJ0utv29aIbX2lAJw60hcMy
r05TotnCNEts/1c/HQtPoNsFRHT4g8T5ODlFENSz6a7iBuXRGU+gCrjeyFGWrnvPZOcO3XYpYi7K
hNzNAxhLMPK9CSmSf8gnaw5YQlc2Rajatg74XS5MXE9lCZAJg5i41lVIkOllgFeK6aaLHUro2m1n
ZssYo7XYgI/EAL5WgaT0kmCs1lg0rWGNtP86MElhkZAU7I0pv/TIvzBjhT/IDS3b4DXsVaMjzowy
/HJckWd+JZpRcvgXavvDqWBrTGNLjSa9ls+D6UZC02bvzNpOhWDCoxI+umdEiOT2e6jviA2Q7kOK
6abjlPRH/vJ9tTgt9Lr3+GvsHuMnU++CnrU5La8pw9FfpleeKZbE7wFAFA5IvQp4WyZTn/KNUSQn
ZJGXSh2sMHhH/llNouab55QnTEFL8SZeTKBoOEKZbG7O7MPfjxhCoQ6A3Sg9+AlfneTOWvOljy8A
GvvMLiQp2ovqf4ueeGA+jEzwwYiCvx+JHM0N0l4eLu6Q7u/z8r1U0xps3DDzb4N48GynIFa7x7g9
9VE0adBhebyKDB7UAh5FgWEj+asYwxSWsbXmlFhxyke/G6XVyj7VUJsh8evPhpxcRgBz4nsSTsnG
bKI2nXLB1WPUe1p2KESbKFH+xvbQA1TPiGjIOtmPZgJJMNxN/AgkkJzaTuPJyBJzX0l5X3+nhOpT
JXlOejNGWI1Bd746079a8JNkXMS8P01MViS7vPwLrWQz8KWb5Ls//J/F7KHKPJbHD+EAkDv06dkj
aHLLPNlWZ123ZM7udjt2KRv2nhyDhZJvHqV1b0MfPc+MRyuFmP2MnaxXnRYJkPwUbiGhntbeMKYN
4pLCzcZ0poUibhfWYg0Bbc4vuhXQeF2BwVG3G1wzyWWvcfppH2/BcSa8ORehVOMV5MmpNmY59dz5
jbwy6HWdrERasdZKZs05/8gb3fLtkYkTzOH5MwG2LjSJyUkyH+U7z4a//nKy7KqkGHhmm6+E9jlK
WvZFXtQTNHmA8/i6k18K2JwpAOmWKBYKvhUgsk4OA/9n3apzmtuBZmj/UI/9EkSV9G1q+oSK3zLu
e4RJCm2F8VrTnexzJYCaGoFzb7hiw7jATNbWaMmKmlhKPIr9Xs/g6Kdo9hveongGFQFJwOmUcGs1
gT96rLI+Cz0rtc+swgn/dsGlMMEEhIs2SSnxfy68PaqacATEvgF0v5Ija/PD7V5k6qkXdUjPzCMk
OMdpKSs8oYPSFNUpVz9LA/JmY+CbpEhNkXB0hNCjyq1qtUKZiH6iLsjyr2+GXfUVKQnNfajTNqJZ
VtzKgpcUF3m4vOELIo9skg5MxKs993KdqIyAx0DqUL2Df/bWUakLPA+i3as2ioWP41XmnU6kBq+R
2pNZVbT2m2nVNKJKtlzC7pA2Pq3jpTOIJdew6dVhe6TBC2ZcV3Yvc371FOAEjtJ4d/bQzmPlUGaC
j6eSb9pY2Nur4mSrnfmN6NXUXF+M6oO5bB6JN74taw8gu1pwFw8NAh7XadXjhY8rME2U2h0N/uVB
sh03YXjCGFdPDMjjMrRjj7MsLbaYFZgN7YeNWnswWrMzKyHcz2GL6J6xSlypkcAIrpXjhhb0Zxq+
74i2YfvjYf4rYoCT9fdFnKg/eMctJmqr7fZv5p1DmUnG2IPtPW4j2O8OgcraPNO118Z39Uoi8/W0
6F8xe6x+FcVWORhK0MrUZTrxLD+P6h5pdXk+N58tiHgxj3/qfR02P9D8e+9LI1kfsxtPhM8ecEgO
/r6I24VmPFcdev1df6qroNTnDcv6P1omCpbopmmWPo2Z1RoCMujOLzRQ9n3FmueO+b7+3t4TM+uL
X92S0YyWJrXGwaJ3CU5Ij6c8iFdl3eX825Q+NrDL7blgC9Q9g5pD8XefqdelnSVXAEIpbtfMNlf1
/7+cRU4FUVNQSHd6wsI14aVBl61ZpQC7AkwYvx8sbLM4jt8KXhY40t2tXVbGF3TR0jQXubAZcnpx
EL9MeR6796AmYgGc59s7OPYORtYxkk0BVavF2Hxpfso+ndyhH66kX+HC5cEPQo+KAupdRsfnkPmO
OZwJsejtZn9jpCQfa9bj54bzNeu/zKugXYpYLu5jPaDVhjkZytqRTjJ+Twcieh9BoQAiTS6eBcn5
tbIGx8h7NCaPGElLfAkx2PKtaLxilRr2z3WuDhpxksUeT6s4kyhGr2hA0d9GyM94NZtFTQapcKyg
Ae1NtZJu9hyVXeULpelm2K7ePI5n9h1FNpqcpodTFu1V2G1hvmJiLt6SkFRn+kFqKZ3JVkiREx9t
YTvHyNspUF8N44nyQVYAHCXE6K88sNLQqdfqGOEqbcdJ9hyX4DRCwsMf4xFbd9zXxjIXMPwxTdRl
H/hpHjNfUKh1YyKxtmvkhCDrEBgEuQkBWh2JwLoBVSS18aSB4UZLJDLMM+Ki6nz3kK60OgWliUuB
LjE4+R3gupPGCMEbOQEp4yVyLW+48zj/fWZV4h5RbjcvKpeaNvIPPxfA4+xU6FGgXBZgAl3N4eiS
WDlQV4TpnUkAZsBWmjqyUV0SrfvQ+WsppV/YaebdnexxURd6J39UrMGvVrqE2aqD2QJa4peP76dt
CrUsjhLlpxoO23meCnhDnchFYa5HP7Q10rqriCGkaK12OTLa5A/Th6WNt1HjdmPDkS/eQwwE0Fbb
oMZaAA/GYMdNTvTWRtUDh3jX03Ao/tyfKwvIAcbZfjLBpD0dUEdPb4FzZzQTtL7ve41DOe21ieWx
V9+gDkDFGBtJYDwECGT5QB3UlmC8Ycbe3q+AcdQvyDeIL8exojlKxwfp/fJ+UvQTKUWV2wL2Oyhk
hYof+dZlVZLjtYUS8OKdcInSGpeZ9jLFXgx2b/6oE0RaEfw+T7k9EaAEpUBaL9zkrFd03E0GIzmk
+4zuMFsCuETbfJ3FkL5Lq5jQVUxZwpRRFKQ7BxcuTnMGXhIMSHoASkYJzErm0x9gGAz9BWbtfifw
WJi9boaidJlXCUQgltAaB1miEeH6Y1wmYIBDLP4sFrAugV5qalbEUj8cTWZmbUDN6ccVPQaC5T5Z
i0uoMANY/C90VQYyromNB5y/i+0w1u5dwuJ3k+ZHYcgaDgEHYFG6p0xcBf4oDgQG0U7niBxzUThX
hrgyoTTgZ0DdExXjDqvjKsbk9zUyLIWdGpWkfmP8Fmgyezen3aUpnRFIbvNt0dR4Uv3EzOMn0U3I
byOpJrtatNOgEzB1g5z14iv6BR01oSJeGZx6+rlwWFPpJXL+yXie2DZLcwwpoboUX4OL+00m8gsD
0zTrOEi6TxcngkLtCELLPSf/tytQC2RCxhaPm4Vtb3O+6XxhmNwLO1QueRHUrP6B02LTJvWKxpnT
i6H51xOPFj8NYkEvhyCCz18P4IX7ilhv79ceB1QkNOVCtTM+mIJ35+J4Fpywf2gnBNSjtyl2ARVT
Qu4O8n7dS5VvTVptPJNK7jgtmtVC9KQak3FUWrA3AF7tQIg4CCjz74y8JKHpfaTEVjCpjW79ROK/
73yV0AN6oKnye6y7yCaWHSRtZizm+48ueWzl0CFIqAsrS7U5NCSjmUaAODX9kJ/0LvnkTqHzJSul
2fnzsd5nEzjSzQJc6G4t7j0VA51+sU15PxJxmuzRAscwYTyZ9vR0fVantX9fAyWtbXEQRrHGMl7D
VibSLQSw68ZPJSa0lv8621iVlJAaDAYPVyEOMT07UyVS+qiffX873jCYownMHdtA9BdXrP7YdXUG
H17LXni3Y0VdYQueRysmR0Sq+jzQBba9D9Vbux/cOCZDqVdsN3ANpuCH+8UrJkOHLpacGMl99L4e
XIeOkxbvtN240+c093kua3qNbVJ4CEqEP2ERnSJ57Ke4xv9UnxPzjB5YfdYcNPQt0QeuBYtjKD04
Ef/nabhVHx+fQA4kgkcG0xEIZirsnsV7LtQSh1UFSqDw+hLGy1Yc+El1NlilPMCB3TcrKFu5FnKn
nYqK7BURDlRazq4pnRoZkDgQUQ6jnMsEbrIgYoa9Bg7hZ/YmqHEbT7w65RcuIoM2LLHzno52tNhs
v9pixyKuj0ZiVPgoIA4sgYZN6kfqj/g9q/MUfL+U7HBeeq9Rlj2lOOpTpcVf5PM6h+IcfHdsxtRS
Zcx4FN9ppjS7As/UVCnAoE/JresX+60i1ocIIzE6nGd2VyrLxGBMng6eGbTXUeEVwO6UOBqfU185
zIV3ig9MjQsGpLulurJe6TNHwwoZKjyK15nrha03t2s3FuLOGQ2GPV5U5FcLxnUihCMF+BPMmvjV
8YsrnktQdZPo9KmxX2HcSyUI4W7aM4yv8oF38/ZhsrzND4fhoOWOzIbCdb3ZSDTLhN1gDLD4hWQF
ygH0O1AkT2lJ47kowBTR5LQRr0MdWUBRIC2E7xnGXd7mikLBUNQdbPGw+/j3ZRIx890fPVKPm8u6
J16n8FpyoxGBppNqy0g+1q7/w6rVD4rP62YNI8BKxNTaZi30tkbb4DjiExvtE2oM+CXf8OxqHi1r
3PGiHwe3NBt8npqYrRQRvD+77H9+XXsv6dS2YwwOwCJrnJN60ciQmbkfM/WyhJhSwPZC+LompKFu
252VNbdV64BAYNo97zzfXkk+ucersEJ4C/6iZKm+Sip4VeARPlDyCGxvMHhbqDSdpdVr17bg31th
yR1fpcTXZbL96V9qpyuV+SlZQI/ZRcgNqZU6yYvJtQ2Ny95Wgfb+RtZqQ6yIXns3M07dSL14aCTK
EyO5YDHrOInwMP7dURxpa5poN+kM88zoM1uIXJ//9hn4cMzgeEi24KCjh4NGSE0F9RaXdiwoyERU
SUSHDmM2Fq86VE5k4+Qw59EUeaShcrwjunNTag9J7NiqMfxK0c1gO2Dzgmui6BQMfqg741eZBLtw
e3OlHKIgbVx7hlkLkrwEcYx4F+xGOcQN61DIxGHmJvGbyyJag5SOL0ETLhklIecMjhI+4uL1ajhK
UTeh9/XKpZv3ypuJzKzs1j+9SeNEq78T8oryRps2UmtoOfWgvLBG1PQ6WTIbYX9zshVO+aku8l4R
yr/2YS2EsW7F5pmV6zOEax13tpMS9uSFPD3wjV8pyhNhmLdmzSkw8lNISg9o/Az9R8Rfsh8IP/QK
nT1X2rn0GAG5uH8Jo6YhkjFjbTyObqX1xnedxoU8V3mE7F5lfwYcLV3ESSPwCbl3u7d9+Eb2KcqY
BFTeSU2cukdv/AVDiQXhIXw0h58gvOYQdwP3put2Duy5e5Gw++QoZbBrmvFmMVDz6rTt6oUqLdDh
WAsGsFkDxdDIQmU0h0QIs2uy4jwOf+Dr+Tm4Uxs1oX930s3ipATjlwslh5sDkuzWwzFb2kL22P7m
g+OI50dnpi1C8F09YRJoQvr73DU9qQpqiKaY5zg66bOptrl+6AGfYmIku5/hNIC7bs72+INtPT6h
0a6mMxWQfwuSu6M9ojE3zvGcW+7CzHSuwQII0ScX38yJaWBmrkFBdh62G7ADV3fJl8BNq+KkgJo9
vIQfrgW1BIm6aEX3Emn3nXv+deVva+anG857Fkc2p3mR2x9J03RFRupyWqJJnAauPYGNUkCQ1qZx
vN2Bg4JdmAXXwJdD+iMyLA5hM/UQWKyGh8SeCBi4abvII27bz1353qgmOq2nJ3YKETamnvq8uV22
DTvGrDoXuJhG5hX2qefLcguPQIvFhMEodzRFNjhR9uC/aLl3ZI1JIChvmi78N/yKAB2Squ75Loeo
n3SqVa+JuCywtUiahOoiU6kYeBK4lGQ4HAG75Vq3qcf6qSGTmnIhmeq63f70V1V5sMrrl5uU6IHt
2dR0W6zuNvcyQ1TWD+d+4g24PsgVZg+BnAoDE9LsPc5JdDJOTCCuuQSGwzDbA56qmKUzXtyRuOL5
QMGsQBhkNi90LUIaeBehy/fBhUE9A0GlUdmTU0fr9sRQesLro3XDxguHL0KwMI8sCEe0oVE31Q3T
AOY2ycGCJX+iNYOkNjkOJqnnA6H3M8QVeAkjguhuBJTTnaBKqpav1Zd8AhhWqDUMUsb0+bfpsIPU
PIpajeRLjCnGYBnHMsj08jjvZpg67Fhuk/aJ2+kQ9SO2rW7mavf8mMkkNaP+E4buwvIEopQfQ+xn
6moLlLCpy8m2gZSjUXDtCK9Cg1BwWL5r7yi0ML0KvSIlLJ0+fIcmTv0SrV8COqJdrnwIX8iolzJv
tmfmD8uPEB6JLaXl5e5ZHmAMMtRTmeMEV9LhkGjVDhNa+s58Qy+izqy8ntOMEuCbojDj/VolInXw
QWOOsSKRzild8KKjuEnaqbpWAH0GJqVqX03b2xDoSsrO3bILTHseZt9+EdKqvrm1u6X8KyxlkQpU
l4roSo7ubR7T6RMC1bt69CxL487agLiSI9b/+WI32p2hT5tczsQTH4UFbnQQsSU7bnrL4DFv88ky
tyAM+Izijw+okVazfRPu02ikJkwv4J3ZLiHA9faC2wTFa4LjalL/li2i8m3h5dTtsRpaB5e4TNn6
ly0X2rM+OlzLbTcRO8ibM9tmUGMJApORIoAsLReXb4GE7dhCQD/ZEhuByHbg3jTjLGOVKNLqKgyC
reVgFyuY3ZKkD827dSp4Xnez/dWP+SF5pT9eKkpCIwDC4mWVhnim8x97EoDTlvjD6dTroSqZXsEC
vBLt93fVWSLECjXOlmFp78Ff/J9aRrEllW+4U4sVhjuUxjIfhkKesQwxfU9bECUm070qQUPf+yie
AWW6dAjFDcL5xAgXPJ2+36BMx1lAtE5rveJ4LfY9lC8WboG1cD4YWP3qi1HmyAaaFTzFfEOXqH2o
tT0KAsHdJS1nMalT/r0Jn+NVNNMBifnJr8EUn/r7xhTihZo7KnbgquayD709ei3aeo+KML2Ta3ct
rNAP/nWKxm3eYfUmBVfBF9EEpxCOpOAplEXJIBhaGFu4W2lQFhGWojnk1Ac5GtKSj4TG5ONaCh1o
o2GwTH4xAgi62pAagsKXQjjfyymhb8xmZfoOVyHr7YDBQBZbawCZPl8Aq4lDgsW3JTdPFZGiJ5qU
xTH1qvspuEbjwlCF3fSHbG/0nTm7ldTwR1lHONr/y++SUMmdvXa09xYQWQHwHiQ6oxPik8edPdq/
7e707eeBZWkqE4IN99Reqynj0TFbEJ7QmOsjna2ng9IweWpTAYgIYdJBj9eO6jDRzBscnENrP65j
8OStu9vCy5HMAgqcAqA6jbi/QrsfXzRfeRBtwbqvAyu5hrsN00HIC+R3zfSefgekx7cV9pcoxzcL
u/E5NDate97qW07bgtbh3mbhmAYpobj+toWeuiSLDCejCOq+DwfHVmYmOqkir/lLEbIfUcu05+i/
id2SqM6DOYhQ9Ys6XOq6N5ED6r3luBXdX1/t+y04pnkK9fyjzvI/F5Co4auIoH/YevaVrcTqh7pc
wMlFDqCxHPKHD6tzehxdzKpb035UJwJH4avhJRE4nDY/lG2xxldibsymGUQyioBbj+L7LsfkSoSB
nKr3Q/m8BgEyRqcwLUku/FueWam7dcseKybgWULXqYFwx+A37bVI6ABsYodBxd2b+StTHXWTHdCS
zp3W+Gg7OQ0uv53/bC2d4UI2BMrhWv4b5oWuzFckN7G1vZQBs+6g7WExlQfhMpK3bxEAtW6biF9U
lEtW1tydT9ISpoQC3oQlddNOjUhok210Z+900KfSZE4xvIWNJ/khcFlNFXDOocpObx7/033jqFQd
3JaOLO0LnDISFrSk/phWyHXISJcyhH2RXg/i7TAkILwNDann6GbtrktA66juU8Nr+nW95cyw9R17
Vh9XiNEC0Wl7IPxhenCz7Mw40dLBwyivfGsqj7Hs+dBmqUA6yfFFLdzd7X/ltHkq/EvcC/d/j1kA
KC5xqhvzZXHWGYLFZ6bwTqUnuB8S2nnsGmC1Pok01DI7jNdgpBWQcfZq0OCybIeiKfkNr+7Cda5s
P2TyM6PMsmIoA9s5ZgZFeBjvaAfAn4ZsZTNn5lGe68iyJ+ZOiqzofygAXGY/i3tVadfgox04aQJK
cGpyfKEMC6n1CkppyeTIZtQovsTkty9blTHVfbBrh0F6Jjol+amjnkO9ZGVNuCtpX+5rOPw7qNlw
G4zqmagrDEW1Umwb+x1N+RQhAzCNZJMU0X5OLyZINld2wRzCji9TQfTzt+mcFSAh0bmlouHD102/
E3gNh+pDcoLEVoL5nivzsgBYzcA1gU9QeVMLZHiOhnK2FwGmIUMOMNbf2MzbTZPAyzzUtw/ciOtQ
D8wQnSG0ai6w90MFybploY1U/ig0j79mwZWNZ4ITAF67vAGN9FAqwHoTPkBMUEAF9ZjtifLPZ+k1
WBeLRw+xEKV6NFrnL0p+x6XtY5PrksVKDK3HHITEkG0wd7VZ4oCheucQzhQyYYj2P1X21hQz9htR
8d8m9nDPieGOOeznlSWMDsCXniyoZnrae4yKk3Qix0sLNgd9xXLBnrqMEv/LecHw25pwHBCuHa5O
8Kdum1IlwuElSn6Q4xmvpKxwBciPiVX88//xPu2MR12qiFOo9xikg73sN7b0yHbl+UeGWkjCh8P8
8R3le9+cY9fRXXu0zyKaJ0m332KA3rBYPdFyulyx6WGr05DAq2MPcFSY/YgilF+4U5Kg6m/Jpzrk
j5qyfNciMEJQjI7LsYm7bjj5A3WlPz3FC90DcNXFMhCcMGpturYI9y1D1FBlAH7170i68YfIsIf2
MfpIqQSk/22pyfblwqrKEC7Hv9UcNmTOC80Z0dOtPRjHqKYLwwKi36eEf+IPThP1j1T6T9uhgsqE
DPtDGdGEX7lTYtYo/GVxFrestPCuMhvgkaJFKWEgNuxHk268nYHxspmRimJeHFJptzZQ3+x8rO0u
MOmspuZFkOqhhFsqcEaS1WvqOu/SbyJQb93+Z2n3Z8XU58LI0UnaV1uwINaFCRCDUAmnAGhRKKx1
p98QzDg2bYOACCGFgM2LmDerkhKgAU3NEbcPqEXCsL0wHbBqofsDZVAyg33s0QSQe2zlqy5K1YVJ
W9JgH3rDqDmSyJqXfL98v6ge81Rwi+98ednN/pLH/wpRJnkaQTTENc5SkkzZhoY0efjwKBNqhg/5
e1PzgeGwz3PaC7Tu3ORyhow5Wwpt7gFn8IZcWw2yuJLLfBJXcKFpSyP7MXw99MiiDCQuA6RAzeBc
yNmBt1mbkVzHZxItzG+mOhzJ2/y4NYetZSu6anUqzE4RIcnYDpuCYtjAA5eyaX7Q1ylENSvFYBAe
faASFawvU2F6ywnzif04iBfcIM94GLtx1ZuvJ2AO3+GvAf4pUn12K4yIYvv4gTYbTnNaxLHswk0E
G8A9GuJHd+w/9Rm+NA9C9c9uohJmtRRHS2uZUsMAta+JNKMK7t4tw30ifazt4axYLd9gQxsjySEC
+n0o7CiapQzrt6+ieOpvT1B60C0+eUYeiHDXunwWw4s2r7nzIyBrEU6846JKhfe/uq6WAwysq5xu
SoHjPPW1UwXpUXB/G6wOythaFJ2MiDh5DAHtou9M0Gxj6ein4e/1DRq6tzMCxDdMU9wtO6nlEoGJ
AnBf8l7+sMmw1rK9WbeEds6BZTJn9HMfLHrDjjPwsnsqgjCELfcM2hhxMfsphTVnKf8CK6MPiOSv
M4cECv/EOCAZZogeDkpFv5bvuKiNfO6WrzxJudaTxVe+5TVSvBp1V2BSexmnFcFWR12iMRz42hpn
4sc5HWcrojDq/aJ0zU1HYMfBGFUWQ83w33i3F27Jz3zP5eBOf122giML5jPgjv4RSUPMjgsX6V0w
5zn24cYxqTklnYJimwNuc1bmod2v8n6sDruT27hAA68/Sac9DkaciGHZLSAHX1Gis7PfEJwo69Ob
kuQkNtAdZ53ZcN73duccTEa/bkz92eQAa3Un7k0Q79x6SjTUGT6fFdra25J6Ki+xKE41ZRAaCPHB
qez2ykcKxQTOwXQBeiBwQ4YDgZkrduPnq0qQv0cG4FUwvdzZw/AlwEkNKeVZlLhMy9/cp9p2Z5xo
DGKqOmw2BlhIXzcuDN31oyGPWddWs0/IBO/jO9jO7GnpSEzanZ36UXxuDYHo6lOvLYr99KFZDi+h
YibjSzyvxUZjdlkxB8PVVHsBlMSVbYeEeuCw/3rcV2LhDUQKrnFaDHxuivYbUxZwqzCGdIUNhEPl
cUanBcwBgmExl8uIgk1NUPxP592RkM/CDygBuYJYF5vZ1SS0OTQTM9kAnioQFh1CtzDylecNZiGG
sYUCSofm4c2kekBtwFisInDVpKsEO1jfA5GiKaTYxfBm4Bb4bmN2hCao3jDZRxoYHzcOE4jEr0EI
/zL1mWjs0BqAnbQ467YH75f9xO64+xFisCAqB4TDEHa9qyhRhlwIZfY38XBrloxWgWeNST2ritto
vQwF0jj11div6zVYcamxXLJNrqe4EuPkUii167bcGCMGeoZsNC6VzSwnZC+2/SUj3xZ9LxxtPzg3
UfcCAiSNmGcXCWa1M/kKbQ4Bj9n4YDRoOEivmMlfza6p2yIsJ4V+o7HcUu7voJRHYntA9H0ihlk7
2a4w5QTyMP2bQ1ET/lbNS31cIl6LXrAPlzEInccQBP8hMNbEGJnDk5gG/Kqo5Qwb1zwvpdy8Ahjp
SoiSITKcL8OvGDQ7z3ByJ9rz6ArP5lj8QOg+Qpo2hoDaMZ8D/oEZ3VXo1tarB0bEYiqo3vZr/lX0
DZdDaEgnl3oLaXbzlEOWERqIbEGwf/VMXDC12UCXENyBcZ6CTcpjmBuEYFSHlkBZyz8Poziby7NQ
yfCAg5DLJZOOANYvYFd1Nh2NCfjs7gPdabETI9uY2a6vuwvoZnrSVzb2W8BgL70gj3Hjdgs0dkHt
AccJhSR/nQ/Y6mkjwSAo4L1aORXQQNl0XYZ8/ohJU2s6VJS0cN3Vy+4sZRxqgCn3lxZLG8mqfk8d
gxCcdNEntfRLAL+bYoYNqH2xdxoGI1C4EiYHeU+PXqYmWdSbXGUdx7gwe0ggzXTrvh8kgUTEE2x0
04YKpLaMBeKTXkLX8J7dYuCEAkECtkvZcAU3GjPDMXJgJ1XPoKT5i7kXPc08z9tZXiFOnZdX6qGn
SdtKn/TMNJ8tckVQ+9MBSaW4jLVVxvVTM/Qt6fmUC+li6tccxJKpX4I6jKB9r/R/MG0rigCuNtaI
G0mvAPCWyAUfjpmtYXAaBXBbT4YRwiFPl+jOm5xKe11WXZvRl6royeCZZxisuA0yGqprMBzgGY8p
5DpPewirle8ZAe0p5KtzBRGL8SNwD1UI7i43Oe9I6/SUATRHsDyS1vS0bOQTv9Tr7oFKTu4pw4+e
UEqbKyhi6Q6QsXK1+ZbyyrHxYAxH9XDKUxKf04DuOxw0h2Np8AP1fxN8OleEsJf9UKnhOaL5lgQ9
AOyhL2GiH8ka5SaGMhP0hf+cgKxGpPMyk35MBt8/IflUifu7RugAHSemhxSCo8UN51HyNajr8fQi
r98mUbB3W4nUW/MndRW5cnmXW5iOiWvRA4tej+kaWNufaTfLalqPb7wyn+4Ypb+AESFr1b6KI70P
eCSBPsooRKV5Gu+j+y0heQFrhFaKqkOenYpYMHEVkL1J3ztfrTCzdGH7t8lMuUZhTp3K42oVJhaG
5wdVjxzmlyN3oOChh0axp4gnNnZ2ICeJk41ixAVYdCy/OYM0Z4w+4bX/mjZ3424ahAKN80IntqXS
7oTMrYAbxsK9HHVxYdWRctyeBeDk3BIAgm84NLhVVVhZBVn0dEuoCn030SGpx2C7v6grhAvds5HG
F4G13qJVMIhRyn3ZVyaiB4meiW0j3IUGb+icfaL9NvRWsEdURKxC522WTlPbfeL+fC2iDe1wub+2
3StbeF2JLBH9jUzrnKBDVin7YVbnX95+1c0SWv04EMaN2xjCvH9XxpZiDWUBKcF9UbIg6j/YTWJw
7vwINLiGWo2JSUcAFsD5fFmFiNNa2AWvEBZUxvWTQsekbXDtrwJwyvT3ZD32+Hge83cHiVjQdpmv
fhyFEeOFA3gCKPqh70fN0ECcKzMiQXI5+Olz8XBGHOOwQ1tfGzdVOujWvn6A1HuBHz3Tu8LGcZ1z
2W8j98wrAh7neWVNN/ihx50ble7Z1tPT89xm3qzYeh7Jel25IKJ2RGA7m1/oCO58eXT6+a7hL/TE
kfdxKxgkOOlv4MNlRSey3592hGxcqqYAf8c2U87zbFVp2Vl/8jnR+RqHMnCNbE3sZ71HV1XgGAst
FlPImaKOOkJqQbAGjLW58nE88/xGxWYAv+cwP7R+CKA62zJGfbqmu0QBZHU4akIQGVzEzwiRLdxq
67P8qP5vnstZpLq9wyYscFkP4n0TR3Xz5qqxBl1dV2/5WQgE6/DS8HaloeZ4ghQ66D++/IdiApwt
jbycQWO/mccWHcMF43iorlp/RRhlBr7kbKBcxGLAZPAcQP474LIMN+h44gtHiLxsarSu6av2Nsvj
WlUn5ESCmAhJtluTvkGZAR+IYmBsrhdX/TAhHmWTUbMHjFgKPkT/XQPaOovt4tukrxfr3CsVhE9V
viJfWEHPDHsS+zRMhAmVza04PSP0Xgda93tOWdvsy1oiwpXPmYN5dvVHuWAujktzKQVwHgulh+s1
6WWzrZe6YrySIk7owvV2VcMkOwyNhtLvMj8WCla9F0cGq13DaoaP6bT1cX/Sm6/aroOf2rNZ0xR0
6/tLQdLI3na7S0Psvau092QW5SsRfySIbi8tz0DMZm8+bmsXeul56jp820vItDoEIiDuzIGvEnDd
WXFXsxK4pSSRugqB1F3yiWW/eM7Issla/s8YolIxWsmcIA2S1e/lmAHYnIDjDmO+Kt+nUSOp5sEt
eYNbvPR68yJ2XsPidwXPYP/7z3IT987ZEAd6PoaZms3hQYsLcs0ZBbaqk+ISmwuqhE+5+lX/haH5
ilhSdVLLv/KqCQ2XCiXjYD6ZcdxaXULoewS0V332juPLIqlnn+h7XMijm4w+gEHBdD2ezkDoT5aY
5F0gs3CoIfRn0LwVf4b+Y64vzcg4dsb7elRP0dQzvW1Sc3l542cQrFM1p8jNnycKhf6O1xw7inO1
y8xU1P+r+EhDMQHloZrVhPNXjFDckbP6xKr7eIHMGo626ivPukXWRHJlNzcA0PY6VaZmI79EZpXj
R9kdX13C4ORXcAzJeFVosM4yEgeQ+qU0O4H5p1cy647OSeNbVpoiq92x0ocMwcU1DHFKHiTW2Rpb
D0qGfMcyOjr0BLtyd7Sc75plEB9mhlj4VKjKvLTC4xXt04mBRku+ZiJJnZ0FphmlFBrP8glsExrc
4FyxrBbDaD/CHblShjIJ8LBI8eZK7AnC6gJVE+15zuh1kweAfaLPaohrZp6PsOhkzCrAApa+eg5r
rE4X+qvnhsP+I0t8AixYutI38rPw1xB0VPzhgPPJHGOg6Ns4LGBr/aJkoEwHahrgchVnaPlt9nWt
ZpSGAUpSDaGOElv3rXW7DEOMQTEXoog1NwCDPI68ZrtgL81w9thQcN0tTLNLP5HWEIDxq62rZ2/u
dopcr31rz1j6FL3wMuARi7tuRR41M1rLwkpYud1R4s3uMwx8O0Vky5TlsdLeOYqYsXUEOT9ApdiF
gx0wLz1FeGECoE0p+qNFDCBUdUl19BRZ89KsuVRHZmotc8CeCZP3bTi4gxeLmBF0sInaCAupSzg/
Zj4S9J2U+ZLmE+HdB1vY/Ea6OHaqHpZKd4azxD/1OiZmU8GX5SobLZWqPtHRpH7oq2Gome3PYUn1
nzCJvjgHsFyYbmckHW/XlalHgC2yJznI+q92dZgxzb2Gz2gLtwhjuTuHKbACxv5bYlVWIPnkx6I+
rxuqIQ1uLAs6nN1DrsBKkXNUr+I1txYkqJ8M6VKyZwiRUR8LXqtsdwjWqcLB82PdEkD7IXxAWvtd
DSIZM7Ooalkub4dedSLCo2koUp1kCG/Rl/PSj/tn3RdfNcuV+YQ/8JwpddCLTBF+fxvVsmgftXjJ
J/cXAFuaSFfHzL4fvk99+uH8/JyNbq82IVdUW5nuVnwoKOwQtaeUrv109b0i4Y7aZoAaL+4D/JYH
B/2piVifE74X1TjMOLzUImFdiF9JoDuaeocG6N8Js/apWESYGLo3OyCXm48iLaYAskpO080jTiz9
nrIvaeQr1+dHdOnwqmrzw6biIIEgangCE3ls1u1rbwHxFC/ULZAwdUx/gX284Vy+g/fn8ZUrNZQE
akAhygWWVGqIW+mpFi2B6t9jUfQaXNbErPZWG+HvcdhN67jpRdxO8g7lsiCgm5d/zrHSL1gARCBz
F6laYzgSuP2lR1ZHj9lfBsIYmEZOSMwsuqD5CDq2Ce1Sx+rbr90jZcKDQuoCqjuH4erENFAaEIwS
UKlmkWj+xppGevvOOZ5K2Jec/sqYEHJ7aP/ROrS0nbATagi8nXA5wx4QS2IiQ7NK/MF0WCjdJ9zC
3/6Y4A5ruhqtjf5yWa/Xo7X92W75hZ5STUEidJ9vkGi14J4Jzc4gerIEiJhqdHOa+KO3xVh85c30
UJExloYUfdH2GT2ZWrlwJqlUtuh2D3qvZC2m6ssBuPc+zdR7e9pHm3eEg2re2sJV44xt7GfKIVuN
4pX/YEDKTugZbkAB+15PZGuwZZY47Kgz2CYEA3Iu/sfpiCHHznOns/FGFzbdCV3PTbq7Eso/TQa4
+Hp+Vnq5u9gig49PAMr/LJ5i2sppc1xsr3ZfjEIb81PWTKYhUqgHbatGwlxKRt7nKz0LIbpEzoiG
05FQsscOf7QCokMfOT7GkWegpwGSlWT1HjmPXEOr+CcCPj0pgaxOq7StYJk0gOynu3Zxw52NuZH6
BwuP13bAHF4P+Gp/zxRZHAi0oKAI37wGoxRfiNnjECrLT95q3NPIHP2EAyhT9dB9UlbgEzzRXxhC
zow9Ojn5kn2ygM3r2Z8DcsEcHkIffQTdoY8da5lfM9GCXPVWR00Mua8Ckv2ZurXew+mGtGPY5mVW
qoPM0u0QDGBDd8viSGF6D3jmgdfF1NTFyAC6Ny94FBLZHFqRUnLTke25wjyHog8mJU5SiA3Wkvhw
+zYp3BJKH1tr2tCY1gjhrli7HmB773yPYBJTsSHQBZYNyVvKO65WnTHUsVBHYZlwDIhqnRof3pwV
FPrKRc5csgCD+ZsF57w6KMN2VaKHubIF+cF+kr9yJD857ECbOQ6Hgt7mYH+Dyk8qxvr2IJAeqafh
rL4oBqedfiz3YQObEgjHSwZ8xWf40cnrAth0YQk9ZuEOjg/ZHNDPA4HCvbf4v/y0S68vqjk0NHxZ
swA/Zq2++xP9SPT5ek6A0QikqA9puqFzNs+v1vN3y9InelaetPphDzyLhcyXjAK+xJdCnBnd0tsv
a6F4gYPI12l8hmYAvIpbPAz0jaFi213sbp/WhnND4d5Ri1JImByLEW20Ox2XGQD9DdK+6/c+4kq8
RPiOTnY+F5e4h0KMXpcTcXvl4L7wSBqa+VZjeaeQBFBsXOkUzqv/KC7vva2TXIDmD3s5OvGPEJ5m
XZmcjTxrakl+cUu/cTYbBuITMUpfV3kS2XmHgJmOLnGNJLfRAq0ZYooAi8yE8mchyYalDr/VVBDF
yI1wjyQwK4x3dkTtgZ9+0om73CnSzjHbAq6Vo9Q6XSM87QICcmVV4/A0p1egp/BH359LTAlfqUht
xC4qG53cTK0hb1xRnjIaLeplhMDE9SPKad21bgjR4+SsqnbZlQmPb2qPSdQygksct3RYIomGXydw
NbfjknUtWulqtpol3oIvokpBhf46hf5KBZmmK8OPYAcoCha/K7tb/PDBK9/sc64DHyJnYcROnUtV
p1exn72xRjAQJoabxWbFSn21DLQI/17n5SehMQUPZIX3Xd+KWl8fR2H30J1P6WEL7sTislKV8gOu
tZvzWN6efbk+c8PtwVguByZ47GN4VNiopdQV+DXVtnF5KDFBNXGBvXlxE7R6dwnF++KKweF9KefV
okUk1d7V3opV8u6nxcQa5D4UNbOzP+Sxu5lSm8ZGmgH9DZMwg9aLpLVMkfrGuz0vNPdmd1mDIyhO
3nFEDBs+TUw2zbBTsDew1+pyaQq354ztD4cRqxMwLU2eKEDE2CsLcsOMmFOp915RFl3+JioAwQvz
fLVJ8h4AQhNL25lpBMkljfuBshLkp5jqhICp1yxfPCuc6JjtQ5yrFELSq1DkOoLUhOLvrqRV43Rh
oIwioR8V8lIVW6RHJaE2dp05ptpNH7S+BJVX5VJnbM6ljOHhUAN8Y6kGBaD63/4nB9nlGDXiHFap
mUytvojbIXnGuePJcdNMdgwAHM24Cw7W9FlG5q0a7ovM0COkrJxDNzW1NzVzHFN6/Dj+LC9wCTTR
BrzrL7eo87Qdfpjortqh40Wwm8TsOcrah65kY7F8zWVHzfMfsm/jB0M7qtoOn2dwBILxRfej1Zyc
vbGeDtbhvNT8nncs6PUHZa2iQCzc4M5z8c02Iqkx4k+4NPD6yAaBEYyBLs5QmBiA7dPp6Be3jDv/
6FZFfY3wmJgzrpNEiTpo6VKuDSAWyp/HpKxJSECfC5YgU2WtlkpIY1QNLesuPkfSd1pdr2TAqYRR
xL0pCClG7tN1xLIOXjv4iQrWldvbPM9Ymzjb8wTV05KY76m3FDDb4eEp5oPzjD6FfuhQ17F0xLOl
D+DbeB8/1Ys63r/zO2Djg9FgwdlrgYM/yAXIfRYP/XmTKXNao5fwFNJKcoe6XWDPl9SD+sARRi06
uBc6rrweF4ndNMdgaaczCTdAHK9+/TBHPjfLhJrAMidQVYywDjmnOJNX6Qx7ju7jN3lKHu85eDwZ
aAHy7heJjC8iPFasqpTA0FRYKusXx9QSQvo7DLAIe5FHJ0YwXsYF5zI9bfiupPrA+b4u9VSkyFhN
kLzQf6CfyBy0Ir0wyj76sizoBs27GPqdDQohojB1D05EneUzUX/XmUvTM2CjHnWiIcBUi+82AB5N
xNncfVUWsO/YlHdqosgLV9rlXTo2+G+tO/tu2odtcY/HeinSvr9EjKhjJoH5TE3z9t97gfKEhXBN
ci4xNLbKD2lOfMewq5QQxJXSNIFyniU7kbUSOkw4y4/pxK66xelroQBGVFPsWCsSWuEXiKV0DQah
2aeOo1ra2xD8T9f8HMJwqUrsXH7d6IeA6u7mU0IAWcRthrAhRjC4CaLoc58Z6hCcOPubFMqFIgpg
XN4ECv7jZ6BM8ZREeqXwTfr3XiAyfYYe9fk44wLRM8CPyn0AlIhiLbwc1Ly00KU7dTslE8tJgZgL
EiHLY6KPcE+5voWD/45sBGhgfbv8PrZVKJaxQn/8U+DKZQ8749tnx2mjWUEJgHXO66NREWFyglVu
3Q5hpcbl3tFpPPEPe6RE6/+NHo6HTR8qGOZif/OSFaVexTCLV9vVQDcheVP1PZP58xe64cDYHZSM
HkJUPTHwPl5FzTalNc+OkFSGi/jGClnAh3rYeAX1Gsr7IFxCDGI2jBs8W4GnRruCdIbk6jUAD+2p
4mThC8UGpu8Vwz/fT3/IxbA/g30pKKEpFzs0C2WWc9W1I5ubvhzbLot5XaHpPTZbyjmmopdfbIGk
VBMNXyR64uT812SsVnBGkV6AoeUJsxbxHmqBY7b5gnSwVLkpOF3dwjdbA8/WLYrhTrUbO3x7CrpJ
zCLDzUBmlvnechIHXZMfUo7raD2c36n6yM+B6dG46VZ8btFDzUPWminlAOLThqA8JkD+tIiGzG0O
eq6gW+Yugz0WoAtyHKBi54Cv6zYzhNf1axUZC8bMAFGSxz3n76/PrLOJ7id6Pnz6inUtMDn4pvxC
zlAu8fypNx02Re22134HHechgGJ6yX1pUPEWcXBVzlb4z44h146oC/2CIViRG0Y/fhZCPTu8rSf3
3zsDsRNy+cwnBREHl2myvMg0CqNJ9IKT4bTQ4k39mIvd/8cnVxYzF/9joATU0FGW6Q3ShQVvV/4o
b08pvFM3HrCLM5T3PK6BjMH8e4wXGEbMGjo8g1EghYnMZ5tF8Hc9KSNr2pU+CiqBSnLYE9rBR8At
5GGtVmAzyfsVujJuEPubCzTwmVMQ5rfVCGdjuqIitszyx6OmLp22VmzT+KpKsyFWrXXhnJ/coy2t
VzweGSKZxtp1xwXE0h5yyqaQzj7zU+QdHAJ+L0LWgRolQKGkqwYsnFE1Ka2rEs78IKSyODtVjiku
ufI9gOOBKyPP6fFmd2mN091WO9KTdSAC9oVdWF2NSo0wOCT4aGAMeZYtwOZaX3nO3Lw2j1VS8AgJ
QOj0lbNghvQJon8bBDSNiNw4pza20eW2Nqizv20g3dZPwJblmgrk+OVCy40loU7ILLfUW4YoQwWb
V4C9nGMUNQ9JsBpql2UR263DzayjVw2RMNiuJ1tQTVeYeSa225F9FHuAbCbdHhx4jXj/3kHDAxXx
2sGZJLp4LOKPn5T6tSTCRwx+OOmNR/Lupisu720ZCP1hmPpq/VRgjEr0vJpSEHlmEKC99tySm+s4
nviss5HC5cTtmKpBHU5ME2vVQKQhF1FTtzWBjsqZMXZ4X72K1e0g39OVDoaB1Rr0aAFIjWtOYgjo
sYrRA4NAh/GFRKFGNuJrpUrB8DIO117ZsPe1YAFNaJmrJXY0qmUwJ3RAJMZ0JEKuW53IZ08y4db2
EqPUhlANnwZxZqAevG+qeXLv4yWzAYdpAn4mocNI6NPRLgk0NksvkU1oAUJdLI+T/UIzdueDEdrb
I4zWnG5CqfNJ7SwAj1Fark8zHlnLbru5lmN2Si9LWoFBYu9TyTQgUyytCzAzyueTI86/uflCvmCc
BcKrYgPm2zT1oqM3fadzUS4T+7AbtIBWXllvfsCrc497t4ZIwa1TlPerhO+v0s5RKKLhY8S222Kg
G8Sjup6WXL9TJGA6/lK2n0gw13neKv/dkmUti3mRXSyNna70wazj13lpubtCqXmMMjPN/lIxEJbY
akTFVf/dtB6QFZslrBhJht7pjH/s5rlhPDjJdV2VwL7ER7STW90zR1bQDZzrIkoIHZgIyyFTf1Nw
LHg2TJ/FrQhfQUcjWbzeHDKws0DMCCA+s2LuEw5QU3P8iSR7miTnoBSngakrD8g6SdJYpUAD86Ig
K2Pm5IaNsPqls1ZQHWHUM0HGopTy9MlHlMGPH7vaKLHEYUwcfHBEDPjRfsjbk0uSF5I5hdZeo8IM
KFfGATUqEM/cPhFj/Uyz4e5Us4/ZoIR+LMBJLZcjrBnT7vfHd6SoZYyNnhLhAKjLEDN0Qf33qSrT
SKZEXtzBXTIKWOUoX4DGbxOcc5nAmmwlvxHdGdOVlqff+FaWCDrXbJMgAhk4AL+MGKv1dHR7/SMK
uIpU4+Obuf3nalrqgJW8Lr+7RH2vdE9xoaTu98bdrnL42gflLC2x0VV/md1ILBwPzmV3SRIpstRA
/1CdGgsr7txdPjd6JydNrlrG6f5S4NWluIrIwCxaO+9iSwOwvUqUaNdQ1XtSJYVawhlkl11gxUoC
qP6Zs633s7YZOdhtxVoaThjnQD17zvUrCe/gDAyz00vcWB9tvlyhhYV9P6XjJgLN5rVVzSODf6+O
ID7GEeIYkHwQor2YCyp6HkLkZzNDzB6rcoc78Ardns6KY//wXKRW/tLtpAbEJHHLQNZQAsJsv8Xe
Xpl6HHDHHCtTbTHLj5zv7azUOVN+RFN30N7daPwOOXb95xNtZ5999F7BbIewtREGatiTe5L83l/A
tmSkCaG5qw1rjHQk10qim9XnwMDwGDMLnHvC1hjnUUmwL2kiXADV5KDRfyjwbOGhz18Y7HrsmoPv
/yDur0s3/nTX8p8Z/mreY6UmVTf3KVwYmSSYFun/Fuxa2ppPu0ENjY7/IqGZPsvo5KIGpBxz3XeF
i/K5BLa8PzGKBkQOWSW8qvUU/ELYGMXJ/guTAO09WPChGNO5Pvo3nKVwL1Frbr+Yf/3yxVblP+PA
sLnI4BVVdRJABmCU/wXDo/vDMW1KT9f2WY9kLC7ZgKnhTT6jD43s1DJwyUmkLuhWGBHyWSjk4OfI
AE+yL9KtQ4zLhE/xL5QJdt6uDw/XGnJuPb7vuv8T1Y+MZ/h5E+GKz5Edfi64yf5KlvndW2gCHdN2
wI712wfpHdN7ISaQ/MUM3Wo/k5lWtGCPX2wkdDvjUnYdey2krAFlE+c2JCW/4/M6QA34xMu9kurY
63AYwGy18CDad9l9Fh6dVVwq3M3Hxgvq+Reo7ohIuIsMl6th+/btPRZeINsCQH3M4IIUH4uZNw1r
vgVPXMR3RdyplDMKN3vEsYn+1/jU9t2nnbRCYSR10VKQ6yZU9tGTUSPRwKLSbTcyRqK+duN8TngN
rFNzd5/vbRoiEyFf5enmmeE/+1UpURm/WUARNF3KnZhglJdX3NtZblwRqor41D9WOF/OntDCYWJT
GhG0cEtTIUwL8pfDBg74SUynxtGPgPPmrnu1NL5Zsc5S5t3FziG6SuXtcY9ZV/aaHqjyIjE9zpEf
hxskWB5AT+ySgqICCdRXt9E/oQAeGoNsa0xf898BrOAHBqxVu0XVaHgLp4TRTzggMEHuYqjMEfmZ
rDXPq8BvBZbvOKWk1C4EI1SzmztDaMG5lRAINNF1ME15Fr+SptSJO3N0Q8F2gV/xgH+1atOLc2RD
XmO6tiD7hBLxfssNnsP6Ce1Jm75zFK9x/26nlDLICqlTcKoypgQrAXdt3u2oGYn/UKalEWcZrAbE
62/joPCH7QH3HV7cD+KSQAcWJwF/KhnsbG8JMAJsDoQZq2GTnptzivZzVrXmlPMRwtbgwB0j4C16
HrV1QTm/4Zasat2LFDIlZEAK9N6iC3HNI0+9INPgWw28dIKh9AWg7BVEeIh1pTqya5NU0FZz66j6
YDgs6x+xrYTWwX1Ubotunh/669MqxfTkqaGpqpaJoBGu09Slnzw7WteOWzrSGPOYI516dwrfQYYX
dA0vswwkETlrtAfs9mDWOgcLPiGCJ+oFI6TsEgtx1bimojPkL2hvCImLrf967AWVsPXwMPzj+nr0
KQiXlC47eqQY6SqGzCvvfJBD5JhXWaOrndAK/52GAf8SzZRZktwxVUt6lu3xD/5aUUGXi9Uewysc
mF+ZiPAP65M18IGmBHECBJkZTIhYo2EAiEiP3yWN1DODYyH5xqeKL72KvdgrGiUwIhMrfkBKvBS/
k3dTPB7nkCRLOpmo1jP8WUWShulkf4GWhT3xS9nRWq4Sh3qzirQXqyU2FRXpYLmDQmoRGbklhk/v
tuQFuE/FvIODgDAZQBjLa/QBPf1FYd+4EUc9pw57D5Mt3Ksm2G9peFKHkf5EGrsS4tOJSJUXAtkj
Aa4OHMNeDzHxZ8dk3wj4X/9b6ZRxHWxBzwsfVrp4BOEElp2hzSUWuxTzSugKgeqY4bnJvqUwvFDS
ouJ5fsHH3fdTj0QOJ7y2U3Vj7fL2dAD6X+a2nrXbay7gXUgjGmkMMqOAzsAmYxMnvx1Sz0YxH4qo
zlEPud/BT8PMJlz8ivdAYE04kCaJrc5pVQvw/6lLxqmn4A44Wosfli6oGDJvOQApApmTQ1bUThyA
YDD8fq44zpKiQGsofv13OmEWINFhBXmh8NeD4xYuqMq8/M501imlvA4qTELSkZ8Kq7E6tN+lLWqF
5+A9y+MV9FbZG/wAm2qSKxUbaXMdmFsfbcrNHG9z2aeUbL/85Imr2pRGA3rnxLWgi8ElsAYU6Zja
c3P9/9wjXiLq6G7N488QmJinyBA/M60Le+wTQVAC/ZqXTb0D78tyh2Cy18c9OrdIhrFZY9rcK04P
vn0ppLcQUO1Lli129/V/e06IgQ1gNkSX7sE8gvj65KJD0G35WMbJHpmMFXrZN07kBY+w0qGY1b3J
vgQIdcSnU56Z3S+AqKRZvnE2dgOWRUMtaGA+3bJ61pUrsTVAX1mnggShACIiclsd4yX1wm6VI0Es
+GdSM46WFQsXGsRoR+QvZC4R7TGggyjCHWGmN+UzGXM00eACflg5eyMVD6+VojmFrkd8wKoNi6hc
kILBkaOy2cTiHQWgvGtQ853MDoSs4dYgxmAt1O0GHQrc3ydIdPvxGDuejGUwtFGobiSYnwjBq34s
i6z/ildKGhfDNstBN+rmYXSQOf/87n2wQ1HKRvtO19vGGxCbjxwV95VgKoOIsseWxD1wiMiLX7D+
Epun/cXJwbMTAjGDbPaRZPeDpeY7SRQqLUPGx0dfjVwi/gdhHc0djnwKsNXaJi649BbhY4HVcC4R
FlBx3qg5PnKip/Lh3nkL0xjbQoxGGzTN1tKa0cT42g8t2OT8GEVeuL8KWJ5hudx2duBabZmhMCF0
Zf0mklJpzXKIz8pE5Bas896YBqUvnf4cfpRXAa/Vo4d77W3qVa/MEBM+PbNbFKzuVr8t2p0DFSAd
uRHzcBgvEbW5nPuDyUxi7FBmFUhU5NeaQ1HOf+JY7U5r7pxR5IcUQ/6Hd5dO3qi0c8ueXukQIqYI
VhX/1bc57Gc9pJCJkSDTlQURrYhBHC5ZAXMENwFJChQNpoVyZwRdDxrZrk2RzbKfSdqz2aKTLn+H
Y2darD0f4qCE5YtyDgogJO4SRRCnR8LIsNYotQLZpEIaUSLVSzk7BomWdoDBDPHEj5yW/40zV17F
Pfr5uCRL8oAGj+bq+acffkQwY6DLgX1nGEm93qUzVlzhQtcXO0PMM1Fl8vsZ2wZkAx9gnDspsmgG
vl1aGnDTJlFkmfYhyMnZCxrUE78ScBflaqe1t+v384bn/lJ0sm46jJteFWfTwzplGa5wSXc0lBc5
S9lhY6WCtyBZNafWH+ztr6yMYOSxh7mLzmzFe+k2UbDtglvE+0Qg+4i3f2vh4zZVDxdo1ng1iIM4
Jb9OczmeFm1r5I5bSfdzGFBmfbIuak0elVaUvkhNEU+BDi45QEWkWJ32idz+fSIIw663+y9u+FPX
Eb3t4Cu0fEGv6zOymiy6UVPoLsEDj4LpjgvPcoaok69wihDWDdoALhNcitQ1TQqSeyOFecrR3KL6
+1MLyJqpFrIdiKVDEkhvR1TLItGuGcCi7HrGgEm1n1UxNJky9mty8AKmHY1h4CEAjxQ91veWbPlB
p2COdeoCJN6wwg0f7m1zhqKEfR/j+MkjA2Xx5qBlfnP8ZW5AqhRRCywDLSeYfvTfQ8yFRQ29iDwf
9RpcUUEOWEDyjuq4mH+4K42BVfirSieH5cVAN5M9Mczyeh4cDyUBWX5spl3gomC7WVc0/OAT/xQV
nN8Ur/DHzxmDMm3YY+Y1LEd56/eXeXZX5obb9Eyns99iih0bV4bdR98Crofju6gbTF9XFkXw7mEb
IvX6w+8FMXc+zQmMjpZJSSZzckkJCnuD8P8asC2or9k/D+0Hi5ZkWrfBJC0r0iXQV1tGLyD3an0q
SETplNxEc2W2N3bMtSlfSu9+xYvnqOCNzEmZda/WvzrNxzM4fekbP82w9eZ7XNLidlxxvQ/Pf/id
wHKayhXCYRBmgB3Q6EgMkxplXImBG2J2LG/hpRvZXTXKQjtmJqej5C5w4vuNwekmmjF80jECvA7W
ku3nIoLMT7a7zKp27+4AwbfUJd47zUa6Ki0i2wymuqPPeVLG+Ul+TlmoGsjXo0VBgKJhyiqNY2Qn
y0cTcq4wDmnmfQISAR/uWlhBri7HbpdoCInMFxe0M8OzdzKYPX0Phqg/RneCYlqF7LSSu1Y2nTNn
MZcZXSsm0HD36bdxNM1Ve+7MbumlqWxYPNh5DN0yYEt3aw7sTX17jChXMfGbqK3PHqjyeK1o0k5Y
4QAZnGidgwNjwxAxCXBbu06VvUIAO9W46wcjAVt54J+Sp294n+O6hT9u7jV/HLNX+lQZJ1IZVcWA
jOugHuDrvs9whsBitaIZDGTSEsb+shEBOIbBKwwveWHhzHqanc3xaMYWe+qt7YKbdkSLpvJC3ITM
T2s+1qoSnHIzNQJAiPEFs3IFajUUk9hLrooUwGVXmsnFmogUJNFBiA2IXzTZ41gdWR7Q7CielyQg
kPkWMpe00vQqr/oIk3r67qS75QgwCH1qefZ88vdlY6TEkV/LYXRdWH+Bk5Af2VsYff8izakMfKWc
BfSrQa+BZXc3kocdZqFWPfJamWD0+nLmlc8wxSs4/2g6L3YvarFakcwTBBWJwv166IFTixKhVcyk
r3mJW6UVGQMH+94E6QX9zdZ7zCDgq66YOUPru7FJxO2gXWc7SxBOt3KffQJzGxyiZxx9sKDVyGV6
en5lgGmZj4KdSb4Pq6nJNnIo3wQ3As/TqwiekcK9F7AP2GMR01PBzvETCvqia+p7zbHTdKFSyuZ2
RMsD7KH1pDlOdtM902Yc/0lMm+nXrTs7jcZlfM8bJR7Ad4JvQLa7yiHOGbWTvxWEhXemDGLgd1bJ
vRWKmMkxdvILef+la4JlOOZ8MEhE+tKOaqEqSn3uKCeGDiVAMjIfN6Mxl+sYP7thNWc7vqlF8+Cl
DHpfheFJKiFoSrpBNF34pO2Lcu1kwsr77vEOx8IVWSJAtyOWrWsYnsUAEABBzkoc9nfWMx/cDgY+
qKV9Ow8Nxljj+X7ficMEQqB7w4/Ro6fKhW3F3jjCDTzTo9UGqbqaEkfwoMjl0bs5xcnrvHMCI9KR
yJa3Qior5bfueoiPaE8TQ6EheiUU1gqo6E3mRgjmxvDtfU/h8089BS/oZCqOJVY41SnZezwM0li1
8muqhDZoVgNQ9Zg1lmNB2y6qRQstLisfgLJoFwm3yBonrFplvcH6asKjSTeT1Za8pmizFbpot5oj
jsH7ZYLyKpNYsnBZ+8nrPdFsc0mwRq7aWqxhmS3tRyeWstdLzEougVa3G5ucuhjoy85fH+ryscHJ
HIv0bnRUQtRWTHVY52CiEthw59kob8CknMs5soUyZe1JPNSvptOtkMc0L2m7IoEqiqZ5CydWs1uS
osUeRInEivOWy2PHL5a2q1UAhsEr+BWZZlUU1NDcMcEQq9BtAJSDNlx5moGnHtYxrxXgFVT/VQgd
7JO/jSt3tO7R19SneKAx3NnvewPcKVHTPSlL+U+vBN2T7tUm4bJlgkQMIpG4M5c9UA4LFR06UuKn
KO+imsBBjoTPifjAU6ip8qbGlXYl9GtbWNdQP7SShVDKyTTdtKzbP6H1iKCJOHB33mhEhVD9qnDB
DwD0do0UI7i4FWdoM0n6k2rynzXcWQmQjN4dSC0DgMz5R9iW3he3HwrkZW9AlxL7cydaRyWCiV7a
KZAXaHUuNWbUhTs43zhqG9vjjpoDX4XX08U9ZeLHpARpriyIE51fewPHvVDukQxD/MULT/6Ztz0r
986rgFoJrQAYIrh9NHFHdMPwRrIuiJ1uANQ1Gc3npReu9Pri/bg2yAAJto0nhXSimQm3TD3unbsT
ScnLmEmTClU2sm+PrbIsmhAkglsuqN7oSwoXHasEbEW0S4VXZCpqsGR21QESAhsyzwQyJssP/jr0
l//MN2bGDcE/pRi4ILSkL2bI4oamCBROrLRmzltERuBB0B95zp95ptB0/jSNjBCUjsrWsnWAwcr9
HYEtJstK+fSewmn1LsM5DktKKVixjw8ZSq5IBL8xJyilPJ+GPF4wp+Z1g6qit562SWXZViXpzwiV
njM1WoKZuMqdYOcZYwXeR9NtSIojJRlyIa84AriSK2Jo4zTSYp/n6b4uLD6Q/Ta4wr2yFIjjQz6N
ooi7XEeP/pCkCDmfJo7r6Js/s7uYrAlwVAlU9IyQ2PZ4gaSqy/ClQgDDThR0ZxSt92oBUJqYf7Ct
bMf3I3x6U/+IyF+ZrFQOVf3sYqqGJ7Coc2lAS4NAjb4dg/vArqSHzsEXQspabMaH8aYkeaHVVWpb
KcuD9tVQE5rMPAfP0KJaFCVWnwvtnq5Km3KfHu+fWXhf5nxZmmRp578Zcx0OSMs2Pj6bZFH7ndIY
ufpA0n0lbqXOBAWH2BuXfPfPJrI6nWBkRuP2HJe6stRdUe/gv6HVUui0Cg3HMaN13lcxv5pgQwye
zArgZeF+eMi+/IzZ2103nH0jKdDpDj/50jEqZO18icdAuKCSwGgsaAE8nHzufuaAYu0uGST/5qki
fuGgu1tXRY8aF3cPLiesxwoiI8I7T931e971Ac/0rbniue9O2PqbDlFKCb4txJYo2XXqUH7IC0ng
C1yPjobsAuj81nzvGRthh1ykBxYHcSSb55o6eZqzd/1dVZ501TjXcoXA7ambsDu2aO4ZxULETnjv
ZQarQz3EAReh2UP8/DJaMGQCEyVs7QtTbAbEULSg+1Uu3OskccCXKbCbZYUBVhlVURCBwyeF85dW
GTiTmkS0U/M5VmZ/qPfCaopyPVaxFLYhCEz/e4H3UNRQXo7ZThRQ+KRPPgyQv8JLGpyzCl1zn01F
OiptXhrfrUO4KgFgUanLbvm8pK06H2WBC22/8UQ5zdMctH/H9NWWTF2pXsHXmDjj1DK7rkx7MC66
VGXkdbOUj4na/s+G48qsOGoTbfDZvcNSc42MOmBlqaW0govMsLXE+NOcm4WdC2V0vi0McnZfA2ht
n3bPqr+xCFNXfufqiGSdn/4sT/lOHC1R/ljXkFHsYtJNqMecx1nVz5iodwW1zPIKfPc+7SRclflv
Ys3CkrUIpQO/Kox5RPBlCXQ1S4SLALCgSwKHIDZxxSnP+RvaHjxcvCbHS8mL8QcrQ4tOsJ2rrgcl
cIgYTOh57kjmPAjI98eqip/0XpmGTT6EA89g+DfecpDQ4gaCWOHCv6K/uSV+a6b8Et2AMdam7hps
mtZ8R9VYh1fmDdQ1cyOObN4/FidR2EPTyQw+dZRktE+zD0oo8lkfVUJrgRlEc+KexVrcXhN9Qa/0
7ePOqwuObmCTUPeRkU4rTXaENYgofmd8ltz2CvLKdI0vUdMUykYqxqr+PpyAr3uoMH5hRVmXOK0X
uEDqp8uf+2rib5AXITj4rpgFC+s1dBkQatAKliYg7dxc/vtMHelKL6uv8ifSaTrwc5A6fswcmFx4
arPLN/hg6r3OlK7srCVXydOpWi7w0gtaCGQK4RDnNb2KaYz2WnbUQ25MP2BJJc5tyFsYb3gDY+/4
jRsX1PVb+A22xyE+RGpAU0+BEWt7LT/eeDZyeXTMPl5kxSNJ6t/Dzcp22ycYBK1iFAyr4FjMoNAs
fNSWlEQ8lo+fOHSrwJL3fAs5oNGfpHNAelLXgwTr8Znys6GGZx+XGsn/w95vOCk4tuogXW/L2OQX
84j+5AIXL8lizYzVCfnK/6tnZHxxE2D0sbF0qzdRucicZ+0NsJpS3gajuV1dQOPeaEU88u/qECb5
/OHJ7W4d6ogE6JIosUcX0TTcKkrXgOAjRVN7bqK6aLtbly0KG3ZV7RNE61+EHNP27FGmZi4eZQ+D
UVV/K8e2r7n7PTM2ktzuWl1RIk6X9RklXvPgzOegYGY9QksGMaoP3IzvvBX6HUw40nFuXGRiJ9jB
BNa3zev1OcJzl4HpfoMo3ICS7haWVurhiftCgBi65vvLCmGFY6laq6QbOMl7Vw3KQsJeR/wXQyXL
+X1oYleKk9UDt7v//O9E1jY2SzDKWq4BdP1f8i53fe5eG+ie+75BKY0uFcnjQCAI90lGyW9dXdhj
M9KOzUxb8RFiSlehF7wuZbY8Rv6Xqzh0oqVfva/durG3kNWanfruMXN6efr4QdAd7SeKS8i69YF/
9/v8q62AF2H+yLBrF5Mh1aP3dnsai2O/EsxWMuiMJQv8rh1VURGtSd1V710KDT4p+kPDKULfAT/Z
dNEMZRKX1f8s4e2FjbgtGsyAuvax8fQr28EA435YXu8EMPdX05w2Tzs5MYXanafZhesun6E2wm/n
JhhR2TakvI2weC+9biFCz2qUoJTeghEoWfOENszcbP3Je1N+xPsUC+02amGyZYTaDaBpFdVVz+6Z
O7HOK2T1KQF6eupjWSDCuXUmoGLsCE5ci5RoBLbOYNT5lOQ55t/U7V9SUJdnWrWrR8Ae9+E+SU95
q06fxwjw4sQt81jhycpu2vWhYOxV4fUVtRknU3eL74sYOmDmEgALQntWIHxU+ZpABzQY1tJ4e5O3
Riq7ipftp8SAk1ZuiytThDslzTktibbDF4ZecL2rUjAk03sH9rUB1rIRkcOnhPWMNSTwxtmsszKz
BRx+sJroQHL5NtCtQw30CsWKnhSyC+/yhFtOMycOYqsgC2cx/RFApzPAdNOi9bALRycYIlg36W9i
OaA9PdKFmJYMu9qDZvyGwoNDPxIF5dXHVTcGkUnsf0WkisLAxsNLEE3PsPdmbpeZZi+XmN8SejNx
vlfZlyPhRmsRARmA+PZZJ7akbdWsTYHtzmw3Vs7hZqDi4548IOGZjD2AQQu2AB+AtCaswxEgjhEd
3+4ToU8U1ox0XT75s9p94ND1XVwiJo3ZfjXHB57kyYsBUjDmyDUp5tIXSv3Dyv+jrZ+bY+/+YFvh
wP6Afe2r73VjyXR3tYftp6nYEFgiwUT+NnE86LObYhUdsSqXv8uRH69b/G4RapHXT8u/Sv6D0I7M
405nJ2wFO9te0x8KJGAsqN8tBe3LDskaqP5Ay5vxQHV0htFVPeP0vy1KNHJroXWA4BsnyyA14KrS
ofYPvMSRRAbKCXte+gSEofhIOa+LZ7jIGYMv02WMtrAfYkKbqaKCKPYJ8LOS1begdYBaD9IsY0A2
5Q7UThb0DV5OKJGaDzlh7fTB+E8Wo4Kj4uV9nUY+tu9LoLMOsDQ1+Ix39+JuQ/IZbMNAvukWV1+2
vAmrKEhHL5zxrvIGV+i22XHEEdbC+sHdA4YbOLYDtGQQIvewix0r9Rxe2BXrF5jzE6WyJXkjMZya
V41iMXpEO5XYddNxaUSbnXniTvnfFR6su0A6BPwZ7I3V++DwNq3vTg5OX46cHTefQ6U/n/9sHxp0
jKIfD19VbffT001Umb9GVaMVk0nz/Aj4ad14kx02QxOoWPvlWJmhySiNCCM3zksdAJImu/RPqwbQ
H8SRi3m2Ekl/FQBTeRO9HlQ/GGQYVzPlYHoMTKkBSB7W2LqQdrTCDAi+Bp9XzaJAdAYogCWteoed
/x7sCRZuRN21g8ZgjOoKt1+yu7UTEHcAYqb1xFU1A2X1RcNY3w2L+AQ3bOwmhZh1mKjWIpTyHsHB
vAb5jW1HBG8AJXWcHGSgR0JdoWEzM3i27uI/gU+KGmu6KYqjghSmR6XuozxMiCz5B2h065NmWqj4
1okVJtqjUBvYIk+xDE0wJ1B3RgAwsCj0G7CTRCLPMWyhiFlQmvYZO/MdzOu7I+pwFv52vanNbVPD
BNWEZzPdJXLR0oXzLg0Vpd/y2CD/um5LA8i10EpMx7zZViUt+ySXQROQSAgbxqTLnmC2PrCTIFJK
u5xnoBRcXZmxZrmSKaoIHP84A+LJ4qVFdXfkXAOTlQrwf4PHrHFkX7si0jOyE72P2yOquQ0Alack
swPD0D+9CvUCYqruaxJVzYPNCjfjDAN7o2fWuYygEy+o4VFOCKSp9L6+mqJ3vIeKFddvtuuVZcjQ
3wgeZxZ8f1Pw45k5WEmgRzJER+KQ0MzDsG9dli5QalpBIXGfsR4nZO9CFb6ZRTXT32F/Pr7F3BDv
pd0RrmoN47exQHqDuy+usyTecE1BiZCcFquqNEsICWAbiarDZK8dRmvoIL4QxVcLW8e6LWEGOTZ+
g6xsskO1GuWXRzyHON4pNzrXeKup93jSbJqVnAnZB6uBMBfsX7PjnHfRNeG4j0eyyzssWPV6KszE
KokRab0SkD4qxn1DXeTgIbSYO/AbSFu3LAu1dVeFop+fU1msroPr4SVrCblzXHFKlSER+C9DZvJL
JTvOxtsuFWmQLtXY0mV/CHUuoiWLblrGB8FjluvmB+HKrMzWefg5CYRfLJurSvJ1T7/v+gINmltG
HsOn4yH/rgTsKu53k/DcSj7OLMKxQjWDLbM6MAHP/JqBvIPHxVNrScQYWOenFDgSGGe5xOIzc2gh
Sz397bp6Hf1uMd/KEAl1ouzyuRJ4+ui2BVHR6Ae5C+XM3qikkS7fdDFk3UfpsHyLFklp29wBKNWC
OomzrchjLFqCpdJGsSWG1CtrhHYg47fiYY8dApZ8p6ZeCjhe5e+0sgssKWxeSxH3UMkV+qWlO91W
cvuGe2+NzjHvc6+d1NRFqVDUdqnmL4W+uBLaBakDMc01Dp0IdOIO7tss0VZwRcA0tyg6x1Ft5Weo
7DHRsGlxCk9sreXsc0RgbZBan0hZLvoRmittbMJ/z7d4I71dNNnTCEkJwJIE/3QS3Jsib9zv4nOd
5a2QeTmPri22g08+IwsPMZDX7TGA2Uje+NVvycVvssnns7Av13qB9BiR/am7kKdvxjSJ89fJv4SH
eCpZWmnsZsXsY5EoiqTi1zv8HOK+PlZSQvEWJEg7+5keeqcy8kKzU+SnaOEGrWeaNbEo6n+RPFU7
Jw4pS+z5Fj7G16Q7biGjRObVnvOVu9HlPoAfIFTQ5VnhjkCN0WhdMDIarw0OVktEAhEXnHUpusS0
q4KnbaNffBHcLEBpfgkCWxCETL7C4amRL9xBk65arOH+DV3p2oDOYzLYS5VjyFoZS62V8GWfug6f
cP1iRABko204oCLjzaYRTojZerWbDposDDWRSM9n9NfPOxpQxnVal1i/fP9SLDkakxdsrxdO2xuu
0gdK6qXP1DDl/zlB/YbwhnVQzdPB7begkenV5NITRb4/WDyxqr0vz5s1jv6moUgZ7VnQR1UeLpJm
4srlr5aMLJbbbsOCzUI5ANVShvbEcjEvix2C74+RGrOxDkLHkIbRpaIQJVkUhnjrsVuf+rJMS+UX
OrYGb612PexdxbtYZQCrwccafRzuNyId/dJyP+ooEXgGSiIyMCtm30rWwOBwFDymwaSqFzkWhZw+
3SKzhnfdbrylUsoITro0HiXpWCVrMKIWHfs8IKSAuaRLGTX8O4diUyz1uUttrb5pf2pNDjL5bitM
fPcP2bCfwonH8nUiGB4wgjDUzcdxrevDXcSn6dlJbsMn4oleNckseE+jKNl+XdrX7BD5B41YTU7t
sEUzaGpD4+Os6yoJTjnhdlnih5o2Bil/bXBKxHqcXbkYo0q9yr98i1YgYcUyZhWvMaqQcHenqIAe
7Nes7Bt8TcWmHkg+5bo2tXAWA9kfvt6lkpsXOIT0bLgvQPbhihhSYFehm0/2MajX9pYvXZZpe0Sc
PdZN0rGxgQ0puITBQdk/kHLNH0rzNqEyUYl3p14eH15ukrFWHs8ileQYfEycPWgPcUvSYg6JepAI
mJG0cNqdAOde6f/vj5rxU+AUINY7z6XByQW31T7YJ4/ztBrZGXDWZrW/3fUejC5+YIYd5oly61VR
VLwMpK4TGhPHS8cu39yzGR4I++ZJPTBWWwz1J8qyMlTFr0mgDx4eaH1D+VeLdUxtQFOwDa0NU4Lg
Nd4UmetldbyvzQf+Gk1XRbYs6OQ1dQwYWXxa4KZoSGs7ZMBU9VaFUiGZhJmZ2hp5K/k7THNSFI4J
PG8WgzSKNMpi7N0C+mRvIGfNiLjQMk6mDwKgH5LajyUw/fpDq/s76tNpRzF/17LYfCBSzix9F3gM
eQSnOTu3HxVLd+cXOYPXgqbhzTI1ofmfLM0gOnOgAYbfrBcj5py5btwCNea2OEIxzEmjKjggfQk+
pKvBBwmSlIaI0IaiYgXvOOuPT55goO6Lalxb89HHhE/67TnC8QecKQh1BdpzImjmaNPmSwQRkZ0N
g0Vp8cVXNLOlyGdItCgI6v88hAD/dUvB55XBXenHUBae1d8hLCVzJCBalKGxsw1YzQM4aBYpuz1w
DuE4N4vdwAgF5dAZFD5LurFJlEfVT3neEiC4YIBD3HH1UhNZVePhnbH9es+D0qO6KQLz3qYe2XKf
1XCDXcUo026/aiLWFfyFbiyJtJh1UBl7VSINVscP5r6hFqwI1vb/NDMDmrdhYiZpcK67LUfXoriw
HXW4pMq2vWcTVztT7rAcXXGuOkNSEhohyeH3DkZkrOd/2lcLss4bqSxuvNNGmVORAq4ZbTtj3Ea2
Zg/2QFE0LD7socfGbOnnRUB1mmCesSVCq9xgS9R9+WlPYIxb5//buEYGyfWznKZWr+PGMwPpFxzA
pR/Cj7eu5EGvBc+o4x6gQ1kOi5CDSonN1apE+R8VLhmD/3sb/ZomhN3SXj7+Vg7wTCtGk49HGI8P
VrrjIGAzOlMSIFzFHenkWCSlQjfW+jyWxpNukcmTPPlJpvltfxtwd6l7mcVio74xGh2DWbfvkSuS
dPZhT+3IbwXDk/zoSalVXr/GyMfFB+RSsvwCkPAmB0iXd1d4cwpa19qm10Td3EdLAcSzKb0DcXDp
Ky/l513JJGyFUZTZQ0NIoIlr57jGrBPpaZCbNAry0J/hTDXXdryudFyKwsuFPUcry0a/HleT8RNQ
Au52xnlksUBfcoxpxWDrEWPBT1hY+gZXPtq0Jp4B/qC7fEVzSO3/92qxsJPcEsBUxqXtkOlmT0X0
kzr8pTnSjZ/oRdPFUURfV+6sYiP9z4fJypZeyivBe5li31zhgW/8sH0ilPDA6iuCcsLEmxSD3sqR
KGMI5hFLjje/Z4zQOCbJMLKOLt/SojCq0bNozow/mGAzqrYe42QQrNb+Yqv7m16/5qHKpsxFi6l4
VeQoVV7yZLVRgsODbDacxkAAblMJ7zX3AzCbB2b0bafLCu5xTF3DKxqOaK2rnxEL91VJOXMCGoYB
PwKTX2X4vRR23Mvn5Eg51CCoNXSNw8wnwm9iVqVKC3CZSCBT4Hju8r8+n25B87YpQyOQXFF0PgD0
7Q6y2Gzp8N3cRLerMWr/t3zCuzMH2EdHAxaEWMjkOUK2+3ZfKiytEbaOpJODoX+3IlNG/1TIqccx
81oRuK21o7O5RRxfbjLYbqz2KcjoqnDdTES4TVuGLVIqx7VgRi2CzlEZ+aSwN6DOWtmcoUBCC9Of
yvb/PZSeykb4z/QdgXe4c7vpZdqQ5qRPswrGW5Tuqu2ZZfvWhviEL7+YG2SieqyPMZ0pnZUQ1UaN
doflLaxQsaK1wsslHR2gdEifUa8XMzH9ttQp7MdaniMVxZh2qZhddIBAXjUHcTZQUZJsF6n6Kh2v
EPXz3E/to71zRQVO28n1rp2qhc7efqb1wmo3YhhKR+LXkxVzEgeB9Obq53SkKeoglQsSHWN5oOmg
9FlDLrcL+XHDpf+cs952XYhgFzWM1TK/ckHhIqAmhj+dpto1hn3/QcwCWr8pbwgRVoFsSXlgHIVt
pEcUFWX/tNUBDYphI9wP6Zh7v8S63rRBJbh7L8I9hi61736pLQrORP5kJ38+jn6hEGRsozJ6rLMD
XYB2npk3xO1B1GGoK1RF3di1JmYdUxlN/hc9WDD1OSu6S1ItpBmtsXWXK4b3BceJ+fjhUHSfni0o
ZNWFD1WgqjGrQ7MQcPId08W5wv0TCJYFbaBfOpOsLqkmbUHsLaLJOZjuebyLIumr1Pd3WuxbkV7v
AU8WakD4dJORBxnIrSeE6PC3HUXzMClNDorqMBOCPwobBUPMgqu3Z3r20Nf6LNFgeWspRUcbZdQs
WIkJBAJ6v6iBR0oGftelT2+s2PTUEkK2sc1CqKv+L2Q46s0VFEZA6D6Enf+mlaVcGB9wcICA5H6a
ZD9hEEISpMTrOy6HH96aSKvV3Xee5SVZrnAAoE5xrMIp8T544+ov9cABHrFsGDHFYYsE/1T/d21r
H1dW3hoc/hgOweWzvi/UHiFpQ/fureFPRbiMS42MchF+bSx43wRu4xfCHSntFUO2Hk9twy5IfbWE
K3TknWQgfU6te5kNvsptixktxh3Klzk9WA/8dq+uhIcxY6t0ky8CBYewD9Gfee58kmhDrv/kgk/P
YNe0daiyn1MT05lYPOw0ENQehxFXYuPwczvw/3kApwIfkmPWJjzQYfFmNDOfW0Ij9gB13ll/wbjl
/F/erRFPpLpn011GXUwL8lP4zDUQfWl/Y6OK93yF121vTVmi046WiwDG3xem4mlUqGEXkwgbYp/N
pYwCBE+n74N68LyoFz+Dy2azPm9Uk0ozffiqE2RQyAgVkIyxXAZoGaNOXzi54QnVox3W0c7iOK0l
ebMA5Zc/+aqXXEXAkg9dDjz5ALgJ8H3fC/OA1Csdv44puk+ZjdssuWB/IAjGShG9pk6IePT2+To1
G5NchOJxWsTmus5+dPukETdD8socqhWIv/lYx9L7k8cgbO5QcbNUSItRP6vh+lCXzOMFXU15JkSM
a0pj9r7HlzzyIprIzlvxY3+qIAkfTEQbzGWMov6FKjDdAeK9yUuBtbzWiTCFeLBCnf0kcJV4+fqh
TJH0IxZnOikdi4nMlj7WLoaU2RMvZoJwaRC9AcMKXcbqNOnVSf8zI2fGam88DuUDfVYKJ77XOKQq
sMbLMh7DPB2B5X0NEH6oErsnakxTzJjFoz+WodXtliVJXmrumfC8ZQHc18bHHDJpnLGuqKTA8BF2
fS0pQ98evhozbPnDiqWv4xC8LUvyxt5tYe0flP3nHC8KIoPR/2HOOQGI6XRAN4xERl6ie/ayYfPx
62t5g0LLjdkekiwcB24ygtCLxcPUZjgMBo8ygNhEVyL0481wUoPGcQoxcqxOpYgcndRsD3KevBBr
YNgOEESRt7d/pjo/qyCwJp0n105ybh1kn7u+qQwFUQR9l/U41ImAGBOEw2OTcbAYm9aOTiQ396zc
qDknCUNB3Ir6BK9iOtrMj7gQnAXiWKh76mEqs7x4o2A/+YAYb4Wzceo5oNgSSBfGmSeWMtMrY/+u
QVWDvteM1EaIgsHsuMpmmTeR2ZMmmc870bERoq5DhlFJ6U/8EEec+/Vn8K9mdZYO5IZqONbESrSa
VETF+gIMlQLUisjwJSxOekgiO1VrNdDu6SmgXXuYxxicbZ/Ol2d7dLD5f5ioyZ0sWmq/AAwO6DJv
5Ou4ogC5fPqjIjAkohxHTfcsMA9Itm/x+jK9o2HMXwVNNDhQjdJ6K3/EewOTYs/hoe8dKodUn2tt
nGsDUfNLKnn9X+fHnKRuZ2boHybZGBW/3RRScDnfoEAJIT26/6/7tSlZMVMEv+puMybmmyLNY/zO
ZbvC6CBHPqHJDjmRyYkJ/UZ3+tH2mN8nw68PSr2wV5PvYiEsMkd1hA/WvFmlyEVxQRiY4bmJur5m
hqMIOOMNedrjeVE1nLsHSxwaYSQS0U7g1qnH2+oHH5T0/scK1b+LedA6kJajYEay+MkZnTYYq8Qe
ZZ9WqV0XOKyB5QJtzFjg6DjDXznX8xCa5D1ZQ7e4PUUuR+6yMrF+JUPkq98GpYwx0XzFx2S1q7AP
w7ySUkdlbobTD0Oy78X6CwxYk14DtdyvqFklWh8EdbU68lfswf5PdujvaSQzBcorB3X+Eu1IoRHl
4jegQuSzQfRKNI4z0wpnVI1ujx7g1bnKPVp2Sgkp3/OBTc6Jya57x+HS9CSQwdbYdYytc7bP91wP
+tG00GESJB6Nf+j4cy8LLQ96pRJdCKM64QvBRCwrzzqFSdwqXQly2nNZaql7kZ9XP+GreZvtpgLN
U8hGiPpRi7R70+7canIZSDps0QcWTGwsHJHBzPjk19iieg/J8YzrJInSd0Ws9gZcmXBcxwxBWLwN
L9gucaB0k2VOcr9/RMVsuQRp4Q5+ToxyZmFKXx6SvskHUj+F57r8TcwgISZF7T4X9wgwjgXJyoyj
wMgvZUAaY6Q0lcJgYwWwrACzGOnX2vK2QOqou71juQQX5PettFvTJBOJmsyrzu2qV88Cw0Rb1sd2
li0QiA2HqLB3J123+8G1P7oJv8TBIx4pI63N14jGYtsb6rsnuYE5r0V99vwMP3eieV3mFH20Rhjx
ut5rbiHPIPhP66SJDi7sc8BV1xPxhBbPaJb3i1xpV/o9cBIQAj5gGj476kwLzNGqr/vxf0Yy+Ih3
P/KZiF74FhEOKYrrHfn8RRy5T16goEMzwoABBFKLZLg6kitm220y7eCxdcc/MMTKygP3jLZxPfoN
EamnmEnAcJGyDFwycUbL5cLYGNn3ekJ++WIjhUxr7HPpn0clvIzPtL/8pmuO4n42kTX9Nk/xOK6i
y2E8nbi0GIkyW+TvTsYqAKeI8hiwHKELjVEJqOGdLfy7DJe74H6Pb3cjyPM7gMJ27I0H1n00scjB
yPty6Y/2svz9HpNSZsbQRUhHwarDujVo9wxn9QQ/z+Z3QI1PWswLyqPMVIOxVrej9moxCz4ErR4Q
UiC11OI1PfjMZt4l7M5xWazPVJx6D/65kNMdPhPF4wlm4zcTeXibYv35F/VAdUbVQx/E7ue7IBTJ
t49FrD1AXNymAflZUX9MCzGLwiXK8ywexjuZLUtZ3pji8+CQe/oiTZOGQdhQW8hpxWpevRs22C93
iG7IjdvvsLzkvcAysl+v2cqAlb+BhG8RYWywjv/7F0bZsl+qdakIYXSx0Gt3G0Db6CfnGZkyyWoa
bEfnf6LS58TmYsi5ZeQ+wjgd3N6n6VZtGOM8u8Vp3BlTcFD2JunA42teyKgeDWtAqUCTEXjGWYAM
P0Frdov5y9fpmN8oYUQhjfKVGI0dkeDoG2JCwVvmG7EcgN1LgIPCjzluuZckS+1D48W3xYnTqHal
PThzgaMwbVTvgeXJkR/IhGz4ebv0ihEFQhjuguolb6Lsa9p+rBUzcDVUACk510YwFrgaJENMN+Lj
5ts6/6CSoU1Y6sdOpe+8HdsARavAfzWAQcltlj/W6VNK+eaB8Gxm9kuTwmExOmyVhiZD1Qth9XuV
FkQ0WjrwXrX2ARz9h94nKkn7YVdn5znfW1MWL5CYN0v6tXDX7EIf2G0erbrcqVoJhD6THbwmKcRP
Ww003/GepTaaHctDfMceGJySkgYb7/Pz3b+MHUny6OVIARRJpqDF+dv4NOOvNZZ6C6q8KclMrb4Y
UBNQ8jLCfk2f4RVAi2ufulQzQAP4DCi8tOYkDlk9ZNNj2sbzY8zZQoQKFXp0TDaoVUH2mb6otLIW
ATdH1vOhmMhhXKGmuE+eSNG3AlzAxDOE3Wv6jl4IiHi/ihdlTQlw/crA/CyyM3jgb3RLrXsvKFnf
mS2rYfl5X9vks6uNitNpcbVhCs70yfVIN2PFGYVoKVdljSSgIvZ573SwtR0CGI8XsXsqdLbcCz/W
y/NvnoW4cigelFVyVgIeUTSNlugrWNArOY7Dq+6UF3BtXd6V/0uooMEmk4j1d0bgA1llXtqvtQ4J
Bs+lHDDjmGZ4TI67QIId24ELw+O9QMb31a3mhQt/gO7TKOPRrCRSUeElyouNC/ru5+CY0xEZppfG
MAMqqJEc2dYNPTUxp+d1HQo81IvJqj8X35BRXqwajuo95k7Shov+Dq6XwzVnHNorqZqEcdEeRE1I
svQ3iPzpbW2Zn8SB24zzSh2e2iPxEYXAjaNWdATA5WFe1J+eeiKqrOFbHHHwuOPMspypSdXkctC9
42B3/5l/isUc4TrLz4th7EePj3+ld/bQY/5VClutZhksyWpb6HREwwOEZHhTjoTItuIMxr+j/q10
OZokYNDnpjLT394tUhz2PneALeCORup2BcV1ywMaIlkdUaPLK+b8gwLcmd3OuOr4z0GO4cBdsm5e
XtJm91oMcqwOfbjoZUfIXo1H3hIukOnv8YsHjV96Q/ll7uXkVZEfOUkuDsKNpMhQ9VQ4ugFZjDFA
nhGlf0psc37N2RUJJC/uuUrl9kp1N5v6GHGgTY6WV/yehbXAfIwok4cUe/ukvcpLBocJBJqlM44n
C4MckOVWcHodKsDyIRdzC7ZLwPcyuFaacBneDMIQvZOZnR21b/m/mTkUcm73yOkh1vbjWp+GERS6
idJIzcQU72+/MzMteIVVPch//yAQCHDXCsdb5ty1YSCdQxCSWpOCk3qE8J9JU8bKR4IDZF8u5fW6
lx0tvs5IFFzZTzVzhwaldFsp7GQsVz0p92Vb4lGdrUoPC3tevemFQ/nrwjq2WA893nDUz1UFVnPE
ioDAeGNjVnNG16Yyopkgi1QpPEKvMnEbo/Ev32hdTJm2shKomIy+L0AD1+MHOLy8fo1Yi3h+v5yH
gy/JO9grZbImFn4sFVG02uU/JNKeUlXp87gE875SRlGTwVSxOJ+oNi3zAQenIFQ2o0v2mGqvuzIH
Qe3Rr8PUAMRdT2N7xFzgoHbfjgtkLczMmlrHurKeGMZtlBIAz7FiDBcsx++O5ZR0UFiz8QjU9GVD
34wTF/YTZIhDMbMDVCRWKXmlLBPGas0sRlxmB3fYzQAOCqvI0CCGFR2N7L3MdT3QvElhmrE7rE+J
jMSv61FntHgEQLVtctA6N9xcmFXc1AiPaDpBIj6IsPrpKG+PauZXaHD+obrz+Q8+c9GNExSlYZPe
KZI72PSKNEIkr4nSwLN7x5ZE9nnaZhLELuI7siddTDto0VJcNDUeC2D3Or7/k7YYMrPVTTc84bH+
tc87THa4Jl+3e6TIUQyRfVKwigsKFYQCxcpn1roYVMJe1sd3ph4FsG7jD/JMoMFkj2P9zHauAdAL
17iTkcUbZfmwXTq/FXhS7y2N2wdZ8gNFyyjXp1L8DFTRjK7QHaIEhZF3ctuDKScRiPP4FSpWu0ov
zjP7KlzEesZwFcj3BcbSlzdpTBrBLnYAaSEfWey3A8M4qRd0v52xySjqwiNY7e3FuaKi7XTD3jz3
AH6s+wI4F5u+lhSMsX+fVUsIVxjRcHxEXcd9Uw/Y2GjG+KztZaDjOgdYrzd0FfIfKuFTF88t2iE7
qYJojDpZiEfaOtSqbmVLnZTTKR7Iu7QTHaioJmc8ZWoKLvuWCfMmKG0Q06R1MtCLBcUAMu4I6bbZ
qNnzNPTCkL9sGHLBjnrkL3uOLRxks0t/xEH09HrB5+WuhlCcM/CPtcvwJTPlNJAXXIVgwK6XrCAE
qvYOMR3a7LYmga0MTH0zS44pDEQ5fz8ZGBQSH4jYpFOz4IpqLsydslNRkvcjWu6Xq9Zo3SMAfneU
5AKLC3H3NXMCFx48nZg9xnlmgtsYpjl3EgXK0zzSUgScurH5+idCIrX2AEXuzQe42mr/0HjhaPSe
BYLQpYLWjOiSogv0lsktuQSdvP1nqWncOWHqtEQkrXjbzC3AMn1PLJ6PEFPkaEdNGV5paxMLlu/s
c7KAa3oQhWQ1m90H1MmcSAwUsmFloue6hDT9ejvleqSEeaUPuhqfMwaTYK158GcIwKeJXpSMCyfa
lb77Uf1oj8K5p0rEOkkQbXBKhCBMn+nGXEUnccVoz+jZnbubDU6CMzW6C0IB9GdvzbLGmqXK1I7y
YNIM+bxrQDciIHTd5cri0uqFsiu4vdFdJirdeeGnuXe/d66a+f6CHLbzdzBZ637wokafZcijCAxD
0XkudpkkB2+QWuXMYWdtqcSye8IX2GpBaCgdDwZhJ2zjQgZ0qE/mhSjS5N+GajHaHbSsYXUDSr8e
xhIq9qob5sj3pHkRq32WaL90ADWpJCpLsh2jNZGK1fJqTkuMfkUkPguVvVHSGS8QWeTKA+uE+Tl3
Dxv/nD38JR+vr170io2r2UAczCsbE5fwU9gDduIGLRH7g8S43I7FMtPC9yVbIiXwsmdNEd709PCm
kVU7Zh5/kev1kV25GUx0zEuqRVK1CryT3xycy7wbyzv+uyiiW4Was+JhZK6Imt3+1Qd4uQZuBvyQ
IO9uJR1tBPH9AGgMuoQoxEPDkdgRfsVFJR5X0hUxhXf2ksMtf4HwVFNvy2W+neniEke6OmLQtAfN
0gHVUgTaE0jdmvaJNDYF61eDSn40pFZLHcJljcSoOLFMMhzlwNnC2mp5szC+v2PhuQx80Ce5UC1q
jpYpuyyi7CNYyluL5gzGAciOyLs32QmlAofxVZnoKkGJFGk+l8CO04wrfUKT88i9m0oXiR2OF7qr
FbPUFIbTZTIq3Yx4DhRtoVqh2Yu4ffdUfSMjd68VPGu85L37leBjnsL22vdXXDsE3c2bku/TUsAI
tvYORJVp5V3IBEup6PMP9/K1smVYS11v9hR+YnguAf79LmYkCFLSYqifEFqz/xLbwbvoL74x2Apz
5Lu91cgKTgvQIf+3KlU2CGXIYHay3EXHqhEziVx1XarYvD81jOa4PGU/fygGy39bS1zD9jhmhq1S
UNNJ1Kikd66jVzIJnBPO5s3XHPu5Q+QjpjPMp0UpnZkGrnZ+kw/VRhG4LYsuBDb3wDHPn5+kxBXj
QS4qIssmKGF9Zvs2j/KNL350RWj0gIWLNlGtiRa+7Cr/ru6xd4g4Xghs+TAKFWW8MBW0+h3T9aQX
c/mKMZUBECqDfW1iX3UPKX0ZqXJljR5RXZPE3mCwBSvQTxR5hokPzPsmp8+B6tM3QYQ3rFe4jHHm
u689ZPISmB0Ol2bjswW/nGipnuNFt894bNjFmuDMRRhNyRfvukRhybfHOnycBEpdmSZIeRH7yrgJ
rd1I6mucwTTARI3ePIVchkQEYYMXOFuKuHDQFiidBgcMjPzAcrz2X/5EJKiWbcD5d/kAT/6PSc75
NvJPsGERRybetOnZC10DW8p5R3UUNuL6rjHA1WFMAru6JdxcS7nuq/DfPgtuKwd011DXcDiHL9nM
kLVKfKIfLIZPvWB1cnLnF7yewXBylwA4TFS6LNyYCl6iafFovczWQFbpMG8s1kQS0lOY2cDe+aOA
WjPMv+lX/OPpdVt9z/j5GCSv9Op9W7Ls1d6X5Rtsiz73/X/2pec6Q2mCxbKaptUMVrWB/XkgmDMj
Rxx8EABzjaW/w9pIkXYAb4aM/vRek/2FVsS7zP9hobTbzR01msTFpfE1wKvqZ/p9MTuQ9rvlUFjQ
4sOLWUFw3KbPpPcNzvskH+/PZtov+4WEhsuyImHWLQ7sBA0mvblxF/+hP/OXm3c4ggasDNuS7ebY
R+w1dPJVZ7wn0uC1cJqgaBrp/ErGK1t1zDQw1hEBPIhaI6l/sBukKLTQbuLYaPaSVOJRsQr8VLh4
x1uI+rzySC92u6f44YLF0bm9VhCSJjtH1bSXx79tMGfuLmWvMbIZVr+xMRgnm+nAAHBYluRj/0vg
Jw4jacv+5Iwu5RDcfim3dFI2aNX6N7ih4RsDPEBzkJ30j5jGGdkImtfo4+/OS14G9MKlWjqgFCre
xmbWZxm1VZ2JTUeNbNTO0KgRoj5IxDSiBFlzlgTou2Trh1tz+2sNhBygdz83HDdApUK0HFUBXhez
SshXHB/tlr1TzagVk6Yjs3DfCNmFuwFCNwTBMPM7ZpvkAjAJeo3rx8/lnBsWErM9FJ51JxZ9UFbd
tP5XUd4xOH2Lde9xA94onRhtedr1Jmm0tVI3uLGfmSdbMFnlyps47jXNCRsn5Gs9CDCL8mjI97jS
tJmASlHXDmY2hD3P6gUPJGPZHNzbuU4g3vt8eWifmVjdCwXV9F11gHOW7yjak2nX0JI3HSXP0mty
lziGunblu62mhpTEu8DGqGXD39fRSWKs6lXVzbn0ZbTpx82gbyaGDzb/51zrr6dhu+12vSBJRjRb
2j0wA60FCxb+Zr4LeOuryTIMme9f3xJv0mDW2112vCh+j+JbAt5/wZrhCpgMt1V70IVoUgaO0RS7
Rr5foafR3DORr/ZVe26SOziksEJffvXyn8ztUHaYy/sVcRj1w/TQtCXf4/yXJdAnt2IwLCb2H8GL
IKht6doWt8ZNK4NddD+Dd07cYXtdUBRsKJUW7em7NBmZPiZv5QAR+q8RbRF6VtBs+LGeH6w8to1+
9WoDWXi8a5uTMgfCvFyP9JdQFmDfNNnUplUTMWAqvGPfBTGWjlmn8D8KlKWm0NaJMIWJf1JH0q+E
Y0LRIOn/yNZoDyfs2tE+QgBfbW9S5gbIqYjNzR0Hb7k6lZbRRHjTEvdvcTELleqkJTglDyJpipgY
kljqGSPaEbDQyp/zdrkwzqcZfrZB6OxBlJsNGtAwsmR/4dgoIjUCtxXUYiAwoLFssZ4u3a+IDmXH
GtHb9uf7rP8dbfKGvWti/R+kEeaS+dw5ocCCvSrNFf8hSq1KvGvcICkGa2aboqNYTITg8E8Zzcv9
3lxYczAbc7I32Z/h9Gt451yMJOvxsVu3/r0UtetnGFRk4jL38b+g8FwtlK0NR+KHHZFsxc2Jk+2/
L2Roih6z7ziEWztahQCz9yF4/3w0eOsiOanbf5ADJlYS2A6RlMIl566P/b/uCNSdlVbMdCp4RHbb
0KkOY9qs+1OTDjUnwQtWJ9Q77bX3Rj8mlK/ADwUREHht61Iwc/heuK01yLMWuW+f8L7oGgykENvN
IifOLvrReFlhs4bBnoDYE66EweqRTr/f/d8o5+7cm++tHAPjuYpXcoG630gdJOWbid2dRLU1TDxo
o+lW+m1zCwNjX5PoPuUvKUtVKgC5jkvl85a8LI1oLRzHQFzsuErcSbS+5C503UmX97mGssTVkd/k
mkzbwM4msJ6cEXVHQeQPBt6x2oJTlFr6ylWHHEc0ecJOk+OR/CtjVjNSmVPHhTyachPH635sR7UJ
7x3mZVIpQL9gViJnBgkvMuAeJ+3lNN7s3KtKW49RL97ofJEkc4QnRHmG22DQq5NFgN/NF53taFqb
nvuC4R6I4B3NyzdH24dmmYPzEMjKtFR6XfPPl5dLAJTmPmWkJK9lD+fE3a3JjGTvQUmKQmf5UOnR
k4oJayR2gqr5u0CXqYWbwzGK/zTOTf7sC3UIBB0IIgEeNNDmrpihrGVVooNlnRssyR9iNz6PY5KN
US4TTcs+Nc84KAdWuM8OgDixnQZa/urll0SwjHLWKKCYBbme5yEnTrnrFvkc6K5GFt2yKYm8vslL
eQdcwjFAFor3BDm20X3WvYefVv0ZClou+EoMCE4/lToD7k01f5a9DxuRzuoTDPuNk+3XzAeVfv6g
jBN20ha09+0O3sqoR0y4F6LAShXjwuxzdjkPDvZRM7RqHh7YjBTSVtx2PdTldZspwZhkuYgEf3Nf
JUQKTYzvhHTn1hek2IiF4+BTEJtMdnUcddwNst9RNFuUYgnfICNcgLdDD0nC6W4KeUJ0g12IeZ8E
WUwhjXNuwQVbCTfSO58JeR8qQN/+yqS+9p2Rql8+sXSiqACWLEvmUhf3tfmo1ksoB4eHYDSCqhQc
7Oougs4oZwlNE8SU4D1Xs10Ls5/kW5UZ6dqrANJN2Ig7hDtRsmAHsDubFBlwaMBr/0d6uEW5Jxu6
5rFzRTOGeH01hVWkGyspRskAIMbKv7x1pCD8S9VRLXB5IWV7QxFQ87KfZhFCvpMQ676osGmjROff
fxBvLXZPkwwxcqCKx7k8bTzT37wQ1pdVncxS9MJ/IexC8QPt1scOHZhIjsRa+zYHQhLvhX7uZoQ+
1bNT6DmNwtzZFdkAifsdNfxTZY6ObV/6dvTRzArfCsRdz454tlQ+F6w/tTImMb0bLyh8NMRu09EK
fmU8oebQZsk0/yS32TEY4z491t3AhTlWndwvngv+ukDjf577e0BMNbp7lcUoLlYD4d67BZCx2l9r
MqPe/jc/RFVCFMXSztglMaI7npza51SCkVf4PwS18jL1KeRFmRQLWrhpbYZpqd0JQPSkQ+f001AM
TKPbsZObdWO6XlGEDpRsdVFqi2hVwLjFvxTHi9bPEq9X9cjYRWY2lTjlD0euyGxvgZ1Ct7SKhJ8D
dR8VfEUWzEYphZ6y2lRSsyKfzhuwH4GU/l9LZSyB6YSPfZiDP+MDgVTDCHnuqliKBJgc8Ase8ZNE
pz5ScwQwQiooaIG9PJJzX0wcVgkubE3YrK68wOwRI65IZ4xCcYE+6noR7zqyIlzPgpRqEfsiAY5N
incwuXCGw0naFRxhjMVNzgJn4yRk+g8W42Q53xkrkKFKid8wRayNjo6adwOnZ7totyjKidQirsST
VZFDM+sW2k3MKfAoUdV/c5Gu/a9/YWU7sgcS+83yeeoSXT+cwyx132jOOtf1zClbLfohr5TICz+N
CuBi5Gx3zRrJXHVG1UO12swvNUvVDGAh2jVQtBmR8AL2MGRXhRuswZwXLh1SlY05ARdS6gxAXRGL
NvhLeaUAuXGHppViSG1WJgVij3jtVRqvWwOYPsMAUHo7EtVCn2sb1EdDngcEn4P+ZmHTBBd+dBlD
cLzOXf61Y3YAOpldXdvZQxzZEK3N9ZHi1bq1kgFSbRUKlRUM1KV8+44Px/T/X7zWW2p71YQ33X9w
urULxfZgunyE2I77kMwnU/75FEKAsEhxzpuZkBuVmj8/LOimgraeistULbft9UOlTo6+mBAcMq7r
72z7BFaZu4FkQ1W5YZh9beUtNabCQ5P/JXCQzRD6mM4+9BIByQTn66jniqTLBdM9BIrASuhrN/iy
eZUaIj4eQZhtDGJkKlfssmRGraRDw1UD2VxeNqct+xXyWMg4HOb9kT1f32soZRjGjkXIX3Nbpl6E
LsY17Cbp6OXRYxfESw1UH0a5vL2+z6LoDKY2W8nR6susuovmHiJBUXbMxNsTvloEGlUsbXgbiEbd
+HIL/20Mha828u0vIgLBbk7s++tSJ/2KEdhclhXKWICVZsTfSKCIXuYTQIdLTGuf59q9dAzXK1us
k95AA/vrJitUHufRCZdMoSi3gsntZAHuB8C1syR09l2LkOw2JqvWOYivLNYQ0Ylxm5D0MSlcr7VR
dHDbk3T/uyM8SfMA9D+2yDxkLvcle5MJiG6JL7GV7R9tPSuutqSL4YAIfdR5tfnHR/Uz6lkGEQ4T
WT+crk2Ar9JiW9XVHhgP9G3HEHdg2jotblnWsDcUhRPNFSoqlAE7mqhesRVbMUOnz6iNHWMutnGr
9+0wp9FQmmcd4UsiDCF30pmWHspUedCce5dB0QjxF7Dm+8xE1lEV0Wht9gIyyMLM1+7vf8B0ErEq
A4Xl4fyCs6dwLCwOiW+mF44pfsgTiS2Qf8HKB9lyFqMMUwhWjp/wgoEdAc/7I0RumPBuqgEzB2lz
LYksLPdGcM+LDz4T4VRHLJUmC1b6ViHvY78iOItMtTe+ND7t593P4JfznfJVsehd92OqHFMj9dzm
ptbIeWPw0olYCh2wCnaFfzvzlrLeVTR7G95KqBiea8cwRlOkrvJEZD2vmbX1k+PvwAtKYgGytSSJ
QWkF36rh95zveWukK+CDV0TmxfLImA6i7KT8HWMHoA3RfD05qMEm2RIOeHc66sFF4EdpnjJeQYEd
q4FUB7EapQyPPoFSdpQb+VSYBLkoBJnELMWRqeaptus7pjlBll/oXANBrBnsXIkh1K0rT5KzJI11
UO9+xKaC/K87QgIqpjzn2my5LQCypaP8uCEz/3BXfQnoAwrrL0/LP81tR09GwsrxCt5I0V5TnxRl
PpB83yxTtaO2AKCiPz07dYLPrTi9wRAHvinUU9wk+ju/z6O17rD4lmtgNaWV9/aXCfMNQpatGche
OFN7D6g82x1znLIelcbTlG0kqBrZ2hrHRzMSGfIeoVdL45BSWB0jY/5/g+/t3RogczkFzSYczleu
CCOdU5t1a2yOVyHcXBWUQ2rPTmEMmJMq9A4j0eDj6vs/AVQ2i3u59xEm22nEufOPTZZMoKimNwF+
/JGEQnhiLo3yTKI9F/8thr1WukYgQOOF1Xih/Zu6SP0esOCW1XWDhvjF+0I4CgVE7JZ+SGXjoRi6
ijMu/nXBQn9ge+7CGi8VZ/WZ36zVUUBOdBRpyqFkJgKZHcLWR0ddi74Z74gFEkaQ1lFI9sRIzHVC
UN1noO9h2sgPfqylErvBTWG8Fnl80X3WhVVSNo4eIsmst0jPiWg4lW4CQsJEoLTpksWEwaFi3bHH
Xr4kFLMcYWndFK74jF7mZQxlwDZZCQ/gKo0tTiSQ+FwXjwcpdYW5GejkcGhGX0qSXWNmDrQ7enZl
xKR0FqWhOhG5YQeMNyasC4ZC98X2atcag4hl8wKeLUbYiHS/lVYeOXSIApupW2Mzk/fKudt3+Ivb
Wfqh62klpIzcSAnDqz99iwiH6uJUpfZ+jjjy9Tvzb736V2vrFfFySGOepfgjJG+COtnt+RDMyuo9
wN36+fN/oB+O739ZcO/iTjZas49rxNnhSlTCaAZV+yKjkVBLSpcJccY0smZZ7lXwjwMgrMizxThj
lAIk3ZqkBQm+xvttU9akXvfFaVPGQtajtU4ztql16FKrBcqtXTk2NEvXBdSza2UKx12E1IQBV2pA
VbW23NKvaDyEQqgFeprEIV7A6p59wS4TAGkGehyWHachqcm1j8OUwW1FK+XjXTRCmAzMcsMqrgDZ
qUcckqcr2+ORJc/j1dlsGA+95FCrG5XLeFF9xRJdOn42ceWx16VAU6snH+5sp7XWhbfq47L33fa1
M9clfaCK90LfstNyLnz5iZWCpatP9YHpEjbUXPUsDJJfxfW4/r7+sVmYfAkvEGj9BfyP5cg4z/MR
BKTYYQCnfLpGIZ00q4EkJ51sYfq+pBx2/GX2w1OU5RWgjup8Y4fcpxghmC9bhe/InNDhKOyRTvuh
PJ+jkbnBC4gtRkF8uy+nbqLyEO4Lv6+siDoesC7UD5Lgwc6xspAzpniLUjYgVCUUoSed2+KJ/xZ+
vEE0bLdI1+qvbPcxVa3ohkMDvKvcFVR7nQL4Cl4WmZyhIW2xLuNsnqwrf1yx9Wo5m8XXMW1vms69
0v6TD7zG2riiz3wATuFYHJiXV6bjNUKVtmHuCPbbr/LXqtk0IInKzahSLzGzS+aCTGWXpjvxU1+L
jLVNzo4ieNCRCfS13EBjqqN117YmTQblmI4vN66Jg4n1U75gItH3/nKNH2PxZ6ja4dNh+y/SBTDX
becY29iwCRT90SREGJJURT/hZqGQKPIxCc+b2XBx6RE+NkEbVQS/H+ASMtNs7hWtqB9Uvo73BAlU
Tj3NMVwfQM7S+8GmqR9ZSKRSpeHfl3LfuTS5rxXRL4vYJA6aDbdHIC6jkhauAro+viA9OCFtbqZv
cWw5mckfQLswTOIY3Os5ikz0yftJcrJnJIheDB4g5Nf2OQ3OsAR4i4XuYoqvyEU6D4CjbYL7aD/u
GrbkfEUd7m9yHA95V0vKQYZ3wpgA9iPU0Ej2CHhm9sCowD1l/q588zRc5O4AWX1fiH9Qf6LWAu6j
qQxOh/S1tBLh6tAP+0vdwZP8zWaAp5nJIX5lQ/QU1fZK9UwDg6MllcXTnbbsnNmpUrdcxCs87x3z
AAZTaHMHuti5WII+g0irxsqWjbrp+X4t6uqS+V+XirYWphRSg6VvS+HpEGsQ4cSOJpaH5uEexdHs
70q78RxhJkrA/UkGZJLeJYxQd+47kyXphP14mhVHI1/vZsVkSROGmD90njU+dwasGE8enXm1z7Xq
wRhsEyluJYwUHn02sQYcFYtaOWX5Sxc010lLo7QG+iqnxh0gTvs7HIy7VAuEc1RnVDGyc4Tgrxg6
3fQQPIEVO5klAwHlV5pOac5X1UDIcSU2rb9RVn/uO5qg7xGAHI5XOsgogRsOlp6sQLxe9m5alyIa
SJnl5KLKk/07Ur2yto7KKfCPesGRA/FPb+lbtnbPH+E/ID9iLUGeugUotmA226lE7JKKlWB6f8sO
qCP6iRF5aeqj3cjfaGiGMqlhUlPaBrtl46LfWKDvqBciIRlqW6XIp/r0TZ6F6k/mWrETMhdllGia
f11CqdzSKE2yN/2At2yyLNt+f7fsOGMVPvoxXIL/s7kYbTnOeLHBcd5y8XqbNaq10w4Xu1H3KMsx
9dfiQF31bzqD5ju3GwmVb5MH57l1M0xYoYLMg05LQdJWiP6TXZvL5N8no6cZQrUoQiTUc77Z36mO
45bAO7BiVW7NtCyLr0ZKdlmN8Ykax/SzewALPEeGt+acwZn4fC9VtQpnqDfDeRASguN7hzYb5Z1o
uZxcqKQv5IoVex31Wtw/Cm5tTBclp30F3v8EyP64i/a6X0WjrbGy10OFTyeZ7lzz/1NayVHUcxo9
BBXtlHU8gFjA39g9eGvp+v1aql/EdNZkhWgTYk8FUgfII/qnT5veuDRs9Sg8ET0JRREkk5lw9qCh
CzyISUlrpzApEjr9XJTFJhmdffNFQ0Qr8HT9cfI895PTPE8Vagk7kphFS61LDwC7aWsD3FB0bkUK
/GXCH6/0a27LvuNZOu4YAUSjCqc25MG5aWq1Vz4ap59hg6hPD5WdEBq18lhU3ZE0r0z2nxPTLYv4
OoXLBJSrFOhHFbjlVcidpv3k3NG2XtBG1cEJKGGLQGznuglOQL8oK28XfY6DkLGInJ2SkeGzs9HV
eP49mn/zVbNrmrEFyN+aLSq7C3kv+sBUwxchAZkZcpJiMElvCjhODCga2DyKLtyn+chyCRmLESoU
yqUj8H8FDH5i1V3Mm8PqBPk9Can6bGVvYQHzyG8+38fS9TjfV5uRnriFL6CRm66MpaJBE6rAhWFI
fOLe/+PK/tIV8jA9pOe4OThHp9/Skw4KYTpuIdBhC0rdVEKi2Qm/6V9ARCYjDeuLgDMEbE41EbVs
n1v7RcSs1WVmROwu7BqNhbW0g3PxLCAjpuwlVtKUsTzISB4xlrbU8mbChOJ0JV/VnlnTgNl6CdoS
T64bi//sfYn0hjsWt4eVVwtWNDMekNe4a6Ijfwg3fS75MxvS/GXC70ZEbrQdcjSKVdqRSd64Jm7c
P8QFW8IZ+cfPxTzkwb3S+t20PBI42DbpTl9BIDJB+bygVOZJJtsjkQfJXOOhbjAJDhn1n1xH3/ba
jaJ2JNhgCjsCc6kDLaEd6/sz9XaExthly1fJ1tM+d0rVn5We5CYBfF0n+MD6cQ7aa6XXklCWncCW
Tl6UMgQYWkfomsucPL1BrtawukhJ4JSa5Z4g+UnomNVrsdnu2FX39P11EZ3dgE4GhuZdbzPFPRVT
28HcyWCIHksPd9XaMuPl+gT/XZI/LOBcUHg9dPt7KXVfHb5XGjqT5yrrSJAAdYCCJf6wYmpjWBnk
JEUxre3fF/+MrAiAOqu7Fq8yYxxknB9/G8Nmx1YwShkcPyNEhFFyEE5iE7zrDq92ZO/lC6dOMhA2
7jAyI5sa9yBaXLQzY8pBzPgSpJp+QRWNqHIOLR9oHjYK5ucIeZOxE2YySJ3+l+37w7IK3pfEg3xY
eTLlNsyUXufFSwJPBp3aPZr74ut7GF006tAIGJa7gzt98WESMJhFjpDjZNhmUeFs1hKgtCxrOEBc
r5vJa6NJCoJC2GS0t9fygWpOCwgjQJnFO/hF1oZF/i1aGpZ05LWgjZB1tNeshz6bSI5UTklkkMr6
lyAcWSh8Q7IgE0KTgUYpIrvu04g71M4aB7SsevbLFVOh6dQVOtQb/sa8OArbBWUzbKWPQMaTzwIL
TyzHcLqRxHjKel3rsmKuNClJ6RfL5vzOFpM32Vv7DWS609k/tV6fjgmsO7ZkKEHcmA9s8Tx7iAMD
/wXM6E6rVxx9HLI9DfVpWbhERWS1tPdT5E/Q5rQ4oeRuDBAvR3Xdrd85Qf9wTrzYGvH0jBSHA/we
5CqXHx1G7sxIU09asqDxfpbQ/YxJwJtkmdKNKiTbeyV1fN4PL3kHFC4H4DosujQmueXLvGMtT0q9
uaf4sF1C9AyqixrCdeodcjRHHJiYeosfQ8QTNTMIBNY4NJiHF4TqdfScDQnEGY0aemfpG4FvHTbb
QW2bSkFejI6zDNHqI05adyAr7O9ki83Cpx6GDaaLmtDRVYgc2gCt1zVJ+sI/XnNkg8iEietsBMaQ
fIBT4HtI8ZEGkE5czrFX3/0e8LOV6eTBjlQC02hzfAlcDK0navNG76E97NGDM/Q+zbARdbMQwUvY
fm8kUqsjftb2SNg6nNCeSJHlmJUNofGsFhaAqVs8eeMWhq+HhI5rw86Box5iFeQjpvo99cei1eZu
a7FQK9CQJODwghROGTiu3OFFN3KvAjkLAHwekBR1bpiVQBx/NrOIBKacU0c+IjWFbhtTKDms8MaR
2e2OVfYgnvpLIZ4xXx+4Lj46bkDU4RLS1cPblOhVBw3SNNUOPoi5xP9r2YBbJ7/mLLf9SV6KNeaE
H05MRAslN3ZOL7cm/njbl3dHfiXwEeDr4zhz0ETPLUURT9TlablRkyvSAyZkkKSsMMa7ovwRXnBp
PyGBwJJJzJPwbqnwRdx1Y766vPGJXB7F8fC+O4XpVDC2Yh+eGoZEaX/LH02A+ohmHrUvpP3LuGXd
XQPHJQ1gG8UNzTGPG5RoHMGe9h3B7THFGO+zgvFrN1HDSriYzmuR3auZTfNDBwdj6i5ZVmIz3+yu
FNoausbUYZtx3Cd/yU6V27P5M7IoHxBYbd5jAafFFeCaySJT/WZGM7BImyZPEBSJEBJFpkTEz/kH
aIlQBFk6F5hZTxbUJ8jTMpbGqWDioaYcYhsmKoZvPA9OcjmOrdBm0hYoICkezcKwOTzAihFMKDi8
OETCtzI1Yy9DpWF9jylwGiq/johOHY/mw64wLCF8fajlJVJc+Re9qcOcyzL9Z7vgrA2KXn9lJoLy
m/hjVJucfLTHv1W055EGfoVJ5HHC11EgU06ykeNaQzIFf6eUUX2m8uGw2ak/8o1bmyct425vpxk/
bmF6j4A60tVvk70dISf0yfKlKM+UpLR7pFRtGMxRqKRQ9oOdRjsD54aDy6wlDvVowj2J634aYg9Y
RGqj5t04B80iqf7TWp5qugkurDYi2bqZ0EzvzRfm9Lg+9KscAuqhiHinnoEymGGE/y/z35oYSPsY
5WNzzeiRmzohE06nbajaovenmuHDueU4Yg73iMEMS7scPWXGEfa9f3O+3MBf7rpmUv061hXzCZbA
08qHvSFiul3B6avAd8VtxHRE3zoKEPiDCUaSEYBMTTha7t21lhnr/gxS9oWv9T7kxM0YIJaBXEXu
0KoVSeC14cppleydNbJHKLt9J8NHtAmPu8B/6l2PuCUj8Q+pByA2RZXEMiBQ7dQIGGwftZ+Q++9e
XpVK+VKcxqIzglPfc/MtRTA08hBZ6b50LdQTY2YMudoTgpq7uZgehl0+bjzTlNfoaZ9LEwlb2IKk
tq5gjWOMtV7V7PNH2njEwPNeipoCPkkNLyzVyruUQVZEDuJAaPaz4PoETrnYw0zuu+SC+ENvhog3
6I3eSci4l9vYst0v+Ytl2cdZOY9VaVh1gRsT8HiSmErrWCys9pu5ruasILjbUQE/Upq4Vgdyb2Fz
akEVu3QPE5/7+sL38Wus4cjrJLzj1kS5kaHJD63sdpoQuD+uJmxSqm0nu8ddfMmsG2KUPTZm5GOQ
wsS4m29Rf1WCSHuwLWiXOurUoLG9I+/5UxdHF3yiTPW8Ugn+nogeP7cxxKerhBPYUgrR1BXGE43p
e2DrtnwVc6Rn1d2uKEP01xMQempjRlvDHrbLhYnOg83XYadD29i7kv4XGyinrr7in/Hiud2uM3BN
mmDr45CO0RkZD8Q1W53FNWjt+PlWLmnMJmb0BCIsDyqcnwxwaNTdA6xkoubJzrFxQV2QqJEeKKvM
Gl27elsdrT8PZ/Ws7HQMP/x5OaFROJOhSii+pBn9B2ojtbDB3ntcE9uWfF/S+AQr+SgTGFDvcV26
U14gWpptlc8oh9IhNXh1OKcdx0y8SJVeIfJFBp2+roorEon9rHVuTkKHTCp5p5amh3zyZ89flfsw
vtU/rCWth6g/3pGsAUpWQcA3HasF5jK36rmJ4++hfZf1MGZBNlPYzpUaKhooCjiQ2AL/rCOJnoiH
MJ7eSWCfkwOChfwIbTjEHMc/KVolbDvVOjNZsfD36njk7SeUMplfG+SE42u+AFhIAqbQCD4z9hJB
o8bhFxQo81JBamSTCpnLw11Qkofm8KsPCOt4I5AUJ1mBsRK9QtkihWd4Zj4zBoClKIdg9W+a06c6
STB0bIiliQBkyBuOxnMLSMqen3le71Ija1YFzMK2mG8biJIQN7WPJqXuSDf4IyBmp0ZUctIYnV9W
c5yquhpLqlh0c07LXh0M1ppHk9R73T9Nx5BCqS0xf1SZgZyajU/W5tYMYVrapQtZ5jX/cvAbOJA1
B8dfjDNqEmWGfPSQuckBAGrPXQUkX9JehRA+ir2W7WmkRsrr47OlwrSyOrpDiuPR5LEZbkqVaecd
uP5Q4uCVyfIE6H+NqFY0RYPPEJygVvfvmVT+j2y1TCF90ICuK7TkI9hR+Lnkcr1sKlldp8gZs5Th
8W+lQhzfugtpjEB/YnWI1eWm1pBgwpg0iUaLU7EXBblxa8DFH5DvZjZOnWWUFW7grJf3MABWN8Jg
DHmo9jUvPc6o4vqjT+lU1GRmmlUOsjntBcYMk979n3YcEBEi3OJn7s9tuHoRlgNi0VThLzYwXSAf
I7FdZtb57CgPEnuFqctxo6zI0sZYz53niFN0zTw4TPDTXG84DErsRu3yeDJ4nfPlTz+ejvFeh6SZ
RNn05KR3SBvYxB0NpD7nwy/FSSu7EQIXxn5rxcb3rpLXU20GtYzDKbG+SHrOCfHEFzRQcApHEMZy
yZ0yj8l2+SWA01Xj5TlRfRj9q2C7J7tSFWY+9xbhnoGYuOoUmpi578o+Lhn+Cm9vLfPwdSAzOSbi
74R9WSYdy1ghw5Q0HDtVYoc9eoFmT+QSMAgI4uTQcnoOYRJEfG582OpllV3T2mqSUKG6PomI3Kfq
Vn9J0Lebkf/igeTq/6uQrmD0fGgd3Q5xvStLZr3fZRGkIFliXb1Mb60F0egXMJTsG1RZwVWBsTuL
8wKKSPe5Da5y27TNC4waY9onToY1dwSAMBTyEKAp5/EGqafGxQiIeQ+wqVpEdJOTvUyJFiOZ7nD9
v9O7y2UpK6hNQ6b6wEZxWXB+W/rpVn+Y0YFm5n9WfSG1iXLU4ODJmCpOBA1O8Cho80vO9JChhtNI
/2KMdySVLGIcuB5TICLOfSpg9oPfeE0nVaIi9eDh7gFJifWbL529Is7RHyyWvE4Q9bKxFp69OTdg
+xvE+Gn4z6u8CkKDaV3lasFnp3VuGNEJ3DLwLFUkW5XEGtfb3VyVH5XYgAhfTT4xvGTMxCdrgobj
513SjIS0p7PRuuY/3DVpTaHsM0TKLsZsyUA2R1Fev9MzXpLM2Nemk15D2dD72FsTkT70t6hcrwCn
KXOHW0gkwCSSLuMCFBg5pXE6C1Oj68mG5rdWMtz55qfqpSS2yHga9dl4CBjOtitoRkTzggx4dpP7
VKBvtz7lFdJSMgosBkzt0VKjHsT6NA/C2eczydjUyLifZibBmsYkT2H8iLwpwYeh5RoOVLq9bhjq
2TRcT1+id8ugdJWt18ehdKcsuk7jsgMU88N5kGyQYjUYcLaagCfrJLcroB2axSb4ZZ/Z9EKgtDq4
+Kl5Q4gVVZVg8PHCFjg599fE+EM/LbrI9zeZHZb5GLH9MUVLJgEPNeYa5tIN/jFRHGaiJRTzzygL
N1LvD4TrHdBTkE66bhUonI5Q33DdDml7shaP6YUUzCdrmgDwOlkWsN5yqKCxXUsFESTX+rpWuDWZ
dcQABWq5numJkIVQGKSGA39iVWAEPHyUpDurgFlJyM1krGrsqpXGBAbHHh5nsV2xcypRWJh9IR6D
JamARzZ5lCneTvCbh8AHQmVUi/Idjy1Tgbc+gX4QNujc05GISsZFd84g8xmiTL6YcT1zTsJkdO7a
EjhkLRqUB3UJPsl8MqMMtL6czzF3vCWEEzwR3FZ+4YemNFToVptmbt/zf+GdcX41AEV937GYjKue
T1awPtOUBJZOx5f4V6YubvMEy6wFUjtYLYt811v6CSdPEh6te/69SRVBvGvjRxtZ9/z066RPS8eN
KsSBb+PIbeCwtiS4GbU46zjmoBeQt0zhTAaGwgxHxoZzYqhVmxlUY5xWcMNahzzraIFPYH9CTZz2
G0IS7PgLZ9Rx7BWxyVvLqTBaB5+0mO6TH7Zib9MgplusaO3/Yn8TRnzgxLTKhNyxgpqmNJHUX869
a+0y6lOHrldZK59Do4/TGPNhdyFf6FOJHM7k9XXOU1bg0fxVsGWoMhgUaSQmLsc3WvHNWlOYodGf
IuCHgGac9Ph7B85JeE2UeNsLgc1QXJrZvi7b1VGCsO9SybfeM2O4cetXXIz0ieksZ1BcYqP/YbrQ
NzJmHyRGuWjNCBZfxbZk4yPPYi24aAFsUXxAkuXr/IPtemO7CrEBnqgrU6x4rwE7izorgpYfR96w
MV8ekQ9BEwLcvOE3SUw2+TsjZBL1K7+f9rool1vEraTMSh0v7P01CTIcxAzyn2rsF0J5HniRuELJ
k7xw0I3Zb68ueWppwet5/4fB8k1oXWvoSSJws7SA4FeA0QyVeaam1deQWW50xLAhHzd2/GWROpVk
tdjO2EsR3wp2Phmw5uM/IjEGAQj/F/Z+MfTUm27lSX91awAYloyfnc7jim2uhniMBRNjdMRh2yEf
QhNbh+7ns7TUWSleWCHtafsqgDbqhTJB340Ib3d6zGXfCwVMlV2mds3n2K/jrBlis9VaO1MUu5iY
gIyLZaybsjA3VUmn2CE6k9t6il6Ys1wBL1ULUR1DdH0Ke3PJDKKSYYTTL4cGMGrOkl8YOwlLadSY
09PVd5tfIlKm+S9Bl+REMXHyGO0xFKvhZpvc5BTqBa/hexrVhK3dEdXGofCakiCCCbv1ZSE6/0cG
S9pmh2Uw3LSeA69npTIvJ2ZdLmxxU7YfAaFM6j86YHlmc3PpkMPA2qsahycrtJ18XITR4H38GZcY
UX6zNBB78C/kspI140cWQeLfgPiqtQVPrfJEVkxy9xThtjbqtV1AWQVAq9XaxZlYP0SPaJawMMSQ
gM1Xm6CCyG4Tkzg2cv77cK7P+il+fO8YZyhUQ/YkPBxDn7hk4Qpy1aUrpQNraWo+tfRkYt9Vf6qq
IPrBDx3nuuvkZJupHz0HTOH+b73C/YFYJKpcaJkLZkJ+lO12PvAhBDvpP0OWhPWZTSyY1LLFzsf1
Kq9wo0gRoa1+SDGWHjlzG3kJULibb27JqKyR892bO5cREQaJIGyFn7Z9HH7iNLA7qa9sh4uUdcQ0
RNHcxubDLvDGN/0oSonuO36QO5V1QAiHyvBUUgll4PjkclXzePjz0wA5puEkIKg7j7wdk/096b+I
VSEkXeyGpP7v3/S3/EybwWw3McnmKWeHpW3d/dFWyTCfIl8+3l8iuej9ExrIYyX6FKRI0H3zne+y
dWcgjG4IoQMQvOEWT/ICUp0x5K1RwkSifT8X0iDwxcqB6UvSF2vD472FvDdB9wdWj+ql3644oRtf
h0dITssrK/Fw/UTSVO4EA7UfxvoD6hvPFZaUaGTNYWxZvV79/Vb12QK4ZDEILzINxJVjZ9CSzsQd
i7bOVWDrU9IpdIbG9N4gjdn6svoIfgjiyQqOkT4W/uLzzIe16wO6PhKpAPxDu+ZTgCoVrPyrxljp
UFbOH1Jzeg6oc9LZgR5qx8V+2dU47GExNj7J5acghsc5JEi/WndFpKQvYdBiHzOqYvcxSKDZabtW
CCqwhFEZjo+HN597+Fi5JvPOkab2rIasi1O4EQYo6uQjmzl/goSthEhFgZThMxL9NyWmMoaj7DR3
05xhSqRR/9KH5x9riZNd6kdosmyBcjmfhcVgjCzvbIVp984IjOHSWn3xyXYeYMoH52lo2c4eb6Sg
kNtOBSYD2hag2lZxr9ByCG6Lu08ixPei4YP7EWatZsN7xtIS8LsyjkL/MToxPsmc6LYEMpRLTLWV
r9WA5/Mm5Pnl/Yp8KijxALU3xsqxqX7e3ML595RXQGXtb2fB8u2pLo6NzteGgBkmvf+RMaOysgWe
x9NoVRJE2JlxnS0rVJPa+7v9oyPyV9tIpjvStA1v8bczDWcNI8nOFh1N0HduWZm61ZfmE/QkegmN
Egjzlvfe+vIlNpZHP+xCKwdIl0bn2dG7Y9TN3zfCETgk+z7+K28bEpRuWXx7z7b13uVvaGGqagbP
GtejjnRDiZzIA2d3jXlumnNbmZw6uoK50snRaO1LxfYS1uzm8jjokR5EmMIV1x4FLCqqdKVT167X
RrgvhNsI2LhcBueW06XaRd+uzi80+FEKqyMzkP0qTjrpWVS2mmVCeeuoCWEF6CpT0WAgIUATdDLz
sB3HpTmM7sjRLjsDW8dzu8h68X3YIeu/hqPaDDObkprl6Di1isITWsQn5NerWClDJxF4CPJsIBIE
Dm73skKU12N+jr38LxoF10/7NAaq933RtNG6QHuUVbvtohdbyP+cKmarU1Agf9ffCyjAJelHPJfO
ydsroimT0/eGX7fkh6V89YIaEm4Ol8iEKlrQqMf8K8QaFnB1un4LJYscBeLPWluxj6moQoeNPcb0
ocaUpb0QERvzqzqqR/BqglTk/iWJqgMngBz+EYW0gFrfLRxTsaxjqhS3NDXtxSVAr/BMITpf+jRB
mlf4Mmgx8+j5lKwKdrG7DPFuH5wG8MkSuuUQyeqFK3XJ8OXVq4xMJMo1wB0TQ4S1DCUf7Te3FnAu
7q/qBWwc/1PjuzfKdbAA8D/GY+ZjfhBFPgta8YgdhjA8zNJFqiKqWT8apB2wDaLuRN34iCFKcJrS
LpTxY4HvVS9Kks+xF/CZnwB4BjRJG8TjP5zlWLJztsT+NJkJVHLeOmdygsfBRlOz8iCcVQap34r5
zW6gZAL6TMDE5T58SK7TozxinRe5HAV4QLOsvRVrBxziqBfKWjzJHq6ExceZJzlv3vH8Rt2eqIbz
KX9DcD+qwzFQ1L6yGCgjKMX3YkRiSuTCcrWosnp1mDSX6ZnJwVBeOHSyGUR1M/WhnOXTShm4WYf2
yFpXRIONtOn9q8IgaVBlOU/qfSvmX4zlZxEPRk09/Zmtndzruwe/4TwjLDkW/nZSpVijrQPkRzE4
z/ZaRks5RXgzqBJeSuo2rI4zHpFCxWkyYlJqbRa+NEZJjYNakOvi0OCAHlRg42khuMhsTP3VuSQw
iYwZ7jyD5XH/zg9WjC5sof5e01AnvuKLbmJHAuqxSl6o3gQw7U5GEk7v/52BvyMyHnoFMzdufYrf
4oba/GW8pKeEyatZp0F9z39u6S6V2G/zNiGuRto/ucwQUtg2RdlfSGHjamR2clIVwsSDImEwBpHY
KMlJn/XYgxXK+7G6o2gCnkUqYW7aIrPu2u5H8L8keMqjkOFQQc4pbB+xXcb/SHjn8kzibISYmHWj
itbesFQ5RYSznD/8s/gr32BSOzI7u6otOaCT/9ecV3qNE0AY9y5CLkFRXf401anecSNxRzXBtZVr
02+RiYCbWWWj21zLZlpY2ehBxjPO7yfQjTmeIkbOjuVPBx48zwyoZdmZ2ymGp6K0R5SaidvwZ+cL
xH/HhYmHpVKYzZXkXux1ose6WzV9s+2yL/o3cq8jTOHa9d1CaePtoqVgy0OXWESjut3BmzpWKK7O
2VG6zVoKBU74xx0Lyq+pHlxTFWIVroqNb6+y1Q93XFjYSVdHGm/jcYKEG9f/lkXTXtqutO/4dR7+
A+ojmGEyY84bZBBwJ6crd3kBumx8whbbj33d+H9HhUR2pNstfPQ3957zmepbt0tMsjB7C9DZrzMP
Lcnv5b1q0HoC2rSUAwKCQqiBJqS9yRr3rXJAo61V8RNdZrmOBmqrpHYdn18rTCeRi0IAPAzRf07F
52s2Gp/H9w4VoiKTax25f2jXE7e7G5lwq9kHv64oAo96hBDTsop3hOvznDs/duI7Q41XpwnDrVtj
yqKpWmm/RN68IUNO4m06T0UVOIkmbtJEUADVCqKpkMfNk5GK0G04su/QEZqRceAvRCIR//yZm5qm
bMriS3F+AgsgdbnoIRoXZY4rkJNXBWHIxOvvUe8UXGYKFHcecVWZgmLlb4oTmPa9KQy7JC7CGNcx
8eSm78oTf7Dj/wYxWtGKaSiFAT3WcH35mO54BXO8EqIZIwmBeh+7lNVQ4Yhw5sfZlX03bVNW/+o1
Tygzbo6qP9b/xTPHlMqZRFXaNhO3AQwh/O3w+b7ZC85ngbHbxAXAZYaaVXJ21KEm87zMA7E2gDmc
vXSFfKDNqNlesYEvF//eeGc1JCTI5tSDOrY8V1APDkFx/lyUj/J5pzePqh07ObK7i7E38AU4RbEU
3Ggen6w00ekMsmc9PCCMEhrV8lH4W3WIbYVil9lwghi0FVEV94MslLEW15L3SC/bAI4a3grScbl9
F3+YfRVmIC0wdwnWeYr9v5IIQvaaaC3Q+nagr9VdD+bG2kP1QjovpOP4YgOwjwMXXfVd7lany+lN
i3GF6/PvzX4r5O8SC7qX1U/9/oqHzzJZ1mHxHwUZONCr0dWrPtkB8Dk9wiFUyHxeD1Cjkr6DhvUQ
oKaTDWeCIWUMUVYRSDFwuX9Cpij+QPBYzVgJ69rTOqYN+oXoTlv5fqgDrb5eX3rZYIYi2oe+gEdF
6ucCaNjR7Q52LwBGYvEhuveynLpnXXCEyCmyOxG5YXK7SWu3uZEXV4LyWYQbSSPv/latOVAaL0Cp
MCOZVf/21QAViWswxQ7B1aIaq2LLp3m/L0OQE0ot/hfSqcDJwyWkC9Kp8/PgdZ5NXNF7tCVUpZbG
M1YZm0ZPRbOVcITlDEGGsulMKyejSi6IszfT2ZTyZCF75stzZaxmdMaBAUDpotovfNOUZ8WNtORg
C3b8LoJCQ1LlvPb6NvdbHfmjBt4A/P6GYMR8eZLoKS2Ltwk8KBITusqTS8+bIx/zScq2ID8irfhV
2E4xWdiBaf97TNGbEZ2wM+oEvgKuFfKIY4DPZb8PnPDoAQwZc/X/c5kxwd6RP99zv/YbJq7iXf43
cFoNuXv0qtFL4JSW96RJsby8+p+ICJqm9oinPU91gDjerzVHiQYA4ZXSoYuSuXiERyftF3rW1IBD
Jf+13oAdipVXVpPA2qNqTXa/G3jy4oE7FmjKOa3S/Yleu/BUNgtqG+Gr0/BVqUaBatbXgpke4MM1
m/ekm3ORKlK2hQe9tMN3E79GZAmSWbJ4SNVUSYWDVkqUE8k6rMyOQXnVyhauO4wWwfGnIzPHwf6f
CXO58vYokTOAElIeOBpuuShQf0cY7/YJ+P7VSikaL17OmF7cochUzaycgFpCJ5tIdD1JwCo15ekW
J7qcZW+sfVITEAO+OelRz+iyxg4BgnSxmwxjlQV/mFtBIKD7Y/mlAgFVXKAlKWTg8rCwS79lnUZP
7Q06cC+9XWdqjhx9NzSWDu58lfKObe90Th46rwIkrXLmn83+O3z5DzvAofqYuYbWe6tNcXsNafTJ
df5Fneq//ASYYmo5jRN1s12shyDFdIN/rtF0ommcvDHZjcgWKjHeN3pEXfwvpK2J94Zfy0CzNCXr
0G0nojxF+262MIaHlDhHQcHJN8P3Y0l6JottmrG0a97ZJOSBcDBbkfUHp7m5r8k/dGC/xvnz/0js
REV4At8kPaA9RbHSaV3DFuN7DNo/4J9yFEXzAdTIZiKxKFnEW99QZpePc6SW2FjqSn5wFqfyXtme
PjWiTiVIyaalxSIfaVLFCNXcXqtP1WMG3BhQV23tdZVJc4ca5POsHP7jnxJSGtNYK4GvXez+QNeg
RStuPHXPIAn4Lf3Z9fjsY8lQnoVQJtjApT7zbFkgCj9TkaJFHISL6+Xy8ogoHwcAG7go9o4XN3LT
o1wx8/c+N8h1tQ0YyhqFQA/TJG32h4WrX7DX6ZJ6ywWAiiEOdyLnxFh6xBu/rh5gX2piLpng9AqB
uHpsywIuUn25OfHnw8Q1X8jaxkili0Xoi3aA8yP6Sfrhmbq5utrTpvY34d9o6z3+Rcxaq3SLW2Oz
jY8O4VZ6ctqGW15p8d7CwQMIWKY1bseuKg0GC4ZOjj3JDflK6sQZNIBVa45V/l4B1d7GklicWeKk
9d/4peaItUBQ8qbDvHqIoon10PPeLrVI1ljwtZTq31YKmcn3zs1GmjK0la0zM8OM2fVy7XzoRfDI
2F+F4Wpo4Op7wxpLCpa23fVr5c9g64xkKPHOmpayknEi+1gyShEWo43k2cvBCA/tY9wV4sKHLcDQ
htNheXc979phDZZ+wJQuhJqxV/iwJ96EDDCuawd3tDToaIJDxh08qkfftk7lBmVSJYwjJDefHPri
ikUr3yvLSzvlZtFhT+ZSrSS30hDSb6qN0ei/XSnkMd4PJSLucmD8Uzqz4q5gZxadXMRUP/i/c0nN
BiSyFsXfZjwa/7PTKDrQYOT4yVDa1YdifHx3Z84ghpyYDUkaqi7iowNwAH+hNRU87e2Tv70Xw4jv
mKby1xyHK5OqRcJTs5c8TS5ar359akxdpAfd0I7AS0lCzyXsUeNWUPisPDZYzX61OXz9hw/1S7C+
Af/m59lvuYFNfMrp0B6O+g65DlsZ/BHKj3yjqFKG+kIXJv3dmOCx+/xGfjhSNPljoDmbWEBqgeQh
bBa49g/v3cCTopZw8dghOyI2NIMH/loOYd9cX0NgMduQ7CSZUGcmzIvDL6GafLEytEhuxeWc3hrP
EJ3LdP06hkGXLcduZhwQTrL4pFlwODfLKArUJ21gKppAw9YCa7DLv7XW25jj/9c8POudmGKV+Eyd
ZRaK2ugO9xgE4gpFUp5BGiwK6URkebiLcBIZ+7g1Md+yCKzQ30EDl6MT/uuPvysZVnPMPJrAeIyH
Nd9vxxWXI3pjXdeJRW/w15MlOCHl8IJO1pX4uEKUQ3Ly0lGyhWBTNIhO39UKK1Lpejyh8sgY7NKR
+zYJSn6OEmy6sVKACqi1NMUCF47qDl+uCfWWoyWennbJFyHjBV90LomXOvl6DdZQY+cjM2GJiROj
8M4CfKoKN9pof0DupZnHnpqa7Mox0shsvwIYeeFvU20Gfciq8VbQUhuzhADQh4Lf7wDJpUz0lh3D
R8aVXFnb7IEsyEcX5OpW4fyRYUyHrpAPeE8o80yMTbc/KinnX4nUfEj5tz/MY9phVhvGo7f8dgWa
G6o/JwnInU8tYzITv0q2pGJGQAtMKuFnIDKkwv+6/dcwoMVToduEHOdVZGyLjMbGvxkH09L2r6hd
6HVXIgTtwjNTL0qsRb+e3e/lvOy34oNZkmt65q4RLzwz7ddw504At8dvlMUDkIE3OcfNyeACtDL5
a1etJyYhdDxPjaeaLgFqdgLVsEa5rxTcEtCpuxzDH89yX8ASoaOL2i+55K1v7Eh8ZMQ0AOFDvFBd
WMbjQIKA5cKP4A+jrkFDfG0ulWndsi3fj+2z8jIDLDDb58GlJQa9T+pwKDrfniZNEw5X7vpNWzfD
ORsLypNGPo9e6rPQdiIpRYgmuAFSIzfBmBW7ChLfzXl2zfKccZ0AUk2j8HvrTTNGfQD53eRkulHR
Zht4O8PIMhAbHryzT5dHdS0CBGdk7TtSzR31sw+HEEzjcPzI2GKisNuVYNbU/IhPlpxG13nRXB1I
i0N1ujRwEkyqQJZfYbryTrqezQJ8BO/nh9bs6Hi/0F4bNvU5hmzjKjYlCrhydR6HE7FWtTJOqhM2
ast8FkqQ9MZGwNA31Xf3T56hAIP+LjQJPWlhced7jKAoiEExkhRT7zJAMobvleONt49MyeP10vYY
bMKmXHIWIwNPs5F9L9rFcLHpQ+EFbyl7qKsfzDh0JvkhOL2JuE43i6JVtwuweChqipYD+UL+N1Fa
qB+FHXTf3QUpH057nwdWZMiuew7e/+3bRNzkCBXyDoqGgGtebOHWNxEJJa8J0MZiggivPyYLqkYA
CfTv1Dg/ZAWJOmUW9W1aLViaNTALFocjFonHmL0Pua/UidZd/Ap7yICMUOyWRNbrxKoey6Ba2SY5
ypqNzAlEgFVoFYAsn0YBLI1tNldpjGqnqReiMaguZma5ayiSXdA1xxo28UQ3FNnZOgIRKDg+3AbF
hg6AIgaySEKcwVa8GF43EMlXrUJMzVOaCurnk6bX4JoSFQvUXBwfMSXS8RL2pxyXiwQEQrJ1TS+w
6Rw7NKH4JuWbT+vs2HtJigsNr+4W/y35+mZgR8paZOce1botaS2l+DAZpOdaZKADBBiLO5dShuh0
wgbGimIqLmIXi4nY0SkuBq7xSZZzvlCn4bWJNDi2qWHLqyHCfoOR8fHIMYJHm5KhDtdpOF0CzDo9
RSdqTQ5Zp3jmgvXHbw5+Q9xRrpZJ3xAG5kMGfiaZfJQQBQAO5TsSwETzsWLRR7/FuZob6X6hCu6y
jKPbdxHVNLRxgSpF7RMScmA9/+MZVqAMUMbP5r3qI5wrCRLwMpkTs+AzOtaSO9kvt1euVWMWRB29
UUpr5c/rcpHgxJ6l7hmW/i3qGI54ovrbeVzeV5d2znyWGhDzoXe/5B+eJE6suaJYN2pVGvgMWXi8
XifURngbU1haN036QUb3ndltE3ffsXQuIepT0G9WRwy95LVColiq6Wkgb3YzaGjvX6oDzATfxul7
fkArJjvBY+IcO9eaZd+HXYLJHiq6cf8M3po43XXYlD/wTDwArW5ccjfFHI0eBPXmTrIE2rXPdqgG
eGUw62qFx+kS+pQqhLkk0zmRxgbtacDH48B9pDK1JbEaqxPjd0ljRCN4hR4UptloBg7GluYURjBH
kjumQR/ym/qrtwY+Gkz1acjBnfrVENj8T2E2LhH8bC6+AkklVFdEo+C8eSpUVAiVxzVIM/iZZRuh
/BPhg/jNr55sRigCA26l+Fc1/lPDoR2+45bn7WWi2snnGEAI4xQ4pKvxVj4ijX2z7VKeZflrtViy
XpX3QhsgP8ubSV/9cQe5WAcXmgpNe4JOso3UTxHmgdayv8wLEzIaQXw340d1tAZaYoDQy/NMhckM
uU573AbDKHTklVolue0iCB4/Z0dewzb2GMw4IcAgs7HBqW+idzwSlD9rJ1DVfa2H8ubrfxQIlsU6
73BaM980zdUW0GkXcrQWZXFtMpnlGIthwOQye0lN8QvyQqt3TdruhL8EDQ4Y7t1f3jzMXxGvA61Z
3VxFXeS1haA8eD3mB8/qGbEzLm46Eth5QEdiHtVPI8gGtRLnq6zSaGPnf69y3pWCX+HU2UppazWd
SKram2dExxK4tEozzXsh8VwR5AaLNe+3TBytXICwOg1XM7d46JKYsi9/dqQf0VIX1rhOtZth2PPM
QeMJ180YRIBnlPQqwMUK7HU9fduSCknIxgYIaljB9exJ9FBwMKEwBSX4LTi9fSL8zR7z3OfS1kT5
JIixDFCO1qi5rIbCYk1ZWd6rKVMrCg/OFecjxKZL7NEdHiCDwxhBLg5coKjpVbbcb9wVCr1g5UWw
erObhu5YIBl3il6c1dNn7jFLtigYd3Sili/TlCJTiyEWS1DZoDu/pfqXu/2HYOerOKlGwhKO0FNc
ZgWWM/y+BiBlLINh6Uup4P4v1vK9YwIndDl3nw8fHHxerSwz1t6Qe+m+nRMI7yW7FmsmTCYKZojY
sCx8s1vKhnjie3rj1Dyz9kQKSsm9B2lhQvV14666gOJWTL5xYwCBSBJ6BL/xcAYaCZMRDaKUFV6i
LKzoNPkoIiM7typ2lcfm7QEMVRyH50S5DtVfncCynUGTe54vGQ9U0qBcLTYef6DsyeFXX/EOFwO5
bUXrhHKIynlCMQaeWvcf/DLtETtCmE/xtCLxnUdHOk43SkpG8ZPeQGR6Q2ca7s3SGVUGC/PSsogH
VODrb1GTipWSDSOjPPJcGokauALqPwx5AD4vlnLuceJV65aUmz0YnnJ2wQ2L2OevWLYzBVQ3SK9X
TzNndvgecY7B2vTQSLnJ4io48dZoSJ337hrVg1tiYbRokr07uTq0Z0Wr16q6/fKS/w5DzNLKM6Ux
t8oYa/SERlVgjuLJH2eM39wqT3wbTgCL99QjwUuQYk0z9SA9o95/v3VRAytfsp5ca4MU6HBYqU1g
kAeA90w08efAILQRhnwHNigO57NJJyFTSvXv8NHl55a7OwmGHwCn9pbxSz0IAPg3/ajx+Ngm/Ppq
LF/7juo2Rgw4O8gEk3xpz8qaIt7yZ2NJ2OAcaMlMzc3413Mz7GIDuqqPtaRg3CEkOeQMjsHBfTnx
sbzTsE2jUqpu6k5yoWTr4UD66LFNEu1Csgrvehvgv775rlUT8gfV7ORNJdTBfX9JM1dwY49aPnZO
V0uLyIGOvo8ktjteYwiTnP0c+Lhqc4PVYYb3ZKZAz9pustCptHrxg3NYvZl9oyF8Zah9BKXOVCLm
DMp8kWWVtUrN4nvZy9HyUXyxw0p56BHH0jd0nd5Wodz+TViYO2zHICBeJr5fkjskSll4gb1yVp26
r74maamCR7CUXDFqr3hDjxDDVa+NvAala2pQUr2rihng1ojJgkAJpfJwgMVsblW+3QuIknST9mdK
c2wbEPALDp2Zkv4TFL+v7Q1HMhdU0k03CXeuJIA8FandD29cdDRP0cA7YNnped8EqyA2h7dFpJ/v
ol/aTLQ2fIqVd4h5CRXvcpeEvSlYVwJDc0/RYkrfctkTN5J21Kt7fwRowZvDogZo3jmborZauELR
ZgQOCusu/ftYtFOWq3jKkJeRkPzfY0TPSZxhr6WZvqKY3+q8irwGLlGFV2xcDAS76HB1XjP7rC50
Jm6HKQ46sdzmSoeMNRvgsBCZwMOHgmF42t7KZwr4q7f0itkRUAJA7lNxmDSB7gMZII8JFzA9PeOG
otPeKgSQgsn3YXFlR7qwz7wN29zcMjo1cKkdv90r15z2a8D6zv7F6RP+iDZ1halzsxzS0PlujNYs
9Z/6KrWbmxKA99Tg1LcRfCUzTYX+3FcrBSq4PPWpF9FP7yX3byltbn6YsNjJCSMDn8wOaEb0TcOE
fIb+7PzxCn8sWLSx2V+wGAG/J7bXXi4jRiWbOzpc84OK1LyFb/S/bbGs4Asd0Yfp/KagLuorkiI+
+e2ERkuOkXkgvFsGkRYf8l+7qowhDyiws7OPfZpFH+F9DC1B2cfnzWvBu7nk4i9PVVGCM72n2yKt
uW5FhWE3XFPGbfc+ceXnJH4ap8GUkofSZUIWV1Z5Pc4CB6WJY/6Si1bGct6x5kTIN0tZAwycN+8d
zO2bD/7iYw40ldCZAziuX1MphyNCvTILViDyrHC27nh8SBSMOmg2vWWYl4VV/T2U+8SOqbwrUJPq
+3Dt481Mxz87jDRytjlmaNAkKexmg1yGbTf+VbS1V8L078j3ND6p5WHL9zXZZe8Pb6ldhYb98zcJ
tBpM47w2WDoTkpA+5viQoL7yXFipE9t1R+T/hW9aq4lGWIc4okXUeuLfrO7l7BhlOK2ctC4jD6A5
4Q12t7yR1l7vk22McPfzjkpr7uLr8nmDFfLiuVTZ3K6ECSvsOoYktK7250mzdyNo0yPVZTHllm7w
Kij/E8CwQBZ8NFM75a0PA4BIFMy1/MCFOgHY1gN7KRQJBo7alWdq/e22HRPYK8wRLZErRSf3U5/i
qRCFDfDWN48WhWVsH/EyTW67p2Q8EsIS65eKyngY7KK+5/BqPnB0a8xQH+gEI/aJb49LVymGC75p
QFZIV7IzBjVr7SN7Y+1bFogHLNEyIT56yTl8u9LZ0VLSPcaIOBP8TyzJP6HxWMnRn/dCUtmFyi6j
HEYoQUe5oFlhxw+78qzgog8t5GIEsO0hL5t8X2tX294JU+2SDC2YEDxZHAm2xIEoFrtgcdotqMIy
PYnUHMZSW0jcQy4z8gPNFtzb+tH0QxypoILkWLWWGFXCcZZGtaSTB/oU/KZzuVhxk2LmtwDBMyOa
JJrQq+/ss7PRCyU8hN+wpHLAHTZmAc/SSr1neweDrkDyy9T0h66aD19bEQxZp4iTG8vSdZFdZ0Ho
XFAvRgK348gNDedu1wyWR87W8vtTXK5fhS9wgbJ4Awu/zUZgQHaDGEmrHerPCmV7cwQCB2k0vVTt
bHhbS5/uZ04Hvhs1WcW5thDozCvxuo6r5OGqxsrPeG0r3mZs5tTXpzaMKPuBGqlnCKN6SPvzbt+r
+H1GUNEmZEgLDmdM+dnxLhPpoDVh+vsM8tGvkp/enluKNeutB+ZzmoV0o+3Ivcj7h7NRDQP9Gr5X
/OTe2CyRlaOhoRju9hiALnQcg5uxUKVPEEd9o35ku/EqrlOY4CW8j46PuUwfucleQm2x1Tzn7U7M
6we27zEXsbctrdfNnhEmJd8H/sjZt/g29UX9xbYyuxSSuk/gHLxdJBdhX/6z+qTvUFUNm5Z9+jXb
VMAzSdmeBanxiGHd/2wwhXmn0sr2kVaTNCtSymML41JbVHvkmM+O7dKxCgx/vdsZNwTvFZUv66wT
oB4ouGgWyorjlo6Xs2M4lGUdYEgiuE9VQ/NMQjFrMI75g6nSUoDxAFwAnAFKlq4Pcjv+iIpJUvSt
ZhxivYxO27RUoYVerto5e7/o986kJgoSToxC/PFHhs3WIi5xxntPIAGiVHcPOKJzlKpWVCU/VXHq
uIDxjJ+2nTad4eNZtNoBTRrYUillRbs529O0ySRamPuZe8WX3ySBgPVxPa6nAuiwR6k+CIjRcoDh
XPRPViJii9gtPisjrWk+I0p51F8qdve1bQOFXnQ6wzOCgqfCgP2SuZn8WodNGop+OhsdiR3W1AkE
OPdmLyNs6i5I7br0SOHxvRvci7Xad9wvNRZZL0TgII8c54D+NKquhe9gdhneYss3l7d2SnvK7uCP
xHyeRtYh5s4Ub+1D7Ne45kYZpRLz7dh0bHQJ7ekuTMzgp3cZCZesV1EGfE27jTA9K9N5AFV5Y+Ja
XTcSVX25l1H7VHPlXEEIHjfOP9YmFZnVKkjLFdQPMFqRnAE7ByUz3xX4YmbIt2hcYyBULoGCI/nI
JWJbAAVc7j7zH5udFFnZfv/I2HIKmbHrF+STaL+zp5v2OsHh+XpOE2MPVD0gof9w1W+aPBLmscQN
1lpUXAPJLNL3WSlZh6zmRH5k4k8XJPoFDP0MGqeel34d/zGEF8pr2iEEko5vyyZUfoXd6t4QPut7
upmc0zc87MxnURfYEGxnXyYT2AE6+nxCG57NezwGCgr9fT1tNzQAwnoK9LI4vTKI5YFjfByCRaNh
srMINfv/BWtSBq3rW7wyDazY+n+inVbp/3qsNcGaoY5kUjmgbmng9c1w1YmvjnAjykr52SvWFGcG
C12JuoZKSpWIc4G9WSYolSQWS/jOWBt0B8+uGaG8OV5YreX+RwHtqaGJx3TgfQryATCrHKbIOmZM
036UaoyEBxq3LsAPgvQ9Zc5qx5VZgGm75JpUaFxQEd98qj56qeyg2Gysb5Giie/2HzKrTGHWIBQn
riUX/M28eCg6Z1jA8iXoqnUhU28yqAqw14VmkuXXByKQDA0BRaxjzgzz4p0p+7lbZ+chDuJDccTv
e5i+brgU65xYlo+IZMrgtK2wTNPCndrh/mltJpPuwaCRWaADwYMgsnx7XTz2+dme1Lzxxd6V5/OF
qM7RmUqGrX3MoyfvJAam+OQHqBiHdmm+77HpNCa2ty2jTN7vbvJ0e68v7Fh+RYCf8rtcUfUp6N4G
zIf2W8OjfrGWWdbwDS16WZb07c1Q5d5ze55lC0jrCJ+alfaudNfi0Vj3VfNmeBM5FV7Az0te3y9A
27PfvS58IsOb0THe82O159nS2d1JQvr41z4b39rUxMcWBZyerdSwekyP5++Rq1egYIP0+Wh8c7J5
0GV96KsLVqSSYyPK06gWlLYRxCwfgvxzUKMPo8ArvBJtCPrqU4XEWu6aqlbdt3026r5zanMTUPzJ
cmnGaYsWcsTlpB7MKabh3/svJQ/h9Wtk83AZzacSEy201VzIkyjllJzSkTK5iIWghTUa6IRBbtHN
2GJZNtEfi3GGNAeTb0AEmO6Ccrsesh97QnNVdNr9A1KlGHUjAg/uRVZtK2AqWmJ2bocduISJoam1
E7kh7bppzd9wvHEbz0hhm4Mmo3wqp3mqqAp3unQTd3Yq5nUeyEHwtN1vmYb8NQkvzzcuW5Sa5+2C
qYWGYqGbV7GkI1dCMEQ6m90ikHLALhdSYZD+DS0CBDLjRBPnC2e9Hz1pfoRd/fB3PivCSmq1JJtI
YK6wqN0QkN6MCGdNmfIF8w/S5uJYLr6brHuSoM8MGqT4MlCXEy3MbJlVmTjTmjRKG0SytN8nXIEX
uR+XA8lVwkb1Poa1fVkacnh6HF4BAtK4TsmRwRJlG1jVLxLRBctOIB301zDIxNYvdw9CIcjmw/b+
Ke1zIkNB17HhDJp/QT0frgPdaHn+2chg0Y7uhU/QjN9ZGk5fst1IM2wLsyCtDDXMtpmF5IshFVJT
QuVvmQH7QMFirPI1cKraxk3K0dmNFb9pNnvdfiBd/7Zd+QMoXpRCXhmvQDD3Kw3Qt+lh8h49YA9P
lHXQtAJD8X3EsVxcL+jcuccMe9sYbPcJAzyK7+JG1G32Sx4XahkezhXnoxUcOE6p5YPBmDhYRw/5
ESH4Rh1SJMMdi/WGFlqrz77hrhi5Csc8kxpkW84ob4OH0CHP0PU/gQ3+wwH3yYb4DtPeVwpUcBEU
TxTaTCHkXQ9yTtj16Uc3Ary8Dkzf7ec2PkhcKwveNQDU/2pHFt7/RTkBXiHL3H1OQonHmIQXMOk9
Ly39zNo/cOlRR2hi0RYNB+uiftmMwFI0o0jyDIYq0I4tA0TZv2myoEzqI9XhnY96AW0McU1ppP1N
70UYbTpY48ZUW6+68HfGi5T0SHHlt6zLnDW6+5hpN6/d/PLBwRBqHQl/ZBFe/YmAnsvaK2xaR5UZ
PeApeVVW6n0U83hM7pp2flJsVLadSNE3HMFN0FmuAeOU+BwDG6bHVWKfNxR+7O+vD9kMPCPGfGO7
QQE/Fr3ChQLY6Sa/jnoUHzjNaeSNlahx09WZLsaXTavC97Kza3a62mPQmFh7cDHuVZWppEHIXDdX
qBLWzG3S9ADgeXPP8KnJ8c2KXMd9t56S1ejMaeT8Ti9/tpj6DD3URUDpJHcKqOKEORibD4i+Poic
z/pEF1eL0RwurS55042U6fB2mApUOoc7Azxr+dKVJEUo/7jZKynxje+k8g1aZpTi9hWw8EY4ligF
v4pJFPEnXjPu9+6vIQap8RcpsRGTYaTdu0azhHqT6xCbK+CFdbI7729QL99VoH9uy+CEYPJhMgov
slhF/AIGEfB4vQVqthtf64uNOEtMaTNs73SLwSyrVFdjVe3xhJ0RsfCSrsc8BFPHNm7GWmi/LK0S
/ttWPuXRztt3G1lfZKJERoPoltUSVo8jMCnuo+L3+/noN+UAIusXGK0Yuv6EoDjPhpOKo24DX1QV
hc71zci+tQE+47iNXhbFEwR2nOCb6OP4b3u3zdlEivfH1D9ARl6ZEUEf/Xm6x+U8CXZJOdvMN3UG
Ljkwk4k8st9LjvXoTQtLtsSVECHfIuGMzm9xbB/YClw0m+VToQflSDtpI9bNcmzH5pdqkZae9js/
uWvcWjekMPP8uST4O7zE859jtvxcw3Ej08KNa7GVSZvnjLP8NVW8+tU5npbUwM22nhtuhR/4NDfA
cBOwE5hx7UUnjfIMeiu9I/lUWnSAuiunUUbCjfj4TZrHRvArVjYlsKeVzr7RUw1wO6Cv70Tp2WZS
5t+BvlSwmBOK3lKkBepPBjuob/ajAe1mJOSmbFwo+m0ywLAs4XGf0JHtL8eLY9qGFA2X2Om9l1sr
/f03qws8VPa8CEuSOUcLvB/o2RBaRHrnYRdDEM00sOZ0aneivs8m4AL0LuEtiEqk7Rl9BZyhyry6
RhE8Y7XvGY8KqtzK2E/zvbhPwe880G6yx6Gb+EzjPb55XRQ16Wfu0ACIEjV5ajsJDBMp0w1DqM0M
dnrdNby/0B9G4qYNYwFH5AOUqC5AvpgCoIBtxHomBdFiVSWLAQPG3NZZKIqx12kSmWEBP/CVobdD
urfRC0eixClWBLKWGIP0E+NNenASdcKd4N+Gr+5vYuctxN05aDyN6k6Mm3Un9A7KnERtWbXZt07x
LivFIVJQ5flA9t+JQBXd82otYk/MiQJEL+AIGUx7NrqpdlKJH2chHO5vd35p5jP7Hv+nQ4Y0kGyF
jFit+zS9QKdVEuEfdurHc4vBxyeR5PzmgqgW6tWqzEQYIhu1io+/B+UONMALDXJdr0fpkRmxQQmq
VTheKxdAfdlM5C14GPKd58PK/ZTq1UijubXZpgFAE7CMakEs11zLCI5lPj1DXWGMibxJgIwVswcl
rzb3hUqbXfv56ycSJo3ddepoWEeKtwyEr3CjO/iTqsEKUWkOQfHtO62WW/IOfVZHpyJ+tBCz88JJ
w/yCS/0ChVLM232K6aIW9ExCUP7yh/bu+jqNTDFqeOEwQ7DrzHUqHm1DUATCd8JZefQuocfv2RkJ
DG/DZ2nqxW/THwmPH4nYuZHFIX++aMR/4ce0Ze7yUean2+GPgaYvaJCaf8SVyOpUlBWeMCGWLw1b
NWaSPnbIaFi9zxiXAH/U7EiSuoWTtxHW9irYFAXcmx+kkdvV9u4Kfa4PBl+klmDF+JQgv6RPluV1
CR7SbTRW/GE1zu6PVSmhV1uhKciVdunMyJwOR6otxex20iSsdo5h9giXzxFyuYSVFLFnV1gq54WV
DEdJd+oIJsWYKFHJYW0QLtl/HnE1qJOCU1xl0RpEbiG/vq2iaBQ6P0UeWYoWskleP7Ly5zgdHKip
q0GwJoN8wGNXZUsgEMM4JVaTEORmRaSrvH68FgsQ1DAWOXj/OWVtui31YSWrBGB8A+BM46C1zkhN
N0zwLX2iqSQybRb+KTTIMTC7w9fXZDj/Xc930Tl9vsgS4numIPm+VEXEwzajacSL0i5PXT5fwQVd
JFYk03JkSmqG8FDvUkiWIqkIoettY3mVfXJ4MakCR7mvJB7t7OS8Boimjjqgy5ISHx91zDQU31yD
vHcl24IEHZfBbDcN3D3c87FqovHTfIKr2lafSAstpi4xSsdckFxlaEwJxhh0PgIB+nFeHr/t0YI6
Rzj3y0GvaWWKzqlJUbtkyCWertkMS41nPeQ3NkV35IfqJ+m2qAZ8Dr6VTExWVxNxu9x/y4V35O+i
EnHLw0mLq5bkofO1rWJ9Y7V1eRGHlMqAQ7gByeS5Fgaf411khrgOAvh1fYcKtYLgvUpnmRGLaVrI
uLUFATm/YDcUTgaOMEsypo+wVCAygrLxmCj9DeyIv3mfXlH9KsQPyg/Xeu/qYXsWdnSSBZ159OCe
5VoP5qQn62dXA1KNNL4PlZo00Eyzn7ewPS3OCiqVrbCYjdjCkVTgRWPlq1n1ckprOjlibwWWCBH4
n1V0tyG7l7e9uokTa8nQiS6io8p6g7tHdIAW8yLjWiEPBKPEiZLs8y9ewHdXSWfQ7NN5sggRPjwK
c3L/0+2SvwcYGl67gQBIee8pfeO1+dUuAhp7UAeGI9zRjP7PEJh+yHyJkCv0odlxEbzv75EJgva2
QEVwjG5TCw5dOgbKs1gFp60tGB+9M6JPQSWvlCndB6Z4krCjZ3Pw+uEaQnnSf9zUEhM87Qz3JulZ
jyaeEaoI/ere8wk84ezTqe8F6vyr07KaplbsQgngdzETSmXGnudgJLnpxKRUbP0fAEOXhWIqSEkv
IGMV+Sw61lUKncWIbVezGWcnMJ2Nb2iZkgz47/+3+k8z1Epwh/Be6kp39zAEpBieAHw6vWYnz8d6
h17V8Apq8erFznbx7KtiburhKvIscXjMFrJmQc3RKZMJZP0SjzYcLqwsuWtsxAQIUX3EPsnkEK+z
ltpaCKZg9NQiFVn6723fbHTLSQGi7ikB3KYvHzQT7f0YhtZNSuzUmRgkuTOPcG1wIINoSbku+qOQ
mC4EVo4XVZq1/JXslYLicK2F35L8zHuF+tQyzlTISoRgvDIn/KX/AvjAFL5ijFvtANtb5uIUz9h5
BWCpqcpdlD1j8cPNn9G6lt92ksAemvM4h67PgbAqishwO27gf0/TPXY9FfKY08knrcfIKrvCyZdt
7NqpAdpaPFuVxCeQLRleXmY8J33sxKOPexixVDzuWzqMRSbJcU7hNqOAB2p7v63W+e8zBLy+xwEd
A7RrR+Ub8VZfquEEGhUW+RyrEzHPVwk0x0mQmvyeDWWg58IPkt3jg50/m6QJRsWIe6BEvRW195mt
nwM2/FD5OvixL33tjau/8DOMawj1HmJUb2KuaONr43wdilBYiWA0KtZU6mRSzRcGaIqxibMc75IY
4dCTnT41Qla1xN5wf3hxrvsVQYH0Zlw9h/l2k9mZd7JcDeo4ZP4MSU93MPk6qvbZnGJi4DSerkZp
/2DM3sjFYPzWCu5I6nM1Aw6d+hDuM7trzt5Lnr5aA4LLvYnGjLZzCPpmDQGxUELkbjiBcml8cI7n
e9ALKKpJo88l7t/7GhlqmvfmYJPTTJAk6FhfeuEWPQ6Yg38lNXwiPUspSwpTAK9dV3/Uw356vfie
VosPtf4oeFcAGm1wJcuNnrWSQfeERWUl/j3VAWriEXtlFn71ZFyL5rEZLMPmdWL417DtGMgqCMwU
opBve1myZOn+H+jcprpYUk9Itubr9veZONhHUvRZSVyz6CcZrcY6A0sXTKbKU0nvheeDxaT745bp
HBafKke4HzIWyhK8gDEUiOyi8WyY7Gm961jMAhMMjs5qN2ag2tohUhDishX3874icULsp+xtTgPg
Jhu63dVIQukJeQIfimyyN89KDPrefq1LE+yRwIVhw/34pgNMooarprYLpzAYZSv+h81/lAiDQBcr
npLqLXHkI/V9WDZ6coKxvHl+RL11LtCpr1uM4Y7s5+0I+j04Ju1F/NzH+V1RoYjNQPpQDR25H9oM
NZfnJ+yQMVUzH6FIWKZAoBk805iPsdSL1NUU2vHMpuxfdN9OoWj5xQprS+KStw2MgwwaW/xSEjnD
3AQPC5pbhMSIyxjBz7SyKpKLuNT1K3GdPlfiJuVQqCYMi406rfgcTt/Dgg70NLd8r98ZSeErcd4/
0oa9/v2oetUFigylunCtgypQnovicvd1Vt4TOfcNPbhvVlwhnAe4lx1wFX6pdDgwTXwHqAWT0VTa
OAUqtWakPRFRyCSJ7XSIHjNQz0Axq93WYe9Z20y3WD/PfuGj9xm2m8k5DKAAzDAczbNMIMjXR8mX
7qOLpHHzZOd5sagoxU7epiJ+AMeu/e73mhKBsctsdQi+9NkG9djrWHQMdF7q1kf7oE6v9kvNU6Tp
GzrXKhHrID0GXLgCjpJjRZFQj+jq09f+OWD664TMQrun1K4EKYnPZ0GfY2uIcO9Ovv5LJwsy/zwu
kWr2iC8mcWltfQ4H9dFvpBf9zDKFMeDyPl5jNkWuSFNEYNTP92aUMA08VB/T928cE/cHo/XHZV38
5/6JHLTQht5B2Jx85LrG+WuexYNhYksbf0SbkhS6GPfw4fwDBGZbSCnSblKnc03FtGUjvO9qxpx0
ki9ovbUZdbEANdbxx3kH2a61fAkE0wRg5oAuL5z7bZ61O/NXzMthstRUmTYQc3SOfr+KuPX8lVtY
EnWwT9VQ4kTFs8iacWXxwKEBYd2ODZLXJAncOkGyI50iTsyND752qayQjmjHKFPw75qiX4fYCnHG
xSM1Hb/rT/f7WT/VZuBQKi1oPlQBdF4tQ9wjORkVRL0F5Zg8twgFPimivnnb/dy20xIEW/Owh4aE
44eL8+0870Fj3fsYN9GnY80nvCvOzn4z7FyDb54ZaB/ulqnDGRY3xDqB3XsfsYuF83Cg9fG36Kft
muJKJsp5qb9o6u2QkSgwoLE+oV6Gy5yanTmeL18mdX6uQTtf2M8oTlo39liuTNhXgr8MYsSloyIW
fw5rgamftZ2rcl6nD/Ixu26ynO0JQezrkO9ugmJZ4Pt+AwehSaUmSro+nI8boPf8z6B52sqxRIVU
yJ9HunLmosi0+yBq0MGLfmUB9NEfO41qzRP+ZfR/ulPsfN+9QC4rkTHXO1SI7VxMzp71HPm8u43N
qM/DpxbBVUSlEF0SH+IUKpecdDBYwdTqQCN+grKxZ8XCkLnqLNk/v8AyPSpHajvputeyGBLrKt5e
USVBlhLa99Kb+p6aHmoWqPeLZs+mWtaLeOIVcwq1OR2YnbYRG4iGySu8cze0H8S88KDB/FV0fv3I
qDeBvBD2oTG6vhN5d/RSVLuz0xuMWAYh6S9URYT1lCWl7Ll9kgiAFU9iE/EvM3+tMzPMej81VAC4
0rNYbXjB/tKEqFYnS5+Y7mNED1GwCm8v73tTY09xwLm7/JAL4IKE4klaAxjTjZkh2oXihDpUnX0s
29nat/ddnIJPIen+ASlvyUyXgZkB+HxhL3WxesFxIRoJEyerKGI9ieTRO1qmHw9QDIgtcHVXUMyD
JFa3WiOa/bmtkSGd76OCXqrXSAulDGLMvHhN30uTuscCYFKMhlnjJBj6g1rHgzWN2z/SS7BbMA0v
enXzS55Zk2DPMiywJdhBoWeU6pFlGk7PYKApO+Kd39qhp48JprsvmC7dLYBPhBRlWBizrqDWVmhR
VGkzA7LH1HH1l563NNSwaic3dBtoyq54qjWzhD2Zy+Q7StN757tduFI7u/TFh1kmCEsJ5gPkh3iu
9VYuLMVRzhdjAszP92FpM/72ccdiWVjMyGbadaXOTR6YbdewOgU6zGke1SiJOx3gtLVo8gxKMOB3
sLFh1bpVHrX61chs0QKBhoabXSGbIG+tMnq1L2hd7BfxBwvjC+wraGLQlFUPYrc0Tz4oRuxI4kjf
SETOXKAA56YW0OFM3G40torlUSEUjQ/9vzmzSR6f2DgOtN4ycOVk0++VGCfGw+fkQrpu/QFlf+E0
M4T/jl4xYR2898dAADMrSCDcYhLJwnX1gpnKnaEEZt5cKqS5GvCXU0EfgmH35yMkRRPBEIuCmnzU
Ip7yW08FsysqX59VoyCUyijItVVzHx/YjVvTFJZbsO3xAf0wOLmr9S7dzMH6QPKBbK44i3n9yZXA
atGQSnonyuAltDMsIb8Qa8bpu1+05WFJYArNbKrVOfG02OYS4nv9TO/MV5Y7r/Ef8/jBlO4hyS++
7owoVS//OTvI2xZnVJ5YoU9ep8qyxTfkaaT1EZ3Kp0vAWtX1XZHASbeD2FyxAiUpgsiNQ4c46bp7
XQF4r3Ib5WaHrLd/YjDv0VLGhYjBwFGlCe4d1/ZgVi9/pKj9BjW+ScBWSYg4r4w5EhKyyjblaHR+
MfdyGls3yj4KQsccedFbtRXdm1MlxhX25mczTS1yPsNK1mmnNpbkQPlNKCZMR2lYG2fbSJ668L34
xOF6mmj1h2a9zJblG2W8Ew2t/YEaPcTcollXruOSxHKQeFamivbZMo8dnLUhM99IYrICB7B9pPVl
8b7k2Qjya+/tysQ8vTwGZHiVBTtnbYzDW8lEWYq1tO2pUxp/KYN5nYLaqWyH0h7L6EOZ2epaSH9P
uKWVf3mQRaViSV+8NhfLBlNd60jvkMRFb83yPwvOO3raPQpXzw4069Ej+/LGj08+O7FYk+7jJ9Jq
UW9kGgwu0me8whuoicst/SULBHwDBm5u26VBlVD5axBZ92A5ug3hZAgQsYg4MxWQ456B8+5s5p77
+LLCZ4+yJHirz6eM5nyGmGPwof6jWcpbio0xdxWZ3mmDlFuPx7400KHld5mSyWMwKQ5YIrlKKg+e
HXFRXSH1XnSNiNB/f85zXBoAX+Mvea4KE+dmK0U2oFbO7DMvvfMYm2Wcl2XCBMhgeVavPPMqXxs2
7RZ29Qu71awvZ5wU1VDBFBenSMh681ZNKamoUI2Y2qtjMvA0QA+MUwzj+ETQx0Dj2o5bKbRTgCqV
T/PNiresfwL85O0lMCMGvaR/dcDBfyQbMII3Sx8eKtdGrwYNNAOD9hLFiV6Jn3jiA13xFxG5GWvP
FhkxAypfV6Sej8Q964ezeBB6fGZHgLKL6GGJ2a6klgWUUEXkLZLrtimjgxR6/Fu9dg7Qz4JiuHMI
0ZtWEtZoSRH9I8BGbbwB0fkMmX3p3SMAqQ2/s9/GQzgodtI5+Eu2+d5M4kraXXBvm6I3fsp8coyy
hWvbfHpQfeSl42HMU2m16zlqBTZUctiGJ937sGz1JcRD+kHR5x16E8zuOVbegy5s91uuafL13+2P
VABRv7+Xuv6agGoQ0MFXir76OtIJDfBoD7p96gJ67gM0FerZ9lEZVDpikIXFKkcFxmJDZzH4j/4B
oS9lZFTg3FS9OKHOx2PT+OfRFEv3s92a7fsmrB2Du975s5DuuA1AEXRXljyi3uclCiP2fHoPtZK0
uxTuxPcDzMS+/3neENgxsfSYDP7NlYtdiLgqd3q5IytAFULVCjQQtpFQr9ZyGlfmZNv4Kafh5mF1
gB+ro+qi2/Ffh2U9lAjqUMbQngkv8exR2vIgyTyxV9nNc/EWSInr3MtYTgNyH50lKt3l5SOZrXGK
A6j9U2pOvVoxWOtcjAVMcrTt/QObrzTxC0smflxJ1r4VSpz+vNSxZAmRKygUSUXW32DvswooiRCx
7r3pyHAea6/fyldi/1fBjAQlw3AXbPoXgvntwxI0019AfwzxLwIbkHZOB7lqu6CytTc4uJGozYuV
gf3lR2ZGWOHPH0K7TIb3negp5oExOlyXx4KepOKZ8KQadcv8I4RdhL3S9fazdUDBIAV9W8/xSiyM
4+h4LtC72xWhvB6gsVdcx8TRmA1kGjRy2Q90c1p0iUMzDaoU1SjiFEBx7MRXbwHhlLXhT/exc611
M9r6zkN+giOww0mDYaNeKxEkBtACFzpkJhtF2BAKXmg6xGc6rXp2BO3h/2vbNFqtCqOYfzVP327y
3vpd+e5+vLHzozpnvg2dtktUcoIaU4DZpCuPmAcF39s8S4RYFlyS0YteRhFy/MemFCV+/kesKd0j
aJRVvvFQJYBrLMwOFTzB4f4CvPtNAVU43PQgddGj4HmCJDye+Bdue8rlEkblbkHa0AztuzZLob5s
9mc1T9izZxsrLccR5Ea26BHoMn/sKxG/0Yblz+G0vf4RGyfUa8o5Ikc9ktcoS3RK2l8tQTd9HAsv
RcBZ1brOQToiUuuLvWLQGjZ0Aa+YYlnOuTJZxpwrvxo7/PCWgXgPtPAAKyHDA0dRw6RtjcXE/Ary
reNiaDb66FbD1NIZAWYWICvd3bry+nT93cj+HKuFsKPEE7YoxQqVVgi3kqWFa2HAnz3S2sIKDpi1
3J6zsf6eKY2flu15gENF7cBybMIPS2/TNATV+UAnoRsIIPdrlQsdg3BDuyyCqbl+wp3sCtDtMtjL
4tE39DJwX+gJlfwcfizAoWjPgfB1vviymKVOU8osWq8nJ0YpUG2r/+p9Wxbl8ZwNa4xxIp1eHhJf
sQkpcwDn5gn3o8xtAH7j0OA7HKjbhtROu7aNY3/q0nIGNC9yzSjI0l1nEFTq/HbRCPRYm8RUKBQO
Mt5SdMV3P6bBapUg77CHJ9y7C2AkpCWiy/R4s/TbsWD4jlbX3e19Yzc5jv2HSgfxhuFtcEVbZ4yg
rJWvVFXih1hMURKgcjrg6MxnJP15MJtkqPL++ZEicuFPFHWIHi60F4w0M+k/TRpSxXHYSnoXO1es
FUm2sdx2tyKV61/kmwN1F40VvI0gRshv2SXK6JPo2USB0v3zAkrpan0mLTKIaqpa8WSDkzEsqyua
9zXPtyvbhbWHmSOjNUqnWBmcWgLr5cgHD1Ks8G/Bxx50JaGtsxIXBgpysI6zTd2M3AAFmGk8nC4H
lAXZjBFmYmQuYWRTdMMfFCiQnXqPrZNnW5TJf9rp4wVOdpzOdcmb04TWTN9N+Ebk7zn68iZpNB/4
XPKOPvARLNIHhRfqWeNAH+n+t8cJN2gqUJ35T9Sx4q3WSjVYz5m8s+LgDymsDqzndJVRIXgqa7To
pskNjH0lNXE6FHjLNk8X+nK36RLdY7V5AU8/ICY+wHpM1vomX4XL6owfL4qevQDQHoBLP1bUj1MB
+eDqOkSrNe14GuxoZxrehqvmbufWLizryqQfwVN4SPlowcgJccQD8TqugvMWORAu0PPNSmn4QVRy
9Krt6v0tkQUSwbdeS0vs60ByzT0CYCfOCtafgv9e1Tl3W8b/RO3p71HJfJS39u7XdOWkwt+16zSx
REuBy93X7V/mD+qT99GulWrhNLh4tURb6ReP00uWKdpLnda9Yvuzu2G4vH7I3nTc3YlEmrBqQtN9
PRk0ZvMgPYGWmhNhl2SGSaaBbRNGgxBczED29o1vbjp21SzlqXXTP90QxsZw9ZzrB9JG9+joymFJ
5v1fGc2jTNN8XZ7ER9MNYRKUG4pCls0N9EDNUkgb4390fFQ9GU9tQnu4kldtNOJtZlNbqj1xgNti
4tbe///rqeOLUCCNvXfH5g15+iL2t70bfeRkOwrGCTR691Z5N3TDHjqSkM0eBhdAWHmzRFppx/hi
HCCjghjtRWYgn/NxL9Mr+YuA7oDZ6q72DlvPfXKp975CIm1QpGDHWS/AYxLB39JP7g3+DwaqtTyR
4D53DR880rZ/jYyl2XKCe1cyo1q6BVYnuFKvdD0pxllujK1WW4wxub4VU3m3fKKfQaTA215m3Mv2
5nbFFkeyRAkg2SP/h/8+n3GdNnsaApYhgjH8xfhLoL8NwoLbx3s/6cQBpLgoGViJLoYnEjRKZzkc
7D+nO/Vc6lnqTvHo8Y1JK0sEYICommskLW7z7pi4+1crKLV4JHj635Zt88vKy8h0V3hfjbY5lVMn
26u9N0aOuQ5FpaIGZMBvYUCQ+loCs9rc/7inAJV1oj+qSLriMvUkJlkp4fdsCxMK90c7sT96Mv8U
t2ah1ZfWsLyMEGZIfrb6zF1neKkhy2w1DiVWWD4TF2hhbR7GiigdIFu5faIpuOe09QZWqJ4SScwG
gFjqShybg6ciNkd3TNSsfe4VPrRLgaGDCRE/4bnt8Z8/bP4H1rk6w2M17LedvmqDwjuZSndsUMbv
LNyJXsTNTOYeVZoUvRjZ0mcMqn+tPBFVV5HOF3DALENsGa7JvMtvBjlrRDBM44FqS4cxleklbcWX
Pm77Wa7N3UReowHo+QRZdj4JchKSniAGBws02RmEPgzul6F2+5P0YmLyizWtN5NihbEMmQ1mslt2
IXGmM+bWRbMLCtxxMr3/Y5THPvg2sBhOOrakYBcb3APZocUdV34BYSdhKGcQIMM2AYWyFcWGxLWb
XQAWlxndmD+dhRrUsg0CvDqROgg/CuPFecOzIIOj+9Wn5RjOnbfuLjRjE8tp2DzO1rHd3eMFwEWa
dqWG3T2Imm2pwrFZF60DIQHqeObLGJVA1VxwQn0WHDogBf+Dx8OlF9r3GuWLDwOO/YtICIOdj2Uh
OZ5eHfSzLdrr+GGr3fh4yf6TV5/aNYRWEMX+Rx5n8wTQZBylWxMbxOK9XXllIz/aSJ6t9j/cHJ+h
gU3CnQyyiZpWT4HHKQz7p8FIUyf1QmwU7PV7dcAm00peDargGsdzuic4Ny/RSJUs0lgSQFjVJ/TN
dJeH6JCqzidWaEcYt/OMFFADZrihG3mArZWEfVaZDfvvxYkdTb1wQ0tKkhIdkp0IHKjLPuUBeKPU
0kiPLtsBG6vDA2faiLksRy3rDz9+s2UwIfNwKpBIOP/mZ6X9lcdxg8GXkoQcfYvpRCkTkl9251Ne
nZLG34iQVb2m8H7peEdOQyejFDQOGeiboRadXGzkai46JClKs49Bcy3LQ4PdUii69jCqpbZLZDVm
Hiz2WYo5TZ6qoRTUOGEZh046rJPcDF0gNMNkv+9l2CC+o+3rNKXE9obX88jQsI6zcStLc3oZpYra
OmsjdrUqaqXWKM+bt6xutMEI12Aehcb/TZRzUvCMXIhDvFOFjhDYikKd0gWUUO9LcEVO3us7hVpK
+eHP3WroU5g3Mk/hsYECOE9C2dasxXar6g58KXiFOSnwmlaytjSr0qDL962QzBjAQlcJZ9Jrswuo
xoFTG/P9pgh+LkEMH8eUWT2L7lteN1ZTl/oUhY3VdIv5D1aFEVmwuoaIkZsDP7MwFIfvgp2WkHpy
k7OOYcMN4G7E3C3S9rPe76rctRu04Ckyg8e6sn0Y6i98bgzP8+CTtTbCQ/TuIuJqXoGm74eioeVD
yQw+U4FVSkjIIz3T0UuUE0DoIX/VDB0Eo06XY6Oo4AgmBFcKyCzCjgf30GeI2BIy4NcK45rSAy7m
tpJywed3ToEArP8sBr4waj3Iq770nkGLDAXneRjDUp14v6qbrOgcmOZGh8ftWLOTdOY+lSCFXdIq
vBpCDssE+wJv40eXbMUXlhc0JwIKttf4Oekdm/SBAzVmJJynhzxoudaOAFM/U8jN7WqI2KgWLKNa
SNXaqcaQPBsIBuY/M2Ft2Xhs22mRHFEA/ovqq16mXGwCWN9+Zhq2rXr3bQ9xG1j917KWykMPGpAc
6ulICvdVD2LYx+r76XUM/xH0EUL9/8YjVllJ4++WWdTjlUbMJlwjMEq7g87LNADPNfU5Q+MKzy0K
bJnrLQYHzX1CGfNRooLfv4olEmmXoc63MPo9uY+as8kd8Ie5GBREQt2AfieZVqBI2SnqNEHkWsOT
btCZiD5/zzdf+ZnQ/QPL8ETOZwZn2uHMqECt/UU0WdyEL7qhkZ5M1kNYklLxErxCfqp1kzqlzcsr
cs8ww8xdyhpkFLwImZdQ35Kwel3kfZF5cJB1V3Fk5pBpxVGcObG3RSwP96H+mUVSPTSwLKF6eHYK
f/+uKssDUTAyw/0u3PJwOLq2KiYncFaijsYgSm/wi40qrTX+4JwZU4H+UaSYiIQoUJas3QRisZ2b
I81l1wgDFa8CRWOzjzP64XAYoJB9w6VgHfqnI7l51irmJNccWV1cOz4ooST90P83PbI+d7v2urj8
5hQMimydLjiJNgyqVqnFIAHYQLep05ce3RRPVNd4G4Gig7dlzD4k8FzVFSb08T9EnxszaSCirYM5
pTIt+c82O9NNvQMxFGrTaBLBeAVzREadvjuogk1UncIpYkR77s6CSw3oj0WiM06uNpuMEFtnEO6J
/wFETou48Hcr9fFQd7kOJ4fizS84vrOxR1BlNKYqVsDQM6K5vvr5Un22uAyqX+ALuoLlGExj4uFb
vt8VLuCD1nA5EOpBJ9KpPu3n3oe0KEBA3z6h71Yd12apZdTpOGASDgvf1RPpoc0Z0iGNnyZHnsj2
pb8QGcPZh/7qKe8THq7vCyA5oHLzZc8gTJBAPz1LYg/LeCfi03L8lLcvylyUZkOKsrIMZYw/J/r5
pR0UlFVbEx/8xgJeZHbAzKHpE0F0hlcgOlPyuC5Rm8uKonj2Fg04aQ8irAHMPWUMnSQ+cV9VlYEp
LmZlbFNqSWaT0C4EmV6aLiW1SMtjIgNMUDQcipZxXGdIrwUuUIuA/dFZdDkv1pcbN9C/Exep1xW+
gfHGeJS9MmaZDB6YNsuD9K9+sI6d6AYRgsfvdDRdOeU3bnEcKJHs5MDqysYBi4diobjjIhqSzGQq
YD2m5HKqdaeIY8Qc4H3VEWrTQPss0ETehwcGm94ZPYxe4qQlzdDht0EFeJmjQrpgt/IhoFMisx0g
c/MsWOWyNf/9glP28JtaUJWWa4JB3TFayqnFhr/bhzCMoDIkUEBB9x2MrENrYbbsxVGPDtJr8j4R
wlXAr05WRy+jnHHi725nGE46m9QEP+rqP8Wf+Cs5fnIwc11hISW6SaAhU9y+9fWQTpzAe3ozy4my
+vEYZYgLUf+IMvlRm1bx8+LN0jz7sMKbXeOiZGJP3s9t5uObKtB9UO5oRTOtv3MNRvRzQ3kYQDoA
pR98sQW7jAOqbmEwtGyEFmUSEeC/BmkuGv89AQEhDLfI/R6evMPPBfFAH47ELc0+bOX40CZ0F3Eg
oNPznVFaSAN6JvUSbxKEjQqDMf8eEDZbwQKubCZCmAL45Hr9UqRIew0qSwiDsIV8CQvlA1ou0TAs
9fQuVkttDkzpHzLnXCH3a0K+s8jpKZ7hSSBc/3WbDSDqYlsXiDhZlzLtcxv2q+/CGyYELjx2wCB3
ARmo91nUnd8m49ZbSIf+iA0ycGx5CywHTyhS/y6mzt0sUmhzHJD3neqbnBB3YQj8gkeihrynNYBm
jK3RapWi04/lzc01VNlFjLmapVQXJc3EdwMSHRsjOn26eDe+cp82eULlJZpbEMlWODisIzH1awUz
ZtsZn2tOoSLSe3pBh0p7UlskvlaRxbI/DW25JXxlqKDJMjnD6hbIE3cohuQW2DO8DMUHa8i0ZwyW
mZ2160Rp4WcSM/sJ8IkarpNr42dV5WryR6hVBSQS4e7M9IsiVasgJmEIj6l8+y1epKsl8JoJzPD1
AQks5Ndpz+hb3brpdxaG1ENOWCHXTZWiF++f8EFNfDc0/9ybPP4euMXhgnCP2f9XAtxW7TdXZjiC
t6FTH6mtugT78tPJJEXotCTgq0bLIfmTMEhFyZTNkzSfXhpY87EfkqR2T/qiwWd2pUwBa+1cZF0h
MpRqrPxU2fcyk5b9LW4ax0OnRNR+h/lFdmHOYEsIqn91+7jNXpvJZNwstoUHbYz5hjLGt1tYgkRa
homLp+tNvFCsH6QP2J58MX03Dk9Xq1sd163R64aaK8qMSs03N856IE+O3996/3lzKEkuQYLzAeLF
VBHzxuz++GZbzqE9Tm9wOrxajRKUyRR/6iYh9KD84WT2jq/5kXaZhVPOtRYjkYAd3p5smr4i/a7t
lhuecaHhmwhExxcZhra6XlmuqXSs5MrIODEdAQ/jPe2SVyAUAYdDfqkmJ4hnfwxkBhe6/vl6osQP
aFOmI7xmrWbUMD2NeLPeBNAoXLsSXvfHSTvUqcCoLdyNAIRUf5gM7RQxEpyCD9GO/79yMBWqvBeE
+DbF52AT0SYQlXOVPgllkUHUctQ4rjeja/J78LVVmsYcpKTZ/mB3UdOlmGX9XjUnnHn7LOzyc+Tc
54eiB1MY8/d+2nQrKHBWxIE/1MVxqhccguYBOZ4O62jRMk3cmI8A5QgnvETLhQb+zOc5NDXUtvrI
qmqmd8vsTEz1+c7Dwk9QhZUcATJfj9mDVKaFD6ubKd7W5BHQrWy1A60mAHd52iDSQkDwRXUgNUlb
NWoPOUcq2L266SZY9lqbS0IeDdOS17feDNeuoEmS1dRksTVosZ8OKiNF8yKSz9+SBr8UHzAePJov
ovBmQxguP6Z+W12qSobWjBiP9CMmtm3ZfJ9/UG1XXKoJVqVfu1syaIt3h6SiGpVc1QD7uO7MRr8b
e67rGnAOaI9jD7uIuObvagTOg5FLWx6ftvY83TBTyte0eJJC3DfErVAIe4lf6Kt+Re+lK8GRPgXQ
mBvAsZt++tX634iCy/LefXZWEkNt5AY9iGVUOaI8A3ARSC7MvV3+xzqB/SLE7HTUvw2qhC3eAQpt
A0tcc+4SiB64OWLCVGEA1QTilIm+yiCEX18GcQi0tAzsCLOjJ8K5r1dbhyuq/sQdhszr1Y0SN5S1
pSK52WlkxBRHtHrin/xnNo2i1wZHXcjc4CgaKuiO75sTip8NzJcy/4oTeffuOBbA1aAC+j/kKfoR
lvFhrE9udXKga4V3PPu8vzJhJ7yPorfpuldCmWcpFXMfEQ+qSTeo0CNLKunzdZ54toCoVGgxPxdZ
JF2n/GaG95KHxyQGEJmRTVbFYWx0PScPgDUzuXbLgKD/6kDZxncBzZm5qVKICRRL419PZYG/73TN
zF5unov2wVe5KyB6Cd7puCxOwRWHVWOT/k6GOR7c5jjlklFmPnAicmILQryq7ap9GqlM+0q8Dnqz
Q4gobVJ0buIQRVCnaqJuEX+L9UNnYl943F0q23RgBgvKX9XoxQ5Ln165ZbjFi2+o5G+zQyMYZR9V
ZNfkh5dbdvdXm0iSW0mgB8DVCX7NkzrpMZ1ZGJpzMsYTgnMqzumhkRGOrdkFgb8H+RzrZAOUVzk+
oU9CL3gUisGGz3DSEWHdOo2XfBy5xbqUmmGgeoHxQiUsMPhvir6HuAT6XSshXY/gf9TGs5Hk+Vxc
He/r+Gdskm9jombPrsRL2PWyC/HAkyaVvAOvq0T2+51LX5P8m/Am2Uqdo4o9u7TS9QP2GHFjudz2
8GJgRIztc+eWupy/fXOu33DN71LIGl/F1IBxi102mIlvv/oYbdYUgPd69soPVgftmjl710hDcJ1K
KfgSbiEkqBvBj9xVhUHFjYqxYuJypVw7xLcGMApuCXMbFTW2DoyuvBJIwC/p7Z7QXJoihsJCMt11
9aJ3ePIPhxUrDri0zxP1U1AjidIvGBg5GhQ4tFCClwrCPMW6auPXO1MLiuTZVNd2WSIir+RjHi9S
+aQ5c2vUMCoRJJ0UOvzxHnKdT21SVZkbpyfVwF0Mw3kRgM0Y0CWu57GKiyzHwmUpYBkAD7cbBnVb
MifMk6WdemYNtZdbsdlMWRmghIl1XbWK6nivCWQXsjfnHsoNxEvTjkWMJQSJuYir8MhghKhg51He
d0PcyBvGwArSuL5QcCi9lT8jSnoL2Ryu1tfHPcDZfj5vYbQfGCuM9wgcP0LIBPhkdJaWHT9UZ/As
AAWz1qDNLfhGiQ6yt0THZ8clUqVZK1R069fjnFPj0Ad3/2KnsccLeN2ej9uEY2SCYu4XTAJy+PKv
BAw9drG1IW032HJhDuBvPUkg51zBOjg4oBmwpve0Wv4GDTJQi7nbeKWo1ciAnft/FHDkoTEHsDhX
OddpF0lkhV01SRYTOiGWCvijpk80zz1V435b9a+kclBAHmUU/+F+uKReRPwVRWu3Xnh14P6nOKot
QKpR1SeDDJWzVdYQVadOjP6utaYGe3xPZFKd7XzjJtoFnmxwdGf3E3cLLHgzi8n9wdrMsp9yDru0
k9SKlzZuEimHelAL6GyWRMlhkQLFH5H2rDGfgzSe0Ff26wvpOwK9+mH0OiXBpRvO6WirW/7RXCU4
V/EB3SZp7CiLa0NjkeX0M9IXSdg+Jlyk7yb82fV7rNHIxA0ZD7tIeUlRIkRmrWlcp194V+L0g1T0
qkEXcNN2dFs5FZrLlYE+yH6H3UqQROWabxGy+qHMTl1cfGRMr7b9DUCerV2957+hyOPXWgbinbs5
zqSs3g4HZu5XMA7bnThPUF3B3zCgZBWfkyXnGh8YFsB9vEq9/3iqIv/qVoJak/y4iQZoTvXX3LP4
x31QyyLLBRlMdX2+lgXimh9gYREE9jc8ZkQZhD4utzlphUgtHV99qu4CQihb1mJSLHD/ClMnegCb
Pz9YLNcKZ00C2c1jSFGHqTkFN/OA/DItpG+jS49zC/cISmO1TCu3hKo0hf792opYBSistqM8Cimx
0tPpwFAyra/DmeABMKtkXVhLohayzpx4HyrjbTdm6qXTxaZJA6Y0f20p0+Qa+P8S+TO0Q88qiXtq
I/II9cOKrrs7ZfP7/RBYxH+yc2urCz4G/3cZ6vxqLwXCBedaqO9iZcv8v0h7M0rYRHFp7tWwVJaw
kgwiJ18pLt+mTrG3yDUBSo6PCB/JCoCCjk+6RV85VChvWDbuBNS79T1PjJ+oRiUArYFjHmcabhdJ
ChyzYmtnBTKpIJ/E/UldU3Lj0crtUrf5jSY8YgtXcB45uUuow9wlL2e2Zv36wNh4bDyipYW7pvXl
my3P+DgAtgaySmGW8arAqQd00Nd5NQOPKWItSdv7F17h0Pf69VipBFuHBespgbArA5WYBAmQi/ae
9MtNAGxrttzYK5VuNQBTeDAyiXanF1BlYY9F8+3h08wdodmXsU2ZMhZx0q/pnjBHzUnPFRFtfj3u
DqzklRhCvwZvgv0RsDbmSvK5q4N2xbwCdOKIY6mx709FsC1TaAcPSSi/MQi/ktURpdWeaKmKrp5r
Wq/NdVVrQu0bZLSOIODK35XpBqwoLb6a3octTH6wvkJPpcluh5BylLukWDr5IcMoTAGSPQUDpUFo
3BsPtT2ssPQ6elltimV4ljJmLAWgmUVzZM87TuQAzz/sjMkjBwbxmv0ZmUllk5BRce4/0YE9UFL0
rHH+C6sG14G4fQQ+jlZeXKiwRNbNcI1PzuOTUiVf50ht3DjiK47oSw4giHpdWGlMeY0gsEvoeycJ
UAdta/Th9OvzIpD7GBcD4xbpucfRoW1zKF6dSqqxASckJLo3awpVolucpg0ms0IpAHUiK8UNwh/S
8kUaCcizDxv4FnMgeEahpo8lahQWtz9f2RKBJN7OCOj8nwKX+XixJ4IFiMFnOjb5C+DMnYszmaHi
O/2ih6C360TztgFA2donxqh5jEaVbbAOHdui56BT/8TBkbyGab8k0ncJO6dP00wam/ImOmayw9lD
co1phRaHLDTnrpq7jBcWyFciWZ59EHGCLvo5grnvmAPMjhhH/T8b2UHHD/M4QpWi8gxSLumLxTxO
KVnQwoqFLG8uiLT/rvqL6VFtICKbmZugsLJ35ZuS0xCeH37Of4/5RuTCuhnSGRXsPXlwBuDdDhCd
gPNIWMlA4Ffee7R1NlJw8kzVH+Sdweugl+QUVPXzTT7I0JSixU4EdSz3clcgkswZa0BLszwZKlXn
fWWTe3v9dIoCL8SDlbpKNlfukO+BRNMSt+5zgcKC/GfLZdSWUP0stpK7Hv9ak8rbBLZdvi7GFZaw
Ve0nUOwBWD9sCFLT3cJgjZTW8u+CPh+H35+hiTb0Lv0imOAYAKTWFKdS17EaXfDMa3YUylFrc1PR
uc7cXns3Wdpgwx1d8GDOJy4KRHDXOt/fbJx2giCrdT9BAXWlt6DlCsXCDPsg9ifME0vQBFkZaMA9
tBchUbj+NWk8TR2uxCiUbhB9ajF4oJ/AtkXf9yuHpgWzrJgVOCLUpLCx+SaJ0tCxu5eNKOIAByAa
KNS44ArPREw8XmGMv2Jgx+73IqkApL0cLQFelQkI6eDgY7p4juYKr9VTlWD0lLzXUOsuzLthlraD
lT65gUsIftmGATKIOpnou3I5FrRvO3i/QKm9/IkjVh/v+4GkLcvcioPS9J4AhOEYpNEInY0brlJg
odwwfTIOg0P8dkdTwAMRlYE8GaDUb2F5fBtoPlLkqS5l45Bnns8uOdVADSu5BLdqWcu5i+nXvxHS
wozAuUggOIiBZ9cm7N7kBJWpOo0WOO6iNMzovht33W9KJ/Nzbr5Uha5jdHZrN7l5XXSXRrfJH8v9
vti4D0guPgt6F2jlXgej2Ovz/JkKBBqhl9JRj/XyOAygV8MEO0c3xzRvjW3K61oQZ4yN+6uGqAZU
bU8NM7oYj0gjX9smiyyfz8bs9Kys74fZRh8T6TyFWZqHWeA6Popuoae6JOMUUvyuH+HiwQABUzHd
Gbf1yIiAjE2SDyeYibL6Hp6y6MnHAYtWCCwyR1BhPWgUNzTIH2Tvk017qpqNrSIByBZ/VzPvGWEe
N3OZlS84HgcotwZg5JzISZ/OTHlp15l7nGQdQU5zCc+0VA5g/o7IqtqH4ysLrKyfqCwa8XKGOIbd
1iwbpPYRctefxm3USpI/KLsueVsI1brUpa39uDy0JJT7MO7liHDWcm74kUo4mG7LGtm4FlqQ4xp9
gfLzxUS0BDg/W9RDBG6KwKOgileAi1jTyULuh0+negqfex+ZthNihE6o/FDNsOFBVZCGKTXcVB1b
UgN3kQS0J8W2aqTK9nKxSD6Fwt/bM4Q9l0hs48mhqxW9rQj+uhNKvBSgayVpx2XLV+exYkstFp1n
6NorJ0Rn6STrpTK++HWtsSMEA6Hrw2HZGkZya/syzCjUk/2WFAq5SpFmCs7o9LLTo+BuFJp5c6SN
Rsvocid/GuydrADLwGePk93a3JnG/DyDr0GrZBplmpz/PQhVPBCg5EcRHBO9K7kAr5tggcv2wmyn
uJIbiXrrKLup5Y8LYuEsRz+mYmU/gN3JGc3ZFeVlyhqaRaAu/dm6BueGDE6bBxJUbmH6w6M53xSK
z8uvkwDqCTy+mYUJuxTsN/fF1R3vbkH6mgSCb3LKX5+R5qXhR5j6xTe8JTmJMEploomjwlXD0m4V
6OkD6Tq22CoLAJVpQemnFendS2H/XavFQ/0zGwOaduLKZ5AGkP8JB91z/Zc56GWQwhrzS8G/1AmG
Q1fDt7b7yMI/jCxURlPp1UOEV2z6zTg0K6UHT133LbK5Jf6s0DrhpUiC91rhNF1mUZkbS3fYOskt
cGbGN0bpk9JyhbAeTLrK37Uuga3loGdjzd33+iOFPAYwNNbgBBi8wHUJENCNEXeXTn1EBmaI/2rz
xHrHwapZP6qwMJ4YQa5+y/ukrI6brw4XHhqgAeuGLDyYhc2EcDVe2Q6nFe5bPEfmM+P0bhsXN+ik
4Yd+2+u+s0Rp79sIZHm0KNnvBc1llsFJAbAFi/oVzq3xPl8OsGdstoyT7OL+GaPR0QpzRgLELDWq
qs6exGKUR3UAzX/DSjwkhooJstpNI696pFmmh1ryk1ki124t/o9VQEuxN6QNaQ+B8GcEQt+a0DCm
qyO4qKtw8cWi5cn/mPlOyuVWpWTN9gebABcHtSJ4Sn0RElJnmQjZZouaW7zzW3C5gxOyiP/8aMwH
Qw2JdZTRn3BeyyMHL/Fxk4RKeW5tDGlGH7k28U3dZrwaaq3yS1EUdKrTrt8zS2tgFtJbO8Mx+kU9
qztSwPKVAhNMFKCh/fAlwtqa5OiEEkr1BBl6TuM9lFouHCvNyyorBolPbQGoGlr+WFjj1wzdIKub
8yrwxMrWg2esuLtzCWzFwoO3QdQCW/jDXBAkq3tHDWptZ7PxKGg9y7tvo4swVWje0sb7Ci2IAglt
m2jU0rs8lUEh4odan+wIRpxIwxDuIW13uFQmf4niVbkCuFRog7/TSyedJ0Q5TGyhLmHiVvLDwjdW
dWdqH+kIc8fueSuhCu6HTCUxfLBaj8s1hzHY6rPq70IzgvGMtDrvLNHMcfAMNGnr74OQLWvY8MKk
/0ZBYCDbhyZsIWXchAdpAinSCvcoRgq0aoNGP/wEECcbhEiqIeKn8fcRpbAbpILwqD8CvSpfjo3L
Q/dqlaQh/YbrNv2a1YmwwEws4v3FJTm6TvAv6ExIzjxYw2Py6RDZSZEHyCwM4H/us5iewGS9N8rQ
wlUYqdCrzBUnNjFHoTlcNMAzjshJSJlawmidXmUK3iZrAddSe6aMVb6Mtw7xjWUMXI7+pi8dfgCk
f8H3Jq4cfj+8oVWFC7BNIO96G9QaMvk3Fq2sCq9XitUGcEKTGcKjK4Q3/aGxKR7jeR//kiKAPwZk
gsoT881VxeE2d1oGwvDyDt/okMguusCOSyMqQYHKqSFCqFwwuk2mnc0czRZtXDQZd7zqnQSTMHJh
aoaO0YVVcc0bafD/QnrdFhOd4RNukUtzVXWUH556JQfJhTH6Q2zgeVGvMJdvK6hI6VnIQwGF8UKO
oPvfzNMFLq6QSrmbTBg1vvvHV07+anmcUhWXoGI/UiqY76id5XLN9DvnpHKt5sgjkxrsfbKlhndj
4lDcYtIcNS92EG1tTuS2aHQ7Lpn9x7oftTU+0i6yB6IQFD6AxaVuLaDxHXDmaGVN4fnKeAwISg8z
2c4iiiBh2Sz5SwntCJAiynpSGSgDsQHoDEgVGCXJVIiTwGIjWBAqS6V0tPSaEXuxcgdNtgEHO17N
AfJ4Y0UQ+83oX6gObQmRlVL/zWOXfe871gnMDEXoavdyvPzi7jz4d680/TaOwKAdzQ6jG+fbwL59
6dXz+zqHXAT1d3ONKzd5uUikALeeQTpULF/wpnKCCB7FebT+lhQuI9AvapfdLpn64DDuAvd6s0M9
FZtnAVAQliCM1MOXCRWZc0XbfokF/9UqpKuTcQtCe9PoocIpwRW5bxa0/pBaNVQg5FcwVJ6G5g4P
F1JgBlpGrOqyxQMrovRxFpwCIEo6UnkDE4ExF4sDOh9bJiQ+QccMyuID/uRh4CHSQm7S0Z+Gi0rY
sXVreA51LqUmuyXFI7oHAZIGlXxdX0/H/9PnyO0I3xEHFfJQ6qC+8arCV/aYHYzY10rqVarekFjs
9P+GVVGiOlGWgZjhzfffXLKUU1QWyp5Qoan+5wQfsHO9OSSJV6zZC62IykBqW4ysQLrl2/EgRil5
0fglzFwDrvohEpPVle92jf7FwPmBvqgmpTEfBzVglG0mh/5CSvNMz8oWZwHqETeILvG5uXRxjtL0
kM6mHdFnfk4j61xNLLWK2hpxl81r4e0YdW6JwCnxUJuEvTJMC9tMCodUYfu62TrA56L4Lkwf5ZjZ
D7P6HQ8It195RhxiHkp+wwhI3d0L6pHNqMsoeU91fPn9DIRT4PkXZwsQqC0VRFxQIetqFpfUM3oN
LFMXLT+ZLu30FQjH6zWqFk0GeIFTEmHaQmgNnLo+g3keNRzFZUccCKagfo8uin0m2ePNqKJXc8+S
XJcDlgrFrx2tPFziSS4W8v/EsmWh2ymuDB/imbCUu6TkMT0g6HI54g3e8fgya92ubykVt0UxJIdz
UGh8M2zbOhthUpg1qXHfhj6xBu4SqwePyLRWLAcCXpED0wom4MdL0/LQzN6aeOehKJBfP//oaZB2
h6uP1WnLiv634ftm12up/V7pARZk1ocgl2I/4cgHU/w/kBcvO0rL7ULVd0/L9JEAT7LYJYyJsdfw
nv2y6tOa2ZWQMFMnKSI/9LN60JnZ9pLkbuzZcrbMDIXsvpAxP6WYw2a600YhO4oEa8kotlQGhO1K
f5d3F+RzVNeXZuqkyZ14ei0jnJ/vURG7NexiZl8xi54YlxcQYeZw1ZjUsg5IzI/Qb+qrbA/OiMsX
zYaZaL0ecWDH/l8gmWw5Ki0bewEJiU0RwkJSiUEuE/dbjSNgohOVkVG2VjMAeSyx7fQc1GgOGTef
IrOFNDJsx4He1efrrd37nwnjonP48SupHuxZ8tXCHAJ9+G4zmdKXtrmIzQrT768iTVV/4UoXYNce
jJDHa5RtrBA3aTinEDJeLgzn6KWXwSeGASIWbJ214gxSeoimpX44VS98dYiGExdMoXachFJihHGl
eWQbMwdhWscRk1UlHG32ghgyN8NuK0zskOacrxu4ZKWMafX07r8zTBU0Kbd3w8QwRJHbbt9Gj1fa
vnGQ9nyVJFe1zNhaO0SXbN+HeFkq9I5b+VCvSw4Z5+7IWAdlrKzUiJ620ekWu6Dnk7m+FhTtXFaA
UUkMRICqYOyYnbDYVQCxUSJ7ZIc9m4u6l6PzCrp4TkFl0HnanU6JkeW2oWNf1HlZ0gzC6o0yVW0P
fCsv6ot7M7lg1a+8p3nZqbmNeRHFLLgKHEkatW6ya1PMWGKxaYtZLZlBbIO+K86BuSI4qI7uXX55
UH1mzwxQ19MbVMDWIvq8vfqDFTW3eqLzM7jKdP2ysiHrUM0x5zgTHhwslO/7wkYxjpKTyVuU7xmi
s7xMy65sP6fjNHAB4+FcEgafpXINEfN9Vi5VTK/0O3Ew1TnkWqiL3lVhUnyZ3WbNXBmhVv1r5Xo5
GpWYA5MFOv0TucU6gwDupNPn6KecsnTu30Ll7mXCNJYftIM5LH43W2oqfP/2k1YQZRV5Kx7J6li8
q+MSAxAf/gdOic3H5eNB1QavDRGlqzFijVt+2TCDEhM/Dlfc8kW3KEATJgOeavPufXwIGBukH2/O
5YAn6CDzGdlkjOhs1Gubjw/fWV4zBSv0QakNblT5vnD88hxqAmr4eyu44BwdsfFz9ay8jTx0Dui7
1QlYwg34Iwj3b1cl1dhfQB7ohuJO3E1XQSXNyIk1uDuGkVVjACfIrmfc11K3qYpQdn16sa5xm/H/
0T4uufGykGOs/n2VXQgs4EkPdt9h223GEIsumW54qhoLB8hH2XuIZa53i8zP59sFKWA9AsPlQy14
d/VpjIi/y3vy7MY8G60KEgrAvrt7Ld1JpRW43cKLI0gMsP9qk3gxxjQ5jD4aUlJHeOv64Ebn3ctS
JBF/o3SvY5dhsx94qqOSndEdeDrSEWelHlSKChJmGRaUTce1IBxQ676QTeKlTtdXsf+5MVbiiGRq
uMgWH4By8jzMBTNB/kTK04PhOjtD6sEJnZNBs4s0ppWYykr8PqLQ3r+5L3viMLFsbAPMl4c2ieeF
nBQwpV9oRpyU/MJnBqqGY6IO8vWWV9bUmE0EP7ZZGVV+Yi+7QXTDqaJoFWaph2Vc+AiZkQL+WRCc
GGr/VgxSQUgd2iYnlzy0PvAzHMywVugVtsJJXbTCV/NLd/npNIvZFehlY8tSceuFWxvV8UZNGTur
6IcIefGILXUHDP8c4AwpKUfhbwNtLFpkJmXqzIo1gkCJhBqFUAlIvV3JvvfISaZfZTb9ZFd/6AEv
ShZIUN8sy5Rz76EOFGnJHEmLA/eoDezarOsFwqEX67va+AcUMM98/qkwCwpHTHGfJqaUWrj1cCqO
BO1amNWbVSZzWmwaoGiadYlpOId456sc6Sgnq10hE27QCAO1ansYn9E6Z2ry2LSDil06VK3GI/dF
Kn0O/2LIFTNaVFc15Qo+A0D5nUN4HatYlBdWuwg17X31vaOtv6kz8pyrZ9nyefOyV0WJVg9IRH9+
vYXnZhDYxo+ULtSAgVsfzmszR5Z65Bg+6ROkqXtP1z+B5FZ8GtPnODV9bx+4N1Hk2nwHleKdHAoY
USaxlYaf/d+KpXkafzOsNGxlwHWmpyZF5oJyqvX+eXsjIboo3RLb+PS+2vkQVR0VfQcc03Ojgim+
sAfxHskO1QKoyoUcWpMhKRvISCE8e9cEHRLRQMv9N98nQDRtuIb0iS3lRzt4ryoDDHHqvDk03j5a
MLDbGddUL96IajnTC9i12I/wxn4VmRKq+byAHuRLkd35WgvUjGtMR3An8HksgL2DyWp4hZBL53CW
Iz4KgXjz9QIyz9S5ycqFtyr4ePsF/H369bEVgAt2ofl8rNsLFN3H01fKXWFt0lnf+d5cLnJbSmNK
uE+qDnVXCbQzzglYXT1XxLXSY9ZX6vIU1ibtmn6lI7eUAjNjZ0cBi+qs9vmwTqY0Sccd1Kvc5kHg
dJQnGburNzeSZEAESeBOFSIRxQ3C62dpIh6NUfE27tJa+vo3CnXYRoweOxDI2j7++3oFMFTU1jOF
r/PiXyzHyeHyFD4xCmGj9B/c6Y47DVmgZo6D+soq8QdtaF0obe5hm8S2PhG3V+LxZiT4thNSJ26Y
E+mTczK40oOfxX3wXdSUasuurwN+jON1hKdWzkhE2bjNaYtWPm8tZmpfdTSf5ySUTvIhTtbOJoMM
W1y552nC1yb9mElB/KRipFUnJBvvopCsF+SlPgYHF9RZphT+HBs8+wzE/qNZsvT5K+xIKekHEvvG
0dhI9B0Z3PV7MXGMATFq/1pbPVDWRMjsguHnpQq0/wIcdJO0R7sdydiTru3nSNbbRAQ+1n9VMSaA
lxz2z9dmGW62x9nrDl+TnomNYjVsfspmLGx3fjJBRp/uculxP015aJ/rNCpK4ICh9ZthDi4L/H66
ZBnzYqmvtetQg4eudwh/qYYO5AzwuuVMjDa+pwpUlcRCIV7BEI1hYmf2su4HNJ5lEU4eETpiLWSt
512CuhBNNUoB/2Q5YA1vqeiS85EiI6hutnNY5J41KU3xfK9XjNnNeCYJ+2NwGd1YhG6cVqhnh2fo
teqx/0mUDxJjzRI4nVoUsEda7yCqrNLVDlPDny5075REG4l6xNoaAa1ms6+3sYwhvtn1AFcONAx4
W2Xxo2hGaZ+sFudUAuv2Q/PCTYS0Z+naYlhDQ7vztrdoRrn1M3inq5rVyDzw8Dgs9U3tot+4Hlux
DKvQlzSlCMYw1+9hQJTc8BJrPvOr5KNkpxAQAdlSOeCc1rZJM9XGnhAfKOxydfuwHYDgsqjgw6Po
qc5HNWBSL/Qj7QGb7UTnmbPA2gWkDDtOzry8u52unTWNdYNlwQ5RErU5BGHEJEFi3bRrcKnHRhUe
t3Eymnmr+1hSRq6BtPUBQGLfMoQqbDcCsXlw36iLVFAWRAkOsODaOAlIEl3C5c3zflAW7eFITrzm
DeqCbskDiwo/pNNvJlXkOwxKWoKj1fbXmeE1/hZBzduMkOBLJlzgWALvNO4WSVs4bP+ouepioPok
TR6XpUGgs2/Qf2GLAHcKzS5I59DuhnRF6AyZOlTTJxsj0qnGQp/DbjejOIU/edSNuHAmCY87QJa1
qM4r7jxWWYZlFa/Mrqjglc+sa5pDMS54A3/nT0R95X/3XwBkzz+yAK6MNGUWfLjG0ZJ9W+47IKY8
8oFGinUk81NXmP18np85b0OHOgmDjss8Y1QBZHK5NtJZe/4Zrs7QwVxCrAn7XXSIwRSdMqjuHKPh
rUT2JX7n4ujI2qXuCAeY9mT8F2c9hXaZchle9tswkglD9npuwWjFfEwXYpG7E3wThKqTk9MrZc6D
27MGNMrmAT1blyavcUX7nAT0HOomJjN3y7W0Aa58RNMel9rHosandcCuJx2LR96rEqPYMW1F4vFR
M0vbQNV8NeliEHv3Da/OkItZpqr7JkUCA1LSIT6nfdIcO1ayDt6dLcJ0BtblGIQJ8rz5s4GS+BVC
q8tySKfaWklNJJRfLica0yCAc+zSj1EMc2Nh23fXVNiJhFRjBlP/wmFq9w3Ln/hPAKEUiWWkhy/8
RSqDW/hT9T12QM/+jAVqB1fIeTqy1rShgutm70ITG7VNY0zKTb4m7tH0H/uaDz+sXgF5DoPpBxxa
U8im4isnUDkrFYj3ktIAC8JDENdPKytAm7U75T8CKRKgq+d2eovFMPx4PDwsaZhWgKHGB0JAwqet
2egooVdqyapg8bw8gYTzoMH0FnlDacB+yi4FTgC8CIh52y1A/XYFvGdTL42rS/2Zc3MqrE/9wU4v
Qw3KWoQgDl1bJJaCliyjJm1drMlZDeoSlZZ9zFj2Uc+FELwujn5pAb/r4/N2ABYoK9bLUeMxdZLA
+OvMqS9Wu5KcMuWjdERe8ZDweIxJe7HdOguBw35EZzyiK/TP9HlXYWfetQggiSj1NXQbf2Abis4l
A4PzgNaBURv5zIKFRxGN25EDEIi9+W9VnZI2dUz5Vu+Xj5a6jHUoQk9d+G8A+Eq2bM9ZAUf8nXYr
0c4uLxewGqlZ6DKyHCbotNJtJCIS4O83zSyF+sMsRGyY+/gIYC2Vk56COCPzCgPGtfrChCtAtEOe
6Jh4ffgXD5lTnXCwh64uPWvKj3xWNxxz4oubLAjDkAD4a+Lwd9GeWF1HMOMVnftVu6ZlD+pWcdJs
tRSLBuLoU/Oj/gLGI7/bDsbo+7NjSxfajZUXBwwefhCPiIkFxVUyhSdXefzQ7DihFUlw9ZT0QReD
g5d0JDw+Bh5qBoBDmSQBNY1pvSl5JSN7DaJga6h7tnwcBiU7DkIfKxVLGvInTYUMKALNOx0KoKYI
aqCuePY8b/CrFtc2ZsghbtMLH+XM3G0Oxd9Yh4h6cb9EcdnGenxgFCSLExjY5+WlLgQ5agLwPqBw
/u8F3cHpLnM1GU2zsc/3uSSHnqbJIZi5hTweorBA8/bJ8Udu/pWEDKvwGQTa/bpijCmbvS9WpnKY
6NVHZFIj7EB+5mfluSvPkYmDwDz3zd8ryMLbgijtFPePIY6NpazLwiuQElAe5tJ7CrmFtxiuI1Mh
Bg+WP3/pxQ5ae2HwThiXMEFQUJOiQEpGmC5SP4e4QYp0n/Dj22Ee0fBRkRYznA+CmoPZV1+PC0rR
p+OwDa4iHKMlf8RwS31FLtd/XBBw7xicGNpybNQ5wAm9bBjoGwyAw1FE+0jZEgCub+SZUDY3CS+f
rXgilTYdJ3RIRjve8coYu2zjAeK8+xjEFpT+ob9C6AzPjaTVAHkVz3SfNC71OYnYCw/z7BYaTKFn
WcdBIAXwVXiS6Nzrz2rrKqSbHEGSPa3TlZiFOIl4QHbohuq6A4cCAOFJleMlmXVMuPVK1eB7w1RD
kHZjcBWTLjx1Qp1f0RI1O9CD42RynTqrIgT/uPk7Noqfp2+eEe7UGSunHVh7XPSC7FuikxhlI5g8
a6rjDVtFoY8iHTFoZmFxqgEJAjCPoKRbqL7UcPpNAH0mM1Kkt+hrOOQRi6MyW3srbYpXuTMI2CfP
1XC/uooOBGSx/hjJWHRvCEVdkBWDmB3ON2OJaoIadj6b8ptFg/mkDsFJrMy9q87A1J8QWaGeOI0b
PP1ItP8xP4Kh3OMNmmsjUDOQX+SOaxI9ef8PCTK+UIjpcAL9dy+FIjaXXw3Kx8o94e7mk4E+bfNe
YCVc7vWpERjUKahJKVx4gKTxc+GmZaQuZ9bjyVwtcYkVtjPmjbp8ACJnR6i88WOtF0fQLTM1sBfJ
eDDzYdGEhzCpCvRj6HTpob6C2NitcwSV6q3Tpu6dZMKXFbq/AbpGJAMs9tGKutn36Yg926O4/nAx
feDuhb79Ycuj6atADjC+CJ8bv1ZGWG6aJ+FrnUStRKcv69CGlpPM/cczgH5kKbxsleSnsR8mH41q
lWuboZkwGUms3YA1/oKk2F8IRVJif1XBRcFrB/ouR/l0xFd5tkKvg33g72rZJi0pTOmebL00VKSn
xvaaMZbZBCI3JG0uzyL6k9mCBzdLIJSsNyfq4vjViQylPjq9NNtBvh30B1e1IRIyK7bJC5AHL+XM
icmnEshHef8V/VY1VuHMubdtac5pqcix6TYFPr7xRQysgVI4VF1yhZmGW4wXYLYtpGCv5nzGkmqz
enG71HDQSpLHzfgL0LmV/UsvLBoDUnEXEH6FPvjCy4OK6TGG8E3qlS/ttWBDJU3ztmJpWKY26wDP
LIImDJIc1Bf7xtbO1F3rGkseEfmevTJHdA/5/GBZ/iV8j1viLebxOyjfsBEtMFjrBOXgM8iiNzFn
1++76hJvnrbJOi1p2k8gV/2Et8FRg2CyNhvoGzhOJ6NZXDtBAiCDLgGzVJ/7cArJDuJJKrWKJODY
e+UsLglaBEv+J8C5ztp7i61dkXFJiRNA5f8ZaTfQrKPGGiTHa3oSyLizvMFkNLp9C9bl6Wq/0oqL
zfkL4lQ2+dFDXTgHRXZZQCF5im7bdouK2X0Szq0xMQlf/q/u23nGPw7Zn1anTDr5d6367X/ws9sr
/69rAN6uMq6YkVEHu+Z6fCKmJCToQ1Xpsz4KuBBaG6c6fmDJbxJyPk5NbFtZaBeYcurGCCP1CqhZ
V9M3lnqJlaoyyw7BENVrpysPq7WT0urr63akFt/FpEDWh0h8MaU5oYsOW30L848l0ztaDVgBr97Z
6axunmPS0zuIRTaCd+TBYku5GgzWzyFMB+iXz5VysUk2e4clgwUvv8w2GHIRe/U+AcjsOETea8ya
JC84OskeXQ9BnS+iHjegRqwX/hZXDEAJSrXt2EWmYq1ElfDh9YQK2pmdHu7iHtC4C5Wq5Yf7CkoM
VtNlEi3zxHcFPGosytyPzrbdtcQDuXuukJ1X6lp2qCHRZZbZKwwe398jsHTx+6l2fDPHE7pkFKBi
0o2xhzWHw9YXeA2iiRbiCNtKqk4Wg0TAVYtY5mw0oaiMD6RUA6n9v6O9+qJoukVMB0mEumEsgNAK
XpBItk+7S65Zwix6QDgsOoztLQ/0BVT2Aa3KNFtlQPccbZ0WPkeyqQp7gsYM1p16KV/IfUOWAIV3
MILksT14GOhMkLa+Fo5dwOpHt4LVL9RZGP6lF0atkWQOXPAqd8xN2P17hsQiaT6i2aHt57XICcgW
5WJMBmBhx9rC3D6w5qr9djjch6aVmEIZ7jojniz/bRp52G18FlcV51Q7Njh/VYL3Z/yh8zBWD9dj
XsWTBdFWZ8JofsKezMJYF+8oxzoM8LrqxbxVepMNJQVttT5Q/zMRYfN8YdZQ+uvEE68EvUvVbfZ1
hK7+JYBORHe1Zzc43PfytZINKEpG4wVtQ2HW0Vt9jzImYR+yGr9g8EDio1/gt1f5IlPamhkQ9paz
Fvn/nI2+2EgSyqtqZUxbMSi/5ZIE8q63XhENv3Jk6F1JSiG/+QbYVMjlZPNH3xjdlH5bHfHfL8g/
GaUZfaN8OfITCbO491wHTBS9G41CFh9KLq5uf2kSG6FAB5tWCpQ5qRAjqN2fVyyFDdPiiGQEl9kT
mURo484SXPe4KphgQf6yFvjId8mu+1JFsbRkxRhMA7KqdCblQQOeO0CauZp7kjEWEJC+1awalUp0
4WOEQgAjHJ0xoQ/mZ/C482Jx3l50+Rws8+dbNjgwayXKUj3YZAsLfifyRuUsaDBmznWmg+FAGsf1
EiXUwaNJoBtAyOWMirankyoxukdI5xV6abb/z+n5YfRUfIXjm2YJDfmkwgDDRbwhBvZOP32vmyS1
aD1WoZZCtXyhBEx6FWuvDmImHrtXznb+hstR2n9Pb2ZLT2S3JiIg23Q+6c7NelU9ET8l1xs4clJU
Dh/hl6SRlBGsS+CffNF+5q1p6optSrJTgMtKRMHde7shaS+XMES7pIKHuf/TcjS1s55W99A82DB+
XJnyIkU98Ie0ObUOEoCbu0VDdT9xjXM6NV8dv3G80JH03bAsOy+KXFZctZxnWtSfxsmXBHgWVVBx
35ZfLzPMday7N163OUWH6W0KJAjyxrnU9M4jZx8UdWNGhwVVlO08nO9RX4P7NQ5vRvl62fM0EIrU
a8sbfZJeJOFCbOSPYIfu+OC4RriLfkR7YxHX5tvjo8x7XJ/+rKTbTcrO6xVnw5azZa3sR5ba8Qzh
TLRdU0d4o1iJLZx3Ic2Vfgzpom7o3kMX1Vm8TMcws5cbkYi7YRSHkS2z2v7QeN4FSrhvvEC+UBbf
eD1lgIhxUYWdQ8NoL0uDuh2h83r4/0wt9BX5YbhGIdmoj4TcTtNLj/6jY0xC3AKqDu44RhZwSKZM
h68K3tCOvPYWO+VJx2nVSiupgRx7xizp+OTHKfZZd4ZYHiaFkBTq5UrZWKyHfaHgBAB51wpB7b/y
NRIpG5QCjHvQ9iBIqVpzoEZIoCaaKVWDkznH7m7NIQ8G53gnGJ6vFGNkOvWZdECeyp6Juzny9/9H
xnt48YwlW0ACUqxJ2flv4fy6A6GUHuxC3tjgRSsbQ2V6Xl6gvgvy5AiplPOYND/Uq+ps2r6qVCIC
JSJm/ibdziu6U/gyJPlcpNAx549PjJQljOaR18szc1SHoZgKpYyW4NMGPvqu+wGW+uFS0FQWUaQm
FjdGacAt2qd+cpnYHo/Xr9crQAAXw/MONtnsqGC/fOznhWxqGJ/L/VcJMS7xyeu183ml2PXqv/Lz
YaDTGgWuCsHnZG/Xx88PuQkkcaD5aFyulPe58T4I3VDlv0SBJPCtMPyzdGuPgCvYTlNNVt6GPd3F
BkoCPQJW+GKXCZUwaoQVYTzCd1qwDOu4CoYFmDn+jXHJmebGf1bq5FJjYmGGPkLoibmOKi4ojywM
k5YGYmgFLYaLkunw3ROqUL0/NjNuwVml1BbPOh1N3HRCsEAbzv0Y7CpgFAp54bbPjpz9Ur5xfjaN
HVm2Xt/h5weZGSAtYzkbTs4CPl/CuOjrlbYZ/J4Oru9/A47EmW6l5VbMrRxqXP5CRNL1ugOSbTym
O0GMckThsrWOxGmgeAA6o0P1UyCcWeBDZFHykb069Trv8r8X0sfYxnE0fyYkXlgNfs4kwE4k3Yo5
26TXGrqVNrzB0weD8Q4xpcOhJcS6mh3LAh72VHbFAqEcFQxxijU9a/bd13JtA6L6IUguCTsYf+8G
45bmy2DKqislCNuUIHYxgUj5KO1n+4kNfanSFAvRVL3dI+wqUoVEEClC7kk4tv3Qi8OMNWNBdPzT
6bgzMa7Ut48sKU4QZnqqIK1RzG2FJiWNiVUXUQOF8HRoZ7uZCDykboJQ64DL3gD3RfntOdZFr+qw
iB/mfVVL3RuyQqMU/QZ54NjCBMFDUmoYYAe8OzKTp0KkHGNQd5/Wv8vh/5jxRggCMpK4l48PChkI
UFF9+WNSGhIhyVFk+ZtjWELHE0WUbNF5C4TQmNwN/tubp2GB+bXYI+x9KV++puny+Wc82BEnXNMn
x8v78AOUhlVkxJd8sbgtSVyV5wzhwYrYNRF3ZfDwcrv2uKedcZTsOjx002Z1K92An4a20/lZ0Yjz
/q8mDiS30/GbxhL/5HWukfd1c4y84qKthKxYduvB6VxKLIexVcnpnxnPXSQnuMWbvtl/XPV+VMvC
D0UdXCOTRM9gaZVpmE5hxjW04waB58sg+E0h1wiaBEHHu8oKole7li6y9AYm7+26xT99Rfq0VieQ
555Snder89JnNMD4skujsft+gcYSlRRAMQfqzmN6XYv5BP90q1eHokkklBmRbfutwLSKWGC4bB3i
2+p9g+lAfdFV+ZoSo5gtom5WH4zVaMV16dKR5E4ADhh5Smm5XGR4RQkNr1yKEYXPhllhGzhYmZ4w
uyzclx1E9qQIPJYvhlBq/IJkuoUcyPtwLCqYP4LNPkAMlzhYsU9+sBVhfFbtMqCrp7OaHmy4Zoel
f+ltm+bbHXzXlY/AJPDuuzepbCfR+f1YSjXn5WXRvBGlS6Gqi8EfBxuN/si8Ar2fEIqpmNnCAr2W
kcWgoj96/s3x0srqw622Vf1slgCoeTwLZoUkIANsK3S7ge5BwcEe0pRNyu4eIeaiH2TRps+J2nss
FMdrRAc2aEuBS72GKTSrqVIMEvo0XR+yHuAlA+AjEwUTsqJWecRWxQbhxPktdTfeTKMeAin4VsJe
x9JpfRpdRuk69KeOKZRDNPa1jf9godGvlory9mehsy//dSCQhpd4aLDGIV3FILUoHKujYFKp8kQi
vqtSJon0+wYYFfXGnrUReySvkkku4ZdQ93ntJU+SLWuRtNFxCR2H6/AqSdStw3UmPf0xyMr7Ttwm
zd/IBZhMsp1/zcAL1sykqU4jXeIgYB9jsWvWW0s8jZHnA9YH2KdYOXvMsExLCNDMWZ89sLjtBNdM
jq9cgT/K/eSMkAO1qyq1r2rgJme494QIolTdgieJPi1iPhnsmxUzkwUEAHIxggfus2a2ymmwGdzR
9v++epFeQApp7JDoJw+gOEl4CSI4r+hBRsd+MBia1p9e+YEjYnSdAwLvhthvZGCE0omuAbNGOyUf
xuIUKathNXrroosEzro/ds100jMkQae1/hC5nH9hgBt0emInB+aw3qN3fiJewOHfgiU0EP8cVO2l
ITdTJPagQbQhTcqAIFr9xXSigJlPijF7YSOj1hLFGWhIBFtPb3bYgiyiotv15cgBTMh4OibylLyH
kzVRaSScmurGm76YDil5rnZ9NvYBR6iNExGLJDS1x85dz1RBGhMH5BvsGzyvprJ00H+mYVAinwHL
hCwYlxna6WPQksZ396rZ50RWbdXGyskt7WZCtLD8DyQfqxAOVEdG7C0rQubdtvKE8rtCQYP9kk0U
WbxDHFxsT3mbeNUQh4U6h6phSEGJrgVgNtNuq95XIXaNfv/sj9xQdy+CDB4abgIrCZEK/B5egtJh
I9QYguiZqt01df9jy2rrKCc4JNjMC77wXmkag6eqA1fvjWDo+mCH95eGPtDsMBfihwc2VaSc/nT+
NDwFFrgX4W4mz3rWMRNwv9qAtwOXX0o5E9m5OXtcTQfwEBj2dec5AH5S5FIR4SRxrFDZf97v/rou
Btoerj8su0TpFyA65DR18ow0V/YlUdgysyw/9p92BTIUMGbQiM8RYJdTmiIHnElZHp/Ee9NppCFb
Q0gYtL4SpahKoHUTv95KxsdR+ITX4BfaX86cOD+469QgYGAO+2d66Agcns3or/D+jMR5Pm7Cd6Zm
jW2bti6MA0XX40wONp8cxyyk4zGgP+88XP+MTADEEH7w0bKvQhSXfFOH0I4foGfn9ergivhIsFn4
E1sgWg7O95GM1pSPHSmIVqelTnGP2i/JFqnFlZuXOPqUa4HJ2ojlbe6W4GzSTAw+8bk3H3UfVSbD
+bOREkKAvERTFWIzZaKmFh6Y7+QujoUewn+pLu5263kOCAhd4OTNPK4FcxrV1bNfmB19nGfInwkR
4Ry6p8IpZCObKlVr9lu8PkoQEA2bmgyYFdK+j03+9fKKSpjiH9xXV/dKXi0Y+dh/1+1wQKRN9ZD2
vVoVQS9cS7RFOJug2tYKf9fM+r9PwlGUUpczU7EiVjLSD6PdhdVs/6SrV8ZNfp0jbW+7Ad/wrKtb
ja+9mKGaEnNeGXD6KshJgQf76ioxcKle//l+gda1Lue3CKtVZ1ic9PYMF9em+IDCuZ05oXtdiNjx
XCzgJwgSuboBQs1LC9Dup4CN5+HCgxHE0LXEuuKs/Giq56t4PvaVBj5zqlXyJFlJ75siz9bB1INb
qqBRCkqIxm82+o6nj7WoEiRbcss/8SRGYIAFxR96z5za3NOxYygvgMkmtD7sm2ukVqsGLU7Eof2b
F0e7jIHpSm0OCRdCeOiedVDfhrjZRKHPdJcSYorhI/25L4Y3i94dMfOSi2oWT/yvuk5e3O14Odj+
Cw2EBiTT+UjVBJPFcTPfuHZVpiVTaAZl1r7cVxr+Hn4Zw8m2IMO0XYqMzAxmqE8/lwXw1w4x0Sl+
PsoiM2CjVyLA+F+BZ7WXdWxd+ZDaOq33mIHetTPFWE4lcoGKQvqhhWySHoNUnPXtyEd5VyGkxTg4
V6Ngmgu/MjjQXXfLzl2WIt4V64AkgrAf87Q1l1gJbWvcMWGWEkaqEHGz2+cZLtwfPNweaXRS0rKc
zJWu3XWqp/R+o1eR7kAvhkvGhBiSaFvyXdPGaHpziOmh0X9DQ/ItxgA7tIAnhFRfPuLysI0L8mSF
c3/TlWYOMZEfnsl+OWG4drWQiGqVQSviIVZ9/43cga9PLzx5p65tcLZUj61Oxk9dv270IbFFxdmo
oSel00bxAfqee6bF8Jsrj/EHEoCQVq61a5ZLWuA9RIv6ErveG4Kz0WKPs8javptxowOhIJeiWqE0
57wV6Qebn3ZnFh+mVT4POzZBTN7bFK9ipRaVa2aQ5et76UGlsBb5lvOVZtVCs0PgXhdt1Y7Jt9NJ
AhG7zvIk2eTAjcvt6/Kis4jgfIT7+zZl7sVNdG4rlJs9zlZ5GMKSz27wox6Cwi6hC0PorgUbQDcw
KURaxp9GPzAA0FhyaHRvOUSDHiumId0VzmWazM+9CvP7qpcijttWBdVj2PO38reOm/jywN9S4jY2
c+gXGGkc11YtPpYhKbV8SsZ5huzoImHxuLKBpGwlQELbylGFbvk7lJwAkWyC7IVcGFPPQrPH6a0X
B7NQePEm0usY6U7akS9PSUkzw76iKuIAMKBjqMOHA+0GuxHA+YTRbt5H4flrWZ71YjCHrqFbjwf+
iNRA4Wr+A/nup0v+yPOzwRGYt6veVbf1GYFwK2dbvraIsFF9wiFvYKZPE3mMxEZQwe5LDnDZrOVE
V8XXCCZLiL2WD5UTtS9QJeo3eeLtZRIQKoU7P6h1jrTxFT3CGRyej6/8IPcsBmILxI+/x2bXt+8a
T5crI6DoAenmvXb5x67zjAfIsFCg/Vu+GgBZlqg++tccA1Y7vHumz1Pru5jPYrPjejtmviSAdDTY
mqGRkcCYzEwpNoks6g+/Bc7KQfy9B7p2xiw53k3fLOMj/4xURiKtbdYHTn29XUp9AVjm/bU7JfLl
vu4wqPFrc644OLyT8bMxrkLM0NqGHe5FcSLmErxzAw4SYgjMctxr8OLznLyuhfofYVWS2a6MEaO6
RdOJPPMHGGIEKJVSyhpXDOAPW9uKSowx3gc8Gs3Bnb8VaADpZdvl0mGRfBV4g0CesXAVGrXnk4fA
xqFcbR71MkBgdNBBHBua1qitxz2LwbZZih9vL6Fmfh3KdCaJDVIbNTCDTzgb7yw0NcXC51vF9IrL
0g1PoRfARcrCHvfU7kKJfuCLff6ojWN70fquqxjGld9uMUfWUEIzjnxKqR3Q0ESJADWkM1VzjS6M
wzE4X4vGVKI6sELfVcvehHijAYukdPmCi1Nt14mMXTUnPYbkY9y3CNolzA0BOuv5/XAym5u79dOZ
urgxN6hZyh+zlOQyNBUE0l0VV+/HyAeK+w9hWb01ifxIHhSFK2UMIKsFePDZxCswXTj10BLbGItS
HmORSaL18SJdrdCLlERO/+QNuRIj1/sw6qVXdkKkVfYJ3HkhFK9+MIus9gs81oqwePEOGhrWX/UY
eiZyI/r8Dsr/o3dkdsHqTS2k58n+Zp6/m06jDso5oYyvVV37qRezraa2KBncvZtZIPDsh8iBM4RI
X4h5MTEfa7JLgey1qxKI72UW2abPKvpDVLR13oiQAvb1HFMjZGioWWRHS8vP/EfCNUtir+EX2fGA
za+EIBLEeeEzd8Oc73S2SY2Y1ftmLBSgTwu07OnzV4hShrZcfUU2kP+T2rITfF/88BpzWWuRHpPV
HCeNqTqneEK1UwUOMyE4fW/mNxZvkMfLagxCe+30tLocFLbT/tOMGxabo5OrcRip8U8E32Zlr3Jr
WYdazF8goIvsAeAU1k3cHBV9bziaL1MUd3n4jtUY5Oe85N0Lbz/qMskApAKLkLAPSpVZsZ0KwI0d
XYnL4UvnFflpjl0KMql0bKajVT79Ej4h+Uu1K88j1tdIvHRepfl8yCwaLdhIhvOdBXRlmPrhkThL
oxXss/x5UERBAAQEV2eQ9QujIkkEkSK/Veai9Z/LMHS8pc5QTyPfLvAYfXc59HOV2n3pzvUTVH5w
PRRxDdnXKthqwWm0WBxFtU+qR0JmfaZDUcNTwrgWJFQcKIEgZAJT7zxq3QabmjwLURVEs0OMfW80
57o6A2xssG3S+2kn/wlKKNnQyzRkoatiBwHIqmWzS4rkPmiDkfuhS2MpmjmFpzeXOTtzh7jKXYqI
f7fJou8U1bivcbBPk1pusGms55GRxBddykIgX1obTt31qb0JLMBkwbx9F83W8UR4EhmCyaB3d0n7
7YGhe0RbueU/HJ7bSQeqeCcGkou/agEfZzodTU++zfcwSaGvgDZB8Zdif/JL6dOsPg/bKm/5yV+W
CBI35g6W+iXXV7VICMWb9ypHp7gfnLJGC8LS5kfh/gUCAGtfhlgPLCZ7MEJGIMe0t1AovpygZ2Ff
7VTqZCk1qdhZtBcnCdI/0JEiBQ5Arefv0y+Vf5w+EBeJHHQD5/bCsTpp4H1t81McCtGlF7auECf+
xzHiJXyi8I6p5KSDBy5zpIsYsB07QYDBzYS9vAfYOoqGX1igNnDfwuq82o9Ty+sHOkDEjYw4Uawe
VAeIfIsYmOcvfyXioxEr4UYklDNa6Lk22Oq272yJ+FiQo5tEV94y2l4tUhZNUiLVv2CuwiQtiCU3
jTngiOQumUdoZ9cb09Ypmg0YcXnO39JQsn2FgWgbTvKrOkmCYUgAZWvuuyC1hjcO6rSBqP+qBCCh
DR8H9l2FxxOUL1zwq8cZO4yR18/D8K30Js49r5osa5OtuVxCsarspBAlZk9EsyJPzeMPy/vCNlcc
MOy2x3J3qCSwJuTsvM34JT7BLBsh4aP4wtye4d95c8Zem3cBUVh6uzfen1YdLYgA0Tq+EZj8s3ck
AZLzsURK/TysqMG4AvRfXirKXsFCkQDeMoeecmFI4sFKcT5bz37tyjwLrlgVTNEm2yDrPkOSf5PR
c4vBGobai0hCRYP55EbRkUCx9YpIYrc71+oRjoYCbxCJ2E4LNfyw/bqKNotB9bi/g0ZXxzN9OiKT
WzZIBd9cGNy/tE9//hSxkzIqujYslysNV9PlcX2kPYgwQQ6ddjQvyeVLOeyLDdW9tKfpU22fZ4lJ
WbKmTeBytnXHN4pVeSsRc3elI/zzh3T5SVmvTB8tqXOPowQ/HgGi9r0jsCFI0XHMW2zPZksHgsNB
VlN/MRXZPyDMhKDPF93FNfjKg+zt/Gj0PUP6NihNpz4dKj864GciL9cn0NIJ2yWr7u4nCEDPAXdb
CISkwF3FJDsyylsXKmHfWpQ2fLGDME00AcEtWFT60faR3zv0lYYcYZiEzI9K6eIR4yLW+ExBh3Ne
pdcHuG+G1lDbnElN28cxefQZZ4+nSGY9rRwgMOvlupZ/BCNaXJJZo5PfZo9C/MJzMUUP72cawPzW
xHB4PsElRKgafsCGs4VxE62L77tKu8g+BEDRfVGETIqfu3sfqU45DSXB1SSp6fknW+HV0/SJoDFA
SmbRtnCoaGaMJAzuEhHvRa2Vm/tZ8WWpzwRz8KTki39hCtBaaeKGLsmGj5Yg8yQ1IHy6PsMmYHFv
kySw9jW4UHJTv7Dxx4SGtCBta6xhJizfSnDJB25FNxD8mdiLOkV2WJndZvm/5PRoODhmZenT+p3+
Lu/NpEvHs3LbEPhTqZYnmMwfL/RmMGhsaLxKgH+mxdayetPfTkHLLHfby2FYj0ax6XTTZ5QYIQBS
TwVc30ULtFq33du7Jol/dvXHqmNGpsKQPoGoxMnphjLq1Peyjz3rAkKE301Tpjsis3NFqyQ/NzN7
HKb2dO+IWiBnoDCUc4kAR38eYO0Zqmmy6s+1aiorpTK2Nz+Cn9oFOqPjXRwr0p3EwHYTbaxn5F8J
vXtyQkzLIYKbRyst7e+J481LnLoabTD9Mk/wZMWs510JIdf4e3iOsUzb662fGIPyzV1Y6Wx7SyL3
xDefwL1LxdfaBTLUEdZi+4cok7A2qQnpjLz02wHEU1FNMq37EiUEI//ZGXKymLikeEQ49gVm35z9
dsEBJlqIaGWGd3LGZlSjb+/ixQ7wZ9BK7ZIaLHMr9DTA274lPuSsXgwKNe3ExoyeRv9hVujE3fbc
elFI9cwtbtUPpdyU5Rl2wGunhyyS6wb6ycp+SATTZ93asDt3Ok9cDKrMaQA+sfNRw6XkZFFAgMjJ
pZMMJMx5MnER8/reft5Xt9UuINdTnGh9e7nP9Kq8owlzqKO3GmOZ2VH5hTuhYp7l9ZtJ1rjaTNH/
Kz31cfX/ET6cqbLs6xvAVUrq7vZvvJYe3dChq4O/Gn8TuIbZdwqPWNvezrv8CTAhjDWLLs3klKTq
8bYBDdORQ+oQqRsfwT0Rly0ZYIAI4O+rqFGgNButq66mXnhZ/GjUHMdLyUzKcpwXozRejlegH6lT
MRPw/kflkygpzLH0CMRpvz+jBhsTycJ2LUiY+OHYXQSqP7fBDILdW3fjf2ONqxo6kqIj9In9fGCS
ffHK6fIiUxI1ojTzZIpYGjRs6QdKlsG47tkxktIxvvbTTGcPs2dgmDIFfUSSnGmrg8AFbvzo1bME
8GI0MaESRXvMZxpTc40me/P7EXLMUOcRtC1p1P/dv0R9c7fRewxFmqIXsZiHOc6Z2t+qbPMHBu3A
nPl9z5hralHKM6CzWMc2EDy0+prwW7aIwlnrgUmSm/ZWKQ7a5lFMgBThxuFjTwta+R0/Bp0W5Poi
M49hZbYKRNOsTo1o5C5aIYJPXmL6ukpA4E9qvIugce1/78/7oHZOH3Sblydt0tcmUz1wSRpHexBP
Wko9GV/g4GPly3Ul853+Avfq3hC5461kxPmaRgEWcMYkcNQFUf4ZQ3XDsayV93x58gyb5f6jobez
8IbrlOyQMX8dQfsx5GXuxYhNE1qoRrgbzBUMuJcmXdiViyX03yZJpXZd9Cp4sAK+s466Z1itSsNU
y4Aw43MhsRTAICUd1xr6n0sdonwciGUG3wFXVKzf+FCVtaU4zC8/37qc2VTvIOKaRe1aJg+01gq/
w11HyiNz1VDkwFgAUSv9QnqmzRMtsPNAxEGlDC0HYji4IZAkN/L0qNn4ANKVHkn7EfQ8KomKkYJz
tZqXGcvrVS11s2Exn0+KLqcvdc+CcrVVLhfbEXFFJ5QDpA+H6KuYkJ1jlvHXrIlx/Li7i40Hak1Y
Yhxgxgz5MQWZFPP481aDioco+70fbsKeC0K5XIJ3ootfZFWjhd5KX97KjTxzoU3ioaRNyg6ujXXW
xG/6ikCJPqWQkdFbXGO/BDt2RvXP1mV6vlLD2+OLG+PDGkZNGhK9NlGzmu0j5nMVZ1ndfEGHUIw1
RJZ6V71x7TqvPb4IfRy7UJ3CHyXAZEILChVHP7Y3FzSg15mkYdvQ1+9xKkJahcd6+3645AeDXNke
kilYW74Gh0pgiL1v1eKYjyfIjORuu6qdzL4+Pi/K09PYIL359RYs1KW77YE3+qM9QmMPWimQHQpI
b5bh4YYzIpZGKzfnB0joW+ebB/cY/kyvreXuS8MGJx4x0GkOsA/IWs2843bcUPleawGkvbqSJB/a
ci6NNXMbFsZDJeWdxlDpr1clahi5ubUOPTg1cG+1/ynRIMNuya7jg6BkfTv32F+kaNu+6lGIpMJa
FReGmsC/YU0P0D1ni5RorS/XeR4/jF/6fqCRhKFUje0rMj75Rpf9KiTzbq0Bm47x8gwa3FE3jiec
nHS6qpoFAv2bilBZnnyYCTiw0OiyBJCJKJ6Mol3EWjp7VKypJwYb2x/eS9UxgoPTqH5sRpB6DI51
mvYT8gNtbv7R1t7LyWT2t/hQMAfnvrEMX8Ut9JO55t3MAe4pYvUwJEUtrnJSnf3VHCba2SVc5G4L
s6Wb/LbK4rsilR7RkoR3IpdHpRg2dHiIYtNFq/ovlzSdBkRak92YbqyPWw5G9WXEYjKoVaZdVbCM
ci0ezKSNffyv24PWg9QuqI1AnvKYm6tqvwZXpZvaGxA0y5ilvbVmFaglnrEDbDsEnTwUGH/QEXu/
CHTqhHyOZUwPzuyT+l9kVxo+3dYMZx6y+XvNp7bwM2mq1swZXRdeGpopkLXR1Mi8Pez8Nq29Oi9G
hcOS6icdMOh2M0kCHQBVg8h8M2BlzDZMHM1Qw4AGBochmHrg/liXImKrJpxhA2Rzq8dL28N2sWNB
Mg05906SwND2VwG8v19DKLVbPVQlwGu4y6bb/kNSdRGV4x2uvhFoq46forgQofYcnLdlBNLaT5WV
KqEZBmxhfC6LfsI5ozHDAZr51OIY9CAFawvOAtNf0o09+BfOEwzkbCccWwoCUam2spsCBKiXOXH6
XoQCL0zfpjH0MqgZXH0AEnrQBZraFLyM6O+0aFj4bwv7EQ9tZkx7Y/jwAc7EJ/E4vKSMPqOY60wa
PNVVlMD7Ys+pc9qH8R+oJMOvt+3G7g2vRFXFdr5geUVVHP7bnM4geDfkzBT+o4HYAA/2Q1q62u3l
aH2LMVGHcD7r04gTTQ/skVgpspL3NKvg50CbC1gOiR15ADOY/gz31/pt9ZhPHTUM9Fny0V7XbLMp
mzEzWKea7EjOoSid3EKR9qP9onmepUE3IxrqMSxWwXpki3wfbnJNNFwgYBl0XcJLG7pQI9NAny1+
DEUa+cMmTFVlAIYI2LMuOg/nIKcugGOctMFG26xANG71PHCyT8DWldjPBBQu0rKPYk//DifbcCwx
r0g85HevRUhR6zSDjc6fxf0tVywaJ9R8zJRB6Jl+ZHwYpPNM+VohrhJPcEEb10HU9wdlIfQV3YeF
suGNX//FrUaw1BnR68lwDxRWidlXC1fD2SMuG7iwryWcvPW1CX1+NSt9kI/4nycNXKEfoIKK0wJZ
qMO4Agj3HtPrS+zTTVN/UQXwPPBQHD2vwbQwy1C+8pU7cIEQOtp4xybyEDtmEEOKYBMsVftQwRMB
pbjzEAeuqoH4ydbY/QXVXa5uW4uMucWpDQq1XkKK+KBliKjDvZv6sn/eSsmCM7H0lOC2C6zKYh+y
i5NZtV1GZgA2M7fV8Et8ByEYJeZXpanG51yvN3TaqNIeD0gL2DIiMiHzByIUn0CYjoTxViClF0hZ
WYnMsSe3291EjGIAjauWkVfVgBw36Mt9k1rPQHGyd5Xg2V1JXnczyyYEqIDL1sL3coP6RKy8kw37
dH5upqO6EEj9PLsbvxxPaxQcHafCUefYlDdkrvKJKHvL2bD5eFr4kM1blf8zlF4NkBPnJE+n3890
0rjYP/d7vrOEO/zWpLhFo6BsNVoPft/V2AR19XogOgoSx5+cY4dZOTA68I2BElcXJ5M36l0PRHtH
zqzbUZcYD+mQG85TmBqcjimot52J4n0Ymh4vk6VZnzfS3ST+QbX8bs6naXClPNqUsZbG/3oM5QDT
18mpUs5dhiJ2QBtsDldKBY/CjA9XcvI3Ths8pB2jmiVI/6U3sIii2O1ZMd2mWK06a1qHZvccLWLp
YrqS8NncMqKOBH0TZSfqe6JcKJilujH0Ztw2DLBQv7WqxSmTeN6K5eIQ+2ssIuvOJYG+9PLKBrXR
y62ZXnJoUeOd4qRaufl1Tp4ZggXBz05dHcVXFjLXMTuQivFF6r1Am3sKQ2on03XC0/lL1c+8Uw2m
zYwJrSMOScP+73VIwlzOHiYZfeNsutkhZNjqYWS+u92sxVjwA8zJxhh5oVQsk4Wg9hu0CycgamnT
UFZUP+H1GpiTZhXic0WjreXReb9/eC7ghrecojaGW6JPLT0qVMS+2Y6E6Mtj7AcLVAaR9vs3hRi9
G5C5D62W5ehYITsFviG4sh+Q+VjmIz72yc8wpiewX7X4vXFgghOByi08N2GkzEzZE38zI7Q/047V
DxNd78k2qORJOYJ236w1uA1NKQXIlBI7Nw0hRNzf7O3XbjKO1A7OKtnNey1ToE99PsaS3IgXXsp4
5ks3uPBKXKJsJKYlOc+nayGh39mN7LJqeHw8gS1bFf8r+ZjYYrISG8XaTB69ueD5Tpxaoazj1EKY
GlIWbTXUqkZKAS8xgrpPn4zInm0HegkYyqNZ1mU8YGLIPy0gTw1aEdUFSVTWLk7YHuZl/NjgP3xg
Tsx+G0wP7J/VFYr39+pE2kkTBDOjzeQHHBGrq5fU/SG8NUCVF8xGyx7HZ2JftTxGLz+PWpcMQql7
paYtPLMfBXMZ7+t4CmZZr53N/YRusNbblijXSKNSKZMtgo9VIObTrhCJPOrHQs4SEMY8G4AeKR5D
g7gwgPfhv12ZFQTkpc4p/czSRHIiiF22JWLoqFy5LKIrGfJkpfrQ5xCiT2vKyCIMAIDyqifkNqeo
KSrgCYLEab+lE1DScA2AStZyguCONOvl4YWglGC8pfveYdBYVHmm9lz5Qswn49b5D+tyupWw4znj
MRBhRXoox2Gtz25CWL5MR75bbYHrVb7KYpIr00DgGorRzyxns5ALZ/+F5rvcIvYWH7nl7ZOlq/VT
5KwYoOIP/jfZ+Zd68BDeldmN8QH+MpEzcxoEtS8rRnozao0srQrnanAXID/P1LCjtERP+6YDXZua
jvmKmMGg/m671fAJDSnxKCoAW3ckkwMC8dBpe+GaV3Clp2d2X8ZkL1RUTvHGo4BiM4BkVyTmq/o2
O8ERn4NDr0zS+yDGsHMt7ytnXqO1ztrolY2RjnUrSnE8VZ9HqxoFhR2tqN/7bEBx0C4T0pkAGIvZ
dMyLzDg8ACn5hXVw7BFcPGgV6FAkUAwzyYJZOQIjpDCL7RdkWlPUmGMOTEzNKik9ZgZT5I1dhS0J
CVL/q1Nl6OzBc/lOXFYYPHcv+098k2Q4yp3L+Jqaw3+7QoEszYi/iUxpzhczcIIevz6XfBOBaO7x
kX094SvowzpCIJ7yGgcA8yRUSFk7PYoox+UBlulsbvOD97YkYCuFKUQcUbK084WxfLHNerMP7Pne
WWn2I6GWd7jiBE0L2o+r7MuZ3FyKzTlrmCx/rs4CN5JdV/dtBmfS74q0qVGX5bYaaAVTDx/JL5/I
fIGNXFpJUKjpB6/yrUGubmuquTJPHp9Sv4esmFnHZfbJ3sdxfd8BuNMmyEPitCW94MNfv6y3Nw9X
QH2Gbc6GbGfi6J2vUnUVxp8edhVxrr8MVPa1ytFL0GL1XnovAJJartg5IoYRyp1/8rzO0E30wMUj
eHCCq34kXk28UdJvvU2mz7QFDuGItONvy6tJGdHAFmyuQ57jEbkDp5IfrlVnvAhNieutDLKCmAs7
IpkJzCsAQvd+eNfe8Rd04BwiM+7RTbyCwzBXqFrh2Tr+5NkZnPWLSf2ew64bmCFIKtYVLda2Z6MP
m/MHHWAh6Gco4rvRQQTbTEV3VY+5WcucaYttPNh2Sfa7YrQJ9qdrys3cDfIZvOEawGipEnNkIF2B
WqpOJXkZRrd8LaXxZMNeGYmMKhAdBgIcSnmZNmSRB4GZ4ciWTKFbeup95kTqWtxHs3NEhJ77xpuh
NTWviSIn1PhG5F8SL3bk67SZrXJDi5DqfIPITB7yWUPdR1ybCHKXBq/XiTZf7vZzQzSyvMz+d4+M
hyvzZBo+Z0X4DhBTY2Yfupij7jn9HcEVwA9gkH5ehPBtEIRaiuXPmohKG/z6k5cZds9Yz+UGFGIJ
radlNTC+K/Caa2znMf96R7VucHE33GCUBy4SblvbzASTfMlkiEXmfvzyPqPrZTEBHwUey9GDR+yE
9RwF2e3d9iQIkA4ZUet2OxseZ5UmrrvhyItNEPXfk2PboJiLF++xsq58EWe0ALyE2pwcVE99qBGF
k025KN5kOzTacMfMk/urDp1Qh8Yid6CMl2G7Ph+yypoJ5EF00SYMdSXHmnVUoAo9tQXVDs4bXF2B
46+XDlWIlQj8qSQ7LEwiDlNM0E/KsQ12nqdt4v33UXKJCMFpdcK5yXjizvWzMriTsEGwAOn4e5o/
JDmPUDvjxKbEHlgDrXdTwLff3sydNUkt4c1+ZrR75JnKrxexan12s9hYMDOCwFQZM03fKyG2o2ha
1OTe6ynImjXGHV7Z/iF74ucxAKYk7S5UGpMruu0+Oa3poyXb8rTcNYf0INsk2ZdCU0Ypx7sOx3p6
RUmN85Xh9sbHBccTiIYiqVhKkUpcoT0e8Urw5ZzTCtP77Gsco2iFyX1dnpqmf2Fbqo0PmuwMpzE7
ZNtp0V6L/JYnFLy4eiLvVVCyqx4j19vVtfZTP1wwepvnkHZgeKZLWpI0oqAYy5u8JKU87/cERjlT
or9lPx/ZVzHu2/jfhv2f+L7LPZp0V2MTzAzNbt0C3XsohaARl9IeLVAF5+5HExEBlidbfTQrqSTQ
WMlum89DB2GdINHj3fCqTEMr+/7kAQhIxhvvSg1H7Z+jhVEA+G/avO4DdUT7qUa6+0H6PPxL543q
Mj+7Z6iXyfDeuq9ZYv89fobWnX9pLYG0bzRkq7ag68F+gCJATtF4XCGktmc9K7N/aBpKgDUktWbN
8ZDU12LepYf8NGZgYIC46tsfits29nYS9VFXtacfbSxfGSl6T9CsKORkk7iyHaGni6UdL4lEtAnu
nc9ECL+M4UMi3dQPYyTFulAd8nbYB8zhN2zU45SPglNgFXquWYV8u79gAK0vwfIyYCQB4UjAeurE
VouoEh5Dq8PIe0Uw4hu4pQnjmhA6GbIfQzw+xR2qQaDoKNB1v/myo9x8+/Pec/MpNpUle6Z5VYuN
4ZvW3HybcMFXUQpv49w4RTy7+hNT1BKIym1EJN1iNgG0tb4jfVwanOK7sCrFcEzXONydVN5GUFVD
HPISb76gaz9ASq4vGeoz3JaFSAHKn+9DHL5ZmMP+BLDonjU3EykqV6co4+kaZsllHkEnCDUkD0Wl
QuA2yo06Duaj/7BBnmWwLGOw90t4dktgzmM9nahf5G8W1AOjWvTvwLqlEjTV4cuf2VlKwS2V9Tvo
/W9x1o7/peL0cnSLBGJw+vfI4YQY31wA0bKBbk984bzBRmgMYX8lz9oiKo4dSSZ/zIdcIW2tl1s4
tjgOkrYIpcdK7xo34rIQ8xxhIqIhPhbPlLQa19kehjWmC9yRP4n6GGePCrrb6ZWAvSpGQe0bgudE
uZlZCSgd5pTJ1i5wav2ztVcUoltCP3MX2J2nphyQLx8vZFhwY25FZgoIU6cwWqlvSk0FhdbM/A6s
MC9fAb5hDdCtKs6xKB5M9VlVJ8DKURTCc9oUxW5Bg+nSad/vFV56BOrC5dPLs+ZKMfX9ilwOPxqa
66NS69B9lJtvjHQGusvZc5zOLrQdepBbIuLaSTA+o+uIFXOMQRiqYu4BaD1KC46VC139/N2Q5Z2p
EnYnqn/TnWUcsHmmuWTqDyqJH0NrjAhiQoNKkOu4X/5mA1W3HZRaULQIPQ8S5/2Vp7/9NfgWNO8r
8BT7jc0jVUSnNIgrjJoIIgRG1jEJglQZSirgMzW9Isam8Oz5Yfsgbq543Kh3nLEu35ZKXqIqS+hr
jzdmkCASZsnO9ErXCYn87ViWiiJDzBbb7s4VeD0I3nCxV6gxdwsQcTLBNxN/b0fG4nkqzGB1nqn4
zqSgSpWSq1qihpOgP9yi6kilVzSH39VJRjTM66gHIt3fU594MCE55ejzJY6YjqW8EkZU8Ggw8fhG
aGcSUIX1Zv4oDWHtJN558DgXfLvX5X2/Bsz4Od8B6+2bz+VkkOTT/F4XC3Fg55fiaBMYXPOjAjVo
aeJ/0jvg2cgpogTu07euTlWAsQgWzWRCtS2HE3EWY5Ri4UKOabAPCw9GjmK2Ax7Zc+V+s23pLDy8
+m23BQeOyO+KOwrzOwXJFHZ5rR5Ua2IYXgE3r3mnZNK6FT0iX1H+aKrGMSf/eeieEDqJi24FRajr
OULSSviSrXQViQGG47zZwuwkNNK2ZApFZeQ/si7Wu57UjvMrwkwZQeUnsai1gPClgMLUOUaglGL6
goWDl9R4SnIPCrySG09IbteTCdT2zhkCc3DgTpAbHFgCm2xVM45GDaxL1YzkbPfBojAFMf21iYAF
V3mQztvhQRSkNg71X0OVemJEt+MvQ+TgWf8GdsSNlQI3A0hWLpKBgE732FJRAR6uEBBDw8kzjUHW
AhGhAaoaFQ7RpvKvonZZe9X9yHtvTioSbklNG8Mor+s0wecQ3PJPkA0ykDtQrG0UHz/+4FMjIYiv
Q6UZ8d6nmghvmiTrteRJ9/ssLhp3ZLtGmKBBXptJgGP6UTo+1hTRVgKA5GGeDRMljkyJq7NJi8DD
QmNzknu13Amqj+8zv3RM3curqH1BVWIVwLTivf+TC34Bhdk+bMx3y/Hi/j+oJBo179u38j1ceALj
7Y1sMn/8jSAVLMQIsyZWUB3C63PkBdT6nVdWLYNwGKeWGZKI5L+TLNFaKsojJa7L9l8LHY9A0ViD
jX9iYOK0dxsYtmme12zlqxtHSKIp8S25cVuxNKv9Rof4zLxHQ+cA6RWV51ahbZC3BWg9Xt0jvp9F
y7K2aOafxi2eCOefovVCXLjjxQXHVwbfk/iRQb78Y7nF7zPpSgjzGeWSVs5FkLKc/yN1w94XlKZA
HB4rSky2iuso8NWBEIooSSGEKL4j7YwG3CMWVmaceA5JeclW5TtfGrsWWixMCTFVR4lFWayn4c96
ppBajcJ17lzPW3iVnLqvWI+0vz4s3lUbtGOC6iFZWUl2v84v/ikEdMs1sraMkpXEGjUIdR9CU2Lq
Ob8w9JJuTBdXFC11rxIiXAMBFC0gfmvK6eAElRdsmPDmIlExaTgaN1WWr7Ct+6Pn2iz4lVhSrEDN
JWMQ7mgTRnR7jhi258CXc+W8fbZNKaqdwt5KNPYH+H57U5z+oMvRRax7jUkSZNBd5mqtjiTxf49i
DOUyR+DrY0MAI89I97ocM3ohgTuXVQVMksdAMtDCH2tJS9n6saxuyRcNtkoxCJx8f1K6gYH9uLs3
1049aScfGvFJeTFy8MfKKe1o+zE3+13iUxr/uLhY8uZ/yK9Um0f5DP3Au2JYBuTcxhV87Xr0Hjv4
elintR2HwVEeB3lquxSu6cE4L27dELP1Q75/6Gr+k4+n6L/I2U0bWgMB5dr4nUH8nYsH/nMzZt/a
ZBk3xkBoWPPF2FPAAGEAkwuI8LP/AR2U3YlAhC8B3emIvWTGLC2T5IuQVI+sYTYWr1qNyIJMepFK
Wr3v8t2ZbJB8ZtJDzrVGwo3KlX8Q66qE+TE2c8g7sMg+XLtEqKpowzr8R277inOKea9JSbio+Ml1
WHHB8mwoenc0PVCUrOFmJDf0+hDZJaXpSBDiSOJY4xuuuuVRLrzr+kPDDzNGLwqLJ/UWDRUU66v5
m59gnVxpXHFzM+28zGNSmLJ12BOINVUEaME+nd0tIq0znVhUKtU2Aj9LY5Q+JvZ8oy9maiFy0RfB
9uvV315pmDDzAheqJxWAZKy0LknocRehUBSAyW3lpMPyPjeCT1zC6WfTeV+LntFkX7C/5MJbMJBW
d4kpanRkIT4YLXAuWrC8TdMycXf6o9qYU0hdmdJmV4mBL2UsBhTaPf/shr18vscizR3KLmaY/Sb1
DX3GlQAI5cZeb++bpY4RhTJXs0ACN03AO11uU473iWCyu9UJz1B+PMh1aHqGnrH8IizsjU403qc6
7Dtia4c54AikuM1lAKECN7rxNivzBfT1LS11PfbBM9Ev/7lDtPs8oytJbK+jp73cZ5OZ6fsFrqDm
f+PMzRoRgHWUpKnHw1oDRv261Jg5SBCQ3iknSyr3wqTLXHFEpwqExttFk1BJihC9H/a5fMg102Mx
X3pLJvTGAueemkBuU21eMzQzGdEwlJw2UIN4UXXHNYELNWys6nLfBHwynEoaPU91MSykkFaxDxSb
QLyf0diAcCrNUpUyxT9ntL1l4CM+ZqOc/U+gPoy8wpATmdgWrD3P+ED4M/QaEPJfKEexxe+nOJvs
5Up09RyDBZVQaHddcV/zov7KKtPycg3IUaJEO8okWx7l9H7LPsaaZSvvi7vtGis+xHkTaBqmdGme
FBlJWJQ2lFnsnFwK9vSvdo+LpDyJxBdvOsU5QQfuc7vioY60XJ2mHI0M7hboNOFV/S+WKeYUUkS+
kQRd48qIcfxmdQgFwQd5xTk0B2arqRs7PkurA4R4bGhZKoEQJnAgAmnN4Vy3jOXDEPrIsCCanWrs
44yL9vwFq2JuEumoL7S2koIQgbzimW+BIJEBf0A1uhGfr3PGBIHfhnOGIEAC1rzPaFwvE7vZqcKd
ptR96LvDu1MWLYIG/A/rTtmAQWh5lZPGdjcCVycUAiFaFcawtoJRogICdEn4k7mkHoDPy8OXd6xp
jnboc1O3G+2g5gy868EI5M5Da46Yk4AzlCH5tI8fOgdSUpEhOu9KJh01Lj8VfykeEbd1HQ/JiktU
MT+7AOselIwpNPqnGxJt/c443X85f45cRNq2AZj32Y9N0JMhJib5ljnX9z0qupoQyFPm8mKN78tZ
8Das96WuXja6sn4XA3QBZzDhk2sD5tBMbNLw1Usz0Ts0m7xRSJI7RxzjC+eNsQsH5KBVg6ubOqp1
Ct5D4I9TEmTaLETcCbi96e2m8EBHg+hQuDYUQ2+8073tyv7NKJ2jA2aRbjMTU5spMC8uXy+68ZDn
i2MTRxNYLIjalZlOecEir+LI+Niy0SGIi4MmDUsX1Scn0oK+Zzch9PLR1Jwlcjk2Iyr9LVsPv6h2
kYSwvwpeHBFdtT2XxFLI5m/Ea9RxxswTgpxSCznwhqGDwaDBLkxlZdE/9gTGsotkDLmByv63JKXN
VtSwujgP8zAldsSMgxv1mVPuJAz8ORi+qTVzK1dC7sQ1KO9SYmfajdIO2ObBB2O1t/080WJz4kjj
wXZysymoQ6A0sMacnSzlTYplyjFwEeuC+oZbhOJWaHk+aaF7adjyuYdWpZJ/mOQwquH4zks0V+ui
mwfQIPrBvnAELrV9ccHXMXGaQGqcQA+GowkGK1PCZVb6FqfkgUcePzDGWeGUuyNSTpSXQNYr8a35
RpQv+7eARVIuBYy1NaExCjnBXdi2C9nGY/izn89yDMKqHbu3AMPjTKibxjBEhNHoCvcYuRBYZC81
VkRfx0XLgt7qulT2KIobGEx9oUlGx0nIkQZadi9bXsegC5nbbpW8A/HrX2cbulYezMRB9lVFHcv1
NiFv+WfIrovEshazURdqAG7iXbagvI4Vv9ucTxmTq5lD9cy5sVI13RdRJen8TC8gBwh6r6rGmdjs
oXEcNGAp8jtLqm32RI8CwKzHS5BusEVDDFQA/weSfuWYujZWNkfRdpb61gFlmfKYagupLNe3QzJo
c9vw+u+C4eAW70W3gZ7w1KyNzbjihZOi84wZCJ64bXSBFqVSX3vJuSnfq21gqnId6o+SwC35YikT
HAUCdxyRVTswF1XGJZ67VmUuGbLi8J1AQwtmZ8fKsCoh7cK3IDa6UFNBUnePTIRFXuKCSwrDCMxk
fbGRSN4up1RDk9gziGJIQxLGr4dYLIzoFr1LQh+Vpgu1Rkmy8tPPCyL1tNgXw8xsl07zD6ttB7LU
GQBo9Iy/U4EeJMRAeasSYhKBdSbTH1KwDM7WrOUp+6Xb/BbUkQOdMzn9cslCBlFpTZModIB+1uO8
tStRKj3oAqLM/CXoxPs0+JXtCaYcv3cMIh+H2kINGzu9U0lRNzBbnW9KgWDqHGyjHdcs9y4BL369
RnI5XfZkQ7lasqJBfxZVRnJlClyB29rX083n/z1V8OjtQG3TfLhJXrf4HzhTDTSodxBADDT/uHwH
XrZ3ZWdIRhdFV4RKYW0l/hDJP4sZo7ZwPlh0Jbu12LFm/AWLo0ev5f7t4onUhRWcU//ooHKFwuq3
KLc4nMLgqjpbqbwqajCP0qhOUMDK/HaIXC+lDmxo1ZyfQwCbD69ud32EJFfmdm7w1PtxgsYqW56M
bTKpfeeFT4zgSh3E1R9hwbHd7kjcy1n5ehk/VhAtRFVCfrHGHHym/08ByTE1r7GcRoEPTIYKYcwv
TIIWAODE8EwfV+OD8up9HJSxlLmPppqZCUe+wqBruzIZVt8zUmjEZeNKcjhw1HFZ4UgdJqgfSHD2
/RK8Ny9umXRKDDeV52sDJK71+nG37Z1psHLjqV+geVPonTFSoR3gkFNSUiiHTeXhu0vxe4TRw9cl
yE0/lC48pit5XKCU1fCUaJ0HE3KpXgTKej/exidoeBJHF0ndcUKMGTbk+0dxZXbhUNT7Wbj+MbdK
W12X0gG6YW8ISgLgBII19RqaG/TcxTvJnYZETPbnuTXPEgtkX41Itte1pdZwlIaQFSPWF6FY5ga+
2I0OH3XEf3pHO9dlpbB/qUQ81QIBw4iaZgLt4d7ud6RVgQ+vcFX0QPkjdYMS4608sE/jqLGq5RC4
JZoo+FXyBgtjlkc2wYDN5xAvtiq9aZ00SWVJDXIOCtaAP12tvFuYWYlVaBdpfb4D+/MG/rIikzDt
eyCYNf/nWlh3nrk4cFCp2CVbtlasrt7io6WasA2mYhxAWaqdUPOiuSglJBywfYj94PqSWbrX9C+G
vUe8euKauUQgQsBiaPHwz63YHIbTZDSBriN2i3lAJrLMsoGLtwJM93gGHPJ8gyiL/7jt8HtEOfre
iC4z9sZqS9nse3bTzOLVyk5SP+nidGQQVpKe/cLzlG6arP/ohKG571FcMXpSZILQH1L4zCauDqAn
K3cIpyG2LlV6LEsMGWTp4RvLzdiPC1v++OMIZb/vMkpibgGFog3ozkQElGNpbQRPU95PMGSH6T+S
Kva3YyvCZrN6t4ONEN4sB5OTA5EiiTMW6jd4OOlcCoQNTdxs5mqUNPF0gG1x2Od7Y4/uiuwfIhSb
UVEqegZyiHYsKAhpwCaPGdX3pRNWFo8mox1gjpMXvgCm9stE6CAgHuTfVUbIPA+oUeql6Y9f27Ss
xBgrRnoNV2s+VPzhWImajSjiEvccUarqlieXjpnso8A0fs4IyEBRMjit9uoXGLOXq1mQ1nI8H7wG
Z/MKBIGdkxzjsY8Q5Lawzy8fyhYig0XNE2FJpxiWj0odAgdpn3UB/YRFb/tuOhuZ1rm86WWrPZ7K
zfxIjeIQdjbAUkl1EQFtnOQHVSdtfTc/FiJUeLZqqF+YOkclBGtY0ptshMUKsKTrrW83K+7vq/pT
xLTW1RnaB7b/arOLoRfRg58JH2+drM795hYPJTKPHUT5xdbGljApsRkETNdOVYqSzOs1hNoxMgrm
hANogl63UBU/w5iAQM9EmWgXn6qpZQzHJ9hcOMadowGEfn2AHrEcf1Z0GGC6C0jGjesOJO574bgK
Bn/cD017xKtiiqCU/UiYaFgRukUIQTKM6D/QGuFtiuvjp66F/ZNP2Ak3yBiuEph1CyDCxD1pKrUQ
7bwfykADEFUGFnazv2kYfNyEj/Ou4u7tbWd8G97Pn3j8yeEsP7AtYKcRVdumZG/Qf8DyJ8WRhI0i
M7f58XTE5cDL1Y4ycNXw4+vmshfPGC/u0N33gSA4WWBeff01KVvAh8kiitNw4R66qcsgQHC+2Cgn
LGDTB3fP/lsE8SbO6RPMS0Pi6TvLC2kdNz6lSCrTtyHrdHwLtjExeGbso3TBp41mTv/ABzISbeNM
3XnvKN9vRLxOnpJ6uMrYmR2bZmbud/DAMqmAmXmIHvVQkQVkq5MuY9/QKYf+c4NX3ZtFwK5MF4Wr
oBPmQmIwikH8TOlOqCTwEv0LSOip0D8Qppxk5GJ1H9JgD5a6bJNz6lMMWAjGqNi3rCJLAKbobLom
q+ZRDf/IggWyZSZT7kmLzSQoCpypERx9Mi4QssIktKZGmji/FONvU5rJLGw6iyFBWJKpP2GOStVo
jN31kKiNs9ozB3vYJ2PvSQxF8luERFaTMU6EqLz06D4peNWI6v49cJHWLbZySH5enGRdP/jtqER9
YrKoDb64YJW93QcSW5+8QnEqCsGRQILrsmTfYfA0jP6yzcO3fONdqGnUPd8pCoyrlzqHY04iUMU+
d+wLGaNrxbXegKDKepWGEk79AWyylen9JmRhWDUertTdxtOIrz8vclcx3yLs6sDPqhYRrGO7ISk6
46tIpqMVzwRzJCR7K9s20MLtLB7jMbfHvZe8VhJNgGJigsd1HrCi35G70eNtOO7XP6vwhcOVRovV
J3RWsHkHIMIakF2mroaahM7QfFQWbM2T1U/lD65HB+yc5oxPB87FVf5CyESFCxJp5GYPMBYuW6Yr
az/P+Rpd14BTwvd6/XV5vOrlU4KZjH9uWEi0fGvIhV3ed4wvsKFSQPKmfTfDvvdywgZuPXl5JVDJ
RsyUJGyiDklHuII6TIYXYA8vzBHEu11jdHzLbjeCrMsXb4iWUfvzdpGalQey0kaRbI9lTSWX0GHq
plM4nhR1ClZeoinBJtW36BD5LCSNeCkMS8uQJc+jSdd3YPbgpSsedRio4o9t41LpGziWUBeAvgCm
Va8zupJUeWsgvGo78cQWFc4yv076d6QbovkEZDVsDFkasiSBUpvBmnU6+NjI25PiO2zp1dERUG0r
NoVqbwDrKxwKdBpSI0qpfbmKjQGFDJj07Q5LwtJR+ZbVDGJeF/zkv3opvDI2t3POpBJLk6q/p7yq
b4+aiIeocHcruN/rKuauqjhXrOX2Z+VBAJXKFK/2H3vRjiBWUoqMH4isTCj46SoMr6TQvJQ9cdOn
kmipl6OQO9RnDr5zOH0MJ3XduFrQ8XuVbU6+cOhYKZLYMqdND+P6WOZnuoZo+128ByqTR4qoshen
8PqhYvkd63SSxwrUVWBHHvxEmW8DAlaNop61CIa5kJwT/Xa8yRxzKiasbbagJ8ikbqotaLHGUng3
/1Z3/4bkc6rrJAIxVfbKk587P9cIRHf033ZKbW6bijYiUxW55m4VQgejr0AfMp1J1dn8LSrRXYO+
Wg95uQNZrgj3kAz4N+fVDv8JI8TlAUA1vE+Kqb3I2oom8dbVjTwQAFZ3rETQu2L5Pqfmq3/9D73z
bo670J1m3tszNp+nxoLC+cxjxGT5QrC6KI6FVM/vxOlQ9QajBbF1Jo2RDozqsStoRrdqarZzR64Z
kPx4ktVd4RGj/rb5KcgPzcCLRPxnGt/+Zx6lbtNyKC1jcHH9ryYf1UEAkiXbkjfSuwLqLzYv/4cO
wBYR68PXRco8vn1jIuAj6iNQuKtgKH4Jv8h/9sDMbddlhEusVIy2LQrRWsDfkhZYO5uV5/w/nDTj
wZI+FKIVwXT5TeU+ysmCy8C3BrD207dDzt9lBBueTTA5a7ycHPTJ92MX1XZpVhFhuUP3Ipv+ZB2M
GMg09Br6822gk3s7M16gQ8HIeb2bH616LQPhCRN/UL0zAcrEHOLkqEvAK10Dzck7vgA8iNeOzt/t
gol08UHU8Tb0WIRd1R2ewaC//vFRGZGCK0+l8QY+uqiUxg9r5AsFwL9B669TqhI3uszX6IUx8gyf
YduX3KYmlFkv9QZacMiiwXXFOKXeMO+u97BfTv88chUcltwWeLxUNdOMK/z45GrHNYzDrxVqHkut
2uqftMkF5tsZ2UO8h2ZqQt6iQeyuqMj2M4HbVrv7GGospIeKp9fXdpyaE7UrJEQd9l4z436SfYY0
dY0wGorizIUuOI8cP4utVx5ZU+jD0eqf+acnanjGttHzEHfBX5Y8EI/rFdhfhxTVcS6HolMJg4j5
1GWsBRr7buVXKJxvleJyoDu9ApYvH1aYYSW1nbL1aGGjA20Zj+y6wIzooUDpvfDJjjPwpnjbqmEu
QYmPdk2UbpPNg5RLkLLeYqKjOO0a4zaKg38bkwnierRI5EVpRKaBjSPe5VjpHmU282z1QdlaTId/
XntbkUaKi7J1kQt+cT4Y79fuAS0bcZKfUmVPqrrfEYuYqPtb+dy43DxbUPbqHUqZuQaux8wTv1cz
3MroFtS9UI+9jiuskfrnTNNhqjYRTR/Us+zFSBklBFegK25GCsE9z/XungT16soRoOvOh6PE26mF
NKxwI+qVmsVufHdbxZ67uzv6zEoo1TbdA2z7bqlCPMOQabtgMdsmDrD3oimazhJK2HunqGesvuYU
LLoEnQjmRbf+U/AfNbxOFw4LZBaM4ohZJdKrQ3xxFNxEdl8Z/4sKnqkBM8OP/8aKaZjcheQ3cGng
dRfXafU71Ldm8nlx5XxKQFwmmflG4KDoXfpy3Gm4S6hd+MfRMmWLwZS8DQN8t2wpZKnoF0YWw2/0
gc0jp2JsTWg0vemeDpxxdJXStpFkT3UuiQ+Af/maZHZ4uIkEXcrVZkzQyLeMuJGeZPoOtWfyZZ4o
WSW9pl5lpeDmpaG1lVFauUhR0wgueh8LXj3pVMZe7u9ESmVdu9pObDQPjC6Ww0jtn8tozLa+ztOG
cZlp7ZftEPC/YBLLiQOkYRFl59SDijE23KF/3bSwolXzjlcKJy8KdQETwA3zkQhYmg1HJQK4To52
K7GtT0fhcBlogPGDECcNG8q8a0S79afYHIDYmaFhxwnXLWGI5SaHVh/YZfT2x9gqKemoh8geMO1i
CEpiyBcI9xZI4tFHpQfsg7tP90EYZu+31sp77Y/owAKB0PnLiOH/n+MXpqwa+ZpkwtCZs8XkP/ga
SQelDPPl00TY8nQ2UciA+GiOGVO8jGj7We9DpKzQFU787c0ATTc5J9JpjqsD9SzjOrcUNXqillBU
OoHfwDhy7lOQMzsBN0VKUYa4H+XHOnKnzgEFzT2vGQwwy1DLcRgNL9F83kNrnhN/weO2Ju6bGTV9
sR6K8BWwuCxVAyKARZ8ULLg1I2pIOBWqRcqcx8xPdkd+DcqdCpVWU4HjztlDZ6vFHQm2BRzjpbZZ
WZIBlBNrmRTaGyXMXxhsF1pD+5SXC6YEc7gkX1Vu0Sl8gscu/0X+5IahXy+6hNVZAejjtcqMRNXi
SyPdAGFGknlhkpVF2l4+2aRT+8Lths1GAKcxekv8RlD5jL/yIKsqU+NunDSZBtSD2x1IhaYwRPNv
T90fdcGNTue71B8lvkuOWHiJZru4yd9C1XN1e2l/FXb4gnzqv2oGM6mQZF2lHJGdlEpxZ1dl/Qgx
88LYXYZGeGWsum1vdy92OKjwdrXaKJwBhcUpVG/QfmgdOHgfHXfGdAtI5UaKMKmLGZ0dlzjK2kZ/
fOsifLNzkmv9dqq/XcbYRfhUAvoiEDSYJUURnMaaDZlfE2A5gok7SSJlm9FPHOvUkKkG1V14AYZK
Q5TiTT6H76bLjDV6IWTrRxHPzOBrfgU06mTPKuuvepjJWppoiJKjEoa7VX+A4Eyl2jwzMvuZE5S7
HNQj3soPRM5qDQGJT6rQNqYQXF3kWYYRBhbz+nOFKgMhRxKpiLoWBAif4YdXdQ4GJIo2pebDQ4w7
l+1yR7wPo6NP9QSK7RiTyP5MjB9b+RWrGH29gBWjAjvljfNRIq6cO1LJeE6M1inz2bkVuNfu/oHG
YwxIJgFXPnPz0caCsYU9C8+RPLhRC8Fwgj0v+OOGVfIzk4Tzb0dCQ0fkIudO/EoOZrSMEXjPn8wL
/APd4EMv54ZnnndhmRJb1MeQwRRovBZXe6jrIMAA3WpyhzWnU4qAjm+g6q0VyPjGgBIowq1FRizo
XbVxvo0GtkxJSTCqMN8/ntIDyw3SOfbP8MaAFYyWLt2s/hu2a32DQ3kjb1hZauwCfcLQKm4QHUqm
po79QPEITW/Bkyw4EDeEO6deeEmC9/zZB5oXxOq9e9IUNZshfkdXMJRdgjpdXpjzdtvBbjg+agfG
QJfWn7sFCKPYZ0MzE2HrKormYAfd3qikgc20n86o6Kr8waJcjFkbqvkujD4jwYenavaTCUvHlDtE
9VSB/N/zmmvrjt0ksa03zrj/HzVwxZ15bqr4+QEVNzRrevvoxDZX/CBAOswW6Q9XN0Pw6tQXs0px
OumG08vZmYJw80YDwVwmTpN9jk15z1uZgu90lvtpKkI3ysg9Krnc0zplAyy+zzt77K9hVc7UpAHA
xJ3L9D7pi4XUt72KLmL+2STUt51TxcRcHuaKw9GI+1xKaaxN5GJzdxVtLBK/UxHqbq0HR/ZiQ/6B
1JEZ9Bi2/Ghw4OWdafx7SrlKoWcPgNn5skUrGUXUP/mwRFHURBlD7/V9LoJophwQUKKhZAL1pDhw
9jGXr0AQ62jOJ31jrpooCTwBYKwy6c0eZohfkAGtlSjlAZ1178nUBkkErbRGZt3qIR9EMA+seTQU
TGQGf7FtfjnycP3am509BRZIxY38OAX45o5evgL1p5UKkZbDPyaJC0pP0vveHlYRjnQBywFkZjU3
O5YtCVRB4iY45PPgJgNtHOB7XMYKJcR7gdiKTCjriLE68zCS3aaNrlRORzUluwD9K80BF991hC6C
n/Alm+YDjU3XtdiYx2tVh7Rk7HoCuMZotMbdizwym/5a0QQTIk9b2mCftrdIVQ9MNw83GtZgHmcb
20RwQWElcRYF/t8zvYAdcDDr2CMq08D8W6aiBO/rTd89nOxt1JwItQSKCGCpvOJ1ln41FvmLJjkh
VTCXWwbebZaksBgC8/yoGXpXL8s9jATHOXNqQ2Ah5EaZJzynqyc38aJJBsr2lJHmXy1BNYHLjsML
H9AVTO9L9T+Pg87TX3zEeTiJj2TFtA/hCJYCWpYPVwvF3QXnrAY0a7NYyoevN2gj2iU4F5dwiaJz
9fMJzPRmsZZj7oRR4IrAV3xaf0y9d0xI90o9Qe94+XgFZYB9yQ9qJMIfA7tMeTMn13ntcABLfZDK
KBhWaTVn8ULW/X2ejb3Gwf2ovffaLEEGj9DjBhz9PJ1jvI/Mr0HVw8M7Z1vXoDoXk3xbqYhW6GJ5
Lm5+XyGSLLkGM/x02zsnVukKHNrjltt2XFFbaSAffrYN5LBHPcQ4e7F32CmNcvpqCNW8tLFYAMUU
FWPmMYpH7FQUCCX1elRqcvf/uSbM5jiVmC2XXgm8yR3zFvjLS9QjAT2nPceFPIcZy/lllRxRzjfp
A0GpvV3KzpaQ3eZgXMtuVuDqXVWGGm5lyXj5vA5OoWwcD5oIWYWZkCZo/c7ZeBCRGFMpJv7qUuEa
NewzymT+tD5o27BMSIC9MJYh8YezEj6ATyRj4xgLGkAqgp8YKva8Nf6nc9pl4jjL1dX7SmGIoCZ1
mhs/bcwtztrYOYfGKsMJLLV0BTR4Vb8Z34ANoUj1J6Le22GTkPyz8iZjMEeupmkCuJkoVyi8cUr1
maYdZPSTcjTcBNIUOg4LBQcxrKnSztyqfft49iPHsh05vi9t2GR5BPjf8rDp02M0nlyy0KuQ7mW7
/N527zhTQvj+GiYFDYDg67liM+/eZDGhUsZXAQsnFeuRHXOH7MAjij2MZwc18l4+tj83MiyQ/68N
NY3uhCIsVeJxMf4gAHO6A77GD/uyPUSmi/FLFgBfryUiJMNyiRscMK1o2ObUA+DTxpi5s0nGki9B
qhqpIP6IhB7nqGbTi04OKuCMfsEuEcNPWVI8DAbh29xkndnSpna6nzO+hDZQ16RrqTRdGQS/sLbK
V8Yjjcrk53nH6XKAdFTCXJRch9bsoMFeNF+Ae03DkBEtNu/MVQU0o6Wzwr7mKgNPSim75n1EgmJr
epmbzp1TgW6BSrt+9rcvMdVsKTaIBFlwrjIt3tqDOc1wW+0CyObU5E3zEEM0zk9B8e6bsmO8m15k
hUUX3pTWoCbs+/NtXSVX/SyMv0zA/Lq/sXgjz1MkAuap/ZrO9uvhATg/fdnpFl5QzX7OIAl85ulI
ucKtI7ftjoGoXKp6Ad6bIvgCWRqBDuylkeCZtDdrSGgHveKh5RM+0NCHhyaMYl2Ml/CYb2wh/Hpu
Sy+3bVjNeJoH4VeJRoAD2zqxbcDwhzL0NEzIMwQ5RbkoupZdl0Di5o7vpXVH2Xsm6TDsPDSP/FEa
n2yi3i7Z2oCXb/E+Wn6YsNAyFWh21xuQHP697JFqOo0+PHGSzSHvNjQO5g3d/9lkVXa1aZL7wtWz
MZTNEOXhgYvtjtxLx76bkLpR12+q4y1KOF9n+C3I3G7xRNYPLVYZBrEWn7t+/UHpoTU7IIYEA9+1
xb8jUMJk67ZndJpeZTeFX7MW++Td8j6wrie33bfVz4+McNTr+5CnbA98fuqNB+r2Tt9RhgsQnvOo
6vULXfop2+rQHF8DAx5z3RpcpG22vBQtl6zv5uEzGVF/PmIOjaYbh0h7j2Yn4HP9HenliH+kztny
y4j95VeGyj8pWwpQqIEaWid/oi2GzMkLcnS3LVaDoVT68TdG8OMYQn6jCB6KIwaR8rb1OMxL/6Qb
8S6WmNCUXTZTqlOl7q6UKrhekSL8pqf8EnRk6NnhJDbA3CqWmdwZN1LcJdq0VK4UoQKe95f75Y1B
hSjNOaatycC1L+dsIRDWxS0zCK6mx++gY5P0nqs2g9RK7ndD0XbazWcyoG9TCH2TbUff7DhK/CYu
gvNYZYGRhmB0TswTV/fCcBMDHiuz2U45usamxy0mPHWs57wkYtRyGtBMr/jcoZ5nGpNX9Y4kFdyx
Z7KpJ/J0/Wv1ntNbcVGlddl/bwYjycjdiMBsJYPC3zrmII11wJUV4tbIY9N3Ncub3NmdeRVzNkw0
4LDhBTiDwsVnB9et6A04J0TkG6xykrlhCycpWxfMGwK0eTXFBqhYEd3XfBmUXodEitDak+lsUVZY
g8jzY2kGe1Q91LRHnUj6+CoOEP2+xc2gXy1oWcwkuQsF78Ah7qUnyt9y8wrXctSB+PGnJsCTSSS1
oMyWEVXljpiDdO2/cYpyaMsnhAR6yXXOIO2qGemd5drRe1QPgEeXaKY+B6V+rOjoPLIn1tU+EjBM
CJnkmw6XdK4B82okBdUOBzK406LJ9KXZm76bMLup69y+toM0HVuAaYcdIOz1yJv9kjPBC/yRRLRj
Iola5Dpzf9jkCCNNLGfuC6gTSmG4j4HKXRFpBEOh9GjQ+G4yzGCPFHErRsVBaqlu5JfbNMfOlEQj
FyU5ne4ZA/ZL9A1J3e/IsiJXfFJ+bN4ZSZd+4gSWdM3eFxC7dZYlFnrPn7VTMhAHyuGkklYjBi+3
uCcdlwspOTuxv1X7b2OXfT9x/LxKQUDGWauVwcELwE8Ff1tKAOCllNUX+iMyTPd6vC1JSZIcIXBw
2zbJ9+AnqCZaaEZv2TalIwiFPgzfapV2/2+OW77Bg+KpXK5hXVlQI+m1yXNM+wIkdvpC/d/Or7p6
DaDG+fZNMeqtzlAYJTlLrimG5WXoHRn/zXL9yCKq957dvGPECmM9A65/xiIV5GBc5XfmQDriX1HY
viRcGcungZdVAsCw7YgKcJVwOjcp+AM7R6lLsae8wcoggM6WiqHF+ST3rLGkleRLY7KUEp8A+i6b
rNV+eqGUAmeeFYlVAeFZBM8hJU/4DPI9Pvlim2TxChcPFQXXgd8sIy71H/zybC7S4MDUfmKcT2aO
DDcNc8ZZFL0C88E1V22ELHA0FDufiYA2q95crw0CIvWnLvtm6+vhO32fgyBCGXF3ZegUdwa5NWkr
1s9OHlyzYJaIgnyEMPldM+r2Yar262LUqnafdeqVQJwNfY6eVqm/XwlzBnVgNXh/v1+OiFxQg2b4
0IFjHbnRhamFITU///8YP6MHvOBAtguLTvBwR59pR+mDtw0w39YfBye5I7k4xLT+L0olZChjfheF
HcPPq8wyRThI58r05GxSah0L2qDdE7ghFMyj2o4IlCQnw3JqExPkx6heGW9+9tSt1lLKHvh72H1Z
f9ob//0MO669/bL/IsMtjwjHjFsb3SiKDZ3R9TSgQ0LdXZ0BgX0Pfko64i2aZBkUgZmrfYNhNdGw
JCjhZsSQVBYMfTv7d5OJwpi2dVXAoQj9bXRXOG4y6/pTpocd9O3MOZ6PQGV+08/EU1KrppEuWVEd
4xeeoKF+dlFJdRZnImSCvZiqRukCBqvz5rc77DLeeepnHET+CXLiLDFdpxO1IGFo972GQvqc+lhD
apVOXxPO4YNn2DYvu3PwLXZEo3juRDes0Qs7sH9tSpeG9BT6BOnyjU0nz9DcSLYT9d1ihR6h2jES
CS/IWAKdk+NnIdsJcH7R8VdTTPLsGAjN+IhCe5RCpVireWz3SaPEOf38hbvEjZioBty+eP3+xNEx
x3SY6gm01Pdp+xrfG55w/Tw1sPoreFx5wIB9m9OEbPmL1FkF+/MVdq18wzao+HY6yFKZWjyB+sFo
FZ0sbmFQy2W+nNL6FU+Y4WJbVdZHXXC95VkzjEjmDSrudj08ibI5TgoCqY5uAM7zfL4+XwItl2NT
DWl/5zoQpdKUA7FP+jxOVa41JqkkdEsQKwHvE+kXX20IxxvOzQ0a8gzhSJebiTP0pGoLGwdlvYuu
jQuRJXVy/aOBPnb2z0wgOK/sl4q9Z8KgILcOdtaFSLckxzLNIrP5ToVzdolT0NNXXbnPZzVLC6c/
/yXW6IuG8ZWS6HuLKgFg/8XdgZZDJG+EDoXhlkqQ2jA8Il++XeOxVDeKr1StZOimPlEyZSt7tph5
Wkvq+yASM1gw8Vqgx7aNSZY6MyJkexhco3QqPTTCAhm+dFJmSYJ+eVeU7SLATgAZ01rZbs6FBFGH
55suE7YeG41vFg+RF0ldWVQuzgZfB+6pRVlWxh8NMNrZlPviR6LtCdxlGs4RuoBtbmOXTYrUREcB
Ra9TPARyFT8dB7HfHTuS9YsCd8q0ibd/JXeykPBeIxsunkRAa15IDckf8BwuUp+DFzPHVbjCZxFH
Vfv4pLC92CEycK+rPPPymh46tW1uHOF/h2zADRroWGRYLhFTJHRcmcDM0s8+4WTL1eyhdOHxB5zF
c/uGxY41idjqIbtsoQz2hv/DW7YP/o5gfWI2ABggeFpINgNP2WMuTC9Xx160Q2JOKwuaHG4gc44S
PVMhhGG7fyA94RL7eA8x73PTvusnYPspMwDIALy0euw7B4H8mBhFMGBI5Rdd6dD4MBSgPUqA3i0U
1SCuVyqLOltFjIqJjv0unpixicBs1aowc1Nw+xrkrXOHizV23Z0zrcATzNgRtToS923Ek9ZTWsYa
oN5Pm9//V+XP/eIewLlvNuOY9whnFenlCHi/SIgVKNoo8WcYc0mV7GwWD3g3sWzkHvfcvracIdnX
uS6SkmE0NU+WDRgAOhd3+VwzzmP09gd23E1FfpcHasYndqxaGUplCd7jZzfrskwqlKmgTc8+pV+T
kCmQTxH+3/+6sqpSN5T7Oh5fzUjZboX+3QuptcG6hO73A8qHmyC7uAfhKSVFXOZgUBFN8pOvL1dE
JOVSKpVJ1czFvX79dxayyLRbPSu5P+nS0jvfb7Jkd4aicUuaPkMVzJ4Vgon6t+2/CaFtJZOL8XnU
XxzrG9TY0sOMrCa7sx0s1wkrwNFTnAqr04V1NEw8tDgmQ1ocJ+wJdjjKxQE9T8z20VDKxKJXeEvB
fRm1tMzwp1puGW1uDPZdH0bTQayIYcuWD2Us2VxxZQ/vt3uzeaQQcg7qQRXrAX+YbqGtBxqz446b
Pd0sH2SWNL+Np+k7UpPVWJRWjYUtjXpsjMPF+f8wFjzBJ1UsZuJwNn4Fq6nMd65bLfuPGqLqFQ3G
Gl3HnvjjUkQooxjOdoDpOinPAHCLyluMkLRmFGsHdTJ0ix5eTGln2x/RNjJNO9eC9Mq5RogGMjdh
BXXgenfFuB+BkJUd0yrCDBL//LBGXJfXjBKU+CMLE6WMAVXFuLbVCPrK6OqMmc2X7NxmT3QW6ES4
dCmtKVHOFm6I14JoC2qDTVJl1ltmFUn/pLeUf1USy4ooZAAjBwT1MxeyBgXChAuhafV2BO6d8xcW
N0EhxNHvi1BXb3kOociXq1XcY+OLi7qAboW4qPCKdb06eJEZXt9CPtu0RlcU6j6kzDNIw52U3Gs2
moDTX1oSannpGg+mAkWUTIKCVccQTirbA8oEVB5v/6ckQPGWtYxOsasThbjgck1VKaeD+ELHON6O
uLo5Etfuwm/V7BrookqM0XRb7eavqztTPReDYL5j2kCn9Gg3LURxHzsRBJ5VE9WTzOujEmdl4rYq
u+GAKSf4J+jtfa1gmtmqdgZCQezuuchlaIls5JiIV53OqGr5mwNolcfGxhgRkUgf7enexME98ZKj
bUuhhmmhPXf+Q2+lpgp/28AMKqfcvONm3YrGwMywjDwMRwoofaJEfxpTTg/XskD5rkWVMKMirl6e
zrENeVXVAAbSQVsPveG73W7VvJKi9DQNOq5z5rHkvWL1ll30Dt1BQLpJ+GQ8W+5gL/7bfq0muQIP
jluZ8LcHqGZDYfUfVNQ9v2Xv04/Y4a7qjwO7MaFDBDG/5Ef2XlePnMN+U5YGbaNIj/4mB9Wc8evC
wVwZu9uZ7V/CgESLtQRjQK9pCOsfAG5czLXE6+xTdQwGaeu93jDZdQ4CZv7i3+UG6nvfv7S091dy
W6B+tWbiR2puKkbrPJEjfIgi+MhTYIyheUxHBjw0l16R9X0KTj/gta/++77bnK5Ita5la+uXNSqL
GJ4G76EfWEUEJhQK2nfa/A5rjpV+kJfXNaW+uRWQV14rk025+7QLNGyWhrKGIkQBhFTpxGI2/Yvm
w/9iUWoIWKCuvQmgk+hoCHlGxS/CfOgJo/m2N7bGVmnJRII6GSm8KzD9tbTJT6evMbIK+bWFwjeN
iE+rFpGXnYg6Tcfo4CCtEG4TZ1im+iCDtlxMLtCUiKSc0gEqQIGJnJQ8m+11Us27DyTeRdWga4/R
Fu6q7kRibqpCjuohSKB4/lwzxxjHgA2zwOwtkHWm55IbVppWhnv7XJXdbLD5rXZk7+9u1B4eCFH/
YYCiBVzWLaCinPM9bb28PiXmlAC5jY6FbN8dsa0OnsZspjFNqza0dKI172YtHUTzQNfCgUqYHhCb
gvnQc1oMlNdBFPx5aV0qsiOw0vQinXjDrihhUwIt/G3Rdn1Z6P3vDJblF6wu8YEiSJDEJqiq0dhU
XS/WOU/hA3V6fzn8Hm3elOQlEQ56J+JlFEIYHZJuD+P3wtqwj91NDB+ck9rsa9PsBU0EI+PJQ6Hz
VhMrU5/RxraQhdPqF3SMy3wFB770kkFz9cSwIJ+vWhDpET/1NMsZlg0UkJcyMrXSRut+i+zRBaJL
nTtGrj2ehkUcjVeVl6N7OhcJX+GGEcco2in18D/e4r6/zgEtiUEoBSniOXK5ewe8nQml+kfLeFsI
+XzobrKJhmbpSqx7s2eqdhfdgPhq4ypKE2TqzYRDXZR5MUDPMCqLqvFApZrAAxzvmlFUJ2h//Uxs
m0E9I8IuzsdPDhmnBiQ5giB24J8rzZWF3PjhxVCgbV+W3H+/RsKTYn1Da0vmMUw91u6HR6ANNwno
Sx68Qycws1dDk5S7QrNZnCVXxIX8xFzwWE3u/AKpSBCle7DFbhQouBBNxDpN0k2pE0bZihUfHsLY
NFqiDeoluaEdWnSIlgqiosy/41h1aYXRsY0cwZt5oEk9jvAWsvxADDex87gM6RZjxbGAmzvpxrx1
IKIT/IlG/70hTY64RBCDRraGZSyFXhWdM06Rixk98I3J+A0AAlccLme1hiF5oUFiEIDfGVH7h/84
SQdCpJWbVi0jq37D7RfR4us2KHyw1wo+1dAml5CYZUhzYEb+5PfG9wk+qTNQfUAuMs0xmDCDovuP
bljDkoJP+uyfEEHd/cwgQSF+UCCrzGiSddPGtYkXZEJx0g20YCItWLLrpbUP3k9LoYKq7tI3QbNH
1ax2yeR7Ftu4EpyigHn6xidA26VUNDoI9R9acZ1me3iSDZKrdcl5s6Ki/w70VsjCl84YLdrrhDge
SDT1US4STTwrgO3Ks8R+6WPV9KJVCApHdSLgjtuMOAPjRNjcwkI15L2olvlyeX0eNR7cj8sYnXTg
df1/kpU8XXggLPQmboVh7vvASxpFLl3Yt4sEf+B4C4gxMGrG9GKqhHgSWTOcx6azsvYxwRFz3xOc
gwrTELnp1PMCNZwn8uAA3a0VBBfJ5+DM8UP0KryrIo6sFqa4mGJuVfI+JU9gA7DFeuNy1zQVNiiw
VOaNxkc5vF2ZOpOe99IED9MM8+3vc2GfFCMMDJOs+hOUwHyYVqFAc4SUWI2p9NxpNEojIqZBT6qE
zeCChD96MeOZekvI33JTXJIP6SjSIU+ASb7acZnKGc1JHTgZBzzAmKmSG1K7YlGbFWczId6S0qQb
+8TMrxrZQ4onG1CqjRTSyr9+2sIwoDr5OEJ7pZ+ULXXdbPu/+Y/1QMis9N68ektvFR2Cz0uTtMxi
6YAmub3acoUI4LZQr/j0V//lYTumBQhuTy3M0GqM1Q1cqlE8ctx93PTDJBC7EUBMMok8ykEtRTDA
tC1bUKo1W9xzKRbv5HF+BtBdDU8xumBFbWa0w0hc6KHxcmuGgNitJr7Ffvy8KXc9RMZHWYwHjU3j
OTjeJOE9N6ugFa100j6E6Gwb+iYD1uPSbBp6uEODgcRX9UWnj7fwidOBdei8hZAmMhgszFg2gu/N
Q3zJuNlTAQywCFTAW43/4r7r1LFV6kR8WNKI6RDlSOPSveIqqiJY9pBpGhExgeOGd+yUDC6LHXGu
6TP18qgiCKhsGYfrVbeDtKKt8sMVJIXUAfUeRBUlEonxeoHGIp9PUtC35uZY2eq5i5AXrXzncL5p
P34mOoJB88MeULKR8eMqC8+4Vz4AsiJ4Y0kRHf+xNnoiCRFrIShZqxoGuwFRqxLQwHLPFsHqSVpo
L0nDwFtYCP9X2Cb1jaVBiCZ5/duq75KcuHj+BmeOEBgNLkgDsYZ2qyTWNDwLMa0HEc8JaUmHGLH9
zh1yXa9j/1OnLk4bt5klV1NvP6cwmXX6GxynM1Dv2pOn6wvAo7HB+FI76uJTFCnBRB1U0XCsZrnm
zbP4RArimi3y5G9GtWaPWSBAw4Q6Zi+kKWIPrO2xif7DHkXNFOSerRRiTdtNXEDkHUl4uDw0b6Iu
L8wFBm/sM520W0PPulldySz8fpBIws8p81emcT3UgxxcDBeN8HumSPCoNIVhOymYhKu2o7WqJg0o
o9Xtt7bYcyIFzowy/AGcwwDf5/RuHZQHLOU0D68cfyIiPnlEXDaYZlLavGjapfzBf+BluA8EE+RM
dMIekJkTxIKDtdBj784JdwhCq0UOKFstEoiNGx0wgZ8JP1lI4JPFL1rk5dL/ssDecKE4wTG3IFKo
MpFPD/aHX3wBbxpps5eQpwpKyxnrVu7sgXGz5X8/aKaIz7L60sNqvyGb9C1QiQ3/mMhl/Oo7QzDC
pE/hrxehLxLjBu9uq/Dw/VmktFLiwRzmatG8Q02rSn4+27Ggrj5nyGu/R1sWMqWgZwG70X0i8Ce8
8OfZBMIAtvh8NOUxidg6XjBamr6Gy/7rfhD1MmQs+8Ii9byGKLEsLDAz4uqdAQ71MeaOTk93tKMG
AYmlw6wJoXIaMqhAV3RCPUU3mPOqHv8IbydmKwM+J41EReDNdaNxfF0kj5XO/dVhDfpb2A99YC2/
3mwr66/XwqmeWtApXHtNu/wwcOBVGJPc1d0zIQDLIUk5HGWpm8bGF1XAF/Lknak4LZZ1G/8tYkUp
VyuYMnrZ+SwT80NkRLexQbmNJRFGlSwRsPNS3HoARZ/DBKdENW0+TPP2B4lQnT9ZFGQANp+ryr0J
kmRvCaKewce6mBccjKXszoPZh5us2B/xQ3QscWdE6p1eoOnBibs6Qdz5dzRtKKdTf1fxmsYRrril
6ALC0VdYvh7yeJ0Fe3EiGe93Rjhfeft5x2QpolqGmbUc76qf1wzy7D47agaWvjAiNJD1R6KqHkRT
19lV5s4duYA3BEw2WAY6B7SyKKZy/6Vlyq2Lol4BLDfl5k/Y9ZE/i83R+LHRjeLNCuJCITxXwml/
gXe4emLTk7b2AMC57eGHVr12QGT2SD0ESaVDgD0e+AiKDXu77pvHCQuGbUQvolDscht90LiYJ2FK
A7pfUSWct8XdN88HArL28zj+G51HoeY4xzf1c0Ar4buPbgZuAbdQmjA/cyBxCUvP/X48QTX2kyrD
HX8n0H3MBk5bryjDGWTMZ/zXIp0+c+aPhwqv+Ih2gjvO2Ua6ant4LsgoustoCUxiFnbe2niqqHJz
J82jYG4dOUJvGHhhGGsr8WWf1A5TXOunlZbQYjQ9YhMW60KFvTDzvN1vXRVBkuSvGIur1lVK4JFI
s4Qa5mTNbd+oz9Ozht5WxAWNygrhE0zSTu7IG6HUiuuCCkNlxW5IwURX5ccaLXakcOolWQxkf8c/
J/5ZPxKgE0GLyxCZHYA1j//x6Tt7le/plLFbb5R07SN/qx81HuA1+5oIVNp+jaSsLWejIOMj3+HF
A/HQ5Ex78kp6Xa84D51v2/kXJr7163ibdEFyTybl/u0z5LFddu6BJRrMhQXFa5pSLYhtvDDYRneW
fqVoUXkrtmkiTa0SdWCDjIi2qIIF3+juBZ86azJdAEAwZ0eRJiQh1pGxYdRKlMv+RO0+jathvP24
So85cmHULGBrtZFnm6Cgxlr5HkggPEuh85flvPj6lMXzdpMeDPSC4Swl6ZfQn4SykfDsOBd8FzHz
jxuSCPbLVEEf36MdwFAuyyCkxdwh3Klnh0gnsEh1atW3bnSmHtg1wozj6jnTVLggGhLFP7EZjNos
n2q+JpB+Sr/XRigg/R2jXpNFDSIyQQbqhjbz3cSHZkvRGsMKj2E+A/s1AonCmQ4v94wgBtw/IMUD
/sqbY6t7kK4L+lff55hObHvmsnHilzMiVDQahHKHRHhuJTuwex53gTbeh00p6awTyuqdqo52KCiH
P7iAqt0e2b/bkHHTsE1UDLluu1DZbinZd79iREwirHwb7iziXkhBUYMY2hWNicaOvUCKQML9yjDR
wsNFYrlR4Fe1EjCAwSUufjYVV3V8gG9vh/kNoR3ZMrkhyzm2YOFLARTKMio882W/yuFSiDtErX5y
ryybAzzFCacC8x5R22LToKwk7TxaSan4riO2Tdxw5kciO7S4Vfof6pZEGQXmD4/k/7CjCSW4fNcj
T3RnjDOtmIbnTkSzVyDSHZK4l9s4aZSMWQ9vWLXw/RAmFeSY2IWx5ruvSyyUCXjQfdKG7XpWZW4x
Tad7rD8tpF/9/TekcwKyFpJbes96phPVeAAw/3MB+H8HJaVEN/oZYTaWRiXH+zNPS/qdH0V4/xVC
TEvVLxIYA0uTHFOjeCzxuXlGCmBrsknJRf352w06J38oM3pWrcilG+QrXpax8DtTxrBKai9x5e/R
Y+yRhK40sKILLeIWwvJ31f71s1uAP6oVqY1+EyAxfrV0KytEYQ1VSaBjlCw7sQlxnRWmTlQZNVY7
B+g0VnEu8KHmsLjFGb/LW0vkKby5IAtEFITbEpA36Deg6Tmwzr8ywK9QqoktqvnYw1Da62pQT3kl
XLjtkTh6Dpfxq2/Eme72aGOuV+PtEXK0eJxUo5CztYkFzAc86e8qwirgS0/IiuCNvqFzh+Sex7G5
nFtD6HiYP43vhziFCF+ri1VffvXo0u1z1uRZb6ShIqIkyZbhz4X2LHSrqukK1cM4rnSsmIaoBlsp
V4yojtKRtXOqlEwlAinyek93KH0Np0ax0gHmmZ6sGwbNTFCdLcbWtM0v9WRNgsIFKWz6eiKfvPGi
bbfw+7E3euDS2DUjHPJE9PWpOoJX+BXy9vff5JLMvxsKhmZUUvDs5VORuYXovp3cs1KQakOCd1Ve
ZTu1L7AAsgJOfGoMqBZpdpt7ZLcqF+0a83y2Swk5lSymMEH5gF8jA5oMrAAo7SD32TVMSxCpjQrn
SkPVwNf24EMv5h8y6K8rBx1p62wptJIVnyMNnBlvdOQjFocDrjGTrI0j9HeXalUYafNv4hYuAd3A
MSYp1P7/fPw5pHFljNul1dkxfxba1LGsOVaIkNVyt3P+Xv/d8YuYZwzBj0D57/uRQCGTVK04QRIP
sRpwPtX0+O6n6dpdOvSoEpomC+Qqhd3xTo8ge8CtuiGJUS7hsj358jmJsCL3UdFpA4bzCXp+4Zo7
EAHQi25CtPX7cIBDkfDypmKL+dPAcAj/4EFhMZCTLH2A/dOVk8TETAVCvQgdatb2FYyVVEOH4Tcs
7lapv8cHr7+OxvJ64sF7gC0HOPHV/yi2vylmiZODWo3oioX9LdPtz31qgKNMa1CGUpdTiUMcMRHs
pTGG+Gz3OAgZCxPP/pMLR8FJsWlz5q6YYfNK00duEqBnkZKc8XfdFfxZ10hn/bPMCa7a9HnZ7I+h
Q1GvHmr5mO+nZoqPfLjqdmrJcxiSEenXGPEbLOeOtvt5ypkkvaViV15VJfTsbELPWqonNNiX0coq
Mpht2NKpphMTnn2SUZRTcNQCEOpHuPubwxNo0I0QJIKDhdMKNC3OZSKVCfNpPvle4VPvp8+89QQj
osiiN9aOmxLTpHnRtYuW0yvKgupfxIVFUe5L8HED6XcsnIhmpOWXEIO2LsJNB/d+AEOO9znKUKMX
0D5DXPEC5CSIw/ZHMQbLzyqFu+07aht1P3blvZXwuRuLMvdBhWpGfV6XpTSdNcdH4m37WfvHjiR0
5GIS0Pl79HQ/a7b8het7EIdGfiT8mUtdq0O7RcVJHbjHrMKWpJiB2WeBjmai5GCJuS1y3hRLxIR6
VOWi9ZiuWtmy1oKrIqgPL0l1znvbssl8/xnBI2z/4d4JyyhNdlwOfQO8T1K9cebCCZJXIdSvb31L
BaqUo0qQv45DiSz7uHaMLmd2f3Ajx7vRIH9z0qtKX5zbfRsKJNcHoJuKANnu8YYC/Genp4UBJOZY
kS1ZETEbjop05n/vzhynEPPxa3NQaupzI8xLibiBHVKeKCtl1VadEBznre0GwmKtUgXt7p6D8VXA
Ob4V9wUdeUMXweIQqyfGEAIKV+Hj6LWVzPYGHLqvPUcU/EzssnGIE84ySf9P6NxAox3tyV8/UekZ
i51/cPTkAOVNFO2265LkA0faBiN2FPmaXaZ5XCj3KroLR6z5GaRFf8L2mAN9x+xXAjE88FsLi2zc
pdHcvPcYTqeZpwoKTw+K9DTUqOtFitd7i6aETSHsh7lw86MJRH7QXRkFqWFK+gqNWcE9/dXjncS3
jT45emnnilz14POa9f9n1z2bOnOeop82olcZP8ruYr4wAoXpqIXDIM0Bb6GaZCv2kFmAqnRbLhVC
8OmjTPU8/aAUWlad28flTIE4bKzK4pGYXEfnB6As4iNitIWqHa3OWEZJgt0ZoVZH80SLZqahA4EO
LL2+Qz05Urftoe7xd3AJODAoDHGD+fdUmvuacmbcsNSN4lWFVSy262yuoqguwVf/JirOkKYOPVBO
yXUtUre79Sdp5b6p4qkH9a6N4jfUGekDW51lZBum0h5hoD9TOjEb+tZjkAlgz281qR2k8Su/y/XK
jRHaccLDMXo4jqIxCyTFyZ/JPw55ctrHpftmmdkvXX8FcqF6H1l+Hxa5o4lszjrKG7TJwUD9DIVE
8S9OI+8KW5hP0l5Ix8CBfgTtapWUT6SSqFhSgDwl7XvfX4f7s9z9WxAm1B6ifP7gl85hVlkizGzo
WT2nnMsnD409cjTeUAceiijANAPdx1R5D6if9czy4wtPXJ9zIVZ5sJQmGFJr0niRyXCOeLy+VnyP
8XBihT8FGmnYcXSW1fossVb51/wRo2bM3Cn0ggSEhSqWJ3aqfIH8e31NOQbVTm7LDos9gDwRpvtR
LZtpR7PL2lZbfxH5qLF2sEBcrr6vDrtmZkX+zcykqq3X9OTIa7e4x8ldM/tX1VM+QjLOovYGOVGR
+tAnm5khZf36oHW0x/e9bjNhGZ5MmSqclFyVqnUIP8MaTA5Fv/Ov58hYsaez6VRXXPRUwJdk+JM2
WNcjd2lMxRnsHsl5kgxNPlzBtizZLcJ6qPt3NJeJ47doQe73J4glkFmEoqYgj3Jal9EIOx220QPo
l9z+NQXvXQfesJ9+W0yEyvttR/aMUAFTG/1tVbtluR6Sx9qkTuy28EcEyNVO3rJ5PbaotQmnDQeh
iuEn1N27aK8xGSZKLLJIoGxa0j0RNzdmTHjf/UMqNYjCdVnaK5R1UPC0SUSJNWZv2Wfjb32NiAUg
BZyp3gt2HdcKIvT6duMZIkyguTlhXYuVgx9JUyDqHfqgmPG6vuGYY56umMo+qcQq2oqZTRRb8j7e
XjCmkVPmPUgTEYi2a0FQrGs81ZkGxj3hn1lMzlIQWlnJ2UoanHWD/2dGsTYNYq08gCb5B8rdHufS
1P0hsSdoNaIc2kxJCJhvbyarWZraumg6JzlIkvkBU49BvPZkMK481ZyU+L4XhTuB3lxPGcS6HUB/
+t0ViClUCiREvuGTRjudeS1Trg3hydf8Ps6h6E9vqbdKEAPzV89HJYOXcdgyswNJbMD5z1HaH6iO
KsaSL4zFCQnK7IC+3hTL+mRptqn1MzOy2XbZNcFnHry7LMLiAVJ3HjVGBf/+0AaDOi0BOUnYxuXK
y3+evEHtR91XnJfa8E3AP1Y5JbZXsNhdkg9sYmHSorxxzEptxUjcZD+dEC0f3cm4JBAviDHYBL80
3BuSlucZSR6xguiiCm1h5Tct2dmLchyIOHJQm/hoe3Wt4EezMxJNHhPYVqYoWut8fB/1jReEpcvh
CyUnTTOpsvhEVtH5QeCbC3USn82baO7Q8kAilIBE7AA4FheXOJ8sT6rjWvlNzeUYRAvaT8outoux
1WFCnuQVDnX3gPBoQxBudW2NFaMkrZv9o7llhTchu9BUm8Zcymm75NNiV6BluYIw3uRMI2SbfcHQ
luEqW4HNByZFzuNS+f9lAFXXIOequI6ItZYB65QVF/X8NHQMViq4zGiYd2tKJGO6ofWXB5fMgOHu
0m2oWAy1BT2DMamcvoHZXADm0lzY6zE0+BKmITOFo/s2LDbZ0/cQRJBEUtX1apcHy2Hr2XFHPEs9
8VxJc5EV2vYiXBDCTCNRHQiXdagnL8a4iB6WOGQ293HFWi5aJjmNNURkwxFIkzBaansEgkOV7SBB
7gkOZF8ny9jFNjDclr/XSVOUHuba0QvA25V/Lqu60yI2zc7YoeGMTwSJP2wY2RezvUqNBJunehO2
Cnulkedcd05AzAy/eRnJ+9G9AB288ziMs5RxsFf24KScnjFr+LfqULaqBY5WGm9teWsI/aBROCx/
aeJZ+2UIJyIVSzj2F5SWTTpp1aOFnWKBXx/H3bmrq8P9qVt/n/FB0esWQ+LUDUoWWVPLsOAl43Wi
DGf2L3bQeYtyEbNFrxYsmMI4zIOmVDVXtXr309BEDieOheE8b8mXLsPYs8OF3nb7M2NYtZPxsDdD
Q2KYuvY/CADoZbDtxbb/gryeCNfj4pADgpPEId0DKcrOv8fcNSKHRedWCVMiq1gAMUPum1VR3sLA
NG9Fqbw/16a93dew3i/xOX23YWdlTakx+jxTdDld+Yfxpi1ClB+yQIoaaz62LwyiJJpQOp6mUpQ1
6NsiIX840StZny2Io+ZuM5QEImLEVdgSQd9y1RFK0tQ7L1ZlnaAAJG31XkegSR9xRGrxEKigXesU
ecvO+jmkgRnwznPtNKIpqO6m9DuK8gPVXiAGbJj5wEJVlR1Cmm/eHcWrL5gnsX5d7/9NKoEiEbkp
Dwd5xGaNw+NUUrwcHBcw7HvaIrGCWZk17l14fd+JBQoIZHHZhVgruzyBpFnRLMFWx5qcXADrWYVl
1a0FNFOHMs4doQP79g4903pFIVpzUgckz1oj0blWuDMc/9Sk+cg6HwM4I3IGeWpIAAbuXbyKjEQx
zkGuEqvyd6LKXJlXq+gOIJ5T4XDLIGA5raZtbk1CWg4ec+QqkQeQ/KzP0osHi0Zj1uoWhioU+NtR
AShc6Et3+4C/t0fyaRmEgZrTTquM/TmtpbwjmdNSMV29LOc1J1Ipy+yYp0QwkafzkBCVIOFOjks/
V/Lvtgd4xw9DsjcTKwy9g0DlzVPMcatA1tUQshdG7AiMO4D528NkXpzjMHIKqwNMWYeeYIuUDG5j
sBI5Hxrsq/2jSGW0iLidSL2nvT4xx+akrvbJ+mx1hKLu5NVP/gvuUR3EsV/FSUxmAf3MT/L/V5wT
yJ8KOTKKzXhmD4830GKm4cLIlGiCHachPt0vMEmPC1YIoFg5j3qftdaIaYZfbwDFV80aw35Npm6v
JGEtWKNM/IfCA82AlRtaHqqczO0BLru1Z+AadXACxv5ZJ1YmPBAyqXbTdIhJnDA62Iue66IBcwYj
49QBbeM6i4z8wxgMgs8FizrvYlogF+h1PzQDVIwj9k38fyOaKbQy7Tv4c3YJIbc1L8a56DsJV1xG
/R7eztEvL1BskDm+LC1GXpq5ByUzIviO1eLAVHvHbWaBo81JdtrDYKmzZLgfFuikn6uEQ6/8WaBI
EyaMUT/Nhs0bXtZ1FDTGGWEsPkugVbgwTyVBLopzxsXHQbkoUePUoLUx97umNi4D1AB2Cq3PxZ6b
87zyAwoyZm/xL27s7PUKDC7saeSMW8MHB9lq8WDu6J2zz7bEfjvKge2WoIESsvwAJijL/+txYz3t
gJuKl2vFdyjC8AzCeWXoXMnJ0on79ex1vo0oVq4pFTHCemhMWloOpcccQSuTJbel2jBN3IeOlQL9
ReaOIVNGRcJzLom19ons40kxX7s4DK71n7MfWZYmcSiYZ6UPqJgh4TpxIeEEDI9tb1qyu7JXaIsw
O7+6ziKyayJrBZzkZW3IfTSP997vRfTJhHsO8R/6xdp0B1B8NOcA5o3TEqe7c4nR5RP8Uun9aaRO
/m7IFdVMmEP7Sb7iFppy1qSYJI/bAuhwgulPyVz7O9Kui3MI2bLQl+mqzOkvx5yY5ImCWBDWjSl+
Vlg7xApUWKZiEkEIv1HvoDqTCU/Rwh2o85UmBJlKzm5E8aO1KJ1Y7rYCfv7+D86OQw4OMkz/bvBr
zx+IH4zIYYy1BGEUq558puB0ija9SGx8SPzUUrnr9yi1nF0b+L+oIZ08fW/v4wiXhKxLEzJH094a
Nh01JuMxpgNmXYXnk7O9pLVlUp/eIhoaZ4dy3dw9BD6Y4miW0t7gcwMzMYMsOblF4vGHtfWy/Xde
Ug0hakRBB7/Yk4OIjs+jzdXVOuCGBMJ4nwSaxv4yeh/T9gMACTmYbVOLzTtBnx0yTNxbSYxbXf9g
i5SDGDOVioECqeGLA/oHzeKe7bKHTTtrT49T5sMW3wiLs2SRDxgZNF6hyhbaVAuRVtbFsPEzlRDv
qUhIHCoiPxAB/exze8T9C/XlhBLMJoYWNLoAFWMikkzHycYlrlsbxsaMeI7VaP/F03C/uMgZ1a5c
mhFXB+7XnKhVl/waijPjLndQ+pyRCAALpANBftMD7ChAkmXKxCdDXzVjqtZ4ylIXd03DD/PPIqeo
f6utk32qjuLGxf3FpJewgYuwO9ecQhOqNt4y6wBvKTv6qQVJ/BJcPRldySZ6e7l+5c/KMaNM4KjS
fbYyM2qUoXq5y9BVwd99v+8fwymmVL4ZytWxVSDM5yNiwhsqEK0PNeyimvNMcdMyuljkvmDfjK1h
wqdYAIgVRbUfVTHm3gj2pohhaOMDMzp+hxWFeFcDcA31ffkDWG1PBPavO4SK09u/ZZO2kB+RuqIf
OJqwEUVj3jB4vPKX+zjEsqINPR8K0qe2SxhtemPxWOajbR9ZHTAtZh+QMJNzuYBvaXz4wN8iM8wW
2cutbFrti+80swEjzRMkF+XkbXPmRw9nBRWkjCKFCAojymrmoTLYeZivl1fHor8RagPsKblBLVCX
sO+45JgiTZE2Pg/NBJs6zpHj8I7pKYPRnSDEkl30JB2HbVjz9fsmsWXXFl8/2l40ajd4USoBhybe
fMAMi5wlonmNa5AAFemAO2h4mYxoNLg+0aMob+51ryAKFaERxcOp6sO71A85BH8TZplyishdo02H
gjhS9oPZkvoFNuX+mhZn21+gMVFYDDYhUSx4QoCm2Sgs8fHtWepa31vQ2QV96K7gVvv0Io4fqknF
iOxmzdL4WVbPcmk9YglWdWYA1jLq0UtZ5GJkD83nkR+S1yaQyHMQyBDAmbuYJH8PHxV1p32X4xf+
p9/rbo4c+euupUbCy6nqP2gXHKR6G3l5jrFFjZFFzloxdgIYr76iw/Tyq6cz66gV/g5d8d9rhuDi
lO1TsI9Svyyiw+G4QVlQKHgNDBUf3jVevVq1Kgeb856RdkK6/23qNqA4wxbXCJFiGxIzvvWVRKHm
e1wqwRgEAVGRB7t/1F2I5VgOrbLKFAp/DOuwlhBKdV3zPHZ+NMvqVjaVmohlGMZJlrqARIdWYssX
Z5aG7cIqmx5nNpnQzlF130apnDAEVbAPhTD89bYm6G+wtmqmgu937SZbzu8aWyZ2Xh3cw0suWRKc
Hkxjg0yj48WzVnjMXMIshas4aszo0G0/eSW14uzOjgkf+LG5fD65W6PdMCPrjCh4gaCzRFPZ618O
JpAcqbcMRKqoQRlBPTV40GABAgBNhFd4bhWGp8XTWt7t2Z58HVbANrUtvJLsgicm9b2HOc8tTXoW
jtUXnaOP3RKQ+gAsxJo0KANVxLzicj1UvqinBLApNx0TwsNEq4L4Q9CmGSqxpIOMX8/0AKAHPO16
BioRs6Tq0enENdFltDfY/rq6KJGr65rbp7uvSiwmC8inGeL442cp/6gcn7B3AkvvZy0H+fXK+p8j
nBUXW2Lu0pOB/OeZlPpBwoWPBn1lDHzbo4Sz3AAIp94TKCoHQRloIJB2DL6KASGrlVftrwU87Fub
Dxs2YoG48rTuuHtJM21px3QA9RXvvHESXF73Rovw59/QzVUYmy58JWjoD082ex6+Dn7/l4RQik3e
++7jQ3w1VuYU6pVRdo2tiO0BMOii2x2ex3G6XwJCCoftfwqe2u5jwdZzZDPdzxnfj7PCPnjyn7NN
Lq76iw+ZIMy9Hbw6jyEAgmA9XJOLhlqiqMGiGa2EPe7WQEniFp/FT4StgSNLWLDNpTr7l3cXtYon
nqsPyCgTh+wVAfqOEt2sH+iUuzhNMZlkRUT/VMH73bY3La6uD/lMWCm0xGlN2OEYrqBfEpzGcvz+
N1zNEcTNLstNSDF7Ner9KkMuE6tsMcn4h4Lr9s7GuMalxz1iYt3fe6Q3aE3WnIhvUmzcHfMNCzrc
9Kz5baf4QAWf/KXcPaGK3h4YR9UEvZUUBB+r3h8N8hl8H5i7e3rrtvGQBh0+WV4dVAHUOZxQANGg
lnFL+XyYtZ9p+84jSZnmG5ynfqt2KK2+1SU/B2lzLguWVKnRbzDQj5mF2jvnhbJCksCAeDRbq6Nw
i2EOza6gHs1WgvbYQwxJrTHZgpqUVNHwu7nTR+fbPaFID8fL6wVBCm8xjb08B/yqu0jDdRem9sUJ
uQO04l8MqZwYKKShpcpx9huXp1Q6G+ddOmK5eGMvqKTMKIKNWkIrfuAjRXeIryJCbRiil6xS5ZSE
A9n5HPxw4kF7sLKlAOrR55oS0R/u8vDtYC0j+pjzk8Xq+B+3WsNV73q6E3T/jwXpvJZefiZL/EZU
gSoVm3RhpbZaCnNt/I8Cigg0dzvtKu65UGsJyHFYUgAflSMg/ibafnU8toatfp3xAgCSZaMj5e2A
4hlil5ZJSFJ0aRkwkOK+nUvCHuY2RCbgp+nIuT1zyisOrmrttgb+T+6DVUg5dEquEmDydesZ1REG
BwyoqYlWdbM6kRrzX9hik9ppLSWeJiUKuc9/Q5UbinymCgzt30lnbsKM1kHjpH2ur2CKdPuPMlyh
No+Ixor6c0bdNKFQsc+0fF6EoNlk+8CKXFupO3XNSy3ermc2ghK7iZN41BG7ooafnySUUZ0cbN8V
pJsfTprAfLjLnVP/DakSe+oARpN+vOTfnMleFQmeuEpvh1dsWbmyPtfpAsqAJYBN7XouZ7j2rCvE
8707fzIXv9mHz1Q14hJ9L+iQxcEuIkwz4zddvoNRS7ErrrLKfWKB/xM2pIigI8+FBvGV1iOkTN5j
Dhnm9YKx3zlpf72hgLWdrLEz4bwFqcKhGGoasshfIzatVMaouc5GX/zeYZewU0+byGCy3bqYhBZv
J92azJOvn+DtPYvVMGgTR3UpjUuxhwyRy+OQlFodjrTZiyQgHduPtRxwiE1ujhf/WymjXIS2yJ9x
K91mfqftmBX9eP+Cd8qIluHTH8oro/XiSOlIXR7ryCNRcU+BVEyb51tAcaJ0A2mU4L8qk00zTbAZ
/jWh07CuvPxFMYiGpWeYvQ1BNzq1h/59mwBjoIr7oOjXrgAQlvivT9Xu2Vwgjxcqv3+FUvoocUXw
DkEAo9OoLZv9NuftS6Ttz6FqpNrBU/1pA4agNcmQ4GQE1EoU2PamXLZ6Q6l0FAff5pOyZbw2Pr4c
kjBnSsVoFO3YNoyGbxFAVIM+sY7rCU5DtLRbkTvvWPgZMRBVisci8E4jbwTGmWsmhMBz3Jm9mLOD
bleCw2UJUQPvyADSVoMn8wIh0xtiSPS7EL7qwu/KxHoNnWEa7tpcYF9C+F2cmWWJRajXYwbg/cTS
FdRMigH8FP93hgtLNj4dQnCJtO/H1wMg2YgUsrTALjsjfYnnryhPWRN6mUoHYUAhZj166NREeLfn
8Ga/wPkwxgArQiziya4hBLTguh1x2sLSrSqd8+rFLETB/bCAC1m4wjfd6OvoS8JynBT3U0l3Hk7L
qfIFQJFXKJHOqy9Av1uWdTEy0MUCvwvgSax6YcrrA876f1v1eUO0vd1oNHtp9epQNPn8QPkTxBsR
LTsJkw27oqcghoRxycjdFHPgVhjFpQNTv+i9qII1QCR0R6X/WtDvGF+wk+j0QWmDqijGC2Y6STbf
KDEJDTY/DR05A8v0U2r5gykpSe5wDpl7En1jMqDz2lM2FBk/9RXzLCHimJ5ONqUBvlw9alZwh7W2
WT6rSVo3qbFYoT2hprlAaPCFuEJYaL0WIHp1pQngCBosCIPTeirt4sktW+ugHukP5Msqol2KFb+p
BOjgzYWpSo4n6SrqbIquZc7LzL4/ApTZU6zyGFDM1yMs1UeXh5E7NWyTNxzM4R0+DM1JPrBYcVLe
Jeyij9WxOxHBl03X7zJhp4sxq/KRx5kTNL8yKIR3okXHf+NzO5SPU5moKL9i2CXvNT47wyxmPN3H
ZyFZgAx3L47TqUVprWPXlO4GEq2nrDT87RjSanN8mjUKyKJHGTidLHp0uwUGDQ1J4YjHBTiL4Hxv
3JuqmkJQaGje44/8qcrc5wKcbC1NjjUZolKLROTPG5xPwGPSR2emTCzQaTiu++CDSt65EwYBKRzU
4dTEionrfcAHbjPPNfi0r6gq/ig3ZLPSXuc7cWK+2ypvjCtMwFWb9WsvnJtkJeaFAYllPhDLhMn5
TcTHOzeIyj8M0+XJjK3nNvNwNFJBez7nQ94FDPslz1YTpUC7HujeRvRwGV+9XHsiAyipKXm5K9RR
E8BjT9gUnZcgk/ySizBbVsPDMCjKVR0j+KgRlnukzmBbjVGH4j7+U/ZZ3csucZqIRqmLeBvAnmRV
jUtg/lHX1jtCSOfrK87m2ZNFHS1/GmmHeZN0F/PEmSw+N35NhllGOv57utzZcP/JRH9nI5YDA8tK
tEDLKGQHt4qQfjnCP9j4zyrJSyPdm7c5dCIAYd01MXIFTVy0G6XHTTH5M6O8e/U+6nV81qjt9sEj
gnr2Uw8WBv7rNHua3UTgZy96k45XC0ZYY8VI5b9hRPz4P2Jhs8oNWsUPqVmQZQ/WMRb0+lcYqlej
9MASW+q5m4MQ0aA9vzoQYik9jXSD+pPyJUkCAGHBmXceeIOMDYXZu3XkKPbLMazzLL79WVOFfrCN
hufZkJ7T0CQv1WdDoa38f7S3uIhsRruEAqX+JTPxqqVHsPkYlGcCXbAKFPF5WbtLdknkEwrAFc8Y
qD16XbdlM66npE+ylmt/1+FTW3VXJCR67CS0PtXsY1DwNk1uNMsN0qwkYUCaloLUOmaEhQ4bvSJh
BT8a+lwyYIAMlEPsugAA18h/jKBmkywsVHOURqLCNKrpRvPG7BbVPwwsI/1CibpVL7LnWU1P7SDo
FAiuLtwlXZNXfbr+tiz39ey4rRRl+/nLFmth9WS7FuIre1ZcO7KJFubH8XxZ1bwuvt8wex/EHQop
S9Ra4qXa39KR+GTQh/yjIx+thLnqqRfxJteddPxGBmotm/4yJlOMPXj4LdJx0C3/flhz4LJ4DFZa
sdI9HEMtfP8BzvFR0dX2lkxKES/Vv0hQSQY1s0b1lToLThUTr2nZ+3QsqIyp80ePUUzfgDdEaYoq
hICKiPdDb4FXlUQKBVxco17/i7bI0y0TPFaTcF1zNdSdR28N5yGvngNO7xgl6CMc5H9NpJszAsE6
K3RwD2tmHpwYi66qU2FG8CuH1bXjT6JHTZL+6krdC4ikHNDBTSMOQXF1MMA9wj4VxfHupplxhG0j
Gv+CyNII7gTbV9lE2s5uPECBVMbfIjxwr8DOvXtpi88fehE5CG7UIUeujYrsEqP3E9Wbz6Xof2RP
YUSN4tWw6XHbxtXpE4MbXiGem5XXJ8nh+3IBj8g8cfRTEeGNWa4EAXWPiffyoJMEVRgwTOvPffCZ
J9fcvwmg3gYGCTHBKtfIsJSjxbc6OWDFfhElOuulgbVwyJcBfK/8DQYzICkra2MvPrGpw9bU34vm
4f/xV8mB3bVTXu+XJj35YDGLkP0yhC51P6r5DFKt7mH0q6kb/08Hv+tn7SbGDGvbdf5CbbSo0sPG
KZ7OSJu32CGCP7sK/HPNxmmQ7hrIRGmh2TU0/relWyTvrQoV12VMisc4ooGKNSQA3VSyJdZ3nwnz
wdGl8CHZ6gJpwcSwBsWxd4aOHeIS3Ulrd0uzXG+/MVfrCmWLBK7i2ReSETWtsxG+LZQ8fbtkI9eu
wqUkYFMgVaFP/NpDH/cFBTa3i2tLCQoS7U4/kC7BTO0XPakKYpHAGALZPVOdbcis5sOTxNYVnew/
WvxAVRwiF6gFTBtb2UJOmrLp0+DK7w8vBj0ncHynVka5bKq3dHbYKpixYZlenSVos771lb5K5n8R
ilSfsAPiMergv9Bu0bdHbrIhCA7ah5nBvlqDvDYm/0dl6ccp+zIAMED8ffRY/H+cKFQtU23xq+yz
S5goNddQhSC6fdJZhJNHhLwGqoZpGdo8t2ENkXLE9yczY3QMpZV6L805VgOwAes0UVT7pUijVe+3
+Jua9f+GqkVD0i6noGAaJca82mGCceRlU+Le07leWRLUUSH3x1ks42QAwGl+e2toIvad9/bHjzWX
rm09kwY0fr8fC3XaxM4grRzbtaj0r4bM7Z7jtNfEyHQiVoqtJLSDXwe+O0Y+KT6VZAjoqqPeOERk
KJSlh4t4Rmh3mSlhHc8caV2Xzb41+zoh5YDCP9q80Gx4CfpibIiUlMD7Z1PLkXenJGGT5EGLOlln
v7hwXmNYNrRbaKXerGzWRlJ7y4SIKgFdnrlsD68DrSvoew9ruWOT+//pK+eTepgCJTuJAzP6yJ6r
RTTTGAbKxrI2D8oKzZd7FUDnOdruZYB05LkdTae9wqY3VmD8MZFh71caXCwJdKbfd/yQuocCrxIL
dW7REFdrMn3k+fCBHpVPtPV7vyz7b1iE+f6pyT5hbPVqhJTWRo0NE+/GCubus3BCuLwdxu8Bw5bv
EGbqsjQK2MxReTD+nz7uIXSPJ4AE874STwCUfG0/gaB6dVWVVgOGRihFnF3u60ic6b8zPnMjVVhN
sUdVYQew1wQiQhn5O4yvI5it1ln/3k01ucuDRsI7h+9xHmCk7NUe0oMXhDfz+eIAx8JDhepfIbNL
AI+ClK6sXaC4XSDpc7saY8ZhacxieOyJLZQOegJw5weg35wAlcPTFNasS7+Vk824S7WmgeYqP0QZ
BPAoZ1QaE0bAzeUPXspovzrViVlrKILtnLz7AjVGw5mpsEQmFPLBI+KiVrysIDj7hgzrSAGNp8jW
XmusR2jBp0gpKYaswzPSOM3o1ivowXbNiio8/qmGQXPOb0EQSyVdHVlpMrRUrgcAm49sS/Lu5S2g
+d+4HxGQrwkORARAbpA8CUBuOEQ733/vMRbC0kxGEETV2nmpxR8Rv/gY65eKdVLC5EIrMthWrkjX
6JtOHDsXXUq6DO6PxoVsOzqdqIwoT3Rcrxnkzi6nt7c5fw/Q+0DtHyIwFg0lAZOJc2SqHlIYi4KO
4FeNqXCx/TEDGaLMHz8kQqA8tBW552M2MmMXF1WcrWAIo33faOM6xhVWnu8M0O+FT3cu30TsNAlG
8lSx1KSy/DPVeuL14X1WBVvzuW+6rvNlk11WEgESIhedZmMo0Mlb4EVGrGyQJ5R/BPD6Y5R13pVl
guArTr/3CDvISGzFhsqSIC19nZFV0nvuTOm74Ca0DNKrl30rUP4mBRGRlMU0Z+U8LMySZxImyJHR
VUhMGEIdTI7juIRKqnDvM5lpB/zup9lJcN5ey7/8f5k9YCtlm/gCW5XiZf8WCV4lZuvCCD+teqZW
GkW0q/J+0Tcp/qFape7laQAQ30EgkBjDKUIKEdJS2Sgguw4qyK8B7f+T0sa+LtUFoeI/JTarXx4v
FK/4X/BentVyFJ8JrvA6sdVWFp+8p9UtyMkQrzrCcOzqcp72IQ4/t45uFwWKk6nwHBBNY2PCis7k
Ulc2Nt5WhY0HUjzV7/QWMobDti5D4y893WbNPi8N7PdHEbc3eEb0o3KIAODuOToRfgcebOzc1BXl
kyV8gRBZx0QeJWluzlOVPGBWLaEroar3RPGnQnv0MaUCDn+hiRaa95hpDopTviH3vpktuVr+d8YV
iyBDAZbc+kOUDUDXiIUWP77WAIJhX4dlVf1tcEsfaZEBk0hrGW2ONkRmD2BAFPwBNGPXODX3PWfM
nIUu7n81ES1vyxDsTQuE/+2TSSxVGXU8YSiIEQMKzi2423KlYpZixFcD/pZ1KjEbsbvCuJGWZKc2
7cjvDjvK72ztgrr9f57sJrHJnc+hrQv3zG4WPgK4CGZ5txxW/6oec2Ri7lipV5AYYIFPbnxv2dM7
I5emvVoGaSdPdeQfIE2voMrHyCUgPWPo72spBeSz61px1EI6Esz10CgELJGPN2hGyO/4lKDNmSpT
rsL4wkuav/ARTZH5tDS2j8h0T1EyNm1Njx6MKtleEPrVORN94kU1re0XdslZZOxxE6v6BXnbCkuu
NJFr1lkP87XTcADhJ81E9008FVLQVll+RQ9eu5UuTLtEE5YB6yfkv3ZqZ2SZGmpbRNKakVOJunTW
DnaOqb2bdgyVH5W1jYwQ2zLGm3f5pJFSFkAwWpCQ2DichIBsJYC18AuuGDAd+/DCAqCjcivA8bj+
WMMy1HY8tgz/kAz292V+5KuyGFb+JICMgzct6IrXCWb/034SP6eRQoaVo25Jx8YgF5sIQaDUovIj
Zqgx3XoZDz4XEk5ndvMd3/l8W7/C0pVXTnC8acnjx31GUfI75Mj//H63YvL9JNpYTLs80lpMnusf
VK1qoHNdUuJVbW1+7OuMHcuTEEUrjeSQGyt0OjUTrrm4qEFxTwuiueBVjyt3ZU+iSzC02FZ8FqpT
y9di071dexkIkFvavZmHXYLpYKpcpNn5FQppTZTAizAg8dgzGyk9muwANVmOiJu7xpGn6u2Gsh40
lo+oFfPJhtLAfUE/9k6BjJ3Kw872FELISgsnWORENw4yL2WfZkgcR8HnFD1FoehVW/ivv5CoyWMm
1jo4YmGPL71VcevkTmMc2UEdAu6mVF8kF/SHIjqcKzrFn00mit8XyWLVaL7q/udbFR2zorKmdlON
gCq72nVF92xI3JKQqAiLMBjspY6HNIM+8IylUxCGcD5S76n7nz72eKh7iG4XncoXmEQUADST1DSb
Vl55AQgQgWS29STlHkDDaI9aiYf37ndw5eJ+lmvlhrqELbDZbR+LdAvZDibDBwnsIfKJRV1vB976
kNH7sEK0RHbknVIyxXpPFaw5eopdZ4JKQquXs3hCCd/674gO45PdSG6S9jCNo1VDAiCBUTjUSsqs
tbSiuSaT7H1ppRuZZd5k6wxIiWo+1UeFEKogP56KHLwcA1XGfHR6KigqNdJtBSehmAym6QfCcsEx
+wZvJXT5V5vFEdIvZO7jp1NW6P5M479kw3m6wJfceVnbcv8nnFUpFHpb/CIRoP3I8/oSrM7uc2xB
Pm8OhQY0Sls38+SajxvnHRIsP2hmXk0b9AaELDzWLHb5hobVaLciyF0XhAQqsqXUWzXLHWnFAMkM
Gz0rBLxp87NJ9yfm1x53rvKcJLEGXO/ULxku8Pdz+fnQX0u/vvGGC4fJdLrByIQI9PJzR0S3ku47
Jib4RFz8l54j0na6Y+6ugIfOdXNdhWIit8tmfy9FkxZfybiJZKTXRUvEX6E1ZpK/KR7DJTHuTuga
kqtYSOGIJQTeJo52MpHfW3dHW0y+K9IhjnqzHOKuZlQA4x1QhAfXx+hY3MVdMLd5jKWkYOFpOnun
VboqFWuTJhT7RVZeUkx9ZnRAY0T9F78NkYS718bMqa/dFgJZNNm1pCA5Lo7v2wxqUD5thnUYRuJ7
ixEmdjwitg4UQJUvjUwJ8/fo2Kcig23gXY4ctQpKwfEUzW3mJQjHZFmAhQ6gSwxRqp8k38LCc+0+
Bnk8EQ0orLZt2o+Tlq344qIXjEnPjdakuf+bB+ueKiP3L/U547iM5QrxlV9NTm4Q9HJ14jj4b6a1
gBlmmHp8AFhEZSFA66b8rYlnmIcMXctFVbvdV4D4s7mcy6hOGKcHZ3ktnN4FOHC6bq5+nbR1kfWd
gMhOnvWQvUB/yFaZhK4h29WGbzAYdZK1Dd3FViqJ/l2cYv3mdaV5flKSoU3KwGPioAU/xl0OFadH
9zOLigjA+xrjfZTXDrxGqOHb60Nf08K8VPcAiaaCdfzxW1gUOwoeGtWZqFF2OqeYGjJcHsNSSht3
2Vz8/pRD6yFyLm+f1AkdXQQsZJQEu8KyNPN0V2HkY7PfHKKm5LMUWcrwe0Gu4sz/0RKaMJfKQZ+w
aDNZ0MTTed7MBaY2UResdBwEfB8RYhksipsFtK0R1QWFpClojRnGkm2YORaVmsZMQjagF+nrTVE0
O7wPNRPi0X2CFzZroKQ4KFAT8zgJuMLXxakzFO2IarmKbTWhYoKqvDXsQviAbjIsQa+7Sy9o3Ggd
NbGTJBzxyypU59sxC3VETX4yDBLb+VFa/6qNeIEUsM1cILpcOIXv+nVqa0sgSMnYMRxqS+Sxyjag
CxIEUQyf8UmlcR3oCmLJtpWwkWut88d7eJB3PAH4sw4zDi3rBmIxoywY3GGa5UrdlJ1l75y591U2
OUZTmvqik1quCf1xGLJZi+imM9QB7958g1i/3eHgJDjmqmi+ePWW5sj1sGfEFgKTh94I5t+D0HbL
qqBP6MGHqcHGXFGvXJtSQZuXT/XCb/2YMHTDVJNSfxUV7yCbt2DnBKRSkP6J9mnVtEGrzBz3h2V6
9SLQdVzmOZjn+NWUagcM93pMdLtwNQEyEtcOU0t9JzuZjlkM7zpc0cIJqQe4hCdesSJI1i5l9h2i
1rwwcdfpNJq+LGYzpFx7p7SO+SvgMAZB/zJd0RlH7xj1vk+WAVMFTw1P5sxZg3brCpMeFjakxS0w
8R4FaTt+ES7Rv+nVmsduvzJbzG/pwPpfQaPlQqo05iaiLuirjOxKtuNSOLHT9lNvQ31ykIK5fiQO
J7XZVbBglxUBVD/u7VqgkN4k7LpD8z7GQ0Npj8uGIz5PRB2aPe6K3EYstjK14AOCWy6zGogdiSvp
ZBRxnJ5e5/AIOQYIYiWE5q51WTunEOL+uSuEAiXXJGh/166QrMle4J1gr6ZpkwmElRk2vo2KGPk/
NIzBzqtcwiMtXrNw9lLtCXiDO34iF7ak4sjb1gSWFFdbL+aPBshq1aNH++8LCghkIoHlq8e8Xv9N
l436B8TbRHpNnRMsUfxCZ4j/SAow20uJol2ORDHjkLMfJ8lacOoaAF14GzYi6la0+1pEAttHEW/P
4wguw3br+tiHXRvyocGt+f3shuVE+hLM2RDMdNLZlJfUnd98FuzSbEAJsiQY7kj5SI9f2gg+kuwM
F4/ItZlaysQ5mn5v/x1UXvjjri//XxC32wVkc3TYoi8DPqGbaxq8n/hviDkhRXi5yFFby8JNgl6J
KwgOVciIlXlZS2/ZTc8iZBwKoU29i6+dghuKYeQ6WWuk4xZ1BajvWU4eFgrAZRs2rnzHX/SFVK8W
iXxulaJG4NiP5RyXUYDbNGHqrtLeCShfyzdjc3FQaLQNvETZLOD/WtL3LGc7z6qp4EBNz0vX7t3j
GKZOfC6Vu2y7B/YOYAPEFRIz0NqtidZBDLqpfKmjPAJ6UCzJS+az9y+2eJwTUvOmOYS8j9BwgEPm
5S9lomvj/5/npZ/v2aUT/VXSP8Caabn5Vxwq/bxEOAQ0QpdC1jXhO5pe48RjJMsUdYIoROuzrpTL
oDH74XMaN3wpMIvPcl73USFp84uqnoB3NO2idcF6Dq/0BoNvwkoxiiLgIIAN5CrMj+YiFLft950u
iEThGzKFnRkhVCURbAUDJ64xz5e62nHHMiINta8defZmieQkJB+aJ11xKSLiIf0kS9sCkY7zUjSv
zV9osO7tzsSdtqhwovR4ynb1It8vziWFUpz9OjFvRIhvnjL2s2UvWmMDznxXmNEOBZcmIzEZseH7
MQALO0qlJUAFYWlMNimjBzKAQf3Gpas0tOCYXqcX53xdySzyK6x7a4qPTjbNBeECBkOIOKxut94q
2Ho1ZKi2osnC/jiHqAxO+nE5d+ecehnqpnGLSXh5zhMNMQ/VxTYLsgl5j+j+WxXayDdTdnOqVxGu
3FzABfS+LU7I7TBoS0Cai50nQpv6K/Sz3JL0g1Edm6JfuokpjaSib5Fx1o9i1be5UjlSnhSjc8SI
z4uZ/y+t8InmpaJOQWdFYBwFL8LuDrJn+Oi6cfshtHROJmfwHD9iDnCXYXZExMaWXjdKJXY6gP2K
jxSk4r2ndhnH7mr3JtsH710zXk7x+jED3zllQL7B+l+4BZqCIcTI5Tl+cQPekRRXBmOx2b8pHRTZ
E6YS3FFpCa2LiylaKudcV/rmBJXMnhdyYFwFWABtcq9ARHriO64G5Xzsl5G3YxstY7+kTwg37JQg
57fQky8jTF31E6GFYGUJxLwg4L1fqq5mXM8FbiqHCFbYShIjIvmhDETsC4rnUHlUHCYLrEWD1fj8
URG0FLV1FGYRBktajCaGYqLYv7fvycGHVOvG9BQyQuekH/HU+ukNX37DmCAws+bCGVEYcArs+Soe
JUAYvVSODZ+yRc3S5ZAsuENze0eLE+GPTe3DqWOKI30IFTnPue9LUreZRtV3lKRKinoi9NxIEQwj
9830xQZUzjzuVsXWnm+jYoTGzk1oZ+ic00gqXMsQNUAUytojB/I4LTPSN8i03dXSHQ8iH6Sxlkoz
y9on+Zv2XKY6I3JGdtP0ZWqbMEGRYz62ip8pIF0z9Zrntp5C4EoG4B7REjhDU9Gvd/NnCtQxWKT4
Z27EN8gGmr9upG7t4oerhDiZlC9J1Rt2+OHnEYgK6qddj3d2ZAJr6WUQ5Y90PklMVfln9E2mGOBI
nPuH0S3cUtiNvw5GoqT7yqYCH7j/kcsQtNlaQOZNoTsAJr/XlX4YN04cLF3VBJaj29378Tnn/nUY
9R49a/m0BFJ10lUun105h99te6+dRq+GCwt9Cl6SNmyzwbVSE6zZiC2zbMmEEzctJVJ+WdJShBcj
giBb4JtJ391++YIBnpLcQMVDzd43Ksuc8jAo/QJEBBHWyg4BSc2l6wfK7BatrcjYFMsXnpBfTUsH
kzwrIYq+NkDSO+LW3Bd5aN/JnhePZZJAhqgbK/1wxfcNrF0hQno8nkSkfqL3fG0hDDlA7Np9LitK
M7Q2XTbxaVH5KdjbH3MIrkw3aTwT5KsOg1874Iss1Kf/d+iUtTh7AT1md2OPo1i9xf2Ls8FQSNtC
W5MtgESetMLDPH+vi2cLTqtGYR6yMMHbK9nN/KkpXCbWjqqN1Q9u1CNWWPYC02p5DNUlytffVPPp
Rcnswbk0BYQlbbxKxaEKoybJvVXJGOOSwa+2/30fB+PJ1MpsBR0E/zKDnV9UCh4xCt26V8UyuQzh
lQBBw5J8bQMxV1i2WjLKddS3n/340dXnFeNKVtiVNUcsWvu0yhvu7IqBtW+54ViNKszHOrGtu8/X
yzctjFStA/nPWnSVnT8QBDc2I30dgFlXDxo3DZCMuJL3m07ZWlqJro8nqW2X4KWU5vXniMRm0gdc
umeZaRz1kOfXabKZ/vMS1CIQh2nxjnqMTzsclR16iFruDyC0BenYLqW1o0vaibaM961pY+JEvp05
nbxYpSENa3VoLuvAKy9iItm9TyMJINJiU/jgNn20e0j6joNVKbjPSt4iPis/zUsrVcWCuaS3MeXe
QqiccKx/bJa0yLX2iDuhLVTTCTaNiAdLxCj00E/Qxa+BakwRZE/Iym21BLE0cdeyPGTg08p0vU2I
ZhIxvEraw6lA4lyku0HCFH3cnTjCQimxoGNWXp1N99sQh/KTvmfsM7HQvtJpHCNLsStAlPjjj5Jk
i8uKd2UPxqRotN/PaAxmTEjurdq9bG9Gjnk+GaPpMIFsU/FA7MPVdERmsPBihWJtN8IGjIyCjccK
3VI35gTm15frOOgYZyy7gxZxPRm/UtwsMYh9h1j4rIRt2v1ZaSI7EQoJaD1hN4r/CQBXX1sthSgy
T+SjzWdW1LV+5pclbJzsGaTev2EsAacNml4bmqrNSfXMT4JJMaNYls1OISAQobmTOC2EdE7HWUqN
ndUWRT03pwvxoEk25UoE71ah9b4EvYjT8/i6J5KChjCgDndwnlYhHJOZJxVU831pGQY2lz6tQRFz
5F8qfQQT8KHjz2CORLtCFPnXQZnTK1YQIITMMgAO77eb5PmvQPzVDOr5fCZQaTC43/4+jqDTEFog
q1T1cm07JykNSwPgsGY8zOcp4AWTUQOHTThvwggKWn2g/quqVMBnT29hchZOdxj0ZZfm1M5l0CiX
8nCkTmqaxeZO5VU9J7OQJ1Y4KCdoibunnMchvSmIMT3mJTzT7bupRjbxljc44JCKmFtIL8jzkSt6
+46w8WVErnv25gqJmzd/J1zQ3yF0jkiVia7+wYI80mvGIEK2BFS/+1h6DXaAAft8PXx9BanKh850
UDxXa4URVCdkXJpEuOmUGvmwY9/4n6Ngg/Cf622gW5CmjRbWhJWBNFKDKwTqQz06jSqN6AIvQKif
3eDEBjPo5PbHy79wm0c75bLbjBaxgpcTimjQhMOmizwx1QxrcrKmFl8fx86vy8TBQiX8yv8vB61j
aRSBhbaOYYjX3FimKfBFCgRMv0E0X/Nb+/YLo+c7uGHYPzOwfrsbEUq2U5xm9wAttt7yw78bCQnz
OfeVOtJtfDFwttoueEpQHKKx3m/LEl0WGFJs8tZZbZbF+RwGJ2XIalzSzkyDD3xiL10OEKgB5FQG
/oDNMmzRLWnD4BsTYLBlLMeDfw8uQBui/vhAdSjnWRr8E/DyEjUycDly7YQ9cGh5B/ZF4Ywqlu/Y
d9lz+qd1bNMmqjKH+mlyZyXf7QnjSEYo8EvyxvrYPqBrXRfGQJcAfArkzbCjIlhxhbipujMA3sG8
U22wd7QYuYl662Xp6O4ehzYpUDHzyNkeDtr2g5DhrEkBvYzn+WFWKMZz6Ow2W4InBqYqbn87CE6B
T3hjAP5fSHc6zSdHuPRoXQRx01KypXp8FaW1zbidhUo7IkcF/rpjLWgniFPfmsc0V8lFLHmnUnEs
gfXL81hNLoGD7n7/YRmna5Xkk7rA/lT9h99BpcoYjiGhaAbuIi3tsSc+28BpZRacEseE6ospE7Xr
HtjonLrHon5ssk89+KErZ7BcTop5Tr1f7CJ33flVnMG6eHscV6k7QTeZYJNu4SN1eoMIJzwmluK1
oHkZcQ65yhKlPstvrKU2SzwmEYZsJc1ZiAyALMQX0X/TKvOAXK1P6AhCDcoMmwtQuaqibkhfpYQd
s8c67koPyYmxUUG1oE3qCEGQlDmsR8S+gtqs2UzVcoboWcOSlX2bFg72JHGvpcwAC7Ao6PlduRID
a7nlDex+qdD95b3q/030BT4hNyfLNaIcDYArFsHrbtzmW6cHX3vIYvb0TofjDRgDbzBM1bMDjfxD
sBpsXZQn5A6vpmcrFu33u64zGmyP840SSJOgOXijy7u2VbUpNUyIFG8Ukvp3TxM9YzMRfTftrW7A
KWZgk1fP4UGlADMMOO63GB7/tu80dqbPlzoU0FLbuLmAZihAVZUJbsQOS8HAtwFd1YzIeZu5mnai
G/ogMDvizKijz3N66A2TaS6Qs6B0AxKjNWwKousELx0YaDu9VYKu1LFedGweELO/Mj4tSeOngiuu
aQS+5LfV99QL38DBQaG1Go68M4OFSePTkWmLMM8Ls/eqRztkjJi4/9dhKQznOVTrOWq+zmFltz92
KVl7y4+NqNzvRoFH5FSnYiie8lr+byA7rE0ruzabP41r1n+8G1x2bZUftOF9mAMxMV9m7prUvmE+
HIE3nwHRKsPquLKmmyAcIb5wF2wBc+3+RYq8ua25i/CoJ8UyxqpKSYcyCD/0mtYNaJzH0XrDwiqH
/TgifQfWtiT0vgP15XoQVOPFmdrInQxBH3XGX3aQHYNplR7llPgYsi6manRsKOAMgEns1Xtkne2G
gFn1u7VT6M/julPGP2hx/ZZeBy3CcJTCk6E8FEkVX/lt6tMxvPeLddoO0ffNz0AwWFwgJrotSlRV
FyJY6OUGav1JO4i/DJzaJ/9i8A23BhtXJgI4vcLCGzIJj+ZP523Zu1JnEGOduoNl3n/A7g+omklC
7ZmnnNpjj9k/sH+7lxZBl1pLECOJxSHInvDLT+8hdpcTx9z/hg1R9L6j4ByDdYXEMhOWtcsDYxD3
N6IAUy0AyxOHyASnE9ZXB+DIisqb2f6T9RV7rFMt+jrWxdYOeOWEPDwdz5vJT8A/dg7eLTH3HzOt
RylmZVLXqXpnHiLRx72QrAaKXX4lzo1ZVtcvIKXcuoFAjhE2b4BT3LcGsh/mCVvI26PbAIZd1MjD
HYVROPh2lzGqB0UafaeZbOIZqXdjpvyBQ9To3uOv/AUhb5mVVbKeJZJIsGSKMsu/GOnfn0ePjH6f
3INSB7AhsMwEhAqGa7ufk2aUIwxEUJO+bWZiFNBb+ej+Y+waUSu1CW6b/l4zjae2Y2rHFLdla93J
aDmW/men0Qt6u+4TKpFKUBJF1CKaQN+F7sP/YibOTljYGc/ZNEso3VZ1ZcF9LXERIavgvLPkEE8Y
NRrj9AP4rHQl3FZJPwMdFqytnEMZQmoVIKqCgkYLv90Mbx0MhYULYRJ8YjPcHsF4tnQdY+P/YXNJ
ZeDNdCTR7BEKYbgriHEwQlk56nVijzGfCFjkHbkkJ6cKBcq9QSVgbTeX/WG6HcrVlpuPdvgZrr3u
VNmZKAUjIsqqn/qjN2PgROwx7SRStLvhYrdiDKh1y5soenr01l+IdkHbIYpFWy+ZAASMVWg6DaHB
gjOBhp967htU0L2Sz2/p/CPKUtTpERLmYLuLrOZi9xTzip8+njzRl4L020/A8dzJdLObff05NjWo
KYrIP/HB63LacYdjlG9WlO4EXiazI4T6BbQBHYgk9grsI7dZTNw3nO64lK9gKwqGMJnqljGQ36tK
ed9dhPDmu6ODVckKQxM8fb0wQ99trAqCrp7gGfnrNhS9AY9D2Q8JsRARacHk9Urn1Sm8obaZv5Jh
9pSIXT7kzltJbNmx489Xvuwohyi4bPDdevpdHtSEA8nepKrwzRc5ThdEHA6tRi8oTcFbIIwkwX2f
whJfGHd6W7J3W4Kr5MiqVm5+vVCgseHljuM7NGgXJ0DvEb0m1Zwv1qn3NSvbzfKn3aODfLGVy5v2
66/vTAnXYWqv5ffHKyM/PdJAW+IIUdEa7c7DDhzlOKuJ2jaCl3dR/0/oAUsFBzJwLgawMMNd4Hlx
xThEEGn81J+Mmf7/xN4ECKGP7lLbHbtAoy1uD3O9fGRrhA/yCDCFZ7MHWPzDQi6DlYp6pfH8YZfX
1AwFR0kH2Vh+ppBnvUUz6YvTy+nyb1+2s6LvSiYxAEeYgOjUApWMy3EXC2jJyA+hNFxYK8cKPVZ0
MK/OWGlzl5whQ63s/ZrbP9kvP7llNL4krbIRHL6ZrUUOWd7WeAq8FzwfDyfPdE628QHklKwmqQj5
FKvIZTsxWSbXf/JxtD4Zf5AK54NegjSzL/+X7qbb3E1dvb9hREOnQRoNgMikavbW8nidp1CKQiaG
+kvWXt3D5HTqkYGgtDOWKbZpF+vJpt/c8Glh18W49F8iKd5HZwhwg/14zFwP160YVlskow1bRzgt
QgLZX4Gb6FiDQxao9mscPkTyzeowlLpR6eej/f0NxBN20JSMhkKxK/nECyW7gmhUODREAutda3gF
It48uB9nuOpkAHuo4RNmMXQe6giE8MAFmffDZLkF9JMse328NVBgOqM8mohhuJbC8ANJE/aBj/tN
fS6N1F456n6KlGsm+jwr3XaIVe1cXAWbqQN5yEP0JCRvEh2rS5Veq9yeoTGGKtEzB68kw/t2AXkC
wqW6LFCQBWY2uSETRwLapEeQznIReqf0ICKKYkUQys1WFAas8Se4UHFh3lF7XfmhFyY++EP0Jqhq
oc30vLlz8tK/FzXlcgmTHZvjSNk1AnpOW2IpXMroaz79rvP8bgOd3KybYqxGB3jm30wmk4jFwtaz
U1bC4xdkRGT3vxGaubbQELqRyjwHPU6kXoHLjN5JlH95vusNWcgOfIq/lw+sPhz1qIWlnKr0qVC1
TS1gMyUWGvfKNr2M9i5o6B9daq3TP67bUQIXUmHMbkRoKJXFmBMtlHXNb6iIU1FOSUTJfqVvXs1c
+IOGLrqkLAnbvcHTG/hNAVgHpo+l/lrFmMyQik/C1CZ96zSc6jgql+UFnTVuJTZT88QCZGhH/WDI
F1vsiotT+1T2KuiZdkhfcAhu1m/7vOLEjisFsUQazcg4iM/lTgjHFW8tLTp+VPwG1Gvw13B0o0IP
/P8YFYlyFNzNWEoiqfQN/lhzZilcwZqBCPl8W5/4EaWiCP2thK9wIHhSKkA0nGjGtVvuOp6LXMLs
HwZKYyoO1s4o4/CC+k9EeOJTcOI4VvVc31pRXNZbvqLLsfMuecCI2VIyna6MfMPt4kJVJcXeN7Gp
00lISJ3FKLpNdSsxyGTJ33OTRvhlHzlOPdaJmGKHBqdnlMksE+jQIzFkND+9Qurzpjbrsds9WRIb
elsofKlcxq3VPxWxckm4dZiZsTfT1Ap+WQCmQ8An4ZlhzXldfFAfDnePyJGbHf+Si7dr1bLX39uB
ZONdboHk/bHOL1SDxNb6k1YepALS7SBRsix6x9c+6J3Rn6CbuuP21RGnKz9zA5HSYdNDO+CQ9QjH
xm3Ldh5MH9CLtTEGwG1Bqlf1JkAYwap81PepMhXBLon95A6fZLOJwELq+LsBsxsne7IMqH6OVQFq
UBPRZuylzeHdQfe17vdF9x0XMnRTeEACazoJwGu3+DiC6nWA7ovlHbltvI6VSPHnMlkAYrfNiEkD
EiopXBC2YXSsWq+k6l6HnT27avnhx+vj0W+kh7TQ7DwLvdAoyn8tKN/Qc4IoGFB0kWP2PxAATGS2
da70n1d9z9YKRycl12Kwvl0XD+h1COdp9DgAZnJtqcYBwCSgpamYOlnw82uu6+zyuXv+Nduud4IU
TMUQBxQCdwzmoYmbnvuQWsY4yhLBtEOxG4Ph40dDrRefoZxcUi1mL71/nPmtb78wVePZcpFUTiAs
waTgoj8H8xSbja7DVGzECpwLX3Ki0WL6B8N1Kx/M/LTLJM5MWlWjFYFwWzQI8Pfd3b5GFrdlWTCO
mvPwSXcp46kwJvNHNHOTxPD2xP/dArKFu9F9XCyyfM+Z/KGTKG3rLu+TxZP46SpkyWsummn3yZ3V
VfwlDUjD754dIyBbHQ0bPEQn+J6S6Yr/jQZDbttqCLelfEqks1MXrwN3YpIs5cIdM3AV/BaaDexs
Cu2ZdzidtbglOcd/dhOpaE/dBJ1wVInAClKw6V9eanFuxq8NJ/grDNsfN2dETfDZDQG6j83twpka
RPIjS/W3l2Q4e8PztnBo3D3rL1yDa/A45Dm+juH7Q+ZYqZ1hePdS3/M0T9IQnhVsL41i1y0tWhiY
kkonLS2f2kSW0pua2pVxf2kzI58eeKj+Oq5mYs6c69XrjZDEBg7akUDVj0NGS5y5rwMHzc5Vy+s9
gZ6ZWUjKQIEotm/oDR5vAr48ipvYFldbSEkN4l696XBKUbqUWGVZHjiFMZ/gTaCswyo9As7UD4Hd
DQX3GJnpF3hL0KSv/wTt+atfQf+sYwNEI4Z8DzZfd9xWSZvmge8IohQpthB0Y4EIu9Tsl7sxd5ib
P20h00IEJG5W0BziR9bIVMGZ+8qUb6Y+28y7vTlpYvWNLzDvaGYSP1FGgNeW0LU3ZEY0bWIIb1sY
clUoqWbUV/YE/j6Wu6uP1Gd462QCLO9Ao+vk8jBjYett0LfN/yds3RKTetTymWniYwF1t5GD1Nvt
PqTfR33xx1v+sjxWfCdcc7ldQMtG80W4BUIcaBeEAAB0GCI/BUWx0KYp2qdSGGUv30x7ye7H+d8D
/mMsP4Ix0nNhUi888XGYOJ8C+rMDl8Yj+fw1I1OGpWvOD33An+2nGvki84X0TvnK4C48cLCxVi+2
1PAVtqf2FoAXju+yEqM2kYRVZqUO/4iQWbDpAciHnPYOtdxQzBEp2frs7u7/ART37z/r8f5E8yoZ
xnpn0cSIHhkoSg7I2k2rDTtlBkkEbRrFdDLPDHJnLK8itsBgrx2odeVyRCHpa0OlY/CytWJRHuEl
Kp6erYYsaSSHLw2XDH63hp5t4m1uUweK9DCLJN9RK/ZN1mzxQ/0eYsQ/zqJhO5zX2Kl9qP7lzJF1
MuI+PS5J/b+yiyzj3TSoptdUtNoJzuMBHlF6lBJdQde0OExBOvHgDr1sFVyN72RugUy/6Afe4hvv
a14V/jBoJZFDMvdHWAFf/OReXZo40Yq0B+jQf0kyUR0ThhQwsK77OUywjLdjhtCS+w8vVC6gBP2T
qD0tjZswQxZA7fpl37i+0I3t2DfQqQf30dc8UWGxT2IFb8F/qQva9grfmgvM9ygqmMnpkmliRHuF
sTI3xpose03net9f2Y19juSoXxs0yNHbhx1onC9dwhNESFU0NpgPFxzUxtdUfl0lZ9qE6uloW5S1
S9TApcTrgyKp09XpvzCR9Y/Xc5tfGK3XBsSMTI/aCmyqYPotZKOaim62swTO/4FyLsiySkP/rR0m
ntpJZWszGgRdNbVh4EvjzrHMksuxlAdStZ6a96v1FIP3FUEoXvhaWFBdXjJhcjtGlsp/gzVLygrg
Ag1NbV0F8+h0KvKJ+Ngwo8mrrGKXOW0dAJaZ0CF8LQOYF/E9d7tAm1i+uXwznK1mCv+nnf7cL8Mh
+6lET6Pq0wiWmf7Ezh80skAe7BN78cL7TLh5ZNadxykzTlktagBb7pWYHtrZGdCzRVY0HDWWyH1I
eYmXE/0x4faTSAgBdG/xsLnwh3VBz8Dn99phqiQdov6j8S6MeCFfAsBvpU6NRvi9WIIDzJE4vUyn
5LfUN9z4Ie5aalvmcf6DRNei19WExFmVVZLP/PVRLCx0ViJoLn1JSz2MqSQ8P7jRun2l0WzKUJ2L
lFmQv/KfV/J5KzKi+TWpzLHquNm1Ek5MThPsfe87+iCvSNEYauBbKnL3CIWgCHXl1og0fOHTbp0s
3qZfyRFAa7lqVzYAcJ5Y7BeQUIOtrY9qSk5LmMAqFJ2moY3y0RQnfckQh7NOz9dbz44M6Bv6ukJ4
d4eC/PQAaxjxgHSSQdwKGU7ijGTQ3B0EHys5n+yPVwKuzzYyJaf+hXAhuo+gd6tFa9+v+sht/E7U
3LwRS3SpA2a0ayNGsM1NwHg00UlvxU7mPgkT4QxQ+vs0hZ+zkAl/z/KUpKd4XTF+CQXjHn9+8a2o
Wk/He5XO4b8qxAF+PMK7BGooJeiCnXabMFCg8o8HMXO2nsN/xlMICulSTYzDdgfewE4C4qA745J7
sR/kou4K/HcvLJoM2vqXr+OjNSr+GqiVluCKESUrtFo/WqHlWmODM0U8eXEMsUrY8Ngj7z6vEIop
bDkAQBN+N9rGuUQNbqY3hx5634KpZgNmxWFhdsbuZRL1fKecDeY0FbMIKjeS+k6YpJN0lH6LN7/m
VwP8mFopjRbHTFE7qY06QYqIvW4+PCc7Fnk2xt1Mc1fYEzFyxUtihsCzekcg+Sl+WpAVIrFW3++N
COXLEbW9if9g+k1JNR+PufgRz5CtVIYX5s3rAVLn9i29/dfErxJ8CFxbRJ8BbhKBWD19rV2UuoLs
PVYXOFClra++q2V/0sP8KQOy0dqgak4NM54dwzf7QNhG4YSHTxfDs/b62IyMn0TwYwDEPj+yi4GU
YidPcJij0yrJL9ApoNor4a45ILpmr4p6a0V2tGDwcLkc1hcCeOp5p0I+IpBAGIFCcqhLc5Q0/iyZ
ICSnVxZe0g4rRs3XEHUOLyTFRH2BaWNxEdMtNqjwqTaJkesFjLU96Meg9Izz65qITLlY4uBonPag
Kp3c2eoSR1+mV3Rrd9LSXz5JyyjrO5up9qXrnT7nt6Gm78zJpBDHvAK3f7hE3ZMAlbmg9oTUvXxj
VC+dZwptiWn5du8HF7k4Qmpfq60kO1815NsaR+s4TsyhEMdk5ibWQvWrW+NPh9gcKxGNP1PedACn
pftcGLM3lOQ8VU7q88vKM5zreiCMG34gV2ScidJ/C5xFwMtqOdIMibXnrDHxP7Jj1XqanMmW/3aN
ORBecvts/pUHtip/jK3o/jDxDuk1IPu7slEk43s5yv5545SLLb1x+9zWRWK4mki3UBuKVMfnGGK+
qUDGn+I8SzUBwoWStX90q31Lk1c6qgspArpbNh6B8Wvt7Iwi3UD3z3mv4OGpJ4xi5VlghMHluuUm
SSY1F3uLRPQD01RqhTzV9zgEdBYF+KwJYwWqVPWgvmPvPZbCsC0oOpZJGt+nd31rEXC5RMrCcRrE
++2t+uPjhODLMuIlPz5jPwkheYOC0LsKxFQYSMrm0C1xmmYr7efxsUNWPjVYuWUAXUpL/BsOEvPI
mZcLzuScNIdkdxBTPoc8YITB2H2P8m7/19YPSPMvN5K8MrwLwNmK89DKym1xwfdpjA3NoRkuVVjI
TvdcJeGrqIE75EMyuiBXAjDRv4CpYw0UopKTWGOFybUb4YDX79jYdB/B52R3TTYbOliUdLcvdUDE
rzqQMd4NidirFg6PBJws6gQh1GspRwPnmUTVAAmrnMeNXf5R3uHdvOgboxlhwIqy+zzivWSBwU//
H84rknD6FeLSv0FA6l104JfoY5RNtbS79mNkdgsP2m/JeCwdgpbnpLSnf5Aq0Qi98o6rmqw8kS1g
JKsd/WtQzHDzKOXN0/Z9RSwDxUz/V4hx0oMh5CyS3kzha0C2zTWm76RYY5VbI0KB2A6dXa5rk7fU
tuZQDKwkWk0y4RUolb4AIaQKxg9OC8VrfNW691eybxC9SAhYehVXZyvBb/A0H/5swaW/vZ9UIik+
pUUVkCgwMeomdiL076B3R0lx9xzeTh579X89OjMDKPRo83T5jj0NF2yF40zdGZBu1Fm2ke8jiS+0
4/L6ifLeut2gHK8p4dz8AASAh0RwsD59cWE65JwWEKkbpvBeBN6DHPvDMuNsBSy6c7agHW73VZOI
K0+jbtpHYBCFmSrY5YqnLODXcIOEgW6blhVQKwHOJmGz/YOe54UDiBYJSHpBuaJJ+MxQ2tWmjNyg
xKcVvj+Lw2x/xhGyBAGDz6Hwh+g81gjutI8jyEKf9/PTFpNQFsCN/e7mD50TAsU5QJeAtfx6VcYW
kG2PHQVlFQnvimqaiP26f2fWPHEeXXNr00jxfpresF/AYYBbHcIfaKon7piOY137egsgtrNlbXIj
yHkXVLRo6pPIFOEz+gtGuLkZW5HJQTKeu01kO1qGmFQ9h/RAetNHcqpKE5til1Qjpql28knu6Q9h
W5rI/MERZd0JxnzPNPxnfl5yDA6UH3bC2A02mGS+DSQf5ylqsjgmOJvXmVKS88ieKNVdSH3lCjXV
xMs8Cf4SbhuzSJ/x3F7wmwGEYbjC5ztu/zG3Dlsm02EGqNeoZY+KJz8icvFZeC9xQDkJW4QDjJfR
nV9ahIDDryb7lSmgFCv4sDHpu4DJt3Qemt77Zf0tJBkRoBup5d2YbHtJ9hPlW/p7hUEeHmPL3RX+
XXKsV2oxVmo8xKXkfOPBFJ30xLqkA6bqoPHC1LTYQ5lEhPg2mo6FUKneEp7o98qc/gML0yKtQl6B
7vJM5/5WUGZYXBgYWU4uJe8FNaY6pnq2b9ETYi1545Qkvfc5u2FtQLzdlbsCgJouvmQ5lkHzhg/o
4owQieLnb47QdBKjCtPSQr5wyYgElu6LCTxWkU+Pbj1ENKq8utr3U0D1hAEcvWHWcySbJXIRCoqo
oP0k2uzFrsTE/gkoMBnRiPlMT1B96txYemnV+cHQc43FuZm05K69G03AesfeOSfrzXzwSY3dguvi
0EPeN382HM3CZxntJR6ldtGEhjj4kIjqA58fN3EdJsYLEMc8ArYEAc/DM+jnKA2PmWdKQAemwPyS
l/VOo5qSCZ4zudEW0QyeY1G7P/0OyuZV3UP2yow3XY4UqfLRn9l3eBLot2G9VdTBOo4CBpqFjbw8
BfKkpfSiZHRpIeLMr6JmCcVnYT8DxQcIrkuFuhC+rBLfIu8EwjHpjzVdXkDOyxW/X0AZwvfC6GD/
Uyw+BkWpj6H7zcQqhZf2hwiYe+cUblRNsaOQmlWs4VVGrHJ0iURq6FHC3VgbRManIplAn+feVpC4
VKjt9krPZRkVvynfbIDeacE4/sOJjCPRBiaY04HIg/hfiiskkieRlj8eTOb10CyKJg9V/RchDXgw
72wbVlYBTBPwuCxaD2+tN/Sw8rV5lOsiT86L278yzQkFD0slfItE5C+FO/znu4CrXj+8R5Wwmpjy
0O+KB9xMW16wpnN5s2xRQOI+b+aCqBR+tvvtjLz5qOjuaGcR5r1zyWts7WZKiDw1Mg31jWdUENLT
5/7WD5NGUcgP/UilbE8mGiW9Gs6QhjHXxXyVVzF3TZL7Dc189e1GkabKi9Pjvjnw1XzWPHcZBrlR
Kd785FWistZHgFKb7N264myE9jug+PlBGSVedBYMm+Cl8cl8luX23vnMxKJraxhL6KXqTcZ+3y87
HW1YH2uKha2beKpmVTEcZ9xGYozMoNkMoOHHYblVZQMN4m0VMpsOeHg0S0F9C392SzDRQF7nvIkT
fBkJp0Ssd73pCva8Du1MSorVmnjKIkngbXE2nGSTevS0fkYwp0urq5Vaq6CGvDUg1Q/jOotDK1En
gY08kJdFv92VbGLuVc7sEzz8gJyz8CSUQHj+8PBTwDm5vyANvDdtShG4fv49CAhBSfTyNGVs+182
vh/dsirVWnKkg1blmdM8K6vu9nvWKlwnt7C2nqBvSvNwrH5OEklFvARJR8aGGyZyHmHgSmeukojw
CCDgwMwAk55GgRoro3wrv4h7absMzwI/qdebElyBgmeOEONF66HjlJNIlvYMx979S0ovFzvtzqGE
+C4hC3P/tnfs1isSxc8ijuVaSgbL1U95TyuiOcHKFqxJ+Xfx42DM+ZVIgqIdjDDkzCPPtyUvYsjZ
FdTIwl4tN7z28qovPaAXiqkflA8avud7q18C994rgKXwP06r7Ox8pL/7yHQDD+ab2KAY4OkNr+0y
tqgv2rKhp+5p7pTGTtcPLwmA7bZjR3WdyNUnE9bD1V0IeHrTHxtGgsVJSvKFaGPqVQTGzOOry6iA
0yoUvfFFwsQyBAcZFBBpGItlIupkk6ofv3FnsdcEKbyOqYaGfBF+523xUBjOpymxrSO3ABmXKEL3
+bXItUMP68EOTWRzXIZrLztZ0fqBMYAH++pgcg6+4GHkiZdoNJtHeZ1YbFx8UYUSlOLUvsYiP7x7
kqhiT6qsR4hwfqNDGG/AkCfwTrjNJQLz/Cvfs44G+J9nzrIswxhWdTEgNd0jvbqYMISyjy99OnFa
WJUukwQls+6sexeDic18BorDkyZEf9XfRPL2lOsVFY2f1KAJV7lbKOuzabIcd5q70wCiUFYXH6lu
N4/I5QFvYhJ73fs+CgpTeEwXnfZJUX6hwzHyuOJlVg2nflxUM3RRmqHXeNz17m3SWzoJUgXOKMbE
+eA/+Z1Ix2QhpDyADIakRy4cUxE/xo2lS9hhmJVZxH5q3+8u5ApTg5UXmh77AR06OXX8gkLTQ6IV
X0qvuy7mjFQgYbGEDMDyuu/oUeDM1QQ2FOzrxXTwxxXUSmC9meIuG6Is07vRVDww2r2r3dCvkrlw
tR2RhP5lnT9MNbuWh6PFC1x/KCrFiXfPb18YcApqVDTPgi1LOM6XisGCoGxDIVE09ktZHuNkZZbE
al3tb+hQtHcnjQEx2GK6Y2YAkECs+yJJlvKofltIH6UhWHcNMtZ98xXp1AvNEPb0C6uVzOsOYw5+
8n8VLH/LgixZcNdvivJiwqMnfu32I1OhywfQ+3vQiL27CRmZDQa5t60FNL8bG52wNDEYGDoW6DLR
Wy9wQNYWsrbxoA8/QZ8Ok35AfpEbeKVIg2xeQ+UF2REDsOsapmXA2nw+1UXYGU+3lkOfgJnLE55A
/wWEisaAB/WOUaTeyhbDeOZ1c+ZiH1bUCpufTZ3kbZTBvP8kU8UWmNiXvoV6hg1WkvczhXlS8rbK
i/Fzv68bKYUCnpHwzsQGVXXDqXq+f9H0teYCTBUZzqzSj3Mn+f2hLGUHEkxWD/mI3HUFvnCmcTNJ
s29SEpYn31PUShTplaktCNAdHfjhCwPhKEncZyN8DNe5JJS2WS/jle5TEhHzKrktYNDFUoMsw7fz
uPhA/nJCGbm7M4l60944/DSM4BwhZ0Mbj7LwnVBJ4TNluukIG+WYg67vbprpa7tIdJ3XG5czNS5p
iv9RwMcZaAhx/qfjm1br3HtlR7jv0S69kIOsoVYFRxQB51z4oAR221keAR6/8XJRauDcbSlf02+D
GPGIlBbpHKS2pPSD95EMYey4fA/dKecngX/XdYqaPHAaRwZVZsNpx1y2FflYIPImrrsOQWTMh+PD
xQUUcjcdSV7yG3WkrksvRVsRptFhGrl6nNGEZEGXsqrVwC0CmBTd5kkURGRH6weu2ZciAKOWOPyU
2YUvFnPVyphqDk/uPrEM448f/GXvfrT54L8A9KzpHxprsqE92Ms7WISK6vwBuizuZb/dpKm+yD+X
69BIhR79t9estipwEABNV1M1+cSuO0GQPdrCQ22EfLp6dbKU8gN6jKpPEa6F0pxJNMTZ+4iF/d8L
slZpMXYKQ3KXgqavGIQ58WuXYoM0PPsoszHEOrwWb+RpmErNPRWUI53TsANhAk3KDYp5AcqLJfRy
I/amXdat/M45D9hcJjnH10QierC8mswR+BxahHM5meinT7+v6hmIyjJolrqEotmANiUbYcyQnazG
xbJW6eV8nhE2pNu16RBg6CJ09zZoycm0lAgltcesH51erusvgtFrzIwi5oTFE/PNZhJyeDBNvtce
jf17Hai2Fp0ViaadXVHu0oKhxCuLzUUAvu4Dp6tS7EAgZ7KmHNKj1h/jMp0nwiBc2iy2n03Ht71l
EQFhY0k2h7pc8ro80NE+u43rg+RvGzL+XjXGp26qpfshlHj9MaEenpTMBkY/EjjDJWgCmw62YXh6
LdDnRGoAYRFC++1rEz1/15m/FwIIJx6XXHd+8ASvnkyBqoes4BxqT7gorCoqzRV1Vk16eXYTC3Q0
OeOjxCWvIaGi+0uQ0lvUT+qYruH/aPOrwPQ89arJeexoKjpyAmC2PY/PmhEMNaw0MAeic8DPEbGp
/6O2aVuUBc2K8KQTeGNWmdBiRwBxqY3K3RohI1ryjCQzaFSRXsy12Wdt1a0zSfwov//tg7T3V59/
A1bNAoyJpnCMh506bvR06QMa0IZlSVQUTV/wJI0fe9zEEr4ObZx2cH/OwKWHgnXGCtvRKKBnNvS6
m4MxHWuIzWx4DJTE3V35WS28EyB17kh+a4WvQ7l4AprippuF2LFdulmvd1tcqEv2P2QC43s40NS7
vkGgpjBZFueUoJlNhXVbBXlSt/4F1lthA6fZeJNNiwl36niOpFd2blcBjLbbqrKPAn6SJ883cgLL
f3xFq7rEPHjFTSEUB9FHjVRdPNoRsuM97bMhUD/Ff6Z+6VubCykPvaphO13p2cswCoPh4axbrPqF
bRVa01z1sU/WDyrVBd+VEUzkzO968wjkTCQb7Jb/1FBmRH6rrbMbVTBaoqyT9gQA9P+yrd0S4Lex
V97Yk49ETE3mPR5xqiG7KRYO27QQs8oHJiqZvNKoz8mLpxdZP5juQFBviiRNM9LI2I1z/H2OvPus
9ULOGVrmb1PjdxL48dVvpSJQS451OQTTr5t+GxJw6BEHBK4uc4suedgClh6FGAa5nfcu3cO0Bvsi
j5uniTrLVVBAwkV9viOy6AK8YfTyDv7LofgnLV7hg6wTqoU3AQoBNJJ94Yze22+K1rJDWgWVG8Lo
7PV9Uu/14uJlUba/LIdTmtCBfGZZgrjvGF4VFqUOIF960c9fRfPyyofEkF+8HCTKHilGNam+9R3j
/6k0IpAAxQBoEJc0UX8KuqEhNRqrgP1fwAkoYCU1lpi9PRpEfiKzQcoIELWCvXd7t3Kw2QWCr/wN
sKSoW8tiyuZdWWo8otFvqBVPoS6F95ckK4ZGOeyjavksIKo+y2FnpJENHt4l0PIyLQc2/R86gkBJ
IcaJixj7J6gz7gPoQOiKj5RRf4xCe20K5GbAP9VkgpvyTpjq/+FlolNH0GRLR1SDCGrQhBYoRPAq
YV04eALp61DGIrLHu9GmzjY7jHErl/8t5ofP8cMuuVtMSTLV60h2/tqHHV+ZsycvEa5WWkK7bxHO
kn0e8Zs2wvYw7qEmEYaGsOLZgD9hs0cMFU0zjOfe6ZN1hls8QFxjwx6cST2E7JY5zP1jMqfVjl5j
2+kjkhU/3Q19yaf0v6FHPmI83Wtv0dIh+5fGGN0O4bb52NpWv3FErMsPKiMtLtNrKrERGaBgbT41
gZ5YqbnTyExmTqqi0xggEzUpSsGhejWXjVUSNgEiF+jZUzVlkPGQOIc67ZztRmGheHxKl8IBSa3R
82b9qWjArEep48I82qunnfzbTgwf2PfDNb5QEnjUs3SPpYwMDarpHYAla7fox+YhCA9f0eQfew1E
8xKkH6UAWnIQHmM4DsXj9jE57JJWVrqRQ2N7VXMu3b1bKQ+PjoOih6VGreFe4MjrB1g92JiApaQv
IuYIEL3vuqwcFLutYDDdtK61Wr30T8EV5o7SoyP4T0MJRUtM31/NtmnalVyWYxGvCnvM0PlEkBrX
WjlqlVeMDFi6hnvoUpJWAH5aQrCPBk145Sd8ug2ZlVeQLC8sAq6j96pLAGVkoEtWkquACr5CL9Fk
Azwf8QELxb7w9duOouhWLf5gJB+yIzeTkw8MlSNoMcpAvbyvPEs28LedyYAICTnziwQcCeoKz4NW
h1iwpwRDP6FWYGWnSWY+6mDQbFeCM2pz4bWbAtKCMli7PA1KDP9cWOlzHntS5HXCI7BCt95buJn+
+8tGjjQMtBXN9fBlsrub3snBJUikw0rpbbnY/TVaD8VDK6fIlpBlP6SiUHJgMK/ILBY96ciBLhv/
9VuL0K/XlMl1Y/qO9XF9oReZsYT1Q4koFca7o8Vmk7UVuqzgr1x1V9JQn6Pg/yJPO/eSiOx3NkeK
8s5cvT8D8NeKOm9lt7DwOl4PnV4g59EOXw0xMh93UCgyZSjuYujSMGWjwtFPm8QqSxqRHPLfdg4b
mbvMBylxAfSDLvQeSvGK6KYYykP7xqjFCS72GI5YXimcx463lftaHxoXpi86xAQu7eveT9nqlwiT
rlHNZWNjIo4usHhljupXzISIls3WlCWtFIFCIUia0mvf8H+AMpgs/wSaz6/T2y/q5S2uindGUn9j
C1XtjUWDmguQOt3gjeQRKsJBzkYN+YsEtlhMdWaRNzpOCZckbPY9AbyI5vSe4zFSlJP+e8mhFcRD
XsEl+b8722ZakLFIumH52uLS0PeV1SEmcPbcJbRI8FeOe7bT8G+22ivfn+xw+gb18C8Kp1dDbLd2
ygKuuk/mQ42BiZsyGSJdouEjS3xpuELSqNCLdaEQxLLKO268OIjPJzZ54AcXH98ggWK3ZYxDBarU
5ov1uyVrL2lWd2X8sR0A9JZ172JN5pWCTTHgE3QSpSw1pvXXREApx0N51PqXnioAr5Ce/6Zfp8w1
MreJLwdnJe13/vEwCNcDNaNG7+Etu4WNByBiaF0P7U16asVxuvhzRea5TG+OrBHc9I9YtTPHTd+Y
MROBfwT3bm/ARc5scGwXI9KzhUXz9YrhbcQ25cp77uyRpAVxiPTsFgcA+12jjlIQofsbf7F/44+3
GAKXqo6OVuBN3LOehxyLercWGajdrfZOtmCtVjBNb/wTWqBLBe+lR1gL1zItDU5go8vnEE9f3H2r
oHyFOpVMlrkcQetfuss0LxxDo9p1j3k1L+txrabKXe2Ncm+V+Z4kX1avWRB+txJJMKIO23aZ4kMe
+t84+ix8Rcr7fAgIsYmIHtD5YOiHkkmGqWcniECntHOlafj9TJzzD9+uk/A4D0EAyQHxuLE16o+8
Ty0LokqdXeM+fXMOjihMtE555ZmKN37M3BMh6Put4cE01pc/MIklAssfoxtrJGBTcfoOyGkfIf5P
goPQlgkqMfkGNzMHsewX5ZDf5bL8yb3cTbUcISnGY9/ugL0tM4+pM88+phPKV03m/a9Go3h9AXOL
/Z6YWw2eF0idqCqAnwSJDLs5fdqdE1DqnZ8Tg1hwjP2sW6MXMjIeWuk/OpnoZBSXlaL6VR5q+HzK
jiulYdkID03DXHNuef/KizApgI+KTfMi/j5e1nWrUWgZ181/2nK5A1iJQwx4kNDSXMtVkM92VjwA
qoeigKmqR3jXbXyp6LuZSl0n6T5/qJVBCA11eOL3C8SC6IN7nCAZ+9IOu61dYyoYPdAOeBMTEfuu
yQk96rQu58RDIXf1YZtmlKGVo2QyEe8nYD1wey2286+ZjazWIBbm6w3as9KiaMkd2VAt1BlhIg3Q
4V0/wT9kT+NpJ36/iRT/90rtPOOW6EQbbNU+EwcHtFxwgPmqgL4aAk2JuyTXhqPrH/Jx/Ofokajh
UdbFwJaTALtw7kotvvRLbiFcoUAmDN3/DhYfudLVXh2LU6uQB2nGVs76Js5J1d7DNCQPKIQEmKX8
YVx+fWEkCk6owFmhZLdGwJJw8OLXtONCB4E/bKhmBdEg7oy3+glqgFVrgr2OsGyMZQ0hx0eZ/4GW
rTIdtqJ+5hkSal8VklZyJfGQMhqFtf3RLZRWuoeFX3hEtptbF1HNVxKMqc40OPTWR298nb0HFqsa
6Mmyj4fYeYpB6FTQFdBou8FfosWXzappSyG3NuyzzIpjBms9msD+llfZyEAoSKmxTtyXFY+/iQmJ
oHChoBeOq9w47qb6VSchQT27X5crTaFdrrcRzxAWU6lC4K+9yzgBsnshpXyCdfkOpo5evjR5H+Ps
VIqE/Uh4WyUZYdwNG9Rcm14W1sws479DRnc6fMzjsZbDgT5Rvkiu1kaGg3I0LaF2a9ESMRflXMQW
kol9RcWwSJHDg5yuExLRX/XST6xBJ/j7FboSXebZrC5rYdgx8vo4iF2Ujl8VOKDdr+fNaUqpEa16
hRUaTTeNTxUmdSWUKGGqtw1bdm1G8wLKZYG1rpGFyPgSu3bka+HqVPCMoheqrKjF0s47CAtNZB8E
sBKahnbzDZ/Zku3GniFDU8TsJtZOwgAT9Byh+BMokFVe6R1sejNaJz1u9fhfI6euxJkCxla6Mlzf
4ys3H66Opj/rECIAMc+zEj9uteLZjd4SwoiRkRc0axOsmLfsAqpnP/o3XKLuHGrubolEY9pOOial
YyxJrXwlhxjGHXaTiw+61jjN9Vw5o6nfm7KX/fayWg+miup9nD4hUhtZaS2SCiJ5zODHFncFZDTx
c7JO3hPkbtWsEBh8ZsQlHVzN7qt+RWWrpTE2SfswrUQYgI6aMJ9X0JgA7aHzQC741J0oBTRbgIin
U5SFY68LLNDf60Jrx9lc0kmZnWnTyhhV3UFQ9hE3Vl0mk4DVAzCilkBCHhNto3cGxHI20LZDeQIb
4K0fnIbHDPiPd+eeaBKSgULorY7U5qcA9rDRtC2oLUKyWVm62lS12m9EC/lq5JuuRpfzHES8I/Lj
ogbiU7FRYSApMvgGx2BNtPjY1FhHQ6lxC8LBHvaXFGK6fjN+p9yspd6R8c0hRy2+hRZhVVcvRqHc
tN9bImk6pOoz53cEBZkCQoa43LSDBNt6z+9XfPAshYgsLjzsgemlCuwoGFEh6bvI0/iE1eE4T455
fZZ6/RGIQhEkLQn8fAFWff6Koo1nc40C3SpuHnC7pmnM0vaM8enoGU06lTHwtkspars1MYK/gRZa
WLUbKO3Qh5DcIRPNn/Uf1HHz3DSXXY5QXoLLMgOU83sU9QlLb2gB1m2Z6tGFhakb+qv9or2GvDUc
4wt9I/rG5hjNhg2eHoSQR7iof36NRfGtBTgA1PQ2LLvp1fIAu34BOBvQpHLCdWm45ZcSh1PpcSrJ
b01xPZVRJF5+uTQ9oo/xCaOp9SrwohFVreCA8gmwihuGpaN9cGMl6Iq/tkFirrZfQCBseXoDuDd8
fw+Oa3615NjTyS+0HvIPa7ggDHAVngJuiR7Pm4MkizicyYXdY4aD0lG084Nfzh8rmi8r+YMk0Ixs
LI7Bqozu2nwHJd6u7ZKOzudUvP4ygeIjHL4YFZkA/2/mbmeUUqnpBsSof4dT6dH2+Fhaic791HYe
fKbV0ERBZFvJXdVwpAg7CDoSYRjekrq6gXnv/1+bgSVsEmgIiCgWGaQQNH8si2eKCruy6MTBZ2a6
Xow+mXZHSAAYxUx06eaKgurtyooUeeoVcpusAFvj2QgGAnlGLrIrW+5psCUjCSxPp+9fkg4vyFvV
6gBSE3XLsR5ggYMGHTvWvabaVL1eGPYLqnHQSgtESwsYP4x+5ngpBXU8Ei9d4/6I35NQ8RCAPWQD
cEVHUW+tssci6MGJpkvC1sKXoX/TUyBB8tD25ZdD7mfMA80QCVRphZnciPVkEhqiUSWeEsfPNF9V
pRuTNnr9VOTYvk3rlBv4UC93QB9lFxvTEzrpRRz7gtmGq6r9UEj0xwJ7bWopUM8y/2HXgM0BhmeF
7g7FIzYJqfLPwqNP4SypajYrsXgDoMF4LUfcWxf3XDR54Nepr3fmCrIJ3+V/E5Q4NudniSUl4TWE
77dMUnMU64v98t5Hov0zPqO1Jywca7PF6BqnTTvSDs5ikzwiT75z34K4J26fNnvdtNEOnquvZedj
bLDG7w+eTKSbWCxzhFmlRCqa3F21n6y4uP37D0rVBI+IAQ+cl3qDFHnorsR2GQwlX+l89Kf3pZIc
EXCgoQCCgr4g0620ciIC4/xLRo+RUINFM0PxbdIn+Uunnrwz0+M/KFxPRaWKx3V3GBHvGjhxkG4N
G2PTHOPPyMEKueg1dMXf41U4kkR0ajucDF+h3ZVDBKjA6qGRJLzejTSWGYzz/qOAJ675GsTQDwFY
LQsFzsGnFzKRi5oYwy2iGJ5XmAm5pqbqb/25bKrmQ5LUK4hDhUFXL++g+LH2Ds4+AqXulAd/l4RL
LtT68GAyAIajGMYVVSAwBP5eekmKKIb8t4Sh61C9KMR/mVoa8H4gRMulc+deAF6ievZg2sl1a6Y/
ZmU2fJSCBuSWaVR3YVVTDKBfeTiHRGoBVR9MOm9J5PXi2LogNH1gQPHNQHk9smsca5Zrf9+md20N
aU2ZZKevBQ4pIZVfelF8kVLWfWwYhPIYkGrKlcIAN11z8kF9rhjD94YvDOcTQDA3EgyPi2flWPNn
Sb3X9VEgApfVp3uFw4fAR7DiFdEoLffwqoqSpA6mg1gezpG7BwCNWxi523GKuc1Ikx4oqTkSkdFq
vxKk0DTMk1CulfnEAL0h46z2z9pNq4ISnS20Y+nMG8Q/VTPzbJv56uKg2OPs9KScBhDjvo4d9sKx
eXVQ4jMqCqCVk/fXfyyx93eMgf5KQQspy8kTtFSD0ZVUjgz8Akx1bRoUy/GCIm3pvX/rCSyqT8xJ
AdzTCTymhwZde0n9M60py/0wrbqrAvVMxgEcXJta1o23GNjRyYs+i9gV+hIFGLiNhzWUNwd4qku6
UgnClpqLszXQtRlUgX5YkimqHI56UQ8wTQd4zIjUeQM1ngb1J1KyYOxrabN0+lhc/8xydfvep5od
tsORutCIo3KR97q2+HY64PAT3cWJIKvGr/ZAsioCZkGLMblo/2/YR7YuJ2K87m6nKB6e8Dj9WZpp
1krxCyJqz5IieP8oNkmtb0vUTJ3M5C4pylY20UQxnGQfASyCKqN2iG+TzJdZXu/8zWakYGCV98oK
ymltJZW0P2YVlSd7jsZznz7PQn/gfeNGBigaG2n0tShxiJNMIRnLVFFpG4LZvAVg5jm/q9wifCHg
hQOyF+/6FQxbz5GNiqv5H9b7d5b1Z7jTj/e5bk+RHLpGlxuotpXT88CPWjtB4/QxuKS4I1yOBFTp
J8yXMJ3yllEqG7ysj2PZezqonw9G2onus2bhWoZvo9nuYraJvIWxIPll5oaR53JwFlD/+fIfWqNG
Wom6J/+6ofuopzJeZnk2BiUnwxa3s0P5y0e2Aa4Oe3h89zlTnwHBHq+yviQx26ii5HoLDz7qSfoV
WVfpPnCbxjsIr9eBHGeF+CS+gFKk2Jae0qeeOxoj9+0xZCR6/+QAXkVIC50/VGViu7HAOEpWcydW
dEJ8DKc5QZkAln5fF6xjThwL0hWwVdA/tb7eQsUMR8UhKMWMcbLSKVEODaVMSJSxI6bmdP4okgPB
DLAdEa7wSnkAwf0kXHWKr8tNKmXjEs0YKEHaiSIl8QryNf5k0PZK3h+ArATp71w5rynrKaoOf6Lr
zNJW3V3NhPG1hoTRwnY3IGY3v/ETA05FJZsq57epHnvwpLaqvN6soL5xx5wgh43f6uLhmaayM4qL
7iliISCfpuYkU+UXwcse3of+Vh4pd11PrGLu5F+ilhpR/k76PEX+jeE6ns3EmV1moQmnxrZ6ODLt
DVhzbNbhk6oQXv7YRgR1ZiJt4rsvWOi4eVsE/e7bSib/WohhSf6qcAGVv12rcvVIrCJIbmPwEZLT
eqrDSiJ6WRvYuW0OUNIGYXwZq51pt3ScxxvQNr8wARjMhrTRLCV19HhLoVkG/nDxHi0HzzCewY3A
JJrqPxKl5u9x3vAW+kL0QjlghE/0ZvD7jDB9WOT1nVaaUKaRje0mg6Xm9JBogv8bbQhxHf7NPhe6
EvLvclj7e59YSv3pnaViYVtfSCuxA5LCT57TKzzTUJeW0b9sQrFvdHEaGijtDVrZkGTAehqePOKr
VblkoZujOqg1IKl/NAQ/7XSxjuM0Lg9+9Z4P2HORHPTQQkZgDYhP+CCNeuCN1wV+CxWCWMmt5eJN
2QRfK39VwT2GOUI9VU0W+YbXK9gz+MEAgX2h+BYtKtPXDSLwE16ltZ1mw29w3admUhh1vn0EiK+t
6DolLavwfC0fv2SmadRkCz8QfellLh8WiWoVNHAbMLoVLF9/9d/B6qlXrPSlR+mldR3368ErLpIc
aQwVByMlI5rv+u+EyQ0mEXGwmU7/GHfTBh40R8JsEtgs/PDZhITKBnC5dEFeRXMSBFpg/6onGZ9w
TqBYXCQLwaD8jyNoofCTdK+JplekxbEDgC+iQhhHU7Cgf5wD4nURPZBytCTjCU5ZXFm5VWpzhKFj
Wwf35irS44JLuqJ087ZCcL4S6uX6/sxYMBCE61KiBaPAJiBDPYk7zOAYgjnaJC+A/+9llgUkzIQn
QaR6ko9bdjNyOlyR8Dm2pBzzCOUVuCrjidXjfgLcc6ZoiNah+mKcrZghaxpv7O156aRaZZiB9Km8
woGytLhhTfj3JZ5i2Rwn9g8Xspcjhhj2WRCU6HHiyvy5c/fQvwGfGAwUAKDpxw5nZ884snmZ3pqf
dajt7BZjTeLyx+hHf0WjViMfz3kj6ayAgBIXgwbGLYScfnYC5a1eNiZANBNOST39uggGaHA6gCFg
iuS4pwfMhQLUUA9o+3EXGjzhC9IieTO6k2rPye4MEpIIl7u66VkmksnrbRn/xIiH1BB5r7BWvsA+
SVAGgk+27qO0XKUDDvv6TDisi+VzvqUeWShG4rowwLKnQ/V/szo4e+Q+yJSQjWHpa1STW4SWyPBO
V2cX0sIofDNouka9byoUd45oPpyIzNC99qmhrwVCfqDnRzQrUVbWDzDglmsDELtHWLBRsqi3jbXv
W3wzW+ce0nv4fWJLvMBmoQEP1hqURGNsJrspPneJQIgrPk8Onu8XmThLeoEUNL4xmIPr/z+Weied
Hfq7RwA85Ids4l8V6NS4UGAclXWa3GTWsuUXPLwF/b13VvyvorWcdm6CW6rSkw7Kkfq6fjMSvI98
EU3GSxiNd3Txzdef8xIMEYZTkTnh3eeyKySmqfwhH/9IntCaFWZrxAtGwOTWAK3zoYqtwHfURfA+
fQXHRfgzhiQh/GS4QAwPkhQLGDZPgpSjh4K2URZAs1IDmvfbCqiiKhD8rShkRvEQmmGZUIc7fMQL
L3DsXccCppllcd9r1tPvchm7Vs9uWyNn5NUADTcePsji5RLi1BzuEe97Cyo7EmTvFGhroDPUA1Zb
SsoZxHUahavEIsw92vRx6w6qg1Bew3HrwHwYKMrQBoL5VbKv5KkcsdDSBVwx8S5RkuvFihlBDh1L
PXEKY61whgXgbIHOpUXL/rEVD4xgfD9Yv9RuLXHmyUe+7/v/NHReda6QM6EGyImhU1V9dODjYiRi
+WFOgY+ipit6BcY7iQSvSo5Z5keOPYfxGHjUyGuw+L0Dib08+Q+FXKHS+Ypt+fIERxwd7TpTQaO8
1Q6KZm919AO+trQeWCTpci/r4z3K+kHBA2GQeLhdbL/ynJDHnQYLQXh3rUeV2Y0hTca0lzZcsNEn
PGUHlB4Vc5ZcdDqNZSG1YLAjVkZLJ8SDkf3uefILESOfpPv8O09n0zNYwxuPyIF1CNXcqMsvJB1b
aJuxX+JbqHTVDZ0tPbmQ2Kov5lNFxrahHGp/NCRin9ygUoTDMFKuQg0Q2hc0Di0/Jx7ekiXnRPYK
AlqFBGRslzZL9lyliO3q7IWw2MXUgLzISpU+fq2IZwV4IIB0c0LsHQPe65MIFqRtiaOvNRxicQyN
+NRtk70fJpM4UN2OXBeh+5Ot4ODZ9cPYGwy9LDuyeSItnlI13bjECQUQ/oHYI48C7j/4ThM0pAgV
lkLzVAllMC48jJfNdiSO9NQJ8cUyYMr/hmLsepE8zMU98DFWCK2A/9X/7nIwr0sNvQ1A+MvdpFLn
TWTEDSGOAuLMqJdujADY8aJDmEtM9eZmPBx5WErMv5681QJG0B/dBDDvO4LZMMs2kovgcAj+jMk1
KIIeK5e0xhhzIP4G9wnZkMOlvCHQ1llKuBlYZDmUp+T0p4/RJd4qzjMweoKxAiU/gaTFdFLTEC19
vBETDApIc0kHnNzyCPBGPhIlzqHEibyhNYbFM9EfoCPsq9pEMv4Utz0sWtJnmoYnTABKQhIrGub7
aMHPiYjWrxsOMtAvvFBQOKRAtAtaFeEEvsYRNthNGibsmL24CcpxjCFcs1A8PtK6upbOZoes+DOU
tJMnb98GMalSzyN1g6ZJf4tNrpZdvG38RvN/80Ta0HorOpvKceIdo4oZDGbnKjiebup6UiD96wXk
H9riiSmxqSX6HAXAc2j/ebbZ+ONwbwFZOHp25Tc48jdKWXXmSq/CaPk1MSnIpmrJpfSmuwoOvDif
whH+WAJVcHoQG1aX5pOSzsuCRB3K1tS+z3HjzX/EjsjnVddBu9UhSW5P830+O6rn8lIuzWUGJc2j
oGXctQGkyWDXMJATQa/rVKmcDljv4QsLu+xl04++etu5Sr5HXQMdWiFVn6yERDWrGc6v0XCRj4M4
zkO5KlQ9kFO4ApfZyoFeC+H6Q/nqw1eJlPwwE6nA7Pm5MmfdqhX3/4pdyW77nxpYWeYGYTs1sQOJ
CUyBzI2jLZbpiYZELnjaWXH1BL2iLEn8FdYW1KEJkFS0KPOg50szSJvuyu0xdXz0oHOzDDOJbY9L
MdAnvnpsJ0daCEnA/Av4vTxPtlZ9n59wiwzYBDLn4JDLM6y27pJTBjalzahM2I1Del4MblmVUzoA
TQWwUeBYmBzKL/qtLpWOY//Y2hvkTqWLnD84LyB3U9DsUS0k4hlyxAPneRA71P+I38f4OIXZt5zV
EnuA7glrEI7JKb6tkLDpLwo0aM+vdZ/a7Cz2lYB/8ndhVx73te3OBv2EfHOASOeqITp7w62DpTuJ
NNqwPtCiu2p9Y5hbiUmEeahw07z94b7c87a71sOQxThI1Q78bkmLo6riB4QDC6nJVzHEdhuo1hXO
sba3fV/2Or5+c7M1+U29TtzGWTMU7ZB4OVW9+IvgsZPli0jbgYadUrkB81aQ+FYV1vRbkeybp6L3
FFBzCegsad1nEkqLXcmvR03dzCjVcxcOxVIZd9Mz9UDYLevTn/SOr0KJbtXnNofVGFIMV7tK2mK1
6NEO26WDByRlKYGLHf+/fAb1uGcSwhqg34CI6fmVYCp9Nq9+P+28KPEm9vm5hXggAi43zQef9GUZ
keVQvL8goimu3b81VnvAelyJlQTqBYfIQs65FYSPuVpvrEZtJbqBE9f5QgvHjStuqrQVuddq5T/c
ONa7lL0H+wQpWzT66GHKqxrRSmMeBtJtR3YPy/lAEKif3RVg82d5Gce9TkoPSZqb6AeAqbnPaXZL
ucwDhZ/jkPcJALcFfkBQC7SaQO7b+izwLbTMdE9MxWL/zHHAG3IX11BmFsA484MAptgTgX4LPoxk
oFo/UI2XpmqnK4ZZzFOTzawirnbHx+A+101hcdMtV6WkZZ0DgkNFnXf/6Wn9E7LiZUL6y5Osld3t
LuiTNmBjaePwOesfy9R9GLdTkziW7lTlCrOKZ6dDxW5glRBWb+dNBoLP9+WeXrvW4IqEldlqJD7+
FxMOd1Hg1Ymrr1iUt2x5AbhX5d97Z4NX4vd1qIQ2ydiWlpPMpIxGobXkzZi5UsR6xxzZYEdIRla9
MGVT8PMFaUmcXy20HI77Dud9Kzblnb5BP6tAH38MXJ5Wy+iE+YmOA/ijy5ZWCJHU82MbWiCwv065
nLMTR3C7l7SNWJD56hJxm/mbdZlET8gyhDvCJtTOr9Vkhj8sQJqjtfQNN8k54y4d2+NcplagubY0
plDrlnbof48EquiDsM2Twd3yPlr7YAizH9AkUFCb/s+BDLqT2wqJQNjol0zYut3r0DRMCzDg6gYd
vYVBTfAIwSmRwhpr4/JBpv7JYMY7j16ymfoCNqnnkRqoZOOZ3O9kxE57XgXbVfbadY+wwH91y76T
ysVhh239OYwUXX93Zjr9cUQzi6xrrcS1Kce0i4hRpwicMzzQhzS/eFIPHspX0z3biJIR897EOQpz
qPWroqberWLDYQ8wmqxjzCPWmtwfp/tFwZL37R6dOsm4A7fOtUtKild308OJ2eXhNEw9ApQAcsbI
tgXKy3va60wDJmZUzCHaLoXR+NfDI1rJVPpD/sdG5CJ4iUpZQrSkxfWSoThicKwpC0ExVUo1sslu
KUgiKW/1M6VTQY/MBM40nXiocpE9LOKzkHzmKXJxdT4buo3Ma1p/957iX1AN/G31tUnDtDZxo0kE
pBrXllDU6/r3A4K/SSHK5nVr7UxnYjutQbkndn38VkYBbbhQNsHiDHtdmdstBV4N7lSK+j+EX2Tr
DI4DMMAdypvE5/qYNAv+zecdeBHbTJogRb8ukcnIDUXJOi0Y/O/00I6BptjMj73THh7KwUzOIjvE
TqRKvhY/+I9ujzuEXEk2H1LsZ6r9m5iCWh3JZM45j3GQJuKWcTt31Fa5pWIseFIGTCtj1wLs9UXC
JqrbgWsI+4l7C7IXJjzANUcJpxq8tXATuyV2R07BUbL2tDnDXgwsrZVB8A7vCrpuFZxkKmW2U+FF
pL4IjbZn8RG0BJ+Ia7bA9Adwt1Xsp1yAWJJaA2xR/cc6vkIYr90tDGaNoBr+5avCGm1vRCD34I7L
7JSBU5W7gp9XBcsU6FaEqKtDwtXUbjo8da49CrKdycOTNmUP2tXtXi8M/ZCJ8XRgQ4OXtrIv5zpn
gp4YPne8rPEMIdr110CZ4LE8N8XwPWhIE7Thd62dtUYCzmI5kxekxcuHmKH9IslK709C5KIZjpc+
hyGO5NABA2uL1TS2S9N75FSRRyik5HfPY16zI6kkQFds0yPoqXjFClzRH7dC/9Od4M0eQdSyv2m/
oLzcpCGTf3bMRPn6ZXmSN6VRIPr8Wo2XId6TZTLRq+vJ73e/HizfS7dGUOdcsuuDU2aeFWUSMest
Kenzo5TwBFfVNP/0hMbr9EPPH8h5eGzb3sEVnVxQoIUUDTM3a6GAlq2OiCbwh2pjjHDGY6f69QeM
s0dQwQguHupFsL1bwp/8tH83w6qz9IGaJ7pX42gaCBZv8NuL5c1GV4CF7FvG0UV1T5ym7W4r/Xdi
8g3zsqiVP5CG8ZT3h1uRmK6H1wEJnK/jmQew4zDYBZkturx3nP+Z0TH+QJX3DsXbzkkV2+qdySYZ
RiKbpdyqm/4DoEvRYBnjEzaDlZCgSzd6xdqVLtmg9UAC0mxzDxoM8kVmVQIb6Db0JoyaaXxswuCZ
ZZaFDsT7QjPbb0Xik0m5+boXfYv/oXgxej3aNf4s88dgFruz62jP2vtSUTmaiW1oYgMAI9FzjrS8
GxONZaNTpo0ZMuRE5b0LMIQx+Iz0CvJ0wB2QsLaF2d/1896gAorqe8kwZjekM6LVhdD1n/0HpM9t
PigXSfEQH1EdcXYonBYyJnjb0h+jRGJ0QY2e24b2plhdRwtSLs+ZO3AZQrPcAFW2UmrsNql+xjkh
y3/Wk3WrBkC7ys6R0gvTIjwdfE24f/Q4BZDFV0rui6EsEd6oNmea/8x4F3q3TE0hfbyJMcqozk0G
BZLgkA8DNyif+Lksmqwmu9B+/j9EHT6tuQeB0pfXpADk0h1sCycRBkCY0WoaFHVEjcUyaq0C3Axm
GPKItZq3pI2DPDmF4Pb1zkfgzNu4FuoldjaUkM6FczUOfjwMwMm9QAopvZmJikXMrDQFKlHNarKe
24T3zuVOP4APfsE3xEEeo/rX31BrCm8xPeBLLfOM+icCnk/NUFD/m6+LY9/cmrYzncVKtrhqH0w1
wvuZ2VhTzOXRkvBR6czEPTxQK0ttEubJkvP6N2iMJs6G8NPAS3FNelo38GQAHzRJzhwEr4/GON4k
k4CDwYDtPavU0B3YFOEHCCYJBnLqsChPB6SHmHK9sezANQSS+/lzezRdYlRqmU86Kvd69BEM4VMM
pHqAYg0CMk6CEPQk9ZNT31/r2ai3Yf/OhpvCCkPQO7L9BOASGI6/N9mH9yiRgJlh6G6GqKfcHAKJ
mkAWwMnYW6OlnGlASnJ66trk7p677uAeZ2uTDBVN3ea4Hz3lN0nWdDYvG0mV+lS5fdDKb/UwVOH1
woDh2ZWP441IhIb6xUGzBGezOYwpUZth0Hr0zcbwWpaRRiIgmn7SoFhjBgE8AgvRNRN/I3brjbet
1I04mDSB10R61P/KrSjJ1rSzpgmO1KqMJn1shiupj4fgXLvZ/KRPohbNPgvNUwS06JkDYMBz7oRs
brgkT3ZBAxrpTwNlexTk6Vzj+28HCGR++JN5saU3Drx5/EUVLAk7NutPPxp8v59MbHn4ImY/MUUT
/1uxXniOgf6qx35WxWRltObxeXYiBzOvz4IwyHxEmqFy57Tl6OqzV3LvjD/WGJ8fmVbBDcW6HmFW
7Y0FJIlrhjXua8Fm8lnNXKXxtaQNXcXcHoqbYF4gXQs6l1C3mNf+zUMcmV6w2Z/jbqZwW/d6TkRm
Dy0iEjaCqSfYM3+0J8C0408yq+wMfe0/n7cj2Us2qT2EjDfNhwdQCePnyDpFIXLKyaAPJvXX4kIE
S5eXL8e5KnNGlRsEfhkNw011siIcBLyH9YzdhdQ2jnLGN/cNMIL5ygiYv2EMBGO01BnJU6anEZN3
F+Tq3armRc4JqBhjb2gsak0zfYhpIw4kS9DTiWvePsS2IE8fB8fM4uqP+XndSy7M92ItPbAgxuER
gndn5s9/xGdMa87EQfe66ZrMSZ80nmaDhcbxn2O46gDAi78GGprCjl7+PU/mYuw6QcIG0BYOXfjM
Uxb6uELB9xRITMRqiIFraHXxJNGPeww6LHT5ryiAe0CDhCW8yK2zA5k0eN3xxHoS6zDRbJXZypLv
KbLpP9DMNhyye44fLIxTNaSOuPazfYm0G1tcHQVuGnmzSPVS/7n9DOtt8v6SytGS4LJrRVcQ0zd1
t6iiC797prMhltWI/3awJ00BPBcFXNFSPHlxl4KCKhyGFiJGXW0WsH/LeD8U9I8ITsibOqdH6Tmh
o+JkyAqJLlroepoITTMH5aekXtVTUmq4yg3ctnqH+GFwxKVz7Srx3W60GIr0OyDq2X0QrQqnJ/q/
qA6craX2HakaZaBP2IWvI4p9e2oe5/ghWu62H6TZo/RwKXOxT3wves10xDxebPulNM/L8Bqhbgss
hOQEJ9q70Re4CjnGQ+dbnkCI7gF0f2nKbCr9pOZVvuKs0+KyBQvNPpGlVZgdCJDSnOLYOwy84IyS
fTWqu/sHkCLQA+v6SEbuzwvraXUZxjVM4YFOeAizyUcXYN8gCbWXMqmYwvE0KpnqwPkYM44NxkNJ
ccwrMY2j6CWoiJYN41Ctg6ACjz/oljS/tpwimlE5ctFs5kVIqZ1sSPvtLT3rQY1SDnjbtO8QIgc4
sFmNsPJR/ldhWfdqAwzUfFO6+H7/lJ8OzkYZMrVbbTqS7pX6zdJeIqgmpN+8aAmiJFL1eF8nBj9I
eW3A7CrOowEl4mTg31UfaKjYqYWiapp01jn0mpbEmvh8Y3A+Tal3YLkUiB5o02GAxcNpD+OYoxoC
+jWQWrPTH+5pdcwalOjO088tPGOEtFRwHRRloTgsGkSio4CNBlKDsZ3vLf3swqYqtkWu23figOYj
IYmPEa9VVfUPXSCiZst2B16ZeQpjjYXVQKNPFO/ot1u7Wi164DBgrfKQsUMv7f/0/VQpDJoIZMge
1FCYTrkpVLsNM38bRuVcKd0PuXiyq8KHyA3c2sNGxaAd6TCL+SyuQRkp+48Of+8iVt7EDOqCIAW9
gYphZhG+6mCIVDoF1KDKdRltemKtbmhHjk3iev/QzgBMK0p2raUEN3EaYdaeyOA3t8u6F8XCHRxy
25qrTJMDlnntnt7DxL/Sjjei4DK76nVwzw6dQlZVe8pjcP7+U1Jh3jFw71ORHTy4Um8YTygHBRo5
d9Jw/Y0OOnUMoGQ2HuBdyw6AuE5RENgVYQGKabyw8CFAYFU4kRYtZ9AU3ORgyHQ/Zhekfzy6FoRQ
3pCBJT/cb1t0Mc2XQVVtFW2KA77DVSU1N58GR+tyo4cr6oolDui5dlk5HQsfnujRRZ8Ba5Dg4C7D
QhyCSxZ/QbTICl2ks80k9LoB8U8FENrkY4TheDvX/sPugXrSrBFJKApCAqqm5JLNmVoBsp4g6tPl
u+1xpQASd+dP9Pb1Lt3yyCHIlCZPoXLIQ+sRObmaDAHzXrGd9HilIvGDamWf4QV6ze07Z2SV9cUg
3BSeAIXDXSjHQ+FnHQ/518lxqc4V8TTp114UkWXVoxTI8fa2czYwWYZ6YxVVYMbFWL0IihjhFs4Q
1Psew0WvAsywe0N+jHrTtcY1mwgZxEDn6kpGk9rFZmvQlm1PDKs+BCnGzgAcohymfrQBUbEyoBfQ
Dd6o9t3LNcOioJERKF3JANxk3vPoI3iDn+NV8obyjzzRwh8KausN6Ys/lG14tFUK/SIOo/MuIBJh
rTq6EfdaEFIRkCjd5cmpFERYQeSgp2iZHHI3yXfXX4LGsfJYvc85OZaWtaY7QnMkLfPHQHqMEJxr
3yXsBDexLTOUpAZhxS0ThPz5Z4Q0ZeNmWUC5kCFxsxne7fw9qeazCEe9nRPxcR6/qsCiy4fbwUSS
uoT802Rt0qobCJRHPTDH6Ep4n+v/2VsahtJaAjYgDBFxn51Q23r1hmQKg74qXe/N4d+BESfAdmMq
mUoikvsJdiW51qViIRkFJo+8dMQhaw3uA7QgafhnmOqOOsMZjgkaHmfpkh02IRJi1+4jmXg2KWGO
gxCgBj7cU+mGO1ZVqSMn92YMNzb/FhpcUYFGodWf1CgmhtNergDxu70DO2JteU2gqpSZIfnEOewr
Ulc4uxGu+MnrbxM6eOT2rHZV+uKrZB80crDfJE9n8fRPH+fOXRhheeGV+MfbRcwYbMMjgrcYLEtX
yMP037Kb2OKEPh8cVF2jTgReBbRf8dQbyMw8FxnNBOTeFNLfgsaKp45KzJQJLoC8vM0rDQ1TWB5a
gj0jF2i6rWWzWUX/wXUbpJmOZOaGn1nysEJubqJdVZRnf/xOqrw7P0SG1dRPzG+lSofKlT2OJ5Ui
loQ6u1vjesDHV7wnsS9FtmkkDLlzWfVsQcHwB8Af7AHBBVt7NL0BcEaL09naTvMbZSdyF9/PZhum
7pGlJ/mWEqG2nSz3k48ZVQv05/Y+zgzLaCepHuPooIiLl4/hHdiuts4E4P10d1FPjKdYPnQismz9
jnXt51g4+xnRP9W4VaP5HLeUTU8qxpZ0enl4yF6TT4HpX62yHqqDBXm7trjH/RWMgiein6odMnlm
RidVgD8/FRsC4rHdbJVowCcBCVFGGO0JWefMnYCTsmVbbCgr5e13Hhxv26/PpYxO/LkB+sFGZwyd
jRkv9yx+M8e5ANDPkVwth6Cu1Tx7CY2CFGOWcxGyzQc8OtVORWVpv/ataAe9G5vISfH3Su3KDeeE
2uaBQ+VTTia8nJDyJ9k53vhIHmy5bYjrSa4DTuc1n3ZtG+3Q7QmvmdF4jcTjzD+t5nEuR0tTfUaM
WHSGXE5FqpXJv8/0CbWT9XWEpjED1rjGiHSRTTicpQZWnUEbYGIpSsrtW0diOhj2sknVNQGVxSMN
yEDWUVP+sS3OCQNGDFu+xhjb7LcEE0fvjAkJDiaLaqLPKqgOXO1z5h0Bb03zDGmsQ5Y+YnlPDdS+
6YxSbcelXgKjpf3sT8ImtU1DsYE+6RD3PNLu9zcehbFXFnhkJnQjwx60/QQmRuoeSs71aY/Cw9O+
hsDK+GtldwSf884Awl36NwWq3KX3Vb0h0ti7p8nt2a20fb0Kc8t5S31DLY/I2BBh3lKQZDZ6XxOi
opCj4cuLag7Yii2A/C8lvZ60731+XZG9V8PTiLLgwTpMIBdcE2Ly5/G6GGPX27EdoHULUjz7f9fe
5vH9zUDTdCYq0Tg4Qqtr0XMLrnDXAYx+wuFkYcnj6iIUiCNRqj2B6Ke6HPcO/T9fhBO7pPPqTjGi
hXsnnZGLLUbVGI2fDFKVha5uYhw97VJP4ToedQHCHq/USrMLJyt+ERPbW4uFDdV6ExYURy6D5mGE
lY/Fq4Sp7cU3uAFFxjZxXOmB3ECWHooV8+WQSfPBsiZLTzIRWmvzAwvWzhmjwz0YkIess8osYUiB
wprQtXy6sWqQlWde19C57iLig/g1AMQoNukFIfsMk4G8dpqnxregJwcgZUwaQp/+jzIZ1VTxdFvF
o63nyLN3duk0NHF0FSvU5c+kplqyk4LIm9PxKr2/1pmHyTe+84MfoWGdNydRlleEjKgsP0G0uHTc
0XBnBrBjGwOZAZxyw76CjYHzZ0ik4Yc+expnlQSrHyyzS0Q3iDkuep5q8P7VbhvEWojHCHDvwyUa
DHv2gQW9A8Whp8/TIpOWReFttp7sc2psDxoxU0UXsimMtA6GgUaaH8znKkcNlUlQi8lueNuneELX
+hPNS661nzN8wCTVV08mQbPM5Q3n3GiSPTDVXaNG+Ud0MNGHLWMhcBTTp2ZquXhQ/jXkRf89o7pv
nnFRqEI2duEzcKz0aMHFVU3XCD0asw7nNfFF6m6vb7335Oop91pDzMXZR5I5JPCwE/MG7ox8VtAg
Bes58bpxpQlxdc6NZGZC5ud8ey9nRxMQJvSbt86gPlotJlLR22ZOUQSJYz4Ft1pdSV2plrG6xne+
mzXKt22mnOVqRoG9DhRMBo1LtvWoUN/1FRn38A9PbJwiuugQSJIFg6RWwbpFVfqgoEWUXldU9m6s
xb0i9oxjHzAeI+I1h313J8rsvbHoi82tcceXsXK6NLjLQ6CaLcp5LB9NTkb7G8zV+aQ7fa1kzPYL
5uh4NCn6Mezu/5P2hRhECJKUH/VuTWSY1zHewTsGL+e/ZOs2HelPn43sEW0i8XY304bk+SxYOs1i
6VDJp+AXAQkr5hGT7cLdc3h3Wdekz/BWNV+a1MnCR/7AxMKyfT5COv0oOPb/EElZN4mY75/6+7xe
BawuFZHxrcoXHKzdkzEq87Xnd5o3uRG3yp2+IwCRr52n1VuQaCxf+bS5iiqELlfM1XnV7o6yDZ0I
TNwvpJb7ua7c5yMlWI3rMZO219CNdA1PG7MLfaI9InIrMR1yfRT3uZFS3+OcJwKBZ+atrXbWCrRB
dO49fZlmJit6wdm8IM72gWsp61ZpwHaOudJoHODbC5IdsYURNs35L3KBaXe7Lerb1LU61I813x3J
PQwYdIbXrKiw16UHsT0JT4eVzsGKFGqmbas0nb+nP3q08vXFOeRgSevkhZfcB76eywB58pPigspZ
3OkgGXA/5BvX2pkdXhudb556tCwqWUCqo+C+mzmIUiYGg3UBzbnS/RFUF93TXTioBGYIF2TjloWH
5AY9bs/ME3KkGNbDFjPSQtLxoPpSCHtUB2YIOS9DCzhyWnyl9R2TKZflx0qcdGHegM1cOm9z3kon
Y1t0qLI6YPZKqc7B7ldkbgzj3AAV4KWZ8O6MBl3j3Sw01fHOOeHB858SOnM9L+L6tUTkR+I16UEb
ySVdxjPt1jkXIOSRGtdzcU/7RvGsFDyBMwFqoCsoOC+fUcc7KRzK2zHiQVIW2LjDs68Y/qYGCK7q
+2ZJmO7G7PDmC0M3XmrWgdPBM9D2ovOlKVWQOBQ2FkSVbnje+5bApDcVBn5Uk755Y9hpCQNo9I3+
QF0qod9ziMlo1uOhf2aFrpsfIZ2BhoUgtKjXk+m4RBCSt+las4s1IkvDOiDqss4U5zvTxsl63B+z
utt0TtfihpmUSyGqzEELor2c2OsVhD2HKxYijeCxANFOrTanwR66O/bPeBrcxLqbqu3JFnZ4IIrc
I5yKDTLZ/DZtHg/th4fWNhjiq5ZNwUfaPQcBz5Q/7EctSFgGgsVfjwss8bwvy37lbqHDb1Pqk/Nf
ktB9I8Xn+rRRreZQ8TSAnnspkEBjVLpkoSKz4sgAprUbuGKx1eUI6PrL5tVuHzGKe7pviBspS8X4
1LF9oJk5X3jTP2zIeIdvNxCwRrnxPzQjlMdOl+4aVz9/4ekiJ39yMOM8juin0i+KDZjuF08rzBzp
PUTXbYArYn9VHruLM3amdJ+f6xU3Get5vCGsThvDosvu7tvFV23PLRtDm4UB1dWssIeB1GgtXB8O
viWGakeha17XEeTz/1z10Knz2fFP7rrgzfFpLk39ncBasGVCD3RgwF6tMRI3NiG5SCRKphmMkPH+
htwROz/ll6NEGhYQAsj43N3P6PH3+fBM1uOIwuG5o9I8Tpn7xY4QKpUwHPdUoqttdoUfVTwYsl3s
Dq6s+7O9ghA8YFsV3s+s3DjT7DCTrYTwr6dgxX9vMjmGilwgo+q6MxG+SXYJ3/qHAUpbo3ym5X7S
AMWEHFJItt2MYdh4MEk4Pz8Hib7iv7koQ2qPqLSuEyys1p/CmK/UxgC/EjzsA/CUkO/RNt2Vh34/
zu7q1uNiuozMP+F/HMM03wXfB5q0rUIa3EgLxENdixv30eufXLh3Is/Z4DQ+o2BFbK8UDi8WwGvM
3F/3jr6ADiwW11xTWsy2kSduNQtRxDK4aFC37Bro6ksAzNCCOCBUWYqO3NHIb/vlW/ezMNd0mSzs
crZgzShKKaK6YUHaV+jo/3P/BCMuy6mZ0QhJCXdMla0gVpMU6VbiNQtSqSP8FI6eVg0e8KO9sP+k
iwYaMNdidrw1/wxOCvmWugxt3BsyMuRnQyQzeBLMAW0kMNm60J5iIX/RvXfxQghOODVjMXsQbL6x
nvn05WzUNDi+3lf5ndxoNy8L1FnZWAQdBI7SjhdwiHLbfscNFWPVbljfr15ETRWa47I81B7XJAQK
reP2GOKd0tO7m1mSF3Bdrt2TH/3GDc+Yn6zp7oQzjWBDcF0fiJ3cMmQk1xdiyZDjmBFK3c0kQ8Ph
Vn1SlM8axk6cBap4J8o7PAAmElLk1rVyfpp9c7tnUgbFBzfs+F6rNVmAP7lcAyR2+1zf07a9uia3
geUbmxXNupKOm2jYZRh2VTMnE+NL4JUyBEiSKFnC00E9HMqk8qyg+Qw0Uf/cTAa2Rpvs3DlthXsj
H9RjCCr/Bqw3Q45anA9GyV5I92C63EIJWmC8yQyX6YiwiI3OUbQYPl3bCHaxdf82QH3AtfkXVWER
YWmaxlvlogsFgzsoiyFr9Afq2cCoTBkCXPN4CkKJTKL9NHRRHUOcRkN2a5bJaUMVwSoKLku3fKSI
YK06ZvmIccrAqEWcaGcE5kpE2aNmRNEljcjRoEgVZ1Q2KZiv78O2Q9iwYx4iSCYmJF614vNfznca
Y6usTnfykDah512SFo2YQUfSY137TLyvB1y4xgQyIltPk33yptimO7JjSMWMzJbadASfnYPJAdnM
VVJiqdjzzh+RfC2swxjRB7hVYhtynib0rTb8PLrMR1/k93bTl3vskbbWbmMGPpGlOSz4ePzZSGV7
T37JPVMLcklZxcE7gWN2U3X5regQSJ2NS2t2w/167cDYLrd+rR4yTwGl8pOZbS8Lj6j/BOTOP4/G
cedXca8u/rr8ajWuIXKs5WBfsCIqp722JkJREWQUZ71IkWu4tZNogtxnfFUfF8gQCm0ryqYDMXF2
JB28mLyWTB310dBUKNilkRVBLvX0PZIno+qjqSminFzr+bjHRqhlJnznw7YARuAfu+o0kYrkRZNM
yaw4XjygmO+noY6j1eF/roZqovqrP75N2AbTG5UCVRcmJWyx3HDCIEuvSSY2PHVFRFcU5cEARslz
HqeucMmJONg2tnQdWqLhi8/xM+ji9bxI1ExjgnhnXlaslYnZVoQnkJ3aP8qkmvCaZi1PO1Ci0+Ix
l1XR82uZ4cZme07qI0E9Sf+1JuJyLB+3fpAczy5UhGecagr5xuldy3eXm0CptpfO/foEUSG0g4ZV
xgjeioVCMMD3JpQ0K3/bc7u430poP9BONkQM1wUsYDccaa1I8vS4nxZL3hDVPZ+afenD5ajnXPsN
U+nnoU/EURMSnwAYItDKUQY2ymV7H41BD9IjV1bO+r9ZpuJNhfORJs6bpeh9h+x5h+umIAoY2pvo
FBqjAvfmtTibgODQ0u1U3ax+HpRvJ4p941uOMEzhb2in7GBGGpYdWWOPy0Oo9gx6LFHLu/ggVcZ7
J/CUV1UbYyEsZNRSCfSMEtn4LA26lWWHvZjr0d6Kefs35FZHtLWEWUvPpMBfQ4oFjTXaSF1vmREZ
8NMJX8H/6M3sTHhzdBl7BGQ9voyL8pk2Jcn+Rv/UFkWJdxHjdnfqkmV4gcON3jZ8fl+ayg9FP+0t
5e9aQ2H3WG5J3gDzfuExFjUl/4ksA+faNJZ+v45Y424RmN7KLXqzq4dVq3NBNGjDAPz1R29BxSFF
Nu1kCbuIzTEFQeHLQ/DY+91anuoQ6a8Nnp4kIAP/nGXoJP/b5HDpRO6g0z7kAXiC5iaAyO6xqVGg
4rbxctnnrLIR6xbySDDt7wX3Of3i2Ad39ioxI/A9xa/YBdex9iT5RhQDOuxC2deJ53SuDKbUdtcz
x4NOrdm97vGXi7n6kmXbZNwGW0sCce65/ULEh+e4VDGqEYC8a5Yn6solws1/oBf6xdT2uunBZDKH
UabFjsu0MIDJ6R6+PAZpKUfHj/oX17vgDHEvEs3qJjLYMzkcAiphMnwkOrww/neyA2IQwi7AOcVQ
/f7wSySaET00lKUziKyTFwjaGwxH6Y9iYlVK6/aKZAVqWO2fCrTHjLk32YFPVLZzcTm19Xiun/Cb
DbvPtb9xPA/2bX17HOeB1bkzNBWG8fbeYfaAQDZhznyeRDCwhZ6WRpL9/W5z+2rXpscGkDwXPKLQ
lVq9vWvrYHTPM1bk/X8Zi8PYUn9iJUaBzeTBM/dch36deSQ3lEsIWu/80makjNYU7qJtwED4qT0H
5QwzTBLtID1OaH7QeKvKRux971ps6oL/zO0MV+NGPHeiGMey5OW0hDCdi1sWWe4xjgNUNdH1R580
hPBPc9Et+SYBRoACVeLfKT/GkQEeIoCfpVg6UA7IctUDo3rQ6LZa6JcFvJ54ACBGvhWVLy+DtUhi
pc6ZRdY6HWJVZFgg0mhRK03sV6MGxXT12YIv2GMUegshB6SFvEBALAfA1h+/H7/q4I3hwaV+iPXE
24X091kkUUNhiK5/KTFNddFrDl6tr/9oKkghqWOnvXIIamkj3l5vfXrNDPZpn5xgwQpqUgOPYKud
0ifbYQX3E0qiJGyr6YrptKFr8ISXerb5m6Znvoo/7Su5OJuAfJ3N5dnC6c8KUNo1i+q7ApdGG9yu
vT1pP3q3vYFsSYQdhi2+nXkNb+jVtKCb8rLM+Qg/YFNUZpGgoFX2RKl9UlszWS0RpYbVnv62WFQl
RiX3lfoFdDjbmfn4AUngcwK/wnxHySpRyaQcVDgFE7JylRvCCTwETTrEczE3tkPZbiuvUDSrMRVk
bSG6PgZ8iIlbo9aUm2w7pwGtdUrH9sM09zVCfO3++htx4+GEgpe4qb33vPOeYrdnew+OImhFQNG0
wFSLeCN2IEq2ShdGU81hW8ozMbNPDWpgSNn+4FPVLJD/gBkX402J29g3OLiJlPd8rCHqjKngqqQu
C8Iq1o7fQ0Hl/wG3y4xBLOh63yLlVcs3vljHOU5qK72VefZ6FrLfldxP1gFZK3wBRvDP4qHGyOkl
SFzs2FxRPxh6CrcQP1xvqExdwrVEb+Mkja3MNDVO3mMPEIMncVeP5FgBSk1Ykymk5aKsQj5mU8Ph
YgyYhNil/esSIeV04f76LgQy9hXItdkGIO+ILPX8tEAYKaCwNwPzU+GiMSKckacy6Q0P0H+THZvW
96Rc4di9r+bR3ukmDS1lUlb78gv00Lk+2x8UklKKO0YVZ3aVwUXkMHnQsESFUWsRHZz9hVzTtmhi
CtWgJGOZq7/N/q5pdn8HLqFAgcFzKnQ13NtgfFlL9yjVta81VlZadlZ9cs+gs70JY3e5rxLilkOJ
NUMwd2qJhyGyi/qTdz2r6ksEKkJKFi9KgEf2QXyArNf1moLgl5xF2xZsVPU1FHpo0WLd430zMXrB
zvyeArz3+tFuoodoVAGr5UZ/ncx1clo6HyFCVGaTkq8ogXG2j8c2wD6MBwKzaOIW/I92nLujlg8w
LupRPcxsG+eGjD2lR5lwofZb3CvHBKxxWV23lHAjBMGfRv9f7rtsiCXd15bx2m57E7mbHl8Ly0Rb
nhtVUeaiTTYB4XKZLnYLrwyGupycDGpI9emYJ6eGAgWD7BzNKhT7pwzFGF0UzvJRRGk8sKXIliYx
ey79fatPTKOQ8Xpn/85+MmGmNRjHYaej0YCzWm643aTe3DWMBtdTeP60YlVgVxToFk+F9ixdyYHu
5J/kkNmy7KENbgjcCBhY1STSCVWB1MY/kvQBV9pmnrL7U6Yxl2HD4K0SUkm/WfdNLR5k39Hgfs77
X8LmYWBNzIqgl8eok96CzjM3KKwORzwe60UU/IHFpgy0omiu38r6YNb5U0JYBw9TOKxkHP9mWTrs
GlUCGx4sb34Bt2OeSAjX57emE4u+/R606nKKsWH5iC11mCy58VARu39mIVLBTHgJLn9l3Uz0lIF+
FI4LwpxdWO8ebXabEDaLwovbSIKWDPxcUf0mNqd/DaH4EmC7LXkI2MoVIIy/M+bd1crSSU1NJTAg
Ow+/sdqgvXqackJGtuiZkqB29ol7+WOkv6rc5d6dLjtl90LmJ/HofAQEmMoDO1VU5nd9rb7SnlpI
3fn9DqkFt55hvGae8U+mG5bJ9FNHHOjULp1Kwlfu27kKrMTYP0djRKuWFZRpuI7ZHto+ce0WjrLg
I9wNMqitkYflFUxOgWL0oVAd09ZymPydYOjsBXvYLyIjP2clhcofkbZj1u+1Ku8z/Nc+zpV04u56
b/jlKDqsAwi9gg/sHmPseyNlcxXiTNeDPIJgpRhnOHIRS0mxb+uVFeGbrJTgiSRdxXU11QTJ6Y6c
yozljikP1Sc0A4RxEIvEB3XD9lOCClQA70Qb4cyp2aMcL7w3sN/dLDQ86uetTrQkf4PynQX7Uhsg
J1Xf7aUhMLx0jpbOtKsOzlPVASVB3sKbau6NnYuGofhefOU0JqW+N/t7vrK7YTdrlpy0IgJW6UkA
+QxfSkXcfxWg+LhjW7JhswWt8Ot/uiwKqesIFXTvMwEX4QpQZ6IHX9zfP2vzZQe47kAbswU3QEFS
1CdPxRqUNtlbXyy1PRsvDUG5a08UB6gREZztFudlbXIYW2wfN9hGKV/fHxQbSgUm0WfMiEcPLPDy
+f1cuKXP85xc5ui0Z19SYAKefNylG0G6x27ZEzd36RGaJLzlsLVxRB9InE/wu7uqIJ1iWmgsa1Dh
Rd16XYMw4iYCUL/VtQA5oVEa/EOX7xGappiyJLfUtCAd7Mvy2PBkp+ir4RtVX6UgZvn8+MbEGgnQ
+3mg7Z+ECEPPymqWuycibLkyvrRiRhXOY2UBeSB3g4xku2B289Echn8EhVlxYH+0yhqNywEr+QZI
pMs7X4VrUyprdFsXpT5kGWW2lqCUqBsiEdCgpYC/J5uLPaoyRSBKIhKiPYqxZJO0gYN5r9vF7zZe
4EABNDuz50ICN10K0YRa2lPY2TRdlJ+F1zI7GHNbyFeyt52uzcasBvbOKR5FnWo8VPDXpuOUh7qB
Uh6pGoWLiAl5ZzwDIZhvnMO3f+3thRhdC2V1B8ZRDrEC+HEaqK3GBoIsmAWdGaomnFtnELuDm8Ko
n2DmSR1+9V531oAVMSExBxRtrioxZPRBCT+8HzfcFwBHBIqKpIM2PAxh4CUxV4DWuk05SACJRHU2
jDS3EKDqGcFgbVebwu76YImgsBQkkQhqceC4AzDmXE44gBt9xXqxYtjpeq+CoK6IAiEddV+JIMQi
Iq84zlAMAw6JXe9bCf+wLpQdyjlAnXHhfe+4ksxAe10xtj64FGgfi06f+wF0jYCD2jnDZMROwhTd
YyGpM5lkD3WTIkpVBwMLhtoTwv5pmPzbjjruzaFvAimovf8CiJXpZ37ibnxg3y1LPCpyz3Z0VWce
ogUDrUxjr3FPiZcVSUOCaTHW//z7uznFtRP/7VIWw+BT5w1fDgkjI8gNk0SwMsOEQijQi1irAwlH
HToXDvjsK5GVnSNnIF+w/TUcvpbBRxXNK1cuk30PZyFdMEkxklALHBVLDj6NpQ2TnpV78m6yZsKb
Oek6YGyaTlDpyUEPzk5w72ztCk+ZVMaaCU30j6rRwoEJeiUfUZh8UctxuuTMeA6v/C4PcZBTVy7t
OT1t0A6t2+Iy89n0UFUoICdy+zEIbrh0OrVTVOrEgKUAL4xN8zPd7yMh3T5nK27x/Xrztzw8rUXO
ZolHXzWn9lpPN0YjjAjrXdjxiaTQXKpwdsxm5UQdjeJBMmAlmoP5KOfkpTrOSEKNtiwLn91acCxX
c9BmDcmp6XguuZwK1IzX3DUWMi2j8uuaWBckdo0yYquDCylZ1OdP5bi9mv0lXpIyovoQp6WkDvlr
Uhq95JAWu6Pmflh1ucKk5GrKl+pvDTd0l2CJXpq2Vvn6cjcMMpPbwdnCW/K7pBMkHi/YI7i+WQcW
PB3DSoTzFfAAWo6QPxfMP6snjLRmsG3qm6RkWgTy4yAAiKhOd4RmAoYSnEythP87mIv/J3eCLogu
gIdJrBlYc0Egj5OtfgiqXFU8oM2gbKQkZ4vSvffsJN29zP0LDw8VV+42SM7Y9+ZE5s97rqQduYnS
4kOMgoDOojkEl5DIcm5sz0Ta++GHJfTDn/6iWCS+/ybBzJf8eoIg0IpbvOJcd39zLb4atrd402hL
Z+l6ngztm/+iGiiV6AJWGWIxvWXvWvpw3sIUN8hdL3Fm4cstye3Ohvs9bPD0rZInVKL3s1Un3Krq
z8W1i2GI6IlM/U5T+46K9l2SNDony+EDuYmQK6YOvBn+PAPJy9RoYMH0md+1NfTYuFFhMTH1Q7Tx
R9kRMl/pEZQZ/2JzShNnNJuw5ZhbpkJp88ZW7l+1FKOuB7xqTpM/3bfp4KfjWa04IQCJ1y1Pm0JO
Mr5yi1Sw5IDL93T8vSFW2MWAgo+ia7AAS/Nxobmm+SUl1YmbSr5uAS9u36TGTeq1gGwrn9Z60Gwp
cokhCLpmBU7xD8ZO6RNTPBY+hXBvuBWvBOr7cxFJAV+eh13S1aFbqiLLCWLIR1/X6PlYUSwbqt76
S7+z7igSZsaWkJAHjBNnLw3SMPk2ORbhiA/Oz5cgNn9t3yHYJKjexEQOtFJw9COGO5hiJqgTsPL9
/kXSRwJDZjEfYBgDPpB+eicp4pqkxQrIhErexX1xF2xVCOUsEHKtrxjgGdiVOMosKGbKjc06dLCD
sWgNk3ZBrmDcmxuTq7r8ieSQ6l03pNuYwTVy3r3FnnNUjxrKsnQ3W53LsX/Njsp+QQguEgZVbWoI
TiQGHI7eaRqB3fyAF5UooSG1AMl1MHbfc5SdgpgOdhae5C0zA7BAAnWcqQawmsTPM5rqs4NCBHuU
6JDxftkrNqIactzKp0u39gtvEUw8wENiZDUNlk0YftyE6iPqklTzmYRQHQpmK2Ps8f9qIxHvDTY+
tTHaq5F/HmcQz1Hg7/GQNTyXB+/K6xDId3ljtlaUUzN72/PTiRkFc6s7/9wH4VmtXNElFPxT1N4K
yCJAzNRT6x82V9+Vv4M7K470WAtnmMi6iPa2wEIIRRk9S7yOoY6sjOH+62crJq7lzqGbI225nNHz
e3qc6KyHSAA9Z1NHe6JaRBxizcWCNI06dya71tcptxd8gsibUgiYO5ofUEJYBs1fXiL/8HAkdf6H
B1p70GlDqXS6MGPrBZ/v/UfyWhHEE0FrGdg2JNhueLZn5nj7V+0gWRK+NF671WfpBjKB9XHZhQbZ
Vvq4nLACInyxAd5k3WMX4UbDUhJyOEaqioYEFNMzK0jVtbrJqGjP1UH5dC5WyVSfQCbjpYmZW7BH
AIxjlU9T1/SBowLcm6qng5t8I2n6Lcm2mIXVlxTu9Hli/0/DFV+TSaRAouL/JpgKliD92D8fTvYc
v7jhtTAxc2lVc43Fv12x2g2zlVck8cvq+AhAZmeJXL8LNvqZ5v+sO2rC0UIHn63K9XIsZGVCfroV
Om8DkV0uFJqdkxrdtr4kZka9G8oDPqlQr95SA+Gr4/bnD+lQYPB+hUaWTRE3r2hPWv15P0PLE1c+
n+zjvKcdvdMSUtCinou4daUEZchWxNhrE4s6lri7dm9VbqEXzZ3LxTouwov+R5pYTA0uiRLIm8K4
zVACxPsBSmxF204VxfmpCKCH0rX5aVErUmTmRLb+Rg4Ir3GoGuStGWH/sFG+vOulcJ/8JZIlL43h
FuCcSzNBUGWlm3eeCV2CKTAf2ulcs29NgfbxFuM7m2wwCei2Rj3Dm4TCWykLPp0NRa3vT+dOOY+2
7t2KejDieUucNJtlfATayG2xB4gtMTcDNqEEnNRf45nbFWOOH0urJE9nK/KuiHaRSNl+QqtuRAfK
5GUlY53F695zno3kNjUp5eyJD95yXhFO+c5DqOizMwHIFK3y69C1rESakJVFri0xzY2XevviDeCq
QRE0x6aUFeyH9SsMYzm+sDphzLRNebxwGv/bTpslpCwyBLLSAyvyXOiYO0dxoEdFc9oY2Q47IXxw
2o0BXR8mvLy8CuA8jsIzRrN0a4Dve6dA6u/iSRRmrUPWdmmrykYrwCj9oIJiAGxe/N0O61A1Ccmv
3oFK/CL5XzQBfSkr+vBuDv6Bb8g9/fSAAF/DLU+gOFIKO7mzRF/cUZhCYTAzEKQeX7JEExptwQcD
ajXxeDp/Qr9hO9wj0VA5RiQSeTWo52qk8cWYCNGh6pm9xZvJk0rkptWeKEod9nB36FSuzsnSlqDl
gyxwPryxU3YM8VY8ng33KC28eAOBsW0ki1So3zTUBeeZ/fgpaCc9CZPmD06kllP5RU50PT5x74l9
EBPG2y29I2KAZA+bY6pZBniuRfLDjiHtWiDGugecXa0akko8GjvmWfPFF0p2ffzEluanbgway7wd
5uNvNEbkEtA9AoGuU0ilB0tGvXVExqZia34O/ndc66uxkeoVLW2w65x073AYhQGViHycEJ27tqUC
gB5XsZyuEZ0rsp1Idw8wov7BaTjRtkguPlcAhIPEy16Ww17JMmtpm9/GQvV8j594QAXydZrH464C
F7fwJKp50kxAVcuDEtCGEtvljDr7h0ghw/T8ctARwue+0PGE+DYFOjDoV2ZuU6SL2dU0IbM7cGmC
PPgYRfuRP/sS2Q9LnZnbdJL7L9XBVwbFcn4sE2PHBOSWgoyASE7+shsIjZjQw6YWCyPr3t5ddoB/
eK9FqP1RJ1/uI3xPH9V0N/SS9iEcO5ou1EnRSeuLezRh1Z6gEYkeRc/MtpVvFubgzlfl33U8ym9m
Go+JCWWpHavzDMHY1+UZ7gf8bi5tq5ZOYa5IciB71MOWhca7oXdCGciEsi02MfQhYWE2OGjQ1uwi
KQ7GawhpOuPA2KHzzcRMcqV9kzrJtb+mc+y09xzsWqM0zlNHduD4OwCK0L+nwQ+NADOTBXP2B3jn
7B5eABm9uHzT0RfK+E0EmkO4FgsrKGb10b+uY/WhEjcQFF/ZWDZcs8miCSorJwl0s3oaAKYeHMgC
JQRkoC92V5X7f0v7CLrTOYutNsJDsRR4F6nxZHkq7zBM91r1SSThTCy86O+lKRjycJVnXog2QHmD
uPDeVlnXQrMIJx7RVM6Z/P62qmBZ32LWPwgfTauvr27qHS8gUBypXWAymNQUaMF8RcEFgpUgHmmB
COIiDDGrxuns8pyyVydWRXEc3f1mTDzcJbWQSovzKBFGsLKajnbYiBryte2Hgpg4+y1HK6V6yNMp
6f9R8vRU4S8Qj7W84DLr0wI1Vxf8GXHvOzYKhdL8rwcq0lGn7TZy2TO4JaYy9elQtS/kgTMtBD8/
aKB1JefcEw8y036ejeb74g/Dmd+ec6oHPyBOI5jDfUFY25VVriK0paZiF6LPIXTqwWZtmA7tGwRT
N3g4/dWz/acyKRrGTzFtrpLCiWpqzs2YbvZjuIfVfPLMsrbcs0IvhNFgtO1DEmrShDICb4S1cwwN
Bht3TIVEOxtyNESMHLHj2p0jz8yTOghio2gr+G+rO/wdybT2ICJPbExGIvBrK42VUVU+u+XfJETP
0gDQbJnC2Kz6vwg64L7LyRPsxxEyc0WaLuwoXLx6248I8f4lw1c9J1Cqs4nZ52fgw0IZ8ERRWIeJ
K+tloS182LGYd164V2w1ezjaVyw/JsoMyRP32e8Vx/RCbo/ZGTJLAPQowH3Ba9ldGaheGRJwPhw/
L5gESWlsPfTMFEDViIUEEoz2Gkh1gku6i1kNLleb0X+Ra+rjRH+pSnQxWg+c+c2u62MS4Fg6Ou36
vMthpvPZUv0PgyN6cuSmOtYi9Otg6ue5h2NID/HmzieLibVjop+Wl04oKlqVg0Jt07snr/Kz5bfo
Q3B/lDPIRPwOOSALWV19Df6izO/GnUUwPYCKE3qmAWhiVlwXnlP7ifDxFeHRS1qxTbTRe4ZFkaLv
xlI99NWZcsPf3r+GvXIfBX1HaqHnbLVS+G8mWzXDx8XnpxI2kZzq8aLpKl3CQhNBuxvXjvl88V9l
6w0u/9ziYipGfhnRGsLuOAUaL6GFrd/EdlqcY6bHZJpaaYpKNFvXjLhilrQaCDa6y4Bg/7yqrArq
8VMfg+OHr+dDUzf+MoDn6/keX5SR/evadz8/kGd4z8EiUETaRNbBewels6lGTquvr0vc+tv2apT2
I+Wxev566F0BwK3aeaO7YAY8urHCu9k5FlBII9RjePRuC2fZf7Vm11SE4iNGg6qNPUBUYLuH8T1O
637pMhhu7sAsKzPvC4aI4icjTjfgV0i3JcvysdkvGFaLDfEa4YnzE15+MaPCe58j98u6LLJbREQI
h7Vg6Y+cu0nTZxwC8ckoTCZh0KVgS03PM2LG+RdGmCgitq5OWknD35C7lstaX5zSrNj0n6DaCqvl
NwZb4Z+72x/8ZP77FPt+i+UFtJaIkBgZTrlqeZ5+yu9uDQYXpmBm7tmFeZf6oqgpHeLhnsw34zQU
LbQyE5sWjy3CekR/efGb9jDln+MOcSBx+YnsCAsjl+b9cK110PoSCd9vBuiEa/2J8L6BayE0gs6U
Z2uj8VOHndOsvrEoKhxUQFoMCK3REQt4nP8WvOeHw/36IQQIZc+7AnlzkAZhb3eHTT+C97GNyCd/
6x7lFrqMenr18342nUM5FAHp6Ucf+bjJLVhnoB6ND86dW+MeHJMrFjQR6k511B96piCYtyQ/BJQ6
b91SCzxEYxxupvS/NHt4eO0UIpv8tDZqchjlLM6V3a03Zm4i8EW7ypRESzfWzTZXz5cxEBKlYEm7
16d1V7T84Bq8FYKS2SVfPHJYM3DgqyvCeAtMniNlYQxph/N3O/UcRpyVKb/ttVLGzSxu4IZtdlPL
I2qQWXtrB25KXhHHIVffEnt8wiHCl5JbW7fTng7H8b0t9USB6TZznVdfuopXTfBQaGNSF28koTv6
3KHkjo2JbiLYRTfS1LtZkq3GJorrFhZfhSTCJ9W8/onOSzqs6/BKQDVPdTPceWwCP1AI7QSM0B+j
XcnF3iRZCq8Ll8e599joSIGNuEGgeiTQ69rgxzJR6E4qR7NreM9oSBQUnZRxOm9imbyuWoarovfW
IFPlI/R2Iv1ud6Re1PzcQtDR+ev0i2kxbZ3ZQU79Ek2Wpjk3R7okO/cfU22gpm11gl1SZYIdySMH
smNU/URx6ysaIJ+9FRNCrqbuobZe+SV4qFDa+XtXfw+y8ksvFidzVqQGkb5pLKSJ22J1IYVGN4O7
6bx08doXacwtoT0IBESRPtu3yVRL4hywHIz7e2XPO5jGrLveceyMxt1t1sbq+5aRNtColJIs8k2J
ESEj1J3RTonTOAzdyKYKydNy/ZXaZDX1u0SxA6xBVTVAhbatPCC0/j8PpRAeoE3UN8GDWD0Kqm4V
L1oQIQbj5ya2gnPraxWFp7a9yFPeOjamJP+UUiFGB1vgTi4JHnk8IKI/lzQVBMoh4p4NXOIBc83V
CZZAovwI69cLVQDY4Iv1Qb88RXIMSC3j/uMb6fBE+YlND1a7K34ha7+QHUJGtiBCX5TMKMUkbcyg
7khOWySyDqD3hoPF+h3t4MNNWrzJimdfPLjmxQjmcij4FDuUUeyn5arC3kze9JnaX6rKWLX6wi6a
dVdv2W/RIwlLNFym3SjC35yEc2wHUmOHSCT+Kk6IJlf3CulQ7zLaCzCf63WU0t0Kv3ttTRwvqIRK
SydK0X+g+Zz/xB5N6Rnt08SMQzV4oNU2+M0WMPsb47I1bhymT7Pzx96p4lBHj3A6iWahgaRmyBTF
Ag+qonWgOSb2dHGbo2v8UQbJ+PMXZSNJuYaeTk5vvkEuwQXjF1OQur4j9Yz+wsRib5MF/KlGog3A
3qWKSWJYe1haDBKvmolB86IDNLI7wjp2bhKNGYc3SSIT2iskjiKjF5ZisSiVyJKUyNeqaWlLOM34
zYwQEfsnyJlFBPIC55Zt4FOUog9DFu+0pSIUQUILW8aZq0kgqEB7iDpN1zvh3CPMqqsSpdojlWxi
UvtcLV3bMqubndjHUVjGQ5ckSDnnfFCiJWUa+feaNgsZVHEUKCHMLe/86i3fP9YLf3pKgpeklDeS
hbYTOkeUNGQzPebnBGfJflzmUjCEsXOARuy7aTwVx2KZY/T5HO3PbUJHjgQOJdLIvrCKxnvK3o/a
BEV94tCbZWt5qvX9vH5EpEY0rtnabtTqbjxXWSl3CtM3ZHfDV9piQE15TpTeo31hwk1hrH6wBqLk
93pZ7QT+tCUh33ok8Qfikq/wu/KEUmHRcFChGNxugj0BoxF/dTgDj0x8ZHcwUmechi+JufHVBGav
F9ww8dJcX3CWizmQJ9Cncy2Ebz6pG4l9Jo7CoTKTCotLCAPH8XnTcbLozEH3C5ppPlsw3Jw94z0a
RsitE3Er7hRNf6AdVgpbs5oMplD6chNMihQQsXgjlW36Xs9aQINhfrm0GjkNrQ+BWncslP8c0T4U
uM8QASEd1vRNuLcRDmnfo0ZnnPaJv1DuRbVO+WEW9jsdIBtblCM7Njy/jJAiyBSK8MCIWR6/QVXb
KVE95imU3w4yGQw6SQlwTeygxL2uMdjks3I3V3ODD4UTPZBfEaxSS/TXND3O3jDEs41R8vadVWjw
XdIKhonqOiz4oSc0k4fPgivZQn5z1G4ByofZbSG5tavc1m+4c40AMep/msEfoPEh97CqKQec/DFV
uJl2NhmnHXwmVmpquATmkvpu7RaVUGtORlhmT0x7CSBfewDe81ExARwV3RI0AY74ODY6xAtBXnpV
9EVOwvQRvcTunQOWtjmcedYM/XbWhzuHAP5WlwFB7yOWBtKS40kRUNbRjtDVQi3qYSZOwz3AbBl/
1jdAXLRe6YxEM5+OAV5Kw8l457z1bOLw8ebpu7mXGQ2r8ln0QUKur+somyYep55am/ufL9EQR8//
772gSoRN58wyhlpdSrJIp+PIwHNoD4jYfnsK6/bKoUUzkY0Jnm4+dLkhgb4Mymizic0+Rxce1lw3
PnNnqozMSfzy6xjvAzN5xMWT4LxAMzbV2dbPBW9dN4dQz869PLjbMo5hi5EKSd5s0+ybfNRvYLfs
Zxad8LWYzPgOcmdiWiItKzFrKOvsGxBGB1nkferAZ0XZvXln49dki3vVVOHEMJm+zMuI1ZLvlCdW
CyVRLHtEH2YBTELqNKz0HmfVKS1HUZtZoJkiEDtyEh7vunQsAK1LlPT8qgPsgpWiIo0zfxIWwate
bY2sxgq78804qIKXPdEcZNLk9ycaTkCSiyNRsn8resZ2PijPzDFlQN+rRHZOtSpUZlJfQrzQFzss
Q/syedBUGJGgimX9SQfj3s9QHS8rjzLS42LJu1v0ugstyzpn9TkUWntlfX2OdrciKpuIpgd5dxNM
OjoQLfKAB9fNuM2MDkZFZ13im01anaH+dP5EI9u8JqT/7N3UlsuyHcWsWHFgchyRFG3Pl+dhdox4
W6pXemtCgWjSlDabFnAfxPg1uIGaRisApSdb40x66kjAebVLuKzE6KyN53UBgC1qTw7yOiSdKp5O
Rc4B27ocEVgt4VwFBQV19HJr/qrGFn+PSDC7ShZYiBHOma3iqhOhuj+Hx6OcYDvCxke0popOlfRc
2jzqT1m7q+lOXytq+nGpdehG/h9DcWfQdwwa7AdIxuQlsodeINYTlbHMEXzAHCPdv8A4oxZk4ZTM
o21FoskuxymLC5Qvs9tDERaEA/pth4v1FXPB4rNcrGJvCEAWqy0rguHZgAHqCWK2io57OdwOfssi
f6vTXF9KNMp/Q1b7sPC/lhSljDhbz/uLvFp4z6l9IfiZd8z+LY1QM074yJ2lB0Om6Ba9YnVmiYtQ
SEaxQMafCNGk65SSoszQ9nl1mbx+ch9/9XU5s6YMGhTZopr33OhmRQD9wdLEZ0kUOi6kGwHncEJA
v4XDUU4WEawOVVqmDBzRLMJOt8jrMTws+WCCT+rxdESMve88w/VeaXkex2RipvFpv1ImtLRjO+xW
glTDAFyZRJY/8XWHHE9OyrDTx8zbqhds1vKXy1blpzNqwScxbOB9we042VXNwfWm3c8ZufuZusd3
4E42TJ+N6EfP5cPRPXhP26V4WtCVJbzROsaslEZVqxv584urUbNBwIXBZpVR7RXyyiASmC77dRb1
eURHsbSjNVuWptNPCo7Km6QfBBNqEd18hTq2Rx3E/7iCu6GyHjTbLXqayOGwRzAqAw5KmCoBYHDm
ujHIIOrd7Iw6sSZCekhZMdEifp6mmlRWyCSF9jByxm0E4EtUIGwOGWRFsvG76tM/HSLSk3dKZa/J
68uFlWLdaQqrbyrcsO6lJkmiybF15rzBjKDtC9iSG/0X/DqQGmswHqFuDAW0eolgMIQ3GJ43GWSC
E+B6d50zmb3pmsSvCSq+lwy4Vxdt3aL006lYiO3sb3AzWICrSigCVnQidRCZYss9JEUIUQSBuNp9
rv7QuhlDpMKz7SHUNtZxib7SCUUZnM2yIUVHVNNAfg4oMWRhVPMqDQWdvL3z2gafmi72rncscZn9
yNiUAIvsO3Uy0T/u+qTfqbqhK13jtwI/vXXLcGpPv6P3i92/21qEHaB1VrTEGcc8gGcIVvnlVS4x
tpOnUlO/JjAVu9flRjuLvSh+AWkrTCl7DIR46ggHt4MWKlx/S/p2F/JOLAxHXKNsVIRfDjePLVqg
L3kosNkHNV4hREkBm0C1q2yP1VKyJxfBxmWeNpjcbZPlkNbiHTM9thgg+TI4gx6dbSXPdp/3Ow3f
4QiQtrrJ990dOWRsOM32n6ic0Hjx/7hoItZamD88aWEvpYEUNbkcB3zPuOfwhZJcKZIB7UJyb7w/
DGq+y+eooZTDFs6jh4DJ1N4awdt883vGAdHfXmUr69zQ9XtEsaKJ0e72v89JKnmHGItXbJhT6jJK
aQO1Axzwxsb/bxcpjS1VORAwQhlgAQWyjNz+kffXlzB7Iuy1wE4dxSoLSIPUAxNZZhLKLspp+eS/
Ao12o323Xlr8aDmF1J/YaVpAOre3F2IGpjni/zg/40rSqCH66tbIZpyIL9w/JKGGqK+ouc4eT8w8
f4Wn6kAY2vqpxlCJjGSU8ogL1t87GWzdF2O+dfVlGB21oOYkL9nQ+ZDhx2yIDr6PinuhCy7DV1Rb
SO63yE32PVV/Q0M4s1WX3VEA74MBkQDadv7+w3/kJfEZOt/OjejU3t8uB6RvWy+MTArVcCnMfcQz
DV+QC9IqQh74PSIHZKzUyTgs6W9oa2UKLX4NEmPITz/i8Wtid7kIfUKrGR8EnR6t5ToUcA/mPAbh
DECpIxYg2XpTJ8jgru6VAMbqA4nScw9ZiL1pMJm5lZjZVSKlMZQVt2ysCzBSMZGCe/omezzXE/xB
b/J9+6gJS1y9jpftTkVqW68qhCGqN82tHpLx/kB/nDN6hcDUO2u3M+Bi+Bb68ncbav8ouvB8LImj
QT6rdhd7EOdCP90sIhaUoPcEmGuQ++7/WKHUAV7iZAfnvHEyF8p/Q71iB947iSkJ6Fh+c/M74mdI
Ag9mjYm2Rf8vW2yJjsX6XEZsvZLPSlTyySbi0V8FkmNk+7iUVL2H8bcOTGdgssZpykQCxiPyeYpH
S0sMrFV8u712nfi1a5MgYatqMKCpFtIoeqqZjxqiwzfBTVIJK5mmG0GYOsELrf//rBiJTRwPEcLz
4+bBre5PwNWwlbGRsASfJmOvEeLFfbPueOtyuNVedl+fFJakAFZe4bC2oCOoIYUYBisz6pAmKHJX
YLq/HVR/xnrwKcOTKV3Pl/VPWokzZOD5nSvjVNkxIiEmsHy3MwH4WZnoz4HmGl+PSCKaO6P9KnLw
nitMIYTNN+Quj9WeZEuS+NtW64MFYA7JtQftuYZTZK5Em8k7B0x9OTqVOy30MyZwg8A1Efx3y2HG
OhwqpUiw3/aSpWV1anAZuuxCmqHloEvaTYlgMcKaKWdHaYB/S5Lcpo3vORZjRutFzR76rPGN+Re9
0xBUdCNuyQISGbWNIkC0iDiOC/5vSC+oDOxXwK0e9Q/VT01SvzTlM8Oc3mISY5HL7OSt764qsV7S
W3uk+3Qy8QV0KTyGbNRgPbgAgOpP7nQVsobbNOz8olUE7iQmPZxYkzaI7g6TRhAKc2jEjmqk3y4o
Qa6c8RGI52YbgHgDOcL/mJPNCgT6dzt6qAlzvGATOqVotw8Eq2qwhRjPakMNMKvBFMtkHw+ahR/s
mouZRYGgnHIz0IgolHjzzFYD+KsyUPyPKbX6WolelZIHa+dkE5gXlScZGjMh6NWtuQfSNBvxu4ue
p4+eJTs2I8+Bg/nVGCpLLVRdTOktFZZEcT8VI4jjVYFJUxF3kY8Rcnq5FUe4lQh56/WB1ZFu41KM
Ygoaw8pfsZ0o0gsxqbRpdNJhs0IiNVp8oHUSSxm9sXJieqEENMsaYIy19B2etIamJ9BDkY3DBUqr
XcrSyMGG3K8pn05OgHJ9wLm2diG3lv26U8fV0KkYGRTJKMSiZb/hLgOmdoW+eLdmHd34Kh43vLXk
MxCfzMzmOQhAQDC79xXoQX29MLuK5Y5U74wsMBApgzylEuHcrO5bKOWyOzvQg2D4wwvWPE7XxNFc
nNZgMjLqJHYQtmRD/zwPt2FimKC6PqMYV5Cfoh6vdgCyw7LoAPMHszQrrZt3b51GHNDkgPN2AvqN
tMaB98u5/r+V6/hQxa+l/+ugxG5spKy7B6g9ywZ5WlYoiUsx2QU3+ZnbIO+uy1814kxoTQBWQheJ
i/kOPkobvLVphW42XPs7a34FMfY/Mvq26E9Fj74csEDcJoRGYRJcsJhBagr3EG2jEBq2Dhj4ulOX
VpttCEdAwnHbVrKg+mxlt4FOzYja+EbDPtkEb/rSj9qnRmamcrxuYNah7+nC3VJESltKoErnLzKr
za1qnilQ9ZBeMaV+WyggDGa/CokJW4OLPSlMfIUiFEjswYFtF3N5/LxZrnhPWr4IjBVEzchkky63
XPDxTvYyh5NFYRSy3U+woLRus0dyVlkVeRbzoV3Nw42t9nMmg2s41BA1XIVSlnL3mOOpMJVjTC8X
12LyzX1QJFuBiEk8iGJ40asllt+FSb15/SSWJKQgsjC+36a7vvohuZQHHU/vKU/4gJz4LbU5YjzQ
ntKrh9Ra+AsKopDggNB7l/VYM0LYTUNNgSuvpTYco6USkpr1Jm2KJEJf7r5ZRAEvYHU8TMMRuPek
T0SN494VY7u2GTpqyYWgBWKZnbX+07MLlBPuxR7+DDaIi+16ZUw+EdfXYqSPe7TmsJC5AjF61Q0y
IOMbwCaLY1mVazemGkbkRZB554YYVNkdDA2QU1Q1LrVe0+6DURxGOFkYMRBzAcqODzN1JEULDCiu
TMLHbW6X1UZUxSS/qmHn9gw4u+XEi0bM2oORP/o+zMJwZ5A+xyKW86ohIoNJCgni/fPEtKFolSRe
prr9du72jCIx31yx6y3dnlZXCT6Ov4b/sDNpqN7tnAvvXQ7PMNz7wIv4uzPISCrGdfjb8m+xFPYj
jT2NF9KylEagKjnknyF03HzNSkZ/NL8xdzCcwHNOV2fGdGfVNGsELQHy62qnEBJdoyHbBZWinlNz
C7wwvpZw8TI6ftY7hyQ5Jk8VqVI99bqH+RLQIzZtQ3vAIynoCtgo38jvzHQs61OxpO2n+mb/uPZc
Vp858EPTNNntKOuIKrGnyM8zk1jdK6ti4QJOjy1j8MUlPLsUk4N+kNKR4R+x1tXmE09Nzdf9FiQs
4mu2vnA49n6Z/uSwpcy3rWmZK0lPnJ0/DiSXMmk9hTlmSW7ekjCz0aqz5rPPaznS1YQl6yML1JEA
BK5L52hmA96SOKXxmtq4Du5R5qKXx+wQPEetilovaLT07iwdtP1X5VKRQydm68NnRgnrRD20GFqu
3nGvr0N6+j5BL0rkaQ9m2JE9G44F7N3ZgkCHGxFnITSGA91dLE2C8qmY2sIzdw3RI3InWNV7eet0
QAgHNmh4nwV8QIqiLk0bx1vama/oraDqw6/Z+8S+f4qMP1iHHwF6NYJl/awG1Fv+yRpd+dfz2kIg
aeLrr1H8GD1NkK+aQWIPL4pzoVOWBqf0F6birXFyzPgTCmmmZKtB/mNuw4Xqw5+kJwiQYBZJP+4F
fg6vsizveYUCck9TBZZhOs4jeKoxH+LGoIxAiyhGxlZF0yitWBb4L3rdetL25BADAIDcWR1biyB0
CL++HbZouvjSlfrSlrEXgg8LHPYDfKcD4vH85f48wwC1SOw4isYpY9bOapSYT7KT3ANxNlfyOsfA
vgerkna5Pbjzeqy280FCXiCeNoxqNMTsLbBOUmB5FQLiiSuPdGj1F1cGH0edLWEBKuthm8Z/gjBs
zW5AYyOPgaxd9IJgibjJz+F4LkHY961FSJ3mS6IHtv0rHaHaKHciNFAOsLqinrCsXwIQXHEix1g6
LuVSdBNrF96kAhXXgCYB4laW44uCp9VdjHL/9R8fjJHQ72V2ItsKm6v1OlRhBWG8R+JidplrNByj
n3j3Y/oOi9wHoEDwkX3M1S1teMP6ceRz2QaCgGtnU6m2Arcblkd2ZMtPuq7tWbaZlAxsgwIkf/9R
n4QHa0OGWGtKIunL3GluQVT2bZkfyX0MPgK9kTA+zHdnmXfJnAoam+YpD3dA7GijwQnvxGOhuv6E
ox4v7S8sDhQsJBNWwwSA1gdZbMu2xw2+zbA5VmQgRCBYLOGxLBOHJafqlsFM3XVCgBaG7EajPyfe
d/CQuFiYqL/bNm7V8L9zmHJyyHM5js81EwdKBNl9M9Jfv0Yi1jny5imqdEl53s1OmzpG44s0Z2W8
wAiIUnnupXmQD0d5uQums4bt46UiJozDKSbC+I3Esk4Mga8ZqiY+n1iN9HicSFeXRE6eBMJRvV0q
QqAAZYhS/6gxrKcvly7w404jG2+KIcV7K4mUtfjEKjP2b7mXVIekdSFwWVnST99CN01C+5HrTeSh
AWkbfQGefdctvfblfMVvXi49Bqc5IO42RIKfn29jnL5l15ui+5arWJQAC2SYPz6aS1EH258ZkL/T
0gi1JOOuqGWCCBX4xzgSD+cf1f7y3bJv72PppyEXI4hjcWgdjCaQwxFUZ5ihHbXzekC7Gaw29V2X
ThuWkKxf2rswjKlqHBuNPWL14dhAyK6lyV5VXrruY8cksfTmuS7lpJOeQzZOLmdqDrHaI8RKN1wc
/DOiHbTPmAL7FBzkVrjKv5YUo1m6HI9MT3yvha9dTwEiGThZ6zusKFfaMu7DhIESVOxO+zmCPsRM
/R3uL1ffhJ663PPyi9vnhmYI6+8/ObTUhjPmmxhO1w6zjIJw/MyMKuRKOs9q5cMmXu7DK01eUUqI
XUF64lbL0TswCYNOslz67nNLmrXK4bQmTV2DgcMR79i8AEs7hIjFD+YO8Jhgh0F6k4ZodR9kudgu
oemg+5jOrGmyVIx6CUbMnkm0ZoWpHHRp+Kz1Dj2YhtSNoO9zLLf9eqgGjLsT0mvOXzR1EGeCkCNy
aBn1VBbJdMKqc9LS+9V3ncW5H3LF5xuRiT28c5IQQq9KbTtuV8vQufJTrgY2R40tAralEhw5mihL
2+Xs++AWwFNMmQTReW46WtApAKMAACXf54v0W7PlHI520jRXROKro4GHI/ziV4TnHHJtZ6mDdqNx
9VxsLhjCmlAPY7Xi/fNjrY04HvVx8ruEBfU0mFCRsjxbdpBsajsl2YLZpLs9DNSUUTU7U3yRk7pc
yNkvJoG5XQG+A7QZjuLqmtToQY+46EGeq8LR8rf3zYat2D1u0HIP/wqH/5O2W2xkwm2MZyXZUw6P
OKv2zV0G65d0mqto8mlZYtN9Wgc7lFUCr+ZJw/WRxv/5SUXAeVK44CnydDq2PUug2xlXsGixXLcP
To7dnydlrhNE2buWXlijwXeBg+ToLfQvJchvoxBluLxX/XG6LBuoFEi3j64Xoc7tUSx0HRtJjAYV
19BxB68j9bOklEnGDBSvE1AI5nPjvDTgvltLvGI/skgkT+H/Hyl1iMjQqGauHdJ1e9KkgOtZCyUN
mEVZ9Exzz5reK3XLQj9Gvy2nbqS6lnsmIRACNDsmHsepx5JMwJKFHBTukSjzF1nHc3y3vgHaa0Xa
lPk4ZLX8oa8qmCeJROgOotMTOlyK4bmHFJ4Dnm6GoQNwVa2WLTrEwyghcXTQwIRDoROf3B7dtlY5
2N61pbpOu8q6/7ASALvD8RV0eHw/QoceX3sJoYr4zR8PdjmXR4ed0IYgs/33QcMCPKOoZg4peIAJ
BcPzFBCcgjaHlI6Pgoy1w0fy1+0B8i8ME4nFUT5aUzZjL3pXwhvLafAi9CwPzfuTlWh5eg6BlcDI
aprWLQoKMYbMlQcxZAQb0FVPZcucWtwXEK1Q5Ms0vtUhLn9ODtBmBTAetHZkqI/GyrwLzW1OxI5V
pWPWKU6KSECm8Z2G3y9cIYmkvWxCLRzrgi4BS5j3p4gvJV2FDRV4rH0PqGJPLlGhYBt/NC3EMKi8
nJ3LVlPtcBW4uatTqzDY8QXTGg3rMZNK7KeKPN67bWwh3SlQnPuSfTPbmNxXA1snVDwsqe6XGcPp
+UtWyyekS3gTaxtN+AwmHBaoREi7HK5G/KPjOy6JzBvGx1XtNQaIB6/ucwAsr49+EVTw7tWAiWL9
hZs/+fge9yKhmS4gWYxU396D2X2iZKW1jSNFhXbqCnBk87NOJtXczJ0F0pZPtx8aI+pRiU9V1IwV
J6Ifu0uDYc98guP8Oe6ovWf9xJBbVODamBsOMD/RBw9BSXsESaCMLoN6R31YPKhe2csxwbZJlqOV
JAlleHlonwGtvPhs27iQRGucQ4jxY1hwvj0r3XyHB4jf2kuZbymCfUwGbVz76hv1pi0lVDyFy7XC
EaUazI0MjMsZuVD0c89Rl4d5UKNDhwSvw4G3RQU2GWB1gEQYi5XrfRC55GarLmj9pA0nR/JlJgbc
KWJ685HnEg9v2LuE7Wmx9bOMjCtBKSXxAVNarbyHzZzgqXLbZ8avzVWrgeTcnGbSsBUu4A5X6IDR
HUrCuY97mE06+vjdjomY6Tn9ONvoVYc4rM8zl4KR/Ra27rdbFPEvhNI8xOFqTr1Rupd1Vjar93N6
b5tx6BoOdSbIerG/WxJ2kgtCeupPClY0eyte9zKNnKN2uYQX1rGYBK9UaA3pWzdPvaZdeWoE2+4R
AsTqVhU2Dc9OUx79+q/9gU2ZnMZOgdtx3+mqkTPVYByRCT9Ybxm3bDMZOV9MYhGyq/8HnSGINhh5
a4yhyOvUa5yp0JXfkqCULpnNxNixdOMPqPPsd8efYfw8VTTEHIZZu+Dz6IIDO8JKKCcNQgko/pSw
F7akn8Y1hDA0Tx4ri75u1FAkATJIaIawsfDRJHUvMjYWEliXhkPiJGg2/PeF1SpsPmKOL5vCd245
JL7s5oTm6MQ0QnHBWhs48dH4adzzeh3smwf71DzlUsnqqeuxf9aXB7QAyjNCVTaleO03ae2Jx6AV
5EMpdwaYsRIe6hz4ETUwNH9ne+gV2kkihxjY6pCtnT6rDZwFVpAdz8yX7qtYFzryG0CyD7hwE+Bi
JLp2gUdpWKkLDHjaAcpCZOH9In+/0gQQtH7GO+zAjBC/eDhJHdQjfr2s4dkVxeTd6UzQiSlJScGt
DBUeHDoWFwtVeDdIfLOQPtFywg3VEL8jEt5S116Ud32ns+A/O5iZp6syuoYhPuaEGbnWPM2+BfsG
Q/EOHDk9DRriTXhPrYcsVxBUfOchYJx/Raj3uBf2IRdZHdEraggWzzp6QqOQn01BWKGWfW7ErRPa
nmCOyuk4CRuK8mo8FjHGy64Uc+rCK2lLvuN2r4YTCdGK03cxeRCBkINSvgPeeh8u7GEU+h3kkZj4
FMZcrOL3+8k5Rk5yhmyhFNwAyifOtkEXfAtj+3wBIiPyPF2Kx2Xi8wah4OwGM0vdROLI5F+z/5OJ
c8ARIMh4bezh1tAn7HDbM5sE+dc64T+rMZqzaDejJsNzOvjS5gxhd3QpQGYfXDKrLOBj1qw4znxh
ENaXyoW2JzgsZeEm00kJvP5/yyp8mSniWracgybBkx/OAz2pXN7v1d1nmlc4aMnb7AqNKMFJqWAg
TM7fKJ+vxMRzdjyFjg1ZE3C2LEpf8xHXGgddwU2gjj7ocoO4Lxd7QIA3xX+sd3oaU41rqcwOTh0Y
3NK+V+mdtjYD1624vBp/bQnQW3a3IbMfctMj+RqoNOQXgkrYnmkw0UzL+TLhZDAhamXNJDKsXRSd
hcTmsZXdf7XBllTId5Uq38CNsKE5CEkJJlsH28Yb1ssYy3WLEmifpZTLxoHWARK2ewCiunpZoxdt
hR9+yywicHw1MDYaRqq49N11FKslmE89EsH7XdQJspm/lipfeX77FOZIRW2/DEowE35kgjYc8dW5
kd21mzazLY67vHETSFRVvHyQkG7znjtZ1yU/PHkU3JipjOokxBRA1SZPXBBwPcjiHzEjCThcYq6+
V7hgECI+RHi0dKsgrF+5HUnw/3CrD3Q5rql0475drpPYj8Kx+di08ReIvU2Ct5TuLkUd3bKoBOj3
FHOG5mQnx7CLHnWQscg5GJKQdj1v5s9BGH0Go5H4i6mjI88qBo2OtoBXF76LaZqnMa7ATrJ33v3U
0XR+iPBU8n00lxn+Hzq2UtbDZMblDQUYDVoEcc/GpP9A33yYbqkltsetWpaVp2Um/EgEQanqrRID
qTMemdMXHliaLSfTFIfWQ9354tlmOsn3YeZ0S4bK9kqQz9/tMTsoUYpW1YDLJkRCsgWs5RUSVq2v
o0n9AsQtFVR2/w0ojtpjWNSTUeB+aC+BN/2tHRGKxSANpHt+T0GucD4DT334RBb2MdBdqtMUgIt6
xqP6an4zDYtTgkyioV+lfwN5r2/CaVi8vcyecg8e0CsSb3oS/Opfd9YO9YlNDRXSmTuTTkHcobeR
MGMhHeWRJyYWiLdLyfcvHLAjMK1FPPQBJ+fnmtC4oerKJi/Ib1rOVMLXFr3Q5mIymWR199ZsNyO5
/d4eEZA+H0Fb9Rx136vvbYJGjocAXXgPCktD2fa8q/U7KUL9941+Z1Yyu7gvGVQOFdapvcgKv0ny
J7lu/+l9VThO3y35qqx/g4e90RlOmmsYUWeMJ0U5iUfcFVkM21MxVyjuGns5teWGv9s+9WXJUCq0
dyaGU4WLXyv5DECNedHRg9jLl9cyreV1epdEaDmPwhXGmXvRFmBbW6vbs7+Ofm6xZ3HRyo9DZz7x
uTmF1+MMUJPg34xHv3F4SeYK8aoClAR49f+wxiIm7XwfDOg11KXkcmtWRQ+QyE1eVkEQfSBQKMVN
pQfqlZEjBrrRnIspqSxvHqKDToLH0izZtFqVLHFW1ESbswhvnxVzL358fA6NAITIq6eaxwZdPpH0
/Q+RoGZ5+SxEg6W2PqeydCDnfvIJfkceh5cSsncS0Yt4IjDsHTXzrKlhqb2KCndC6jh61cv+aLZM
CqpKvblZZXiRChS+vvTWVoiksGKYH3wRjW6cbl9n7r1CXInQf0MfDm4J1zioRQyBJIyxXza5zMBi
xnvZk/w9WDKbyyapeTTzvC7VSFxv7LE/BaELPTHNPqQs0ayWXaUk+y7X0nIw6eJ/P+tEohWO7/7O
gldOKbUIt+PNVPUCyQGxtEVkEuKbW2tZxG5X9TkTL8kIluEN8SnquUKGoCrulFnTu3Uj0n/Li83h
y3bbpktLljicEMrpCO+Qlt10DxlT+BFytXWX/GQYotBJEsFieo5WfgD5xE2x3AjvmUAV1DFFIc6Q
bP52OD2yd+5TxzTD8Dma6lT90sXsab7nFaK1/FLWzfoNkEHWDlgEslowEHgFD8V5Iz0GhgSqgoZV
H9/vBq2e9x1Bm5DdMzb45tPcMxgVjme64QtPQaUTUfUr0ALyG/lmDOYFzb9aCBpZ/mDsOMM0Vlej
N28i2F8xiyvsy9CyHuQfYy63oGCiOm9bJDV6AgmRYbG7d5a2zsL7dY5lUf041BVQg+m+8FEe3Caq
27yWdq+nDdTs237+UemeNf7eS+mKpsylOOfKb6wcfPJNTxFCU0iGyfWKNcZvTxu0mvDvndiVKTu2
CQQ1a5PeD56Y3vY3BL/xBVf/oM21finsFemCl7ojYj5XNNQyPBmy1S3aIeO24uFrM32H1fKlnqlc
ksHymv9iPkYxUeZCnnTA7viGsRRDEMAkwDlRIIt4v+2cVs0ZRcqjgJiOMkEFKPLIZHd1qfBzNdxX
8KBy31SVbD8GaMPSt5cETjSzr2v7hrRtfKCN2SDVuXZGlND7+nPifMrThIYWCKX5Wj0KS9UQ3ERk
G+oDp86V0i0NXf9broQDkzED/3OuQ75SvMOGRD1Ca5iK8NDzdhinPCIdIuogVqq3uINmavrikA56
dtPvaKm0zV1zug5o4uSiUspf3qfOSeZifYakTFVWbxkFpOMPafQjHc9i7w23OzKcKIEj57Z/tVkh
zGQwR6ileqIpm/KAasAVnJTmxr7bA6A01NXXYZJL0jP0OJoCIe5AelyBvHFbZKurA4p9KZYUMOeb
nCXNT7bywJuzmE7ec6ziSZAtb4NFO0UYTAO6NYrS4X6Uo7h1zqSooQHieVzyVM3GYNX8psDphXgL
Yqza8jj3wKr5nkwevzxRWo9qI1cz0yaPLvMihg67t3qfeTl6BapdDtu4k76kQdOjeT9qmW2vpe1T
XrBeL4IEAPRTmnSlwNEMqaUyjoLQ+0/oF1xPZODXc+0ZIEXpAUKuXVhLJ7M4tFOtGuShLiDic+22
U1Me/9SdVBiF0d69QUiQyMP7uoOHqsFQR66Q33cW8PwHfgDxaa4o4pDOSVH1x7dRjolETVhXReoG
QQIstlCpwps2NvMaXGYFFPhUA4IBZJhYTCv9BnekI0EI3VWELERhPGsPwhdffxds5o/59s3Z3/Ou
jY9XVuwST7XgqIen9DWXfWAAPdeLfdgXAKvT/UQ11W1C3roQ9dmFgD4mYeWz3DU4WdaR6sPdz8xk
VdZ3BS6CBwABM/WKbRzgJ9hNTgdMApuGUsAK4D5ee117mAaXovfzdbPiJe+/YzZEt5itGMi+QXvO
epVpxq+rklp22wiaIBQpFRm+rGs8cR7CmjVshyGeBbk8ffUB75K/b0GSg6xcm+r1tIkzCGHrQWgS
lfDbmk7YVcdvRrNGgd00qfPpM2gVThvNCZDRBzxH39pEi4za4VLFDr5FYv+YttUHxgZAT5YK8Tis
my2P7kByiR5mX4+vYgngKwHZ3mFeavFFPxttmh3BFJgcQDzjyDuzFqI7nSIKI3Dxq65TnIwdozoe
6OVfKceok3qwARiteSeD/YarMuslOLcB7P9zn2o/HegWITCUjAKPMkc7cbnWbRaByHM6cp0NX/w5
seAoB+70EKy5LWtbT3rh2P6iKiqR0xYGNEb0nEoH7qYGah8/Icpj7FyRoZ3JTTTTIZqUJUmYIa/s
qi11va8mT251Mlkuuq1N7q+I7vW7fFWwungWmkeZHDSnF/xzR+aoQMdGTI17l6EkXEwv4Mee+mfj
EeZFB94nPszGPJ6E7QTl3Rtx779gHidiyqvkZGm3pKVF+MYO5p7bkHFlNKa3xjoNPKgRuK/yEYGr
28PZDQ85L2Zznvr3r1MD0aHB4wPknFKxFnTRJAD6jGmlNrIxFM2oR6mnObogyjUm9BOZQlF+Tewu
UMWkeFxT45kBIrY8Ndh3U7nDDCt6bxT3PEKNlvC9tUIQr0RX5A/RNo5Tf8GrbxN1OnEw8Dfa8AwU
sJ9yP2tmG6R08Ej5LqswEGXL5+zA/TVG0J7vjlS9OJ0i885vD8mUDy18kG9ougU/CnqCTV30YtQ/
BeRIL9sS3IcG6ZYXh5oSap5HFSiN2Wml8oj7JiVZeN/h8GbItNS8HMDqhBV2sipqwHIc27VEZny1
EIOZy1ZpFGPdtQ7dl/nrLDPQSm0IVeRyx1reYrgo8kX0fUlpRng1fKvlc96Fmze9aRRKEjfp7NkJ
T9S6Hu7RD53jq8Na/3Fc+2ek/sU0sJXyYzhUP78XyCkZELjmOjXif+JgnLIlKkcbGEzlvsYDJ4zK
cZfbSlAPM2YO1OYNYKB2IqogxEdKe1jS7U3l4LRpeBt4CKw8QLkBqrhfAgRYBlme6J7YZ9M4c+v/
omdfTzpJhkzBjjO7dgmT7lOvUZ1Apj3YX3KbQ/OcX2A0OPWcYT6yr5ajH60uHoTBLhAynKEOp5XM
On8lmObvJqvxJZzS83YB2ftqSM5Z7Xdyw0ytNWSZB5jmdIa49iysxQvszNjAUWpxo8IbXdXyn02b
dy3bO2coMrMkQnS82JkRVOzXUv0PlXoZ4EWYsDC9x1llX/yrqkRimd0vzNf5ulvqwlsFzvl1JABB
mGqiRUtF//yhOhqknSsTull4HVswP9IuNIfQEM9fXUSgwlKgGo7WL0LQNkET5d/EOlLRFp+pzjRz
uKvJDARl8siswZzB/NW0aE0xg9Q/dyCYFAb+J2PKNG2QXmz9QwtZsBL2jxSyaI6ThZ2dUzkGaj9g
2odDC8nJ4gqj5F+tKP+5AsTUR3COaSNASy/6s+QTmWX9TgpkzzH9VwlnA0Pog3GezEcmD2IYaMRx
q0OELKTOrPCWZHkdecqzuUKwLH7vWV6Nq6c5/zimraR9SG7XqdcLojc6aI2SAjU6oxV71n437+Ln
Vd5P64wpoSGWXLDubh0QhGqCjZakTLyFiQ6zWHAgywMHbKII8yHX30KfHdJnM1y26iQW2vZOU1qA
/635OnVLlaY620Msx6x8guyhmpky6tyYikujxo5PimhIlbe4rtH2un29u4iY191EaC8RD2n2sPnf
un6k7ykCtXU/Hp2XfEUZ49z3mmpl+df/WTcsnVBRXfNvEpbtcNL0CtGYmTdNfamx0JI1QJyeL31o
XtXK0U3fDhoe6Fv6gZrsZNaPGLd9R5uBx6M9cJwlHNqBXbC2vLqo6pV2u8fx+sM+CfWQwjE2udWr
1YH9+zKKP74yHYMOWJkPRXBtZNMYVeDJdDWN21s11PJUiGa4g98u0y4Y5mroRe9oG6Q6XbOhjZNK
F/3YxA5V0nQ4zTBq/nEV+i7IVD68+1T1jYb8Q5jByC2gtFRmaCGC8PK8Vc3jx2mVBbzGOi1pMPH8
kQdQEAPLb7Kb17rHlCJXEi0mWlFQ/piXxf/UE/dM56R6cEJAt3f6ixNbBBZilw9v5A2WHJT7mcsj
tYvgn6rurBMoPM50adduroa7CI7uZKzfT9FAX8ezcefLjQSceVqwGBprzsteHL3fQvoyS9aeX3l9
upgl0GEGFTncmNDTmXDGYJW8PkUTPQ/12yVk8rL85aQdRtKzhBQM09+PWo/RDhRrDTnxlxxoK5wB
sv41rV/jGiEnsSSXPbiZWtj8XSn7BXRIcXX/7StnTBPbPZ64cOoqCjKJ1NLDSOc7d4AICzzj6x9a
i4e1o8SShWihgqd4rSGDaOkwx6qDZZZNPQc7wGRPx0fXQub/Y5Tl+orkbHDlLl7KsxxoMuiOLRim
KE+j14cxy1pF1IL74x+ApVGr+NLood4SxNf6sdfjvTWy2VlQhbgKhJfM+EMMc8e/XQj2ufkoBJR2
YiZX3gims7JUrc9vtUQ8mGz0crX6kzUQHSmuElvGn1wBdCWVvpJ0GlIGP+mUIFN6WbPNf7rnw9Ln
Y/s4hnoVHtYyCX/AnHrujXkkIJi8/UoyVEp73rGCGbP7/qz4XEnDOc3WuCAJO66UPltfqzEHIzfA
GbayW4aV2CKexF+umD8B0SLrgZUdgMggDaMGOvTyIP96C6XnXZzztrGbuweJynM2z1pOl+a0IEiD
QNbYC69LSe7PiTueDLso6WrCotPBQmrd4fc6ji8Oi2/EdfTkHjH9BOdJh7ecE2qx6rOhtS1sk8kZ
925cUG20+IniAOyPW1SEbPx0cD9o5+Fkfq/ZVXlJVfgZy11YHytsItrLEbhh2Oz89BKv1ehRSvYq
fqPvV9Eq8GGm0g4czFgtE4Eu2oFM7N/2tkC0uRNm8lJOl+Z7ZU1xa81uLTKNP/0vRLc+SMh8kbwR
zv1JmkVp5qVIkon+SIl5bY5FNyk1Pnb1bkY+bVQkonspgKw/6VZx6sSwIkzgs0mAWwfU3U42TagX
PHgHXS/tuEEEA7gq2q8DrLcfYnROIjRFBWiFET+3x1wxNv4fsFy4nBs1oeGWU5yHtHrtltKzNdM/
01zlS+Dxhkxx23DF9yHEsybtM1xQgYTfxbolwzJRc+6QHFpVCuwlFbjwuFTADoUd4dnEv8boxOOm
QhWiy4jMDzdUdKOwsMQ45hH/iVlYSywyFxNy4dymQADja3/4dTUaKuDR+YikmNhbP0Nk3yNBoluo
YSRL4TzXjMGaIaLu8P1S2M062hn5nEdDVRaGMl/j4fHFZYMm8W8APnk5cz2P9wKVlyuGYMTLrFkm
4/m//Ezs0jlYClD0R/zwZV+oSZJPJL3gnd1t8U/doeofPMJ5uOMJYPfortk6WG8RAJRUSpoghFNo
rT01qdzXJxLlNgiiqSZjHTLibZSnm2KkpQNZofjLlkwYr5zRLU7KTq+vzJkcNt0DQmqYEIRZqmLe
+3KdiPScm1VlIkLbkBtSDDN1iFVBo8TDj11jUenTX70S8yiCNBmROPg5lV2PZi4y+1SakcNAiycL
a0H7g5uSliE6z4P9B2a4AkrOzzeBAKSwuWrwjXqQcos/jmFltTUYqLr69Gla5QwH6ZWe+0ldeV9s
ioDfFXHzQGAkZJIdPzmukuyz+xQfXbFqt+IqllG9Gq5KOh20apDlhFHqFBxx7JSssR6kKLK/NcJo
5yx2Fublg7+VTUzKRUADYZnAkSiL5f0ZJ2RFBdLgcgafM4pJOtVCBvibcnamXoz1EeNwH22j2Gug
diU/FwVuzbzKrrcMb34fKMbzphhKzqF/w685sxXy5rXaa/9TETV/VjGkiBbae0AA5PJnnUEJ3yQa
jTE8oXEcq3io7EXVFQp9+c8z3JlUDVb+YgYyO4SUnO5GJ8yiRREO7wQzqdbOxs7xMnoMaYMw/Ebj
myJQny6LyDqVX9SgHK9qFrMF4iGaVrYaUMtsKhwK0xpDEaWW61WRjp0qUcmY/zE+jCrCiDO/tyie
nT+AgVe7cPyVuYvweTKZDt+bksHBtp2bcrbWFswP2gPONVcwtLKoiau+LaLV5T9sJ+iRB/LMchZ9
t4S18IbcGX8m/pfTp0CdamgK0q+rEYF9JcIOGntODNSc2f3r5lRpxM70DXB/hLSHBHSQF1MGPpdp
67lVdpZqFuhm/FJS3/zE+gtJny0AjHc4RnN+iMhfTOr4ti5eoiVixn59ZEHm6sQ4RQCRPYJL75Dw
GMLle5besevfove36CL00kDfw0hILh+1YKK7UOsRQKyfkc4KCy+pAzOU0vJp5QKfCrtf7E6zhBXq
zH6lfnXpdI+8LIeKZxJBc+cX1xRTINdqtNQFroYyDOO62RcK9cCK8T93Ob13R0TzQh5m898G2mpG
pPYUCm3oDSsRCaXKZrbo5U2W7tLjP/OIe0Z+9AsaD8q+TyFAyUlBcanIJ0o0pg4dqd3enoABf30T
wtlVW/aflT+VH1IQWszwTaK0z02fP8DAkMiwSYD7PBghtGzxztV7A3/+MpwogqtHz29XDVidZrTP
ng9w5AjFvThi7SyvTXU6CApxXQAjJfDZYjbxZnQ1nkMOclnzA10kG1ngHTPkw83mBZMwAlsoqbey
vJ2ZGC+2jq4aelWN3GoarfIC87784Pp0QSi/m3b9LGE3Gh43YuIlUZireiqZCxo51Ked1zTVi2wp
LG1Mlkf52TUSVNEm7BJdnkaX5kJ0Df/L23i86piuTZIjekRN9J8u1Ir7mawzfFvALCfy1ErU6ITL
UR3ikSTAydL/TigBMNwgYYyvKIPv5deHT2r9N+IqX4CETHrwlkQujc8sOcm52kRKV3sjMS0jSkny
M/+vsLC3U4QC8gJY7cp5GFEpfq2St7ugWQgs9XnWVF5VG+c2oK0X10r4vPma3LYU16mIL1TJIKOK
FcsDA6AfvBsXiOwClZ9G82u2zR1cG8LEcInsWt29FLiqfTqxQkHOqy0KIHXY/vtEamYaz4w080+q
tyW/F1qNPdpAyorulXQYPyYPkTzocXikX5Ns2LeRFx9nHUv0xnh3ub0yQuoX6O4M4zQUW1VcCJg5
eX9tt15jSHozt4fV/aUD05mLwuhTFv+Jp1MFEb9+cIhEn6VlwKxFiWq+uPcJnCHl5MtM8C3mjfuD
6+hgTJDa+JxMogNUETqy2Vz641aj4XD2ME4WmXavPm3ejuU7KuCHdpRQaA72wOOs4C4oClVLqbkG
mzoV7ufBLF24v62zq+qwwS+6fGrLCpc0cE+2II++HKEHjPdiAHw3lq3TmybzY2EzS3Uelb7q6FCd
yFhMb/1f28KQMv0hNxE8x8XBOuTvPKD3NkGPtVv78I6Yy0FZeCSHaXxhB3wVw2ZuLV64/YapA+Im
9YXvxtNc53FDj7i1JHZpYd1SA3zJq6fzdTixseyqGgkwzd5S+10TDrI3xvraoJFtmd4nxHVsFes7
u8qUf8QmyjtnkePvr90w0iB0wNPFtWSRo/fXH+rcw6xHetWOF3dal//kdjyi1tZGVeAqns9kXjHn
Wz0CAs8/F2QcWex75fVXScFNCT5voAK5vuyB0varpXLu3doH5IzP7ifXjT5WhmCRTGhWs+ZBMXj4
w8SnWQX3wdiXxZ1oHQzo1eoIRgs5H/9dDBOA4VHSLeGSaKYU6G2kKrt2M4ksQvvs6Mn1EZirqTUy
4RInBZKygODh6XYkQHMgvEyLDTdfuq7ZaMGzKUAEKXUIGG9yEFeg9vpG6UManlnGSpfvPvx57+5G
yepwX17w39WOyddeI8QiRwYCYhtEciOzUu51p0gtsT7Yn/ozlicZQbzGH0prCyye5bNgRTTjnWOA
8VFphRE4ypis5sWS1yhD/30nvCweWV9xEVkBpdjHp2pK9f9aFMczqknBlhMoYmx4XLzcA4xxRvwn
Wg0BH3XdH0YShSZ2RTbcgd2AWNvAHHN/sm/ra4LqVXBsVX+vYostNK4gUFeyitQiag9tuh/Cq8gd
FQdQFHF2oDaJOD40xV+QCNe29iFOam9sYUmzk3abXZ5YKKeSRIauB3rudtyBJclvyO4ZzpAAerwi
WyJO9Ibbo2ZOfi2XRQDQBA2j15rD1O6AxX2KuA2EvQ/JIikDiz+9mr5Zkl7XA13iTcU1/qfpnf1f
l9QRr4Zm38TBZBdJRY162NzqPFLqtnXq+EzE3PL3HVOWJNdBnZgN4TkqpRsW3Zhkc4Cc1Ktcek3N
IMEswt/X67rSldOy8cA4gtE6uZtDh14pNl/jUayfRn59ioAn5o+7tPwm1KUm+AEJzaLuWr18Th2O
/U+R7qBtv8JtYMiq+C4AfAGr3nFfQCm6SqaUL3DXzXwQ2d97hJc/ZnLwnQZLgb6XLSflC1vXvqHa
UxBOqYCX3KtuJryBnPRd6HI3xYqapV0dex9RmQs8jitr+SpeZQvGPQ61+qMvrg0A04WvR48oUuvr
/2ljXabNtpN5RY7FBN3uqJSWWlGgTywAk13vSkF6qMP+fGcEzfwJuycTkrPM/K0woxpwa2WO4U1J
/VIe1kuhozpCp3T9mfBEVUBxEQMPkpA1pLK5OfE6Jn8w2iVtYpyVIR/p3pxn3AYADcEEEW5+Lm26
MJH5u7yIm+C+BtKW/vOIN52OLxgwSeHkkCxoXCqD8J2Rlx/E3XbRjk4jNNHERdEB8r3l5AFDwurj
68yS+zYys0pLIfJFQbu7DsbdLiOEloD14xst0Bkod38y6HQVYzga8eNhOCUK+vM4/X2gpBjOrHFl
oWr1BVOYHTcsfTecEWVd1LFxrMjUqRuLCOxQ3AZFtZd57nem56HW3b3KTSocy24+D+keY109Mu5K
iITYAi085kdv+LX6xVEuz6b2GODY6o/7dYE05hPkXaIQVwE0AMn2Jq1pkCStUjyzLpnoltvdeP1Z
YpT3wtIdt6wnhX/P7YjpbY3JNFlmRzh/0uKu3YIeBWNXhR5QMXY+gbZrvGJLZWD2JFtf0kh7fJ86
qYIZdJ6KaH3fWP/Ew2HGg5HNh3I/g7CkNGQe8rw4SjvYTfgLy2RNmXgf45QVXP9Ediz+Mmp5O1sn
on/yD+H+jty/qrIgOcmWXSkvETYb3dAnxqzHEVGowVqgEL4o+J2N9MwdxdL3QoFQRMhSXaGMRqnw
n1lRle3BXdFkUDsSpKWUNF/Mnn4nFbJ/Y2i94mj4nu7toIQBqs2a6Qf1tXK5alJmqj76fkVV4w5w
janFQ/B4Qq229GXO3AFhtMr8AkcTeAGGlIHlBsZeHXyLBIbjZaoZHYOd3QBmFZEkntTB/pSkyqIl
sYkjZfLRRkgiYDXk99sbF3f6tzgTfsk4GakrpLK7kBTvgUNY1IJyxD1Z6oPEDkMlyKtRh4JbYize
362ocU5dRRdOV/XD3a6bbVsPiC7lbxFnshjPN974xRleNrhxOR/NZzmSylcM7l/lsBlu1u+Azd9x
NOUWS6Yfn5C3jFbN32fdj5BJzfDvimFVAHTqPb4cRo8qqEvKwAeyCvi12/OOcIXTOsj83Zx0NA05
ds3aOmEuKHCowMLR2B6mFOhlw0ulN66qNOEuixquAQ2HdCqIpWrztp2LtYVbcwHBH9tZijVRCgCw
gcjwWSJa/U+5v0/jjLKOgsUqlaJssj2kxlEqk+o2hixXjfBQ/Hx/XhthOOUOZ0AMlVCMcKRiJOKG
eJ9VUDlcZDRPuDIg/FOdZktvJ1L66hVrLwNGFdAar8OBbl4Rp7JsZLo17HFv+Oovxstwi+efharI
AEKdiWMc5CKIcnTP9J8pkbYCZ1GjwC+2XV5wink+sicGU9ERPa8qfFTnSdm20SYm9xj8OGL0GzoT
UJyqxDfEGa4IXg0hKRE1kH6JGGxb9FmA/5qidv3HzhLw/tNp5c8zB/BTOlNuBIYsgjUxyIPUvViv
AbfvST2p8/zCfnAqtx6WNligX5YQayDkVtrXwC8KpcWKbvvGh9EbK61z9aRIaKTnxy9Wt2r+3WvE
gozEjbSsrdrq0OTp+IPAXTPpF63ZoYLONNyZ/GBo8z+530bnVAh0sLhhU9d1Pgj1fgkWKx4mUZkU
1+WMWWeL3GX9va5/gcn8Ci+RbGKnWjaB9i6a8GJbDh1F9AoG2F1yMzHp5JldSrsY1rNfi02e+EcP
w3bx1YTIXK3Ti4AZbaISwI1JMwxSFjoc/4nmUmVt1IoFsUVz95hh6j0rBb6zAct3chvRMrscAcTA
SVemxjDolAGIqTwViTR0iGBbP8p9Yhqam4XF2d+3YqrtTNYr6WmTJoOpNgnm4On0t5zxP0gaaF/6
A5lYkor0XLecimt86uxBj2hnHQ9F2Efa6LM/MhWmYmgY3kSjoUd1sb1jhQEtELL2l0N6vQkQtIY8
QR+J+zl3VeAOsLzK+uTQxHuId5IKdUn5NcXrkyIluAW/26rfS6PWk6hlRK02yz9fe+799DkhtagZ
nv89+bpB0HSCtFPozaju0rQWEYmrehVYUDHWhyLLdCJWTm6gl61ca0XE4TMMsKxW8tTw7TNqS0q3
Uuk985O3csy7gIKPV4PjondgaNieKp+ps/mXR/IpWnzKDIDVfrY7DOu7n11HrK1zoT7Jcr+/WPj+
YAH0go+nN0bQTDGBh0YvUwy8cAVJfedebv58gtYjKzxk/ECIPlPEFUGG/isADm/dkGtzqVhKik9q
qmycY1vcWfjQY4BiIIfJpeib9YsswpJjDG7Jn8bjjVQGhYKKpk26kTFFLJvgL6RgnlA3WqOMDE15
4zxFX5cVHE75zCj9HJGyLFvSScewHa0DRPiTz3UJQ8M84+g4Wdqyitcm16fQHVnqXyWCz3Mor56G
SxeWWWrrFedC1zPaaZrnBiBo2outtwrzkf/YdKilwAQlW0Q5vpYA3CuCHRneVnM8kFSBkZyVkmvX
1H8Dyc7z2wJCfLn4SOUuRVFCVBEKFBfnk/EKchVYy8hPe1idVf1KdZD/NrcL7zs1yqaxTMT/sDgf
a+tNw7uMZ8dnKbBsBKGiIC/ctETKAvtyX5OOQd0sN38W9cE0CloKrq3VqeK2XgjLEEA7Y81LCsG2
/xFeSdnGe86ksHccBEV1Pd9V/R+Xp5/YEF+KZq0xnAyJOcpb8TMGS6qmVqaMpgRg5D0EeA3t6VO1
ZTATtpBTqzbMF0sdkGB2WU2+o1Av4O6XhxoFjTX2GUAUhy/59KJZ9HlkgYDr8blevK56tZcwDKOt
tsAHz3Na30a/XdDesmCfLu2dxoEcR57J8zi77bRc5O4wJ8QDCSdnOOr9X2LzKH/DFKQajOQCFKKx
J1TKri0cenmOs6Ed8V0wX6vWUkVTKq9Dl6owsqtSId4gu/QXYyXJFglvqH0oogg+Uu+4KqZVRQ24
CloV/biRq5hYhYiipgU0qzKyhTjUAtPRY3JEFYhUZqNnTNfEmlRU/lY4b108eq3ZxaGJHqxYgHIO
8ESZIUSEV2S1UEu+JMnAFEb1tQ7+l6zYLhZIBJc+3ZGrfGuJJj8sSvVjy0zIfZmQFTtJv0OlSt5+
owjMPVETYZlw88wLTu9dPRKjKGQK6+mUYR62jNSlTgriI31r3O/BGKDLrUm6DtFV7IkXtCrIVbKC
M//RZN4mqSXN3XNvrahmm6807O0wiHN2ZJt7pUxumtZ2h6OKHK+7jD3htUjHvin5FngXBgIv3Lca
Cu8MQ9hhA7wgwUXTAXFu7nEOro+Y3vK/xo+wOhITD0iMSvPkHMK21+7J577w1iiFYKCPs35MqWi1
OyoZULZvpBX9g9B5eL6ml/ggObt05YIsHUgqoorWD+xMxg3nhNYFSU3BityLC3OcoXcGtCci9sPC
BykH4q2lLIJV0dEr1+aQX5/gjewvERCmpfMQGYxyOsPGkWQ8FyrohFyiIoOlFQFSBzJEGtJwUFdH
/ZpXIBs64GU5RPNISICJDtl+O96nF7mXyG4FOnBmblXbvRn1BvE58nQgQ8X9xSbBQYNWFR5Yw1CJ
WTbTq7hloBTLbFdyeEiwcEas+evl8soJW/Etja4B5ZfjlZMmxaNpQkyUqihyfl+k+UghXIC7ywYe
ay+0/BXkSyXkS1mYgiEMGJCu60n0k8yZaK7OBfXk7KZ2/laj8xkV3p1aOnSnI+zRMTVDarR0FE3o
zQb/L6QYSZlIaGUBNRG8ulv8Xtj0mmRJZdIDQD0v/8lLQO2asMeaxGLvPExrb05Z9m/h9cC3+lev
WSGp6wgLTiaL45c+XjKVc8+bVhEaBQnsW5ApUxW8bnIWDFxyXlom4oSWv2bQtU/XRFmgkVq/4EpB
n39G6vmtJi+nEQ5GjAQmR8EXDmc214oDJwaGOOGk7m9pqV7+ln/LXJxrLoGSeggPDPphDOaQZacf
QS3spmlrir5KGxEcBq2Rpl8gQOuN8pGiZOME+dgAEtPzGj4MuF2oIS6dEiHQYjRnlDow8VfMxciJ
fR3jsXyitCwBpQqHhGHxBJScQushTfWKHiQHUWAdDTbDdOTmcVloJIP5R2giP2941y9Dyr7MkEkL
1Wi/IP9Zo9YSVNLIzf/eazeGBjW+Yvn0YNYwScCUwmfAZO4StE/sTIGa6E10ql686tgaSkMI7rub
06nYC6YlKb9/5zYmPuNGHYnJsOvItKto7xk6cRh4NtIYCctumGlftph8xwY3lfdoea/sCjMffZxA
qPxAgZZCDjslBBbW2ywEEdTv7cJTC6+tldjHl/16IEZy+x+UF6SVIr74mUm13KQJBd0JTJoZPvQO
Uf3DMX7iLoX3HqefPIt7a4OS3nnVUkjjxBwY8camutOWDxHVqkAxbsuSZs6NZ/1WixO1ZnsL33tK
aFliSKKbGyymIWHZFUSQlFTN+D155P8++7Hhi2d7FdZu2ekC6FxpGFsm4NaKm0FqPiaMG5hrt90R
aeoQzjBhWHFO+Ho/RqEi+kFYJEdvFS8wFSC6GebLzCf11On7PX+uoJ0P4vZTFcM8S+Tt/7aAMUkc
tnFgh7kc3LEZ0W+i5pb4aFCmGzZWVOWuJCWimlJoL0xcbxlvuE2BjL5m3wz7rpnr106o8meoDzvm
180NQNfhbXGoaiF7Sgi5FoElx2DCW0vH8hVZFTWeVuLIglyY+4SS+YHnxCCbrGgGPJH5TVM0Txax
KYev9HrA2fbnrDYOLfmnPCVrRJrhv3YASc4TKNGwxvL7EkgNxx6CgL6BjH1HxukJI/ctaC/JCK1P
3vHUhajWcE0her+lA5z1PX0HMokJBX47vSFf1cQDJfvynXBSO2F2SmwbBS/aRLQCicDaXtyn5GgV
088sarS6uxJIWurSR3RTb/pPsaaZdkHNz2CxrnP467PzaNxX+8aJ796aryNJTyZL1vfL49YDwOpY
3oGEOLQEDRL2p4aKI60eyUhdu9aKaJ+ZP0uMYlAV+t3yhhxH0NkUamaATVfviT5weD7f+o5L5dDH
2IBAnyeOvPMDaoB2dftzmmlxbkWpk1COfTNQIiz/wzZuxaClOnZc2+4doH9AXihQFSnTdk1zEB0s
IEGNjGDTGK+asIjX0M7F/tLzCQGTx3Rz+hAKKzy99TVzkoM6CLOAJ7yi4rtRdxm2FOa+7Rn1+6ne
Dycqx4+stDvlgbAUKFW93M2KxVDjly65ynD+vozYoo5XftetvydISxMEgSqP+pJ3PzM0m00sRjVc
yMOd3wX4ebj5XbilBHlbJeOU6kv9Zx/iK1aR+c41c874h6RJkACFtdJobIBbmxtu3J9pCJKi9szt
pPaIT/06WJCB6macvUB+cqqy67N+UicPJSpAVpM/inZrmUENyHT/iXEYJGfLxCnWoJYj/7KjaGrb
CfxJzGkA8UsTzfdyV26IlAbskKI2ymiJGhWYLTWB1gsLvmmX0i5Fwrr51BWV2o/MN8d201D5DvZ7
Q8sT2hbh3UUXXi0W/T9J+EA14ZyKB+BcEnbPEka+K6HmJfTHwZolwIBrVe6jQ/wS+WU63pvnbr4m
HqTObBZQ5ER0magJ4U8UppJD/p4NzIXyTkjLM0ta3Yd4UaSnnAaWu1LohB+6o70b96WNtbwYV2ZI
1gKc/yMVkEFfNrLspG3KVdMkXXfvvpzDx9XAkjr3Q2q7IT2KPLFeexIPk5zDnypPHY51Zgjcho3r
nHMPSkWhV54he/R/eu7eQTsVfx+n5SCFfxXmItxa1xFQ+d3PTNsHVdbhDQUsfobVxyh5ac3xRs8g
MpwDpiKlai7tTsVx6GpdYNC810fPWc6qlPKABzk23KNvE30HcQhv3prY3W8VPEhRXhvITKkstR/R
CJ0CCMmQxhnVXyrj9EUIq17ymYWLbCVg+4nY2E7E+dXJCgZojbIvpU4R8iiSP3WccMWWq/eZog+Q
HORpp0nSFEfBa/1ZhdgAduYjnNDw59f3woCADyv7NYYI2VGHI/8xo5nXdmSd5A/bIMefBUqel9rb
29umyCR0EZEB96tb8VYhGzgJC6FmLMO4067ZJYGN8NxGAUi0KNRrBvX4xVKenTKHhqcstYlWQkeV
y0l6+sZ+WNjKkY5Oo0XsX78Ld0qny4eVOoFFCRfqI3rmMNMulbbCc7jtZYgoaTuNoHZmBND8tkFg
I2ie9iSLJSW+iNke1f53U/tHvfZyrC+dJxAustXZKQYoWQlTWe2VegJGSMNLX6my7hE2zrGUPU5K
PnZtL30yC3a+7EcHKQr6xg75TRgVewz2YYhIY6U/dB4PxoliGkXNO9o7+iAO7ipKuM6E3gZGl2nM
5Yz846GarpyPPqQPUEwV3iA1MPJWwHNruT91lnqbuxPo85HU2ZM1H4vlDSSz0JRM6IrTfAj7rzGC
diyJuwwMo5AhKZA4U02UJgKwGH+ijuoQg7mPJxtxkv/ofuOIHhdIDms3vBxRYrrFWCUOYrcw4Ow3
LdD600pwaFTSm/EQ7uORVjkGqDhXnrNq7Mi7bvKxkA+1msQq7XOwQ2tsb35gXiuX7vwmsvlrS16F
a0Iq5hHcYuohksJllt5m8wN3e1cu7vO7l30s7xsD7UZYcI4a8u+Nv/JJGzjeUShCCDSIMD1SO2Gt
bZD6+ME30hTGdOQTTZ4+fdq8Nn5h3jGGb/DGiStfJsbKNgaZLHC6ogn0XRZ9dcsNn2Fo0xKTyRij
PTm+dTW6R5j7iWSH160Yn4ntbv09BcrEvnjVt1q1ZHV2xqN6WFf8Jga7d2w/sm6SQ1SUcxiHiLkU
BqYwuFQM68VIW/IWEB/JPXc67LR3ddFbvWWOdkFR7FVxG9JdExwLmhsA3cIGGdVx8Ns9ZAb2k6vk
e5DfbfDKd3wQRBzSZ/RFC0LhAifeSXYxSxPrAElfP51IpOUzs/CFLrdI4YK6dtDuUQOquzh244Wb
MFCSwLdtTom5zD0xZLQ1EH2O/02wbIWgivGnXj7TUnjQxyM50oQk6QcDEHtdKpZ2lJ/LYhN07TI2
rF5t9ak0HV4WLrcji3pIorMJ+XhCgoFt2jRJ3GKk7pEW0oIBU/uaLGHQzzacafhUnaiNaF3rvWQP
7IUiwVbHyjRtekRlBHfPmb4uqeRdJEtVBxhd5x24fcT9Fa45ShbUqqPms1po+03fJSw+Tock53e5
qQ9yg2W6eqE3c7AQV7vRrL2OvC1sKDfvGEeaLa40sP/S3sWV5tJg2wErDYpM0j2O/+ybaH7LNn8G
twgV+AroJZA7ksiUXlUzuJQbWxsPhUuD+0Y5AE2eCQLcQf9lW3kbaPrdI67vc2FRNlLAeYMzYURB
9+Yur9ndKmXL8IH/uWnZg5msPKHgi88WTEks8dTgqSNJc7ib0OyePYZWN2ytax5zqa8XrrNZ4/lm
XXrGoqJi9bpbqZLV/CYkp2Sd5V072yX7BkfCnurlwYA/3FN9bD2sOg+JWxlShhfwG6MseNewUJPO
4Sv0j/cwVjf2S7xifiSj6gVV8Wu01ynGHaQygjXti1bbBBAhcycXc3eYHxe6tyGPt0+IGEjlLu6A
7CO96zbW7ErPwgpiNk4F77o4uqAg+KKKpcbYJqgxqSzbR6qVQGPhSc/fl4uhmULh3YO4jFM5vmmF
VtetMDLdiFxEx40Zpw/I/dxQ8aUhNzUvPQEXQv+1vE7Hup08vNSIrSDDCKK+iiudj+S/1JbKZtmX
V/fbs1COIS/bHdrPurPLIxdvA3P6h3xV1GdC6sidTXyILJhIgSDs3fF1r1BpvEMnVAh4TkYCnrVY
vF9EdW3pOkwmSxuQM326uITPlj3sPL1dnjZXoIzaWZG+BfZhpI3Yhntx56hutHrRUFRrNtGK8b+L
raT910LQ+58owQy70IFdqErnPWXTqw0kJ0nn3/StVehu6g6r/4Cgu9yCX9yJyCNcvmVXyIBA3xAG
J1KZ5iHxs+LYnxWHRi4tzIsv9zi3cGeLFHg4UMfPUrz/s00rt939T3O7GJN54lh4akOCpLl0nVzr
7oiKJIdim8WhnU/+EbTrOY42DHbMWoO+bE4IXDhhLCRjHmjRHHxnDZWhpPuM7tNicY/NxhSUYvq4
YMUoS+I0AQlyUlIt9sfaHcWvJqdykPJw7M9JRfRSK6xzPuSkYb0bycZWVO2uf588Duuqm26waeeX
3Miv+eqCVQoqNkmZocI9pqYaBMXD/Iw3v52+jm3vR7yVjD/lp4Xs8bXfzXsyaaO3kgHSlJrhRUQe
s8hSdYFD9pf96zbmWQIxRLatYBBroZh+eRVSP6YbtUdTq3SXCIwix56OWcwImHtqAdhTYO+RFwjA
6SBg733SEjWlvVAxteueTJTuzEtYRe+sf4aJz4sgW2qwqZgqQxX59vBxVKGq9YwwPMnlPFhKzZct
+yixLiHxEYBwGTVyZxZlhm3robP5vRV4EfooP+ZOouAuGjfIGaRh9lVO2ekl9GxKBRYLp+llrj6t
h20sd86KMMOZpbA7mEXfJlmP3zW/reNeqswOPivphHDxhbG4HoGeFgYwdt4q//vz69a1lRS028u9
IseUf+wvWw7q19Njz+4JoYkp+S2pqQTWQ9h1Y35BFS6K0f0ISdkJ4HaZrfagfhAszwLhDoD5vUrC
inhOTYej7s6rXfiFW4XVQ1lTzpQYjokrxW1Iy2pTcQXuE+FuT3WSDFpNurDqxVefSyYmUQ4foyQD
D5nez5yNh4lXI1RJxo125cnVqvcv/UcMiLwzrL2L2qXBwlcbaFvgtJgGIenGVOE2v7I+uOyz1WVH
AfBcZpkJgrYyjtK4Ez9D31SXbOzSHIjkYKgwCWwNDgsdZ94EjFMNeXykIAeDPKobXc84Fe8ScJ0u
Met2vG87N7bGWwJ43Rhp6sEEH+Iwq0reoB/zu6JUoYuA7sN5nydQd9nkD7/kvOWVbBb4wsmxOW9D
9GIjkO42vG1qBMVsfFCjhEo3p+3hjYOtof+fRFgiBGbzdwFCefw/DJAlo/spFE4gw9haIKE9Ay/y
0dyKWoUdn91eNVi7eLHGuHRibo284FR7RUrQewtz2/TmP7HTUyuk/KnFSx55bcIeHNfiQFiqYrza
y3zopSpMD/b3Z7/iJc2f7/0BYUp6MCGCzSTUGzy7aKs5YLnUnTM3rdA9zft0I3bhMu/FGwjAZPs/
9A2uVZQ3n9TlnO0k2FpCP75Z5ZQxW6wMMyDJpRZxN1C+IDiCSKbFYPRLvRrGRCeNt6iu035219vD
uMgEoaZkeDtF+QlfRNugVo5Uf/bQLCr9Jjj9mkLpSSff0LdYjcYvlLT4q/j9q4XL8LEZmhgjCz7j
ygAwCZPCYA8uBlG8REjyTRdNhZE0ws+QNqW7w4AfjQ+5fy35H9oJjgE9n7tbxdrv8HDGDrAJsAw1
D4NKiyOvPsVag9EZI83cRPn9Lt3WFkuz6r92dcwKUWc8j74uVthpojeOYLcHqqCxmDTm5dURIfGs
+wQP+qNKvHXP+adBxP1HZy1T1n8bnRWS40g4a6akWcRTMb5RqUr+KV5h+8y8lASZsFgQJfBP07Pr
YU0rl4qugVZyvt42IyEzKLBWd/A5mWomhl6hPHiglFugQt7rtQMcZ9a2Pa0hO4RlgCaE24rRMASK
TYZ1mkSDPURKcv2eHFm4Y9/SBeDZHfGZ4TQ9IdwON4+DpAX/WLBmS3VH8FmG+04GBdRrRzNX2+jt
xbSZVuHzjaFLmc7S5ok+Imv4elEiQ6YY/FK4WTMx16vYLF0s9J8qOJPC9TscmL2emL7dP/E1Cmqd
Re6eX8Nkr6Hj82BSOope4SbYa2Q5qbm3RKM43Gbq8tjS2TwyEi48hmaDWRsKSqaZOd6HVcXS7c+Q
O83NNdIOectknlOuB/ce3Y++WWW3webMvuZMSjHQzqFRFLiveAc6AXitOE7YfZpYW6vpZgcsG0+k
sSYGYzBCPkdXvfxTmCJIld8/u2YaGSY2t6ZSyKCFXXQ+Nw0AKuiqnBVfDJZWOg8fpK1MplpFuIjO
YHwdUARTnv/dZEcxExA3NbMflfLD1iGikq155uIt/xPcsg8DWCPiFbTvMVlum+cW3qyZ49UBVhpA
Y24rtyBoT8HugfnjjPzrMEevAa1H0A0Q0JsfIEnRgf0A0xN0breg5oSIYECu/tpN5g4mUl8CgiAL
gQ8V70p4jvJInnyr/Z44fpaY4qFjwGn2MPnLldal79B3Xga/m9u8lDR05ZUki7nIpsjP4sW8ef8o
1qIpOTEPCqtU4hKgVjsf+bvdeuz100ybtfFlVQgHkYN6a7j9ythbkfB/TJb4A4IU7yHuNAIhf97T
ZH7Zp356EFTY+BCwtdBlJIrr1KBrnBW8bl89pb1R6YBrrKuLO5tgL2yiSR1vyJWRMsjqH/8ec7YX
FibxrvlXJMYwxQVxxF9nEy9WG/lQKzZi/8xIfd9gts3YlgUYha6ih2054Z0KutX4C05zGGQntUZT
Mtt3VeBbo87VWXJvsRm+ibSzSkiblOKkUlcI5A1O0/8S5y0mWjaTttqshdCaEwc1wJc3g457Zk1S
3+7lt1FuLzmi8oJce/eE4oW5ffuDN3jAn9dwoVQmaMc8xg0KsJeOUmE42O3Dfwv1JtzkZgZr+h+B
xdl8CuGpNagmsi7OeRn92KgOKsx68qVI1X1rU8+dHcGGfl1s7Noo63HCDuo8+TebwWTugj1vAVI2
Zfk4FlQ1RpObzWxsV+KXDO3L1UfsyapptgeRxqbk5XCxeqjM3wgyzhtSjXBpWmt8pgES1+qLpuLj
rQ545CPv110//n8n6/+jcaA3wGRycm4x+zCPh5lTGH4wNNyEUecqTsAS/VUARwvalndiq0+qHAeR
ZRM9AcxBXnyQzhYrXAPVw/0E0QvO6/kie16ufBAICAabFlP+ZIIFY/kga0xtSWx/V+KzaZDlmEJO
MC9uR8zvffoO1W3owPfHcUDmU5USHFRl5y6u4ZN6hnjdiZfs8w9lzZ2xRNct4v9AN2345xzILcXW
/b/Ng59jzit10cnNhBLW0Af71EKOsHPHN/WRFInYcB0FYf0Bx1DzbmEjWYHKuAbB5cpzhkChqaP0
uVu1rX13qt9ro5+pHNnmJ03ohV7MwX/QRaidyGhR14DFu31PtyXzpm2n4HYjf5KM1KpeoZttNszk
GbE+LvMn30LyP+M4bm3dBKeoSZNbWqrR2LacQXcl0ZDKFx0LJHS0AQYzoFaO+yXZgbV7yW0Rgv/L
CJrFUUKYSgDGj+s85ed+zor4vIiALSATBnZvTNuX2g/IYHxBeByLNsWrlnlYeqUFLyFASrYQXedL
YkqQNPJUPGeXYQyej6NWEoMVU44h5mo2oRiuHY2wYSTAoWZ866Z7hZa2kHNyZK/JTUfyGduG8XXO
mqkvxlpL3u4cx9Xjbk/3rMCL0k3h/R2c2BpXcsFvtPJuM0IhPFloy++08TSY+/6oEi5/vdklHHG+
+Hlw1u4xV0OivuUzIQDJk8BKJMsG6YWWN+uptaXOU0TyI9kgxXBRg+TPlIXu0sQ2JL1/a/x2ZZti
Zm80eITM7wd+wF7QaUFYXt5eK/AerOnEFAqrBzxkS3GONs/vIhd8RhQx+he1b9j47wqSVrEhFV/w
2mg5PP69rn4WHkym59aFQrl0XqSVpV6cs071T2T+z4QkjUJ8XDnQj8+Py2Vq33IjVtQ8HxYzBYVS
aJbPhce99ijqnQ5TGQV2MtCzPYxC9XGVeW7MMTpQr0wBc9gqNhowwWNkNmJmoZZBtGA6XTXSJ0va
gip5I8yDCqO4z0k+NMYRDVLIPVhzIu8fUF2DhJFnvYJqYJmhhjr2Zy4Z/8j9vTb09Idfmir0g/1l
vMxB59mrD1wDfdSj/dZkfnyGaLy6jPfJP3v7GuzHyYY8qW3Ako7axJEk/e2gNw82QXCoC+9s/7Bn
RKJ1w4mAC1ZkK7Ab1mXUzqn8rVOIQo4HkLXTo6UCsWX08k47TTyvUqZecPvhsfMg3XXmQyiGH8TG
tC4RCC7QNlMUbaLY0bgArhV4TutLQeayGS4ObN2OhJNH89dTqwrjv67j/91hwB2IVprQnZA85X+d
aid8TKw90fCOMf326ztzJrcE1No9HepOcCPOLdbUMzL31avBAHFkrx205PGQT3q6uwfjegfbn+ku
7qSVzZSUDSrcj1IFXmNHvy1DgBLThDNi8gBvvwvJ5EYUzqtuaWiWqYYcUmz9dqzm2+CU1Cpv1vxG
lcbjHY7yufZrrQ6hI8+C5CCoAJdZRu5Lo+gWHQkrWAewJU4BAH9ZX9VV7krcjWu+R8eTRjkPIjd9
XyQ5L69O/gJE20Xp/etKtk5rzB9f2jRbAuzBok7PICuTS65ynDYw8nYsqiWltTqbTyq9/7srnU/3
gBNWdGFTBOrkJLfYUHKFK18JosrZMPoAt5mkDJK6Oa3TiXjPxt27ZIZCDIsYjTqnLf/vuDGQIERd
ACZcOlNk4rVesMRNMa+VlNRKjRiemhsHpHufX6+np6lQHUcR3QuCPMO7tlHQjQy46AVlm7+HSoO8
Dxc5vf+5nVOcNM9afERq8DyTbLUp3iYOEIjtU7YawbIU0UTRSa+Aq/J+5yThlwN/3tYFJyf3u/89
wRKhvqYOqhlE6+ABijIwmMQPtt7Fimhz2gIKarmBKy5EMooUytt3t0EFPF8LgbPC/+WLGK8VFTYt
yx7RMm4425rkYOb/uRh0vvV3m7N10cmjE8jv7RlLzDyj4tuRUL8QuuKT8wb/o4YLb+/Gy2q2dhJ1
fAsOU4jwRYQcfzuf5LnFxo/skw/Xm672YSx3DLqfj3N/SP6uAY0uUwJVadAScVwq5XMmkmc6eFsZ
lgQQl7trWR5Xanm1vFXyOeMJTmyJ0zgC8nlOix74XFMA0cQjbO6/hh11IatTT9Swr39OB/Y3TF3/
MBkrDTyUXxvmozQaOycN7qvY0hPxfrsIP//9Neap5UlbX3vWN+53X2w2CnR7vsfcXe6I/N06hnSd
X55aMMwVBmVYj9x9akiJug+LbrTSH3Zg0VLtsD6w7L8HyproL4dpRRC8FJvzLhYyGryqbPu/c+Qf
Wu64yFsQ8G6Roi6s/LcpZ0Hf/CWiR7SEivHmxAPW3yj+sa634Sk0kJ0vQxF3SdGDNCyry+em1x3T
qn9qWG2OvD/FMgQrn3zW0EWtrHwI8zRFdbOEWNrj+l2D9DUishROX/oRiAc1fxBafRSA+2zCsK5/
n0K2ngB90/yIDAsC79LZOHQ5AYY1KFytFVA7HtfSa1h7LqLi1U+1x2zfE7/whf/bpJmKCAYT6R/I
cwbB3ytPVXMOEuPcl5fPADFiTrKKu6tfeEunRk3ykrxR1UmFVRrhWdvnPbuAjPUs4DDmt79C6wbD
fvQdz15Z4I+WiKtmt1deo8O7C9QpxRYcehFDVTbjIwzXt8HMg/V08LYfmRcmR6/zopvRJkjHp9uW
SHKSTPEWPTk3kl6uDJkhVHZPMpb+pa/1RfJGmeW2t917laRVYAhHGk5EuE4Y0aX+DOhrCKRO1pDo
MPOwWb2GLeakHok3Zcptz0M0ZIKuWuKdWEPjwZaPI66mNvB/mJh9X+CYu+X3vrJdVorsXHh8Pvi6
YEYkfyv0iw84+NzubIJu/tLlhwapTB67/E1ULottrj9r+nisRdXjA3fAquN4yVkBPkpIrv8hOPvf
KSbqmYiZdHwGm0tuZ7/dTqS5c8u0M4l+vIi3nuYj3lVz9xT+TdcZ6wqTc8hgA3SftcQYp0+LlDXL
uLCZ7hvwsT4uXRNZosMA5GUQatBbYuvBwwtB7zgOho0287YPairCWEYnWeuZ34k4I4JTKHnljI7s
23kO63O9zoADbR/gbIZM7+dj99+e1+7pbjTYZIMtpVJpzLubX/pX+P23XhcHzsN2fl/dKp19KIph
U9cSfq1dYLT9F+WAzudxr+o30hV18eveA/NQqDBUBEBMlrW1hkksfbrQRhkecEYzlNbh4xGR3ilV
rbOD63yH+gUXEuSS+a5R2bbnnJzTqjd0uqk8gTP0sqPSHxxMHGdi2Jxo5ctgQLkSA9/Jt5P7T3A6
/r9nQ6eMDsh3hFkH1wCYczw7kvWgyH+X+q+WfhEwpWv9B8iAi7wpKTl1Mg7Hi7L/0hJCnjmvvoa8
4yqxQ2hCiWISSjN0dZGnmJjVQACLg9GAjarRmgJFHQxg7ABEfYFJiUXcOadGCue/4F3gkLTfoRWI
5/VDfr5PxCXwNOuzacaPuaCCbfP2y3FpY0PlNqRxftLDY1DUJwUWs008YlfpWaoFOp3iWr9hA6TC
1SiZg0fQqj92XiP/kW8rMGf+0aZN6yrcFxFUqI0a32Xk5/ZGSiTpIWLsPIAw9oSzp1e4eJJ+D6P1
hFcLRWW3n27bZs8olsfRpF4oP45NePLlDIx14Qu3KQdn1XTO81rMyMpycl7c7703SXJOWT+MVAKN
ocv1S/OJmg1Gl4d9gQ61eZV5XKZIDLxzHE4Hm2WrToxDlOnlsXFiBcx0ozAxwl1+WR1NnOifGNUU
uWB7hnEU4nR8330MuiQEcmPPXTh706g7UW1+48xjcXvkSvs99gI5oDdOtZNcqWB/0lFAiSR2zUJk
M98PCiizBPdq59bIxO4fyNz11Ixut28fem5+2owX6Eimdbu4NafNYArDQi05O97QHQAgRm2IugzZ
fsx9Wy2qcrnHyZvGydOSN/aG/wEFuREtGtgwVNsFClN77EmVB+zFiN75rkXDXhXY5luKLddf/QTQ
ZAPl/RG75f3RdA9Ev9yQs4mBWCGMOkl7mB1rgqLFrH4MCLXzOYBMuov7P2tRcZwKUgv2KFCFSYTk
VAk85IXfM9s0eltwoqmivb80cZbHCxVfktr8Stb3GVDpUsFBEfQkvEozpuN0GAdXUmLqsDppo7s2
svW7tmyW/QJPHUtLDlJXiVoY3yLiaCrftXDtxvOzZQbVAFA7JbgzNcbcyPkTB2bC3FWVT33AAMlJ
k1/rYK894LH8/ptmjpnxDhhLyTYFkCl5CR8GfxtQwOEKyvhKVOzlhAXqUyCLgT6dSRNGYsIiD4nB
RUX+Fpex5EDaQYXVxUvL86BQizguuJADPjNr2A9M8rauWh/QmzHGfeYR308PBssFqj4cGc0+1jkc
n14LB03NuChWETD9h0FFaaPlGRlWSbJHD+6wItOgFSv0oNhhvBVs9u6Mqxg5qAbfrJWZxFVNMwxf
zUXO7uDRKq849iv6EM57B5QmYVWonb+h2MIHURtHn0iszDG5r7cDqPPCEnSPDzze6h07iKNsD0wT
CY7jVjq6dFD6rDhjciWt8H4EnnZbdgzOlOYNyDPQ1EQft7BNeAjMQd6hC1M2w/lZTlNaWzdXpUce
G9I5HXmZmP48FAeV7gM3pb8qoGLLFbLuaJ84+pv/w7Gqv6KTCq9SXuuNYo/RwTV5wFJ/lULgAK8m
Yi0tovCD1NUAnftdahEjbLQcKb+4p+Yu3XF2w/1cTejFzlI9GD4c1p0Pk9VjAHgISeL0a+o6vZk7
MCIcuXPjGUa7b1/m96FmvxfxLtX+yu7Z2tOMAfiR0ebZmPln5ixcmeJU5MQoEG38hPQyQNp2NTtH
XzvqhixIgXEc6b+l9lGRR81sgSrFP3U8hJCF1I44kqlhENeNMmXyVh4ZhGmWd+HrKCGvO5+symRN
BQKhJFrd1daL3wZHsKWPAg+3LWTO6nuOwY4s/YQ5gUw3Eg/oPCiWN4WliprLapaKOQEa3ipoV2k0
Xl6+f4ZocnYefuznzWMaqdjus3Ds9BYaimVXrwr/LxT2LHXxBgTMiUA9Qfe1kDwIRxg7MaHz2g/h
LNKEOQaTY1TJvXOaV7v3MVLYOuGe/fY6Jj5NFCkpNLb76mBgtkpeALaPzgC5HNE1I2CTeH0OHW7z
Tu2nhe4f0/RXx+NNYvJwYdFE0G2p3hNJisqEYwFOnzdB+zuvwhO3QAsaak6Fzan3FymX6TBdBC/g
nRYu/yySzXlPCb3PmK2aAiVpItUBOs2/yor2NOJsCyDOckyD4dZpzV51clFn+DmAH8jb1HYg3z+a
rmVqt04ytZZI46qMpAMhLSuryNCJErqZCZ59Lv9r8eZz/x5ykeQLCYlR/byiM6OpgwiKQ9/gaLRU
3LWUDVD3BSdEpcG0VI9GlmkULfUW57JjrxmRlx/8QscQzr+ByeEcZ5/PXGD+rCfpFuoC74KRfweM
jNKag2nBApj+Au4L4uCmPryq2kkNP/aSz/yajU4jsJyZ+5BzHY7ADlyj9HVxbuNED2iXe4rduyJP
AfkQAgjNCbh/gynKRLln094ggppm31uqwS5li1f9a6gDLvBRWk5BI7BninBVS5oG/U4iQFR0Z3ru
M7Z//2kRrNIs99wHwuzDQ9ns8ePEkCabb0z0q+nI81r5HojRZ9KPkvxNfvCdUnbqhwKfAVBChKMc
lAgPL+vXTIlM9pIsl3MgSaJOHoTcRv9hfFrbZs3+0xC2vag3HfdJV1tuILrKZTFrKtYre0Uo1xAv
It+i7BCRcbpysJEGqoQ+agld7MLii3lt3md/fNZQO5wGIPRrJcShgyT4E+3GLDoeLnEJbtH3MWO1
U7FzIpfc7RO81lrZLolRhUtYAmlpoh7zUMHpyMUZHzlRiObq4/xBd4lNvEMCyfYAJG4egYsxG0uF
pFcbWhbAfrJv+lBHCDjEDRBAP00vxL2gjD/D0aKL1v8J74KXL78hbrkIXL4Lgpq7VG9s86x48tU/
2Q0Lgeopu4AdTWk4OuCxVQg7yHlG/LEYs2LdhIvetPn2pcAfc1laZHhBDFU2FTQg6V/E2HtGgFON
EEGs9d0TExQU6gh9uIT/kWNx9rOCq11JVdm7wbBlamnlQPUbNSTDCsJmc2UJfzK7GlQ3O+zB+dzn
YpZdz6VzIQSXcprG1FzMGGEZMVyDUbWROSKLYA3K4HIU1NyJA0aumbBv97Sx9t212K3rva6ss6qv
6lm+4Q6toxALSF90tyxvOvfcX9FZg8ZGeZnETCiAmPPI5zssMCO2m52MdTXlwowhUJ9jpmcwvK/p
UjZYbsqIWz7wWz+Tb5fPUasV9BqA4+7wvdcze4UJ/ba1OUffxT7qYCGUuOW00QPgMzyrsb9N9anC
LwoHJu3m5qkbRBXDoeAzrUigSHZKtXMbYdCZ3zGdSETqIoDWH1I12USdyNAtA3kNADonWnV8EdMS
21+WnOj6aVHB4NKdGCRVdZTma3YHHioHbjQabrJcPW5WeonqOquywZZH5yzvPaTKTOJ+cXyZvvdH
kD974iurblUMF0J+3y2MnK5ytqik4s94iFXNptR7YYrWXGKRG/f3eQ6AUGtpDa8W9VVSbx6ALYqD
sAPBXzPf8sOzuXzIE0xZCPGyOVqThVjZXU59sZHjKgZlg5iPxR1BX1shnhars4GjKQvYsjLwuXhm
6cHeBKCalbDxW8enlyxOx/dYNdMZ62hE/8/SXepANxE5IML41aS3Ec3aN081N2BiuCjP16CL4OTr
vH6FlMwO9vYn++cqxdw4L91FNQTIHN7Zb67XE5IUyVNiusdScrT4ELZTi3GjoBWyXNsL4aabTdWK
84PoVvrlMQ9JvnmTmi+M8fzQPcgU1nhejneb7/vibkv08I//wZbObtHbcuq0F0uZqjuiauBA8mRy
coBSNFyBhInfCTKlC42mCbcZj310QEc26KvIwFskgMeutk0eofsdwYxL+Jh30hq7BuUSA/Adif0c
B5+AfpWWfZC+HucJq/ht3WsXktP+plQ39tTiaim+/MohqUO+DZsbyXvYLpfwb5l5iHgODe+ox0B+
WHYGLdxGOfEM/v5aAaXBUxLzNw8ej/k01VKUYMQ7I2OwiJn56TbWBiE0dbvJl4HtLgA3Kg8BDvlE
2lGrUWSddb6K73GwiHAYODkO6rZOwDm+2slAdOyEcTc++IV6DmU+v2o9NNO17aeM1uFjocE5xB5F
liAjsdp2pIfFz6zUZYH34YXrQu05az2EkfF7JUWS++eJGcq/7RX1e6Voni2+VG1VuM6989srI6ku
qnGdjyAhjjpw5zrg1c1RF3bOL2MvZvGzzR5Xqkoz4dXpAriNIBNZodr0NP91PRstqhaIe/RspOFl
vZRd6ae5iKEAAzH4GqbIkjkYsHZfRwDgcQJ/m3awQoCp9lxSKY3B2MQtWQ3zd5CkrZnoEtSzLgVu
x93qtYGkFafDlXCX6mA9H25ZCDO3Ps3ZabSq3rNk1BuvXKkpJqrWVW63Um3w25HKs31DD2CPhLgZ
z0mO6n/OVGyKmHevORhoRStgM8stel/pGnbN695meClLnB9FYPBY72QopMYLLotjHgSkCZtpS7T1
KBb7yyWQHSUoFLAFgDb0HDtqxomaAGN/41VkylG89S9n+GKxFMVGXagI4WVj0FDXLyQvcXJGW5zi
+RzXDmlC3q/TirOr8unVi56pY71/TkY04xCfHwIWUGSGtz1V1Cs+zP1Os8jhb5MZchtOxQnbZpBo
YapkWrQBvIJvpi6DKOJ8g9lLllQvaJ7Jxg8HbmbNRZz6n81PYKz0pT24s64HW2DaYijqtYwGMmtt
eZD3iAAxE4jO1yzUVSZbd5V9mLSEQd+q2i8qsjLf+DgI9/0F+elMu51zcdjv7d6eCPT754fWGw7u
XAviZbpFTBkmprWIqEyvRFf0qcjZlOwMrOlwbg16m5MFKwD+r0bE9bzrWYjPsQPEJa5k1OUvw5lR
j2pSoc0ex6RQnC6tDmGPbFbnC/EyT5dhV/1559o87eqGsLuaYgiixg/dS2B2jbUrrA4fueFH9Lje
nnXr4OoTiAIWhzM0aeeKV/lIPQ1FSGQ3Y7C9kdTCIERsnlnWE3Ip9eWCk2wBXWC+0EP5I1w69bQk
i3Mri/f1rENeHyZ6LTwbRDSevXiqQTD113zl46X+X2bT83r1lw2VIyisgdz/32NAlenm9vSf6QfG
+U01i80DVdbfarTwVx90NDCyeXBe5eoKZAeB5CzBwzSxGbkRZRNph+s2QE0PizNX45SZ088AePRt
M9TEt5UH6WaOBgj7X9tgr/i/ja53vNxS6O6UDM5fQmPwsqE6NfxKpsFwLlMWOfZthUdW9b47i+2m
YsD/R6CtBPHrFqUtS+oFmQ6gK0+I5ki2D1YnlgRbxevGAEBRMUWK1siCReNiJUK2hlVOZn9vnzs/
fMLA6BVLffJ409dtTnao5VT0XryXB24zWnnUl2YVOUoN4Q+tuwkpXT3jwf3jC4FswjZZYGKdma8T
A6rYfqjJCObtWRFcR0d9FMbAsiEbYjN3lxoPpFD2fFF4TvGLmb90o2zXBScSZrz6pu+KITOCeKTw
iphMHOBi7lxWvpvafW2+GqygauKyYcbEF8zPoHh2ese/63QB7U+KtwHyweA4SkWti/g7uWVvF3b+
6+s0NNtDhCtyK7Bx+yGAxHOILDoQ0F8djfQGrkOM6+q7Wnt7S3BYVq9oP9NmSAtHNdh9pmpeRsQ8
vl3Ny8c+9qdX/xIQEnevMINqYSBmQZUglUVZ4+ukJJvFlFzs34tc0FM5TnJVTYp39lyNNdi7a6BC
TXEmJOMQPkgyMY63Anjuw6+PMX9XemQT5NBti9ewJLCUlBCuhGXCix0o8zjWEy0l5PxNNKlCY9/2
0bSKbCuG/B3YGCLl7FGJw7EqF3BQStdEN3YCjW5SqAIV8AgSkuPq8g37NlJoVDlUdxqXBU2pHgq0
lkviKDFekOFDgdygLCrVSDpk8IrOQAdLV4jyABrV0dwUQKMFinW4yZF4Ef7Stw6epEyoBGfMgF+/
5mtK3VBMUYE2qLY7ZXuaL6cLa5pBcrO85buA74M/9yB1Ib8y7vJVFUaHxA1tc4aHPjawGACT0uPy
hUtXHSiPdwmceRTH5kGOQyrj6sL4uBz/6YOBZ0lxKkDfyekPI1nRYEHmoe53uretk7/35WFSMN4z
g76rtSQ7D9Su0eXJJkqUJ9owmU4ZnlZjL9Y0YYfjwgFGtff/TeIPqzBAPQiinb9hehGHUypSKpxe
xrCjlXO/8nJ0b/pIAKAksX3wOjscg1AhIGSXmrAGN5EwUSmg7jJdyieILY+iGAQj/8U3E5Mo7rJv
owkC0zJuyBaihweJGoXtaTyfJZbszSIJcwLGyx5vPNqGMukWNlPOqVrT4VIr7YPbw1BIuok8OcTu
qOSU8bDNeTpWj6XrBOi/CtrncFsh0ZJNzmW7Fo813tyWuDBUaqzmkar0MlEv/QzbnQTYSpiDjvIb
Vl45tNrxdjrDTuvtFGBKZb2DZHkofuwZbD7fcr8/4N9q4uWugWI7HXre47+emVDkrKgDQtJzh4Ez
zYDxvdhi7/Urd18YX3/D3v1ip3T2E/5p1gS1dxl69XnO2EaG1gfrAp5bn+0mj1KmEGPax6LRTPdd
FHgNmvPTZMauhlYljo90I+S20TLi3sUg4TKQYzZYIis5u6wk4J3KmN3Mk64zy4j7ODmHl6vwAAOv
N8PpklUZ2y684DtDcet6H5Jh48lxLkLA+1DhVgX1i2P3IPBb4s8ECmeIC+RUVs7Rv4keRzEuwSGx
cmZcgO7RNtsDNqWkiTUWE4q46CYiylHMBEdY+5W2hf8rIravVh6+CiL0ZjuoQAyngWxxQ5X+pFZW
dj6TZF5wSqd622Ldv7oXwcyziVy4Of3XdkVbUvr5KYnn2oI/Bjj6qOTFWwBWBSOJaZZw+Y4QXTOB
jL3kLP5c3oIDmkpAGW7l44MmSrJufGkymwhlTFSWXlZS+tt5QY2RZElJ2b5XTrYRBkO5aqpsw5eL
i3J3CHEpcvWKk649gCwI4BsQbc9aQQeJ28qnUGU11B8KV/1fKOYdCtpbg36fNcr1zP6dIQtxMOyT
bhlPEX6VbYEqUTkod7sKhz0X2dGcwCIr8E3jfscLdK62XHmpCAa3oFOb6o9nkvFAe1FMvO0N5M3O
AFnvTNdcW0GnkNPe/sn1N1gLGVQ/AmnNANRu0VTCaZoAZEvTtpEHVIZKo43nbj5ttwKM8UxSPfHP
w6NCuQgKOtiCxzk7CFnkCyU/q5ASmO04z9qwJOcLXb/Q52kpmRfWQ6FOLsTXWBL5qOW85T2NthMD
+BKmFfWejV4zHP/+UhORq925jJ1c0eX1thSG4nnTY2VbjZwKDIqJeUmVYINpu0tMvhoInIetwyQe
CM0uK85SpMxiuqchUxDSO+Q/OP5K4VtKAI3//bDKfUVVaULOLMXNxDUxXPrLlcl9oYRu+3xjHeZq
u0A1OJKo0sRh3YYXYJipXJCWRDGTaWUGOWv8qnskjcWa9lY6qFcCIyOsJy1tf4Ursv/NIkv/RNcr
5lxDluxPJD+XOZb81985aCcqYG7dV2jGvu78OmlLdUAOmrNRPIHTTgNW28eiismnoXkWQyRDc2L8
7nP+1jCngHbdd+uSXToW1k96RaHs+4u5JBU/hdlMnaXCn8zcmZLV2V/3zGSnpk5RXW6W5zu07Do4
3zzlA14Euuvvpele7QO08DOoDCgGgAnGLHd00+BKDfj4ajTz2PNLbu/4bQRGww8iReOl0Ig/KlSJ
JwBwhX45ngx3K/Mqz3qk/jqEXNJQKRCMpS/C+o4LkeZZGxa7fbVRhIwTXg9iSCCvD12IiHeLGGuS
DKM712EcApQBDKRVgwgsHnZlUGRWZirgCoL6Kk4PAQY3cQWtH4xpT7nosLXwBuSgSWxVsf6Aiwjq
SfmGtxREOyBSTB8ZC1gDxTLLI3K4MC/sCwTMCzBFqIzNIItFK5QMHHGZZmO1PHd6K/4y1+GI3C8l
UD4Li4LpbG3lER8ivprDeasVpbIytHZkHnkTLcd4g/LCF7VqzXpihm0V0CF6mcfquQLnozmWN+BM
/tIDeDlKzdLLnM6xRMe+LeyrsZkGsisS7y0IYhbLVGJdaGCakOoqoBAgkTK25Gmg2YuOsLmcxK3m
/m/E4llS/AOOntAVZgVaZmYqXNmDtL/oGTe3Q999qqm7kxoTHv4NwiJRklJZO7mUJCIil8zgjDEl
beCr56qMF3g3MB5mIHi6z5YspEAbZlwkzT+HfQobSvRd74w5j4rprM/JF12oJKHOr6zAN4/XJtee
h4QDTtfzUzfFbUkyXA4ROBvqHbhIevFzcs+4/8hNpajkrmXWkxjOGrAn5sXm3yhvu7etCd5XLhaB
H97VyuK9y9GwblWBaNA6ulxISxXFL1CbIWNzpw71n2JbbtsN4o6Km9lKQsoID2Q46ZXl56d+W+cC
Sn5TxipdyHzRgJamHkR13I6pYcFBhc8PvbY60I4qBYh1HRJ7jAMygZN3mLbsIrwuCksIiz7DcA9N
iYP+uWuUIiP+baaCUfWUK3XkpTKv5afaI98U1tbSvSqg+fQczRkI1UwS71m1zRbQBdz7JcgzER/D
/AyrPtk/tpKMTV4rKO/NfQ83fgoisQgfLFCOv6oUZ6UfhFyZgUVN0p9d/yVz/mTbe+er/Iepg+GM
x9kQ/bq6/I4UNvfinCmdg96L1SqwVZtgIH9aAD5kIKdj0D17SuNAY0oszOJ9X3I+hM7/LMm2Dl0Y
z+31YLKhEi+NDrkhjP3+u+Azohj39eqdnzNkwr8/g+rPW5ELvla32By+dktmcgpEUb3X4NImX7Ah
tB2GUEVhcdlq5WwXl7SFB1jzEwN3n1EV9OJ2cG4wHCR0iNts3s/iWl0RLMWjKkrAPMeml5tcyKaE
q34OO+Q/cYBk77fI/9f/ADpDYffOa69/nLpoVTyvTDQxyOm6wd5L5D6pteYPjxY1WWhD6PdvzUBi
THCRieMrg1cvgl0N9S+ETUcsn1fDVS3v1wLaVjrCaEuHQ84cTHCrzLDM8q7PR5fk2+zhYtoMDTdb
d9otkVjNZ71dwBaOKQid72FfQ1kGvDir+ungQkH3N7UDhaCMe9afx5erBYxWZXTzownYKSQ/cwgz
Ng4zekForzRsC4fVUzSUzlOOKXMpqz+lhbBK1QUKcZu6b3HtwpZJfHfB0b+TyJF4Ta6NesSDaOEw
YQ19sirB2cqgoxG28tfiCRWtI53NGFAKWkvMuqA3FdQS3VLWA/fQbUPuIjR/TZ6OjQQm1yI0VGBL
js1OBch4iu6cEfUwZBLbMeVHCfIHn2BUsEqPKgcnApWQ1HWZVysscTNXLe7lwfMqlIaPtIzbvbnZ
psO11GjIxAiZs+hCJb3vqnA1vDBrfVAkWeaBfvl0j17Px1Z8ufK3dXENtmXa71bvzJzMxFlemFjg
/ehaw98rGQbzNlAKkjuM6KnrfcWyFWQh0pmlSltR64NthR8fPcV2sZNFijUVWKgzvNSVkK7dV3y+
ssWtHdtn/O6VFCfOJvDdS40JfTTpL0KV5wWGxeOW4h5+mJ3bf8GsRAMyl5WsOMYAQSoQmRL7i7o0
v4ZoeegzDLSzrGHYNqki1zvHDz3+ZCeELt8e+Zr/DTesHFrpmW8pEOWGk8rIwdNgC8XhFjcSscIo
W3YDuXRFHxBHn9QvU7zxj7OIkBVmqpBX2Z5aHiYeGkcwSG0j/Xw5tDm6iSQHYLAkf2FU82LGOAal
ISBB2bkBldRskLD9MzbpTobk/RDb1TZ8lT2L4M30CaJkFlqTQhiZHCCWmKZWDKt1hZpzBVshxWRw
jMDDqNeaxiL+16or5DGLSsuTGOgSm9f+CYgnPagK1ivHekyjdyF8HWpmHlP7X5uSsF17D5aA8511
LPBN2d0NUtY0MmUqv+tWYBJb/TS/NwziofnxVgH1RhBi2/HdxkQbP3MWq9+LJaAMFzUjPjyZ8Vab
zrK3hTxqNnSiDIkkX3Fa9JcWIH2kNwodT6oBpMf8pSSUpXfpGiXp0qU6YdGRgnqUionE7ftyfpzr
m34blDuQQdtc8Jaa+IMR19j9RwO5vF8lZZFTd8wjaw9IO1q3BVOE1BOSR66gc0ccQmpXm6eXLrRs
qP4VwQWt6ikjXrwVe3+CGTknjlUTFvixjMbUORsFdWZhXewOctCgOCjVnUO0UtBeqiQJBlp3Pri1
VL+l7g/PyH1nEZCBUTCsHU1Xw1b1GthqEDYkzaq5E6zf+AEH72S+6AJT5s31VYTbmA/zl1vrZSzy
Iz7Z/JIUAs/bUZM7wh1TGr4DyVyx/oUL7OHEjYuy6kx0F2/krcmleDrB0FarNq3N87qvpcB7dbC6
e8JAwEQ0oJNU7fTsInWEjZHaOltVEuVt9qbf+ZlfMUoNR5+NPMNK9g6ncIbsinyjmnkoxk5DK/J3
SedqW8BxEEuDVGIjtr2ht0kI/Y4+VAoQSMQhz21lEFkfAGMFGelWLXX9C0Qd6+u597/sYfhMyBai
xlWrCfBX0JDFz+hRrVjsOPyUBD8osD2J5vemS83fPnebatgg6/mOjh/uhb9URCnAr77Ji9vzjflQ
QCmKMf+2zDYeFWnGGITYKjw3FeAQqEhCDxciOWLh6q5UJnFxUd0CiB79eXmhAXxIrGahlZ3AC1Lm
RXJ9kcm/83uDLcaq2r3BrRw1zmHIrFpJ6qCWE5hOYBzXkc7wcQJK2dHLWInyn9uAJMPwpEq69Dtz
Mc4e35URhv15Y6RTrHVNGJkF4Puam5bSc1F6VGGVQYIqDDdkCvjcjzM33yvUo/IdWS/RQI65C2MG
whmzBy7QZ5inDMowJfY+/oT/5LoR7X+fNd4+D2ryWZFwO+F68nUxxaJa6F6oQaYDMXTjARkmIYT7
Ce1QjviPYTO0QuqiMc1fJyWjH3L/XLabJOkkbGP2S5ho9ZSz/01b1n3FrzH7D0AK09Rnd5+i2aNK
SfWsya0y+wI9gSNBCVXdCf+cmIOMn5GWEJIjengupLnQa6p8ciLTx6wisCxPEl95q3NJv8O1Q8bO
GKMtihKlWio5WBasHXGBlo+aX1K6vevaGZs80pcrFw3Gb351RrWPYjGu370lSxogQZpjii/xZL2x
ElZufyCoFieuB82GMXnN4DcVBVwD8Zjf/tDL2NxZk58PJG4ukxxLgJTmTRjbrBILFpj1nCAiIWC7
r22yCwSNSFwjG2+tghHOff9DMEJm5jX+7zeWPlIUU6IKSXGMYXQMbZt4GRC6uubEHI7csGuF+gik
VkyXXTUSy7MmO9YFFrbURLtjxWN7gV2b+D9rY3/fxHyXJGQZLutwGd2Vuibgps0G33inRFdeK0zG
nwoLjeFc+r/5o55wTXXRrzPkO2a30spXHCylvKOQUIbD1iTPeu+7NeRNj28lITbmAPjribpkWvTn
nDDu9jOxbd2Lf5hgcUpxbzqK5NqQ606EIp4qvaXbsnkVkJJgmYQ0pjdwVGSuU7yEMZ/LgutqUenn
nHTZT8k7v0IcnZ/oFeV76UBPifbIuEvhRN75eAwKx5hEUCiqnogR+KzP53tj58CwYkX4mVCzczTE
mVOFAFEq/dOeH43VWdNvSD3KspZ9WzaMSVrtacyOlndCnL7xZmQSuSPlZceU7tFnye+rQij/i3yM
3q9cVorVEvJYm8LGK13ScRNbUMLgEUetaSrP3/fiUc5q8hYiUpIO06dTbgCZT/pg80LMFE52mwm0
FZRKzBUo3O180T17/wsrJvPzBeqLCGjreMKdcbmYOGGx8p0iwJBUiKAYtusaGaThpnKuhL7WkH7m
8xRYJAjnvE0F8xs3eYvJc/aZcWhcWykQuYdPDbsjrHjTQVUk5pCXMe6I6955cfXzQb94N/YOouE1
Z8AY8d6+xmW2z6x9gVxqPLz3+ZPZYO2MIsawxKFf+jpstoDQjAywkus9uZi4fJaiGo+Np3c8wrXh
8aYhf9ponMT/Nr1axUMgVTkJV0xSa6rIAZ/COXWKH20AHNb8T1gqq0rFvtVws0Elo1xfQrgWN8ls
CuplYgJ6TuODn+XNRsCnlK1XWPw2ZMitPK09H6kVGTPsbD4QUuxH+SfF7b2C2tWbh43gl7CGah4p
JLZ+XGiq+GNZVCP19WnZ8zpB07Md9LRg13N23dmmtyqqygTJWsJ+ptajyuOtzxe9EjAij+kwvoRi
htq71UMoV37cTdzZHwtDb2z4vWzj1LBdzp+qSM2tXALI8a0EliHZ/nkBf3N3MMIjJrzcZtPhOkxw
TS6aasXwRPN5LAeCJN2GL6WiRExS79GkaXIo4j9DrYxgYz2YFeNcGp9EyNa11QkWQTdEhNDDnE6z
vOiE+PbamvlrMDJzWqyAjWBZ3tq9ATY/eXsidDcsNGqwJepXFAkU3xXwkNsI2nNjnjk40iLCAtPm
AFN/MdGV4YJStrnl9ihAB7/Kli7nldrnpTzviqH1rbU4xZOJhWWOrf63gwCuZdVKqbNgCFBoBxH2
/EQw3U725GOK6QuBsdYM+KsHqnW99XDcbay+Bqq+2a8S0JYukA7+rf4SvCzhOBvJ3VBdr1wz93+Z
x6fYyKWbFlbe7XD7o7QMrmb9tGfDJTmAgzhnrBMfldyTJqhW23/1XMzs1uLS0Y7KUD/DOgxSVpof
DNIGWfweOFPA1FYuZKF+CCertUq13LtCuNpSj61h79dlLzYI5N1NW2FWzjE7BSz4NBrKPH56JoVb
ALu2VA3woNEbcwWUeS+Zlvxprjho/6eFZk8xWoHrXkH9YAs2bX8NC7FgQ/pfzYeOkbdD4XMsd4GC
BnznfbK+E6vIakFV8JQDEJz2emjH3tRgUSg/1OxNUvjLqZBP01uRzTekJ9Clvpx9kLA7HwnWSBOd
W7mB7TkTodjcxsYDRVAgZux9pjCRptX/Qxks5l4MCBdQaHhy7AGTytjE0uZHU57g+YOJjOVApK8N
qzHf+oO/eBft3km3UxOwGj4Tq+zpeWPG0p9bcd8Hgc0eXNL33KB6aWtJIlsolMEuTWS76wRo5a/E
VrAR102DdMS3AdTbstOCi/8nH5VC6l5fWhk4hynAu+UpouzmJLriBSxqHtF/Vewryl2VyN6+FsMI
JE5BvwCzf15XIo/5RBDxOdBHI1zGly/TZ9+vhRK2AYppLp1CbKPwAiRdkFnT9P+VdElch/jJ5vgh
OYT6b8Lzfrcc0LmdLcVxP71ei3hdQM9s9LxJylfyaVT40lAFLT69uq2gZcDsfwJhPrb0lVlK7M6Y
q/ZrXMODqCPjAlfdGI8MrkZ4q+ZSPgZBa9Gr/JWwKwUWDGJ42dzccKiWJRXd+w61RwDEbSJAonqj
jFL+7HKY7SQu5gmiK11GcX3OqAMi7rlH4SMqq91e5+B/uVKMqOmCsFOGmG9cnPWJMrrbABiu+MuE
w00B2UpfdNaemhYwHK9rcP3IyqdavNANB0uyZ27iSU6xQArm0qekEyC3R8bu/vsKgw69W7tQdDfs
OwcrwK4XRWAzaucYpLFkjo61Uu7A+1QLawIpNg9ZsKUy+3qlMpEU0911uZAct4LAx032ezUxM3io
iZC/B/X5V33rlOPpY05gtEO4igaY4Temzj3upEtI415R0JfD/Ey5HD5puSMvaVTETFd4MbxbLe2R
dt/D0mdI4+OQDiuMbxYr3BALCd3jnlUIg5vHHwyS0iK6ew2099l7vpx4HhHOXAaAcL7b54pAI4i1
dn76n/w7q3Ae/Z0P3ZRBaQMOSGTJl2+K6EKC1Kz1qI1eersHziN5HcKbPkPNBesn9GmeuQnoJqfu
0gYHtSgcnBFf+2pe1WSiCJWQKcGkPmfjim/ZfCwPRTphBiKTpY+iWcjFvYy5NuCy9OKzk0K2uSUb
I9c9sfYTPPaqeHPUX3RkKXOcsboBFl3Chgz9MjQtDSwnWRDFzYcH3GKT7DXpENvVgYcZTXyGuX4I
he3h9vQw9/7uu0QtWhublIpXLlGQfxQXkEOs7dpSTv+X9AQ4vMaeIjhHFmcupHb7MI2lbbpDTlOV
xVDD1Jv59DBtoyRRX1C9Fh52Prina//bWyEIzDX1RpnngqIVFQmtGhyeM0uCg6qd0CtVi8TfwmCC
ampTs7GNeTaWrt4FRsUZuE1Nz9N9zBaXIrBOcxkjDkz5iiBzSE9Hv2jjrhbc4YRTiXF6TrndVxUT
rOyPUXRUMvC9HT/4qcD5slARtzut+pGTZ6Dp9j5X7Y9VdFq7be7hKaYbfflDeY2mrjfCadEVyAsA
3AeX+peFuuljQ0xgNzatMLLkF7j+CjqtBpxPiZ2uDfOLnmG5674nG5ssRNVPqxp2xO/t3OtCqaKI
31lYARQlx5UXUS0Lv8SIGJOWXWFRngk4a00U2dq5vDAdgsS9CwJgUTqTTmYggk9rVc7GVg76Whk8
PmkTPFjDAQ0P4CSAZiP11v/WtGI69ONa0G3ZrlktEaS011/JCdl4Inq3JdZ/apN3akYRbFmjWkA4
PwHqcsqDurCI9hRhCCNeP0StpY6n3ToqPxYVlpGkX2NxWMPn9tCPR+wi192OVYafyDbCoxfBDsl2
eNbvLdIzVV36kCTcwjPaXLxhEwGuh6o3Rs54a0vgBQQE2e/84VOV5FM/P+QdvP09R/6mxUVyAfvu
2YcdNZ0IudWScD/sC60qp6st0qps47DbpzDO5ntXt8KaXFqnS5Me0Dp9CizAcxmstr8du5Rv4Qlv
JmmoEkah1mf9maJTx5zuD/F7CTUty/KsqyuhCJHazBnNy1j3NKmjIwus9LxFXe3aT+Wvd5VXy9jZ
bxRAPtjb3aPJ4ep/GSvcBf6LD7XYQNujEThxjlSCLs180s7p+BBVQCs278Sdlzr6HbYet+APhgVl
I2R/tq/doAOjTePHQQ/Me1B4bkc+KbTEWYoZLxVlQGX6DMXcFoP7it0Il8FvcSQXMv3O/EfuKIYp
osENHVbQbWSnzFORPGCCdsDXrNUx5lco8x+OixY2gzUNrFL5YJ++43T9Q9jnjBIBopb0UR8mm309
vi/M/FXY+mOS4syXVnBT4p7ElKNY3auNK39c1UiWK446SAJKLfyxBoVjHqEVB0q2DiJHhW3uGN97
iu+Nrfqq7WsioClV3lcZsqyHaTU2bXHGptJaF1M0raH83MkD6IiiEBftQm1ziUKSa4swHtDxhyHk
3DTES3dwiWUqXoHgB/uawteF2OH+Oy0DNaeMkFnhhpQzauvlD8FqxJkXLy6qKRPYWyCwKse+DWtD
Jm3RSoUdQAuaUCTrN7bvephXguxmK0ZGrUYg8Z0XghUZleSuFwu6SqTOj6dk6IrtCvqgJhJ/5krW
zTtbJQ/Kta6Lykabc7ZkS6WTpUufgjwF8qgFmooC0oOUwUIUQQuJc4FnHGSs0GkSPcDTtlX9UDfM
12UXYpBJsz8thVF8oDz6CjBtyXvn8cnk59iLGz1Bn1R1WgkX2tWKlG1FmGtnoPTt3RoLBB1ANPYj
3w/ywJhgnw+02pDr/7nWizgyiENf0QhLtdmAU+jU5VsVDxlWcMbk+DztUU/xbSvoWaN7br1ygfWo
XYNsugMQINaoiN1fi+SkNaXdRIVEuNICqpefvseeBGZUN9I+0YrDbTOTaXV2Oe46ETNAwX+hM5Sl
edPX56TnMC+WyZniOynQw7sKlbQCgFDtjLwaYIcOLJ09sbQfeJuU7+XIWqrs50OCqng6pnmMcVEb
B8b9ENULIEaozENwpGFfuoehrp+aXlBlPtNZLRZUotPcl/2A62FaE1hKOqmgv3dVvlMZqtPpGHBX
ACPQC4P5PBzRXPEWeY72JTcqHxr8xi1UGQy3BqmtWb6zVP/lK0nB0VdAOCSoKDnDsJoRuGAofUVt
/f+HTSK5gkU9vvl1iWfdqg9teOBjzFQ+83Envqo1Lo8hSi/E6DL7Z8aHgGEgqR9b+oaaTug2CFHv
WFCw/+n1xLs/MirHFf4CPlEljHFnaRf8hUONIwVCiux5doPGoD2ZZg+0dSI56gj2R5ZEPWHouE0Z
F4sxlSQS/yaUb4msw5C0OuMaouKkeZO2tFDf7ud/9xWYzE0rUdqFYM7y88B0EcN5UwgkpKxfhZBw
DCj7250BjBeaF/Azc4BZhtVLdSuTAb8PBTvgURaKmxYn6Xkb+9sfaymg8vMR0LGM+l9fibkTm0qG
ygqf8ugZDIA/7fhR6vjFj4xmbUnx5hox+XBrgg+7C3CPjOk88Aq5HxV5OlRVgsFlNxZ/nNAUNKTZ
FFOSyX0tet+fayD9to5Wt/DU5iRTgH/H/v9MDUp/zYZRRteZr2PZuxwW1StUBXfvWIirXnvxFzv2
JaMl2zyZZYy4FsdESsByKbGWu3z2/k0NtPI6m6TLBXijqdpc3BQRR3hLFnAQwcSBoHn0rAbJlYLX
kfc3OXJ+J316MWuiHerjBz06C9y7XuFejSAmxeNqIfcNDXhCVsKcuvUTjwC2GrdJLjcI5UoBPEzW
dmk0Ui85VZXX8TPm/6C8LUUj1ITIAF0PhKbb92aY4ZR8vydJP44GLjqpfUnMM0OcBiI3BNwuKOUI
MLaFNoYHOB5RfW7S8NL/q+Ktxt+7y7MoVVdKQgFCkdpDWN8Oqeg1zO32yucoQTGYHXiqZJUxmapE
TilAIfYg9ffDJCKYARh5l2H/vu5MB0fBPKfeycpICr5yxtPk4dE3nKHl0xTw7Xa64MNNg7+f7C41
ZbD9d1k049HFQqulPv9j+waGpSu1xoWx8S98tLWRv2g7/oR01Qz8sjiixTtTmeMUa3MhMgORItIo
PNHRliiKZpGBw1DF0H0hkmqP8jZWHSnhEV5b4Ekd497VK9kgdQj0xVPkenMCa8Z61uyoH5AJFC2l
K5b+gWwCxNEAQ9iBYYfBMy0sHuPcAoRlYNV3KuP5dskQPqnrV53AeB/yG7Y7CDR0CGYHbmupj+CK
rwak60r9h6a09Q4HnJ0iV87YtyRnbFkiWK9LbXE93vVUU/rizYu8tsmAVYUJQr3z5oqVgXM3/ULy
exWutJyOXe+nCQJHLeWm10qhiCqswYamfbodfSA7OAUBNzuCVVrnNbLC9k02HYpCcXF28ij4fzRx
d+jvjoLuhEEotVkU8olTyViIbs/+cR35Wmm9KwYiVQyCL/hgxjufRiQlWPRHGGLILAuGdmpeP3ps
LZ9hfyrvwyD8ijzcx2X6G5ab45MYIyXgXyFySHwJP6lXQBS3b12yV5xiNwSfPdb/aje/khUOW2b4
fs1wGjC370f6YgCSrb312XAdlDFPhivcxyAMqd2Rjy9hMoPS0n4WvFCZCoGwnWfvGQb1wCZl54jT
MTp2HxgQiu7PKuPpq7YRWkYnsp6hkee4juiVgdUWNFlrj9LeGjy25XTUVigbAlRcwmNnw4yQi+Jg
rW2gBTFcj6uIrH0jXbZxC8DyQHH1E4cAPhDhHfneP2jZFCkDX1Hi9o0vf42SPTHt5ba5IVXfL9mW
/uvHWsIdUfBAYHgerHEgF1QgmzI/7VwUGzC8r5H8smoAe54M52w2sDhAggwuVSNP+x2Pq7jTNIYI
Z3yjew2NaZZu72xhfUCd2Vxpd6TD3l7shdYmJ4O221s61z+x0G+yaQg6nNn9MpqU+qZlzIxbNs+A
dEqVugTgjcgeh4EaOvPTMWnnQyeBL6sYDsaJ7/G/NHpi6E+qYttZVpZ2F3YaDM4a6Bv9f6521w1t
cBijMWJo+GmZD37NruV0FQZzWtk6uVTncs11Yb9WD9WFjfhBKCFpOLwT13NY3Paqrk2TLTNwXEDd
iCZPv1b1gcIfzPPdWkQpq33wRHs3JBVb/Y2HjGVBy8ejOP08I3YkAjUUngLtZ513Khv5S/B/3ub6
aLYRBU9KwoYSPj+J+mZVEdm9JjypZas28wt2YTp1O8hP3VlpHG/hNsE392xUyi/ZiYu4NB7YWwjm
P0KZcmjivQBfRWzH1LSg2YPUwKMqy+KpHsdCIIaVXSMDKz5J4k48dhUAzYM5l2OpvSqmTrpqHJ5Z
m7KUpb2I32XpGSKei0gxFsOkvDuwT0LHsfSrg9jrv+pfN1QkH/swpdEZLRbdEZoTKhbjHSatzvDA
yDl0JwfRtnTmhJvS9yPx8r6DAMVCuZ7lJqisLwX8zCzKMFQI21SIvv6pURlov33Yall7G6A/A///
roDSPQXQmPcg84BTO9SSqwHfdtnnZGNbm/VpE9j7b68BDmGEh0yYEwQxe2LyFL6KbxBZv6N4C2a8
jjHS26+eeLiTVXwVnJ9q/1LIrmZQmV0w4FZyDlSpp7BTxG1so9PAwVwJqMizxqrKDlx6D1dmf8sv
+Wu5wBiduGkpcex9ZnRPwxoU86EzM7LrtTTJvN9JgT0T7GMMIUx+Vfl1g6KmYRdrgkW20f0Ysg7A
l8N7PQtV1cI7SvZ1Q08vr7kyaEMejHdofWNRNFQx1oW+2Q04Be7bmD8o5n/IBzftvjmpemEmnCGf
WgY+q71Na8VOOVZ1phsychCLKn4JObPlThhUF1OsMoRApCMdhSdzq7sjK8fvRm8mo7fA/0lRU6fi
LLBGupziOXY4tLzgFjs4VCPdu/6f25p6MtQDLjElr3PzrPL66H8pD9yzarBRUoJlhMFpeMNoLtmh
LYFpBp6G1+F/0LLWqUgqic+YuDuY4mhAd4JILcTM0yxCjhCcWP2Pu7xfN+liUEOxKaVaeo7K4dSJ
wjtwKl9VNIVZn0EpuZdXFHx5ogB7QPp6GZFsmKKFDh5iNIseOeQ8LuMPqhCFnV5iikCg/KcAMNOx
ReIL/tXSe3j7FCAEZoIgkolmH7Kng0pAfYTdPsbxHhmjk7vcP8k9e8RjLR82WSIF2x2zGXZqXLxQ
c5nCy4Km0dccsCQ9va2sNTT6jJSKZ/NOT+yNuYPXU0DV0FThSPlRlJio26tnV4A4x8SCMcSDGgkh
QyUj+jpXvwzDEk42/NvR6k2rZkbQWcWhbd/4/LdbOnf7P/lV5b5f7OT9LHH1YDzzeTeyHGHIecU7
3sfRf8FeYrq3oZDjPNKVshwZIpoY0vxK6j1Mzia5KmPss0E7NQkhZ6p5ahEHgltYNn4paCgiAAzf
J04dD7RrFWTbng3TWCcqoKoTvn3hwNQsfxrKGlI54Av/zutaXSzL2FpnH86rpd/Bx303AYjFujMI
NKQjO/3QKt3p9shtqkbZl3ONQvm04TmbZ/Kbxakk1KI7R5S1f48QNKKnFI/nAfjFeYbQxs5cp15E
U6l7v9uPPXMSAQKnnM7WQ1qZlfgioOFCPNlZaOiIK++chRQL8/5bEUAjlw+MiLLrAFpFNIbQf08o
DVLPkW7wkhA+2wT7r/3+lwv35sLhfS4daywUHalZyB8I0U5RZLkS7Wy4vyNWlFy5yRXPiJQ55Wyz
SQcEhjBNEtdByDnogxSpFi5N+jFnkAdh0c0J+VB4x+8iDMrVcwHJjaoDXUCTdvoJevgUdqqVhzBe
PDwl8RAxH4DLgdVH3fCstxd7cpwHXP9+az+GL1FVsSJqyJfkSnn77xezKoW6eq8YVt7hJZhy22in
uBlZZKsqTPpzaYIuI5ohR5/bU2A1QPsIOQBCGss8iYqsr2EKqJNxAY+lth/Cg0m0HKUi1WTUsBUN
1cxNmy002wGwIUS7SMwy9TFuzhz5+BJa78OW3e+kr9DCWcttsDavvjzlFei6ktVRxPbwY8UxBwlN
gi3j76A1s3TkMatPSNewJJxNfVC8/WI6HzXsKb4yzwh01+ZcFP356F7t1GP54vy0voybqLtEG2IA
p+NAtT2PGnHzq4+hNQAUAcYtvu4L+V1dmx/ECeavT7MXWZIx950UIk8G1gtrc+Mdxr6rs4tKAV0c
LJkDE2eG87ypsmhkE6ODZGpcj5SI7mn56XeF3y9WIb61B19zfuFFZPEt8aeGigPaJ/CPx1gPj/tq
8cQgJuLNJF0aPZSnwY2/mw4mHvZPEJTBV8iPITbaN85+SagVPIm0jcSooDWhp9yePxF/z+w+Gb1l
QfTJU+0oI09ZKk/pIa+COgZ+kqc/QAbYwgWvXA5lNz40fTFyBe03HckD3+oBGvRqORYH7HcjawBg
PGynPl5Qm/qHnIrYlbz3FNkedrYCBRkg+CaNr3kpIQiRTC6WL2LaSHgu9pXT3oN9h9v/aPtUQWar
tSNSpRZ0jdrxLPy0MlA/PPgfKHI7tktXj+u9W6SvtuPjKcVU1T23M40oJjcoSfJ+x531ERnRZMHr
w0Iz8X4qOASsAom6OzQxeGMkibVUvwatXlYNNZGi2NAcEC2o9A3fY2Yemzt3+v2pYcuJC+uLW/xf
pj2twdRRuL807SEJ/AFZ1UrMI47xDAgQ8ep7qjms3lYvIXOVcKU6Ly/X4QXnQwMZHi3Xwn8/tDTO
/s4vFF+MvtixwQPEGoJvbH99zCfeUbo9ETWyQH9ZQv9bs8kOztpf2GfQ8IgkuCizQxGUJ+91+w45
bBOdCBQ/wEnEm/6B+GeQz0iOeoBSevaZbbr6Yf0NmrHw/yWug9+DHQ0c+2XcjjBJkdIxhCTZkJ1r
VATYeeaNow8OjM3YkljpXoHx4Ki68kkna/YaPnZoqCaV4+JQnQ0xifJAItEogIIpxPAA370vwplg
bY/18DzMYMfmikbRbrWDtvrZFXbol0HkId/SPOfpkqzZyedcRDmbwtg0w6Ie59Mclw2ps4qomTqj
EGqX0aLpYKwOOHCVh/UjyPv2lF0q54dPd+eqV0b1CSxD0mY7lqjVPUfsKj5EeCr33K+Af7iy60mx
qADKnWSDX/o+wxkaEcDAmVkL1y7JDNtnQJEwvk8tdhJHd00b9/VHDrh5XCiuos+ZYDbu3Jq3IN2U
H7OWpf9ISOMnCiSoagrZhiXzEwD7KxvJUENgGDpkcXBsYgmDvH/3elgIHdL95O2WBAuhIZR7tS/X
+U2pl40gUKGY+d970iOmfGvwNuOi70ufIQVhXfqpD9eCxcxAD7v03OzBsC0ynVx9LlArRlMEaeA3
kTiCV9e//sY9eUH8a/+5ncxcYQmButgbiJWlxTjpGpHTDmfnTqx094Nfz+LpfObpXjmilpXPXvBb
mbT9hkoiGAP6YOwsQsTXvyNVE3fIWFjuUrSoQu18IhhC/aTnWevNXNHUhG/zCIcvufqVhuAfPX66
Kl6pSF0v8woFqEjhnm+ZPazmkwhFVCMZWKQVHj5DL6xnfwXBKxrjO/yIXUDErbXo/GRUaOyXSV92
jdk52p/M6dfb3UWYy6h43wHDW4t7b9bFf3zm0RHwJ8REuk8s+b2V5rkZdhOrXhL1LuDzuvdC+Pl5
aHCkQBzRVF09AJPGYDs7IwzvjIxorozlpVrGw7yJ15b5sm0G1aPWUen3wBwLLZpOIIttJ5wleDQo
8hgGLMtIbJig7Rr+yYICPVjImgUwMh4FwcqHMhgDOGn4FcC4gw7KfaYwJ0T3FCKakE5qc5h1PZgU
C6VOobYQyMZu3J1poIYmZd/gnNINwnpYpaLZOqOT68ivfVhfkeJ9QNNC4XHUK5yKkhuT+5D/c6v+
Ex2iJDYlT0xXIq7lEUpsRIElg2s3odRgry9YOHkkXlJLAdUvXXrI3L45JimXz84cLRvR7LVZ6+Ww
EujiCcp5uymUJ6OtqIuzvHhM5yqhJx0tmnzgpzmZHB3LNF+XlQZAbCAcUlig+62/w5LwJWLDOGsh
6+UZhAOTjqbomVRUH+iCZCNqwJZW/shhVoZE7IVhU80In5bj9z77U5dYyQzs+Uoa//ECmXOBpQhd
ib7EaEMj/Tv1KJnqmDMhVkRldtJr1bR9aLlITVSd5yx7mX1YU1cO+QOYEIBIZZiJvE1gAP0jsUwI
tMiGml6gko5M5hXtaJGsICZ1Y+5MIth0ho2BMx/GGNMxGU+XDaVMW53lK/F7oH3Tcz2OP2kDztpm
Eu8HvLYcxhR7qYZsup4aAZcB3RPmk5OVIU+tXe3SWH369aE2xtBNSGf9EMR7m0nL0Yw6leT+yx4q
6TyTu5ktEBXYQIlgTsAUsZ0PGyFDnqR4JSD3ltJBC3Spp6t5Lt3i/3zXYw5xAn1llCpgmewOmMLd
DGG6BtHep9Yf7SbDw3s//POGcsdMArun2v2ePHIC+PDdp4jQTFTijnd8a2o6t56FCAqz2jc9eGFp
SXSBDctbK0vwgVYDnbZnI/7QcRGaLPWeSMmsB7AY3efnD3RgWuf5iFGSIz3MOzoC5cydDkVIocft
kU3YsT5UjK1NatZtjOawR8X8phvG0bHZ5m/LTZMuE/bZ17NOCJcTdz0QqmIz9ctL9JxodtlNulVC
FAh5N8EZ15lcs0d7WGKX7jZN+H0G+gDa+tX7u9jpp7Z7U3NpIaPFEpJrB1CKYravO1zVhfRZBSPF
OXOGCE68R1yU91aDYfz83EETE9oAYf5Zt421KN5ESfZAYLhtiJO1N5NbITFw3IGmP11FAj7AuweO
xtgxVSGZ87qnGMgt42OABmT9WvGFXYAW3im7Jg4x18X2K82EXQ+Dafc5CAVOVd3+O5TqW36n3D16
YKb+Y/E7bT7hfU17CNKPquvAS2qNgrHln1wp8u+Vt+Hqbl2LfiI1wqGV4uz++jQsskObEydQ2MxO
FifR9TjBbKLxTj1ZYKBY9W35Q/R6aQhw1xtd5kbp44umOSZ83IVQejEZir5VP80rB48eQou3rMvU
fJqo1+rf9bOAb4v5DIZNd3hVa0S6uFjcNyceXhKaGFNWrKpVIDqdXAWQVSsvGTJDx620EUva/+Li
JWtEens9zQnIFQJ5cRaXr27bj30dTf5p70fIFqUHdsZD5+I7nWHZI1jZ8vEimPFfFffP/EvVpcUy
QwYNA9iP6AySUiyhuUA2J3LaC85vLc8bfmd7usKjSu6sh5w5pEb/KDORzFM0S1u9JS3fCsDtfwKh
X28amE1NDsJGg5WAUP+KzM/11yTa0D4EynPCHDwUrg+H73EALfjKk0s3qPsfOJqP5CrshH96utjP
xySOr4lzi8GGBo/bUXD7L+LCJJVmHFjn9JBR20Q342rcqNubxx92kVY+Ux0r0Pg6knyCEe2Bteqx
yP2aILIH8xa0NOlrBobQfzAzWrGVF+yOPmDhqt4VbZyTOdKYlH+5HRD6dCAch9xngzacz3qsFKG/
T7mLNlmDWpWKhxI3TLUe+LSMFvcLfLiNSnE9ZaaRoZTEP/jHcDjgP1a+7ctRqLbJ47cpcCQTxiNE
aPyClxShTC31K1L5b91i0iYdU+qZBO48mXO0+LxzuuQOmXtTKgDnl6CWu/AgZpvsEsiGiIo+GU7t
jCy/qKZvYiCSz0HDI/thbuvYQVWCsnS5xuicTcbPRWeldHGfIBu9qGXtoTBAOa+x7fjRxtd5b5tA
RVm7lI05JE0b1nO0EqwyLt8w8XRrhq/1ogom0As1C/hPsog2PgkenaIjpylca6dhO29fqCKU5NXf
zV9OVvLh/XGRmO2zOLULTG3+xUnZowMFapgMirSJQOjqtSPbz7552Ea3+jX0P6032NbvzYCU5feB
5Wu5GaX1of+srFw3Csf7LHUvb0p2e3HfuPfY17wrIPUYqVMBUD9ZoHDcsHsVVis9XOSj473YMY3J
D8KNexjUdmb80fh25MFyEe43j52BzQRoV9iTaV9X/F7wdANlW6t38M7xKtAoBbVq0OrUBtk83TD3
eq826nyDNI0fu6Miv3PmkKvxPqhnKdhBf1Qv8ptTmmPwTDwch31w4fa3ScLJ8GJLQHpcfPzAMzos
s8CI+tbl8vQGQHjPac/g/PklvZs1pC9amRvp8wWtyFxNkANJ2hZAQIq+QgjSkjvhfZNAtqS/e7+A
gH0ZIwlqhYI+UhGVPKcHZq4u0ZVixVORPDui7/4BU8La6I2kOsJ34q8F0xDoB2cdx6VYwTq0hEDz
wjhIb+Eh3VvT+/MaoAgQe0RyAGkoiH4Z4sutVTPx2/2THIox/Mkq31kUOUWK794CsFExkOYM2BE3
s+DE4nLOpaEMr2rqyPUq0ZoXbdY5vpDKxa0O6JOYXYin34RTbbkCqRB118vi7NI7CZQ/m7WRrJvi
psB3ML0EXk9hGcVJNXJCo9tJ8OSbZpaqbYgQzdaULzcR2h2Owe/s1mYiLCF9QqGnWkjC0TU2+8TI
HmLaYgMvLzSypsloYDVsx1/LSHHiEDBYJGhgwKyiMoqxUwVe3BPq2sFU93ul4qR6S+1nK11/XsO7
QL+RAGOcA5Im7DhRlk63DV+vIKQJT/TD8KHrzAxPDmdn02fbLHs109ESGU3NWeCS9x4T6Np2CnEI
JNAln8sGL4m/4096m6ASWJSxPJ/TnRisLRlpr75p1kEjFp+7DreB2N3xuaSx413vSWDUUbsNNo87
jl/pxfXj1Nl/vNdiU7qXnM4+xNM6fru2D8/5U6eIPJoBFIv2+9ldrIpj+g+gS3ljI53EgTDlVXj1
vcV+gvlINCBA7Sh/EPtvQJjxRUqMR7LezM5Y34G7bTnQ89itIfCrVbcI4NdzFvtLsuoQ3jle78F9
yOGVDSn3AdysC0d/Bvuk8VtedPxntgoVNC7veL2b5tx18wF/qzf74M5EjQu2U5zJie546G1tA3v0
OHk3ly2GK622c8ARTg1QIn9J7xxYBOyptu2w+WGjmFz4gq4hoGT3dzGXsj+7l1SS7o/kEMdqszHE
zA8/o3CSkV2eTB8piXOeD3yUqnAmp53vyr1RcLLHXFkggfm2TpHq350XMDA7dWW1rtX3YynfUG3t
4lVwxklYlBIXV4qTU9OFO4Y+p8jRihy2ClmhF1/oafQg5c8C6FP6YsqrunsQfZHa9ReM7jzbTVET
RfgvTTDlvpZZYacG5TlqlBHA63+mkm5FjS6uF0CAwqkNPjrUB90bvQqRnbnEPzhoOcSC59dUXrda
0trz+/qHPkB9lZTDTV4g5qutUWMWxWIZwfnV9SDJ5wkiYJEyI5n2pm7EkkKx8BN4yDdDjihGO/e+
UdSxHTMatGB36kgzK4gOfc7OYurOJXrlaRXEz4r9iiJ3z+jsCiJojqAFghQc/FB8HjVmUZyX2m60
r9BN7KM2dm/OzY2NrCIuvYzwQwuaPDIXAJCsS4wZsOP3Jzngfow8/hhA5BwLf3qVabt5Qmh7xCBh
HBlZ3p6EcdGMskzZJmSrCOqAfj3lW0nd0IeH0GtePbSnJNunTHdQ7VKcNzhymypyQ1SkziW7JaOR
bU6z3Q0jLnsP2oOnb+91zhtk8aw4EE3uYo+GPjqKRKDmA1JRqz5bBAYnUUV/ZKx8G7erNVKmr0tb
n6kvWqrx2UVkOwmmBy35J54muzSeJCzs8TY1E03KUZ99YnCZ8md0pOX6Zug6S26fsW8oxztTUafj
uErZstyHjAAqt9WxIXJQXqMj6AxPEwKU34rHHI68ex4xscPAgkL8uOpRp64T8U991g7ngrM2Uti8
Cp+O3jAxb0LfAwavaE1tQQYUF1DoQgQhXdbT1d3jgk9MxTTSQCOvFrPd54nL9iQpciktmNk3RnfP
bjkQ0Oh26rIWDh/YiHShiwfam51WzxqrAanQYOafNptcgSx/8EzMrUxfQW0E7s8mlBlXzRgoLEkw
HVoCJ+O+xc8FUSDlBgimkcPcan5oUdx2kDG9ojti86tcHbh3lXRCK4Hv8Bjk5QwmuUt4PSz1Gm9d
Kg93NW9Sb3rpUKpwv7rEtEsjs+hnsPiJlwu0kEzvrgX9lvRJLszqZYqtU1E328FKtUChx2I40XIh
NIxVlX4yKj6/y33ggNRJ9mdqqOHIkJ7l1redbicAP3Uh/+gl+G390MSzNDzKq22BA0qUl7r2zmjh
X8Xv/ETJDqHwtalrujcR6br93WV4ZDLhAG4dTgYJ4Jqwm5vruwlPncd4VviZtxCu6C99CgLAbqjW
sScNgfclqpZtXvMDklApPclaVU/hEXYF31sOVdX3MPaPXCVdILRQwUeOiADmFJLNpAaeH10SdSLY
hJDsU/BCajUeZSjllENRc2lBL7ZM+ucXIXiSwK7Oh6F5Trbr/D5ZDwoLimTm5sCqsfKB63bEpjg+
3Ily522vKjV6EHth3j1WfoaGRWyzS0YrVbXv0ViuvCBtjQTAOlBGz/A0ujsl5WZ7odSP07PFnweN
JnOZkNvyhysdNziQRysCGFQ3EAqURXRoQFTfYLcNT9trMl6dPqdG0bsfO0Yo59l+ZOS4VGSDr/TK
zm93caIRdWgFAWOLEvZwqi8IMxeNvXtGGWKlzyXWJiqLRiaETj755T8KK2kqk5YDTpjy8uICW/Im
TbXYTgMqiUy5UGHWnGLQuRIaXk1jfcKg8Qra36DKnxHmbpM3D+PqyUmuIxy0Jijdvk1XfIZ1jE87
jvJsVxoRYlMZoNKHnpiWrqlagdnPBxobNeBi0Xi6bXOjBk0uUjVzkeJ8XezvvRkGuINBTkCxRUq0
QvM5dOg3YVnExu2SnwwQ6rtcxIJf5DersYDEvdH5dBv9TnAA5U0G8GgFULPb6i2ln83ojRYlvpVX
mh6kibSyh5IICXU4BDmOB7no2/sdk4LeMoe62wBRqypUa9y/XKRfvbkWu/TAfnwYlQtmxr03lv66
zteY1lJhzXyHy7nY9CZBJT1spFleu3LTNXHwHTj7nQCIqjakl8AC7k3waHgdpYVZ5JTsGHJ4wRwo
cPA6tLWOrfpbVcvPeL22Tl67Y3eC+WTRMP6T4rW16xgYH0YTEUuasVf5fuYK9cyMH0AJB+vZHhxN
bJGYItkO3lMjyNoyNvawynHaVLj9J3u8rXrYfGYOcRmLtweJNbkSlhjpim5ZfpoqJkQucGZWgRsP
xUKc9WAxBrnSohoIBgv612wOInP5MFXuSdDjggL328G8BUXnV2yuCh+58mYsu2uehgxB1u15SofZ
WcSCAgGzdZS+dWOPYZrRLeRRa7qPm2wpr3+HP5JeaPF5P1PZpVao9uibm+0e6wNOBvvUYjqf2//5
TbjEzIFWHOB7/ot9Gl1WJ0uSBpJG6pSxiBu8VBn0ojqqSsfeaJFH7fBuoG7K9Kt2+WC6FtuZjne/
U2+jkfxfUR+CxaeWwx6BD87jlMjcsdb7pv30KIiJ1Sy5VAdWDIvPXntJNDnGmjKueF1ZC0mAr47G
MB4RmKLs8DeGi0YHNrppgatry0Wuj8lvhwJgLFou9Yv4WagGbWga6pWwr3cGt0yeK0eDw/Bf6sj6
GTyYsKDRc/etVaRh1HsULvQ0hkO9R9ZV9VQ/isIdrmQBKr0ljEzqJ4BfeMWuvUKwRWlQK6JneY2D
0yQZUnAz1KkOi6SsyYv5f4R2hhfJX3jV6M2ih/xbcq2XoeCGgN0avWruBL7cvtmD6dNWUXBslUMX
PkPO3otZNeHxQ+/rfaCM1vjL1/zpVx9iQXJG9teSfxYtiw3lfomvYo5Th+XVuJMPZqPjzKNkvhWS
tHJBVyswN0rBpJJGNmvnfHQgGaUAJ0zFEyoOUPqRg+tJuu9gbCrBcNEY7NNKKu0gE8M+PkrNzw6d
GuaZpsHmCbUwixct/UA3YqIKO6M7OLBu2ABhSQDyBwzf4oybmTuNXK6ocRHNrWXlsEgpp0MyB/4M
KhyPj6uhxqZPvtnDvcpyamddVbpZmZioHkNqZri+xEXTFLKzbMQ71UJjO/cCXu01OxGaD9BlNbIe
BEqdSE6X2ZssTnScEl5L3G3rv57nJSXZSbRaECWOkrDQRkh55mRSFXwUmP1PGQosvayGpsx4wHcE
JZmg9bZyu8wPOzpDsX5bgqDL3jHSqBJZ7PPCXcicknFVrFJ5RqavqKNpXmNMf1yOdRyWMXaUXz80
ik0i7TAT4vZrLKtUpRuuAa0ilcVZVcU+ReG2KsCz60p/BdtOJ9fkaVuGN4O/OZk7POsDMbRiM2Qm
MaJv57asMjIZBO2oZDXT4r1Ck2IXG46p46xWdvuLx9mTZD45bcjH8O+NNZ5vne/F5w4+BFavNFgq
1sUWnnt2QfBEZr8yDH2SKobjm25yPK0cF+kxTBwFYBxKhMKIkZoXYmYFJuf5/tl5KmNdB2HvKsUc
Gbmobb5b6z7g5IZM73jwuD7cDQQmtuQfs6PEf2eYGuds+lkRKCLv3AiUIu7HU1/yBkhE7cDZ5C7z
dStdbfdiVv5VWwoM3Q05e75fI+AxWbqXssF1SpYnsg/umEghB8SSVT9LHw74ogFbtvxLqR49MP+B
JAei1Yp86eRjtiEf+oiLXDfU0ZBYwyfObZPlhyNjnRxemhR/u4RP+uVYhPPH9gY7e9mr5Bxkv1au
BlVhFRP3EnEb7Mn7wHq2TUasLKJWpiiIgSCk1LhZWeB28PHwpca37waYv2i+RNtt8YVF6HL+mHLX
e1IEtL6GC7rfnU89IHU9N4Y+1GzwgfLLnYZchzkC6lt7I8AqtVgT9F365ZuP6zb78qbQVtjLGfFT
N4GwQi5xOJjwJsmKOPUIDsvKBQA1pZXoRLJtdGZoWo42nh1i7amFUYnUguTmvySEu13NX9nWOgcP
rJrT+UrboyWOC/M3Cwx1wqWBweI0xqZPmZSSgM7RkjsGQ4JjjklSrv7e9sLwbaIzMfhgpoI9Q8ds
vUOqMjgpiUUkRDNR0Uqzv90PvpcMUHaECxBTJAttNDrBNuyF2smSOQh6TFricJmu+zf3uCaQU6BF
XjbO+gWqmgOK2oDOwssiO14d2d9TrbyOh3RCwc7pnhZ3X1aZHHDOpH9bf+WJM8k45nwCabKLQeEd
ZiUuN/aLFBqA0JqVjewnA1RF9tA51MoN/zymAKBRqzwZVezKGwgeKxktWPaITyl65p1qKwHX3Ue6
eHrGSbEP0+0Cg2F/VjKJXREtYDYaW0/kQNGkvvQdG+UkhNqZhEC+KJc8BtSCRnpfRTguxWkRfgKR
ge/87bJrwSywn0iVfX7+k2lO22IWMSYCGpSZOVd/HGMJ0VO7bRkPwWPAoU7crs+oErH18Ercymkk
BzIsyzc0qqEDuhH8cB40iSneM6rCwmkDLaoYGRAzbFiF9VyPRpH+ttYlnn9NZhcdMqKB8EYig6KP
myOeOPVYKGn4E5thSLpdJrOpYM4pxIyXRVxQx8UPI8DRTHbGr25q5bnfkUZzeZBjZfU3GRm2Vt7u
0HokmE8FNd9MDAa/ZV70xWB8WhD3lthO14Vh5EXCEqA6njT5tcqh3YzGjmG3+X2dSh3obd35y0Ug
5OwW8CWrynLejzej8zvwedEX3FkM4uISuUVrcfl5iZZIhGpBclDJu4Nvjm94Kek0Q+l2+0vxCfM7
6omQpkx2frU6xpXQV4UHLhR69vGjS0nrjiHKnAKZ55TuwnK3R9x6lqu4445uMcbTkshVtO1lwHPq
lbfRbUtaM+eebeyD6OreMC5Foluj42CecfMfwAPX3Kor/Om18BkvgYBHxhj3ci6isvDpUMXvVGnp
UiiFuIUtdN24JEJZ2Duz/LP9EI00fj63K3Q8imxKiDz+TU4rQ+4L5SK3/DTS9qpnT01/CfbeTnCu
KPcj8luUaOiYzZqtBEF7+QX6eAZoRDrSzauE2SY3iuxQ2zyDroKo7UT6mNXqoRpT+Vgc4mXeriPK
opEGNlzkpYBXIzlPMHlXNAcsXZ+/7+MqcyMSsTtvPJseo/Ep0Ue66wv83m/ztYG0M79BVA6Oj5Qg
WTh2lOB65D/5wju+puphUFLgBOAh2HHBfoHQJyzqMkqUPd4tBotOmEtB/4+Nn41+93ZD10cNJEpJ
RvMQuMYBFQvrpLVNNdXqhWrAmH/d4XqpK5JjexKY9wYGXRd2BJzHnYGjr2fnic6dyKjtlzwW1aR5
j94Nx/PNNS9RjShtT9eEoIr0eHmfsSsOSFIIlbSMjUfe4REfvtdZ+3QRsBxCrDy+JryJKTcqLclR
wueBPQZW4PgYLXGClY866N8K4FShSMcOmq7ne3OGUOWq00ehBv7MdJ2tEy5UedVN1J2dHm8aPVkl
FC7gZVUEXXV4GNU6bO1PMlkGMki3N4mErrtzD8Ov83wCTy5rX3NSShvFoLgeXpH7NCJMnu3mCIx8
9SWG6E+i7AHIMjf5c/LUZ5paMzsbmlWJpM4ZYYCEcBv2YorF9HeK4fOmtcVyWLfcXGlVhkB8vY1U
OPh6su9u0NGqcdxV5BprBqPOkchDFIY8H4Q0+3+uBoHZZ33nXGXQ1aTunxDXwm27Bwlf5MPKSwsX
FgyOB0t0jpFYWxgVX/VAfquoDP2N0SM+CGw6RCU00XIQdTh9YFII3lcgT4U+0mP/11vGRro93qP0
sD/s57v+4qSA5XyMu2AokZaXyDHoIubjSt/6xJepSjCE9odqOh8drsN9C9UdramelDuplChLUTZV
jyOXbXivwTSiPL9g1RuxnB1i2tOERNQQiYMUp+KkyDbSKFkMcvdvMmQ3zkMd+x1jY///dPsC5Pmf
pXIOhKAQauhEVL5bD5XZaoxwTfbFG6M2eDg07mhT7fD9xWDRQ2unsz5Q1bAFx3141SawCnNYBIs8
rixr7W5vR+uPPftEediOz+bbQ1nom4cUTLiG7HYyRq/Cxdwrv3SxBO6WBDenPM0eYtqk9LMxOA5y
QGezsj+EiBJfvPZpli0kgA1isWygwtxiY3FgMxZje2uNjg62NdzUbsTAp5Rs9kx4E1AUegjf61VH
4K7TdoUeuXkVoyYpcYnKEfJ9CCssGjDOWTqx7yxDG7UzA2WKMjxd8Hu/OqMHDcOOEuXNqTVxxSwZ
CYZCqEVeUk+iQ4SuqrAcZUJW4WsHYrkpGFPuUpDq+mgMDRLPQfEQvROX8iCYT251AuHCnLdEpK0b
WT6jtkIwZYsswx9Bc33NhO6i1cwXuBSPJDfn5kp+51e+BHmvsVf7Fo9IlPNYVcLoFY0x4ygZzbSx
5klzIW9QOL3gYN/RPxZB9klW6inhE9DshCht6SpJxNA+xM7WpUxRIyvz3f1lchZf5A0TWAfCcckn
65LEdsqnjJqN6eah7/SulNOgtEiXo1BSBuPYWsAsNJjRAAyy9TN1nRfYQiCI1WGL9a0VQA6X8k/h
IXoiad3gbQaXHEnFmynrTeZYOOa2zxz+OuKqgrRJC9USL5YFPYVQUOo5FGaY2b5oAKH96+kLRXU4
9tuYxZrYCwmw4anvR80t4H47NY1hDcQt+MxlQW3/kgDHLtxWm9azRtoCBOHXJF8jS1iVZT/R2ZGp
evUai175pDDQ4nDTpFhozLZQ1/rQvljzbXPcarTbukzCBBORgnTuYL+1NAsDNqhmA9dkZhLftjs5
rj57H7/+QVaesh/YKlNasS0M3jYL/FrMfSy8rXnQAJcprcH9F2w19sxcrSbxBWFXE4+BOBtL6qcs
a0R3FD8kLlWTRysH43RBy78ABliuuZ3RF71l7jn7zb+8E0Ueu7gAx5DAsX7KN2cE4x/C6sycTMXd
qj5aFQJfnIOUWppmWAB646Se2POLYkl9Xe4yO91pzAgwxGadxGfBs4Y/c0X6tLv4vLiTo4AB7YP8
2jCJ7L/loG7mPbeOpxPCNLGQDmlIREUgys6VipphOM2/3AJblVyBsG3IlibQQk9FDFgjod0NhhKc
t8zEBajRNh8ujVZWYN7yUsqmtZrBqwtPUwtd5W4hR9CyWzvgilgkl3kJgy7KuuUPx0hgckDrfuTp
efqO+T5X/E31EX9o6vO20DxIIgOP0UgSnzexRBkc2OlUnKpRnN2T+NBZfV+dDrSJAGxwwoscv7y8
VNyfqh52wKpNtVP2H0fYpPveM1Qfrw5okhLU7m0+EfiDfoBZKNV6x4umM+A7E7WNQFVFu3gahOhO
91S488ZwOZJHaBy3seSFMYdJr7Zd8+XxC+tMCe9aHOzWK/TQKM06mDxsHai9OgSIa0/P5wuqn/mL
tQ7BlMWZPruoNdp9/sRQNpCdV52v5XC0YwBO49qOe3ly13tOgenub0d9BFyOAnu3LqMjGWpNpQya
9T5e5ma3PmwfM61gCwFBcDHR66Q4MeezoT0iGyUGn9c+Ch4fsRiFPW3qh0jiUNK71836K1Pkrf2W
KeTXBeTFWD9JvLB9Juc0RrqXfMhsBXkFkVxMHibhr4dDvhorqJqTyUoh12SkTEjfRYjbcdDe+8Ve
5R4d1qsszJCb7PVFBpy+2oZki33kb/kx8OF/jjZ431pVwVQ4N3izC4bNLDfA4SXjArnf4nnCNLL2
5qjrCHrn1g5xuK3vu/Ps8E38q8DXXLoXfQX515Sc4pgpEJHnfdyV7thqQ878Mmfj+OfI2pZ+zlsH
ZnS51JXT8OrKrxFbLk82iEa7vhbmBj/PG2I6zlnBCdf5C66G9psvBhAnnjgWYuNfJMn754zjTr4A
pFatGuoKwwTjINy32dkBTNQrqkG3oE28m/ELn+vMgUOcn1XcFwBEWJQWhmZJJHfAD8dq+xlax1HX
KAkCL77DThN2QVsQTUYMWXYGB7wqleeRz8VUFT8PrjDHQHrgF9Pr5+CPcoed8SriQHHJI+5xVX3n
4fDDJL4qOnzfsEbpjj5Vn+OrcaxreivPOE7L7ctc+PuK8OYuPdHWw3tBjPpzsb2NAa1D1TTPxcw8
av4of+y01B0r6bJ5kerHBdnEjcExFA3Am4PxyVQQzzy7i3Ti68LudK5U+22ep5VrnBg3lDzH7udT
I9ohIRDsiT+nVR1Fdz80aUF1M6v++A+SGgg5aEZHJyMJguPSuNTFI6Fbb+spowObU7HFHgRhkcLZ
f9PQVuHNnJasSH4CcAGPyOE9aW8crn64NPqUFTBrgZRHvgaQ17X7WAVsTNOwnu8b7Rswrhs89fCV
VgVkOtI0vh8jL8+/0eDz6r8Mt74ek0NynY5OwWwdKxHKuypoqGPUOiYcqRB4OKpB15O3U7QhYldR
K3x6j2RjcSmBG97+D3lHgIa403fib4dSsPDNE2IMZ96f/NW0gqOnVia+p3STLT1OlRbCIm9BDPHg
8rdBDT5BKNWOvRU1GqZ1b3I9XI3+Qek1ip4mYxgvCgeAzJFMT0n2AeDvHJ5i/IxHp22FuDRyAxz+
lmzhVCQ53T9DEyfKCJgRf3YhjvZh0nPKOxf5QKtw58EUAtHjcIVX79DInfiLXrc1XPQ3od9RjzOW
63LjH27wGpSoWX198llurur7mLPfFLoxo/YfLWKGdCY7JHMnLkEvr10wlQK2Hqd3gH4yNjcCnLcZ
iuZPurURf23Y1zws6gN+1+SGiYPWrH2gv7X351fBxzVZM8+syJZXsnUXRBxBjju8Dr3myHYP0Blh
XMPs+9zy8Mc7SD5GCwdzj10yHAfkg43EIBTVJ9gHDgwOAFivzVH7GwlNztNMSkR/LdmwUwN/Ont2
L5onbWEeLKlqJ2scmzWWC9OgJ2DSEFY+2A9Te5rQCBMNQulf85OkAJ9yUZVoLzq5SsZeq0Lk3erc
KDXYwxt0OZeGAmgGUBWrmuahsFC0xhO+d8aA0o2BaMsl9kCLswSTS0dAfGFPrpOx5nrgAf1tkNEV
W0q4UzDSDLLo8SBl0V1VYrhnwFzscJ70YkEhaH4TXyfwhf8h5P2UtjmN9kkWn9LTnOTJ22/xxA2L
exdPZ29Q6+49CJE5D5jZkTv/Y//4XOT2h9a3wybWNXUXZI4k/Z3z4R1wOLPBnz7gFnw7I7KcS8Ff
747np8kpTW4IS6YYo2hci7vUGGxN6n6/zdoS0jb6NkmCqeC54uFASuah98zhPwfnSQyCDEXiACfe
+1yY1pw17FTcqDtwQbpxOZFdAMeN6SzmanJAvxzvfMVclRqRub7+2QaGSFVqc1G0KRXr9O1/skLp
93vBmcHbMtgTxx4fmMUv7pjVwF5cnQnmY3gRQ4gNQnmmn0fyd9zwnxohnVYBppk8QzJxjTa822Lg
AfkSpQEA1ZeWJ1HG2OHRtrdY2cV6uDOX8dGhQhHja8XnBbOHUwV0wgKTUvZ701KJcEigWqPMlYgC
zBDcw4wlp3J7DDybMP9tR6/ElcFIzrhr8VqaKWJYoHoQE0aEUCYj6uHxIowO4nbGhvAUPwVY81+E
8HwVMmFuIKwee4VshR0V4B20XyLll5prd1iYJsZ9EXCwc5JTNys4uoXwmFJdZ5HllTrHmETCv+UO
Fu+uzbNzG32dSGajhgYT4bnHzge+JLO37Or06C5mROBogu2NmdWk9yR/xC77RE+K0gtn/XEUk3Z4
mzRJ1bObjkHMLG6jpmdFyELKrXE0XmvdLhxJCUJJ44Qlg3TO39zIy8SSdhL7iq0Gc3aShoeTizHV
DZTJZYgAh2RqSqjZnmd1TGyS7KXCSN+2vng0pTNuEeaqoch9xza6BcagjW4+xUfA97C7DcXOobQB
MwHFJMkURyxKSb/qW3iyJhaHkTMFcGqulzaThXVyun+Z6izVb5wFjpjkTDZqvPDFRrNmaC32epTd
MQeeXi5cHhNzcjL9kY7kViHup0+9axW4q9Xyq61daB04mbAhzipeiHhMgKt+b41Pk+jOMg3CYI6h
J6rANCoCenCopZGTmcbwPVlt4NSw+di+ISujYSVgEHo/cr+7bMcS3MVNzBYBdRZp3Snoxey6BZMc
DEhoCjnl6JvHCa4K9X5czmrQcdYgoxknh6wqDginztKGZsjRIwfbf3jWWkVL/VeTi7hYCEG0xrsd
p/jY27t4+DVijpn2vdigzDouw/TVrMooli0fefTkiViX7DeqK7VvAL4gq4mYXYzPIKhgqoyiAKQK
gpFnz7zR6nJMtllf0Sz7Aukh8DqKqgMVNzClLbdXr5gA98PrBqxWxOxby96ZRakfBNsdzynjyCQz
AIdyyS9buj/h+4r+bWnYok2g0cZCQ1+yP+4zGFUZcMiOauJA6cQc3aGchnH2qd/1qaftZgxdmKOG
QekfEPyk1BpeFeH0/d/xrpapN0fUSWvAMislHjme9vAiwQmDFoEhZGnt8/pEGzprmppecReVUwl8
C07XyHm/GozOeVwac3pyKH4zwe9VNTd2YdlCA3RatLYwKiF5ANlyd1vCQ5M59dMdt46093QhFx9S
Y61qmbOSkKJkCHskZOKurftVDyhs0U+5xuyTvQKcGRNSj9DjKWEfU3WXd6EIyQ0HcnnR+2q7ofcK
M2fAOM0MKJNEIRcamTaLOqVll1wBuo1dy/LR8aezgE+oiBe0dwHCDUurdwZbbYCJ/odv64vqRwVp
+ma7hO/Xkp+38NdGk3Qq714KwRkQk2C/BrxF7oJxrKA7kIjcDf9glHvMOvoFnuSxnaI2bkS8dfC9
KTW08/hQNP6ZpJ59kUf4NIYvSsgxCMs2nVQJ0+X2dnaQce87G6myPnoy/BQLB8ya902igYPjyAuU
4Twwkegc7FNh1Z+OpEaMcRnWxM5vmZdgMRaLFPLzyRDXPN7+3uCnKfIAa//6FI2QlYlPDOBQS+L9
1H0YsIKIC0fqoI/Akd7zc2D8GS761AinWqVqyh0wD3qHQ6fe2a/SOCBROzVQPfIEpA06CZGeRgze
NJeKuuXUohTVZItjo2OHPfwTSkueyH2s3hxwjwYR5T1mMIZsbzqVoG6BN/mlg2II4PRVMyIa3Hwa
6sOeqrrWQ+/Sz2KgsyXJ8VorgF74t5Cfk4sN+kxSvRlH80j+mEICX5ijPgcdc7vmU2efwUntHFSs
ONhm+XB380IRuWZ6fJAnQwg3Fj8ZvZWr/qhC4f75U0ZStKXyY3laap1JwBZquu1J8om0u+JhWeWa
uls/XFneKgVER+npIuQkEVj9aQ6d1Fw2R5p5O0j9AGpacBEgdFCap3VJ5ngW99bHc/IvltF5kHFl
CP0bwRg/j4FRxS81stHAvmzDStwSJmH33Rp5lMriuc4/V3ugl9+E+6eV9gQjV1no4JB3Ps547/cw
ViwzhmEX/hzoiSBQy/M8LEh6Vi8NTiMRaT9OvVJr/It865elj1rUzNvJSzmoOwZh9X/S51jTiGWT
KkpjfYhxJd6G569ClzaB4UYNadMRjtBCSGHiOHRwZ3IU2b58BOQrW7/r5mjHN8d7uIP42e5Euola
t5h3aBOLJ6QVQu/8dyDZKYFoRYgbMi5EcJyME/tuhPP1BAMMRwQ7xt5E432PNrm2/ElYo0KrZkkW
f7gN5VaY8oHk4udNdoBp89MtUDl7rkNt0sPhqlVjpsn5CPIj+fbDEr23HLSFbGhCdla0AYNc+Aie
w16Wk+artlxS0FiZ3vyasZZwOtlLJTtvMRgpgM/BpzppU6wVIsKz+viowoyprOU17uIAUJkQ/e+T
Z/IPlliusddRUfVv8oE65pTqD3OPZJnUOLyIo8Jp3KphVDB5TX2L5sP0U8pK0iMhf+8fRAsCHEWQ
1+ML5AH9R4jZDxskMJkYJAODofC15tWE06KASIvNTRSti8pppfMOrzS8T93s7LSLpwgWlowpKSjb
J7eWMRNWO54t8HysRReiqtaNVO2t5ghjOZNrdAnhXQeVTx0TH1PS6OXSviamvwyoRKr2cdfe0eNP
UfaliPWtdsSFvE0sDN0w8/t0xfTW+kX7GD+H8njJxMpgHeu8vbOeHP1Kv3c7VJB15qmGI9msqOVC
5TtBRodRRjXtRD2DTfCSveDCCFr3PH34Zm0RaPX1MbWQS+/YHQCzLYWl02/qbQgpDqsldS8bVj5U
ohscupoKmrCvLIopRQ01KU0lD4dlOLMpU3Om0V91JQS5KLvdF4CkGbh34XyqgstHDZ55eLw3o/RJ
ilMRXiQNAYw+efw84JKhI6K+l1/BeyLmU/zR5d0BDLBYaKADvqWP8Hkwue49gAvoLIQcOzrClhdk
VkptslyP8Wy5lm7nfxkzx989A5ijT8E61SVxbvu8eGQRdC7ZAIbr61U4LenxB1qibbVvF5MKz5rP
tqgFmh1bS92shXOlfB/sfMAc11XyTlqD5ZBx3TbSw6DxnVuynxuzygk90fw5r4L3HFeAJQAtMj6g
zMvGzYnKJE8h72/DUm1sdQPu4JqrpxfE/TNBaSbnlTvVJ/TiFAS6soiAy5r6WE2uEG8wuzlDqJtU
hxY23VmNH326fYGomF70UBA0mzZHeSOf8lnjvzDM4sKN8wrtKEWciSVOAw7xRcbP7fEe91XcL6fH
3VNwROk2k19SZBUPdHivYMdzInuImKz+CFKQjudUPEl4qyrMMhzDU5HK2WTfiKNmwCyt9aT2GeQ/
uxFY6UKeXBE5r6tFjZ/i213j3wSxoTwONilYmuWWYrrlkVDKSkouQ+O0C8KpnSUc8NZijWwvlbuN
f6hzrPMYoz6pj7OCsyDi0RGSFU61MntwZD1vVcMzH54DLyuT7QsGKOVbJkZ0JsqJAInwoHweegb8
2qPUCJMNryihcVv1BZIyLTBwq5ZW+EGcd/gFJHFx9nUFqvE51CRQt+WExnviwPi4ME/ItLF5OS5O
P0gswIi1GdjWAd3lvZjEa03V9cVHn6RE8BSMbtTIaV2/ErzSdzkGdnb3t4Ht3Mf9+GXgAxBqLfSe
JWbIkpl4BqO6awIy5CUHSzkevvcJIWDPxfjVldnn/eKbcvEd2sklA4OSwVorrS67nLXAQGv1ahqK
DA3XuquPTFV9gAqnaqbfubNf7kd/U0Lq50ehs5ZzHEAYHL68HY0qEzqVEagYDmRbcAma+qgiKBfL
9FfR4tlOXLZ7RV77U1XbMfrcEBfeULBhs81VMbvcL6kopM++J1AVcDycb5hLuY9njBLXnZZxj/Hx
AL3IgLls5J4FcD56fwLL9/2TenkGKFyjN5UIru27OJ1H9OpYnSBsTSpJpc9zOBMLEkKtINVLQdZO
S1oxwRMro3YyVeOur+zXcym9ByF3BgKt5aYXwJwY+rvUk5O8exrA1WLNpj7m8JUIeouFm0ACAc0N
xmqrYoyiYqU/eHaNHyr216QSVGdKjoVlcNoz8LdkRbV+2Mvb3Lg/taV73+YcdDxgpIfq6Q8nunSl
sio6xctO+PdgQnt1QnIEl/1vX1MEywvmR+MGeyXlcNg8uzr3Kv8MNbERkX84/obNSj+cAVbRu1CU
wxFGuAkMRtcWw7ywnDlPPNaXcNxwD1x8yYt/x8DuMz4LCIcXQ5PYkn6CphCYiyPO287OLXwHyJWu
2VIDpsaL1rQQ6RuRZwUPDzS6mi6cNPKoZR+GRhjtARInJxx6qSyglS3Vxhh761AZ6cm8KBHlZYH8
XnBlLkNfj6v1QR01HII8Fgg2X8l0nlyIMrtmmu7io7IrawnYghmSkiyXjharemcXfZqn1nOkw2cm
kKaogr4MqsYKhhGulE/TD7BkDUhU6gJ42gRarX8CZo3kLfXy0FBsSP/gzocEdLqYKQNO18Qcnbmw
j9/LfgLdnotu6M70RqoFTFzvJJH4r5qiC6zP1guLzBL/QEVxBLUD7WPucIV1Yd4ERSrtQbfj6jC4
0XuRjN397ioH1nQI7oWrZ/saHvrCX0PNTM5NXJEfdIGC5vIsD5ySVoLOOx4T/UWGpycAC8OrQtl3
jIkP2iHbGO3o2NDm+dRrk31ALraPpdPbnccDP+FDckFus7aibVAcR7AVIaAAhPhnY4cR4Cx0sym8
Fz3uGNkBT1QpMSB6GyzavIBlhnDlej+V+NxbF6U7FzqvZN2eVa6YFNv0ZAYeD7fDS9zKl9QCGMfy
l0FZu7hHVo8YsMd/vAPBtUxrmv5/TT28iy2uDczh8Kcr9XfnOAHQU+xDI8LPMXnMmzrG5mLEzaNT
0/ZHWw3gqOOANrkuRyUof0Y2jkz07GmIi7ckt4u8icjLiTwCPrNHfUeDmuXKv4Kw/oA3zzWUkU76
6ZpzJ6vxa8QcTFUulLbKCBMPnEb252RZlfb+846AkomIzWV58YeQuq4eBQrlO8zO/8a7ruIlxb8j
fZ3MKFSvs6VaL/hCcdGXrkDcBtoGcCLSvu2QOOkz7boptKu8MrC0hftsx4sZ6pJLoj4QsCHXB0sR
nCdXdosZTvSN3rteb3/JXYzdMvQ9JFCqXIYqOMg0Zr0n3AcqMcfuSwYaRkv58jXRx/bMn66zqOYf
lG5oyTkwiInM5nx/QzhpuktSRmSdsRKyjWXA9KXb7GzlTLPKgt6lHIZnnrwUdSM+k9cTdE3xlviG
i0Wx+7g0wPzjlOPxOry9tLF/LIsn+ikDE0EYhO1+HrGpkd1s501uhwfVehejlehcLkEvBR96MXK7
A0LQzCGR5gDXl0ogFIuSGI0GopeR4IYjEoTgpd+t9iW7v8AghWeSKBd32S7ai1ML/289CfV6CFPd
dlfyqFpXYPGPrApus8SGK450ufxB1cFFTAK9NyX008enb4p+K80WxErIn8GMdqqIG419CPaDD6DS
j/b3F975bwW8K5ORfykgm8HKgBdPD7QTJrr128H20JiC23CowOn8N4HnCyRxUcwGl1VrX38Xo0+P
QRdSv7Swan83wTeDEte7S0PzhI9mL5n6bYxPOfNlakdndIaOvWWyqfcL1yr4wiKw3tnylol6FMml
+u8DJrvkKT3x98GMaCrPhS41zsk3jPL4aDCAaEoiJE1AHtjG5PRAtXLzwkMLeK2sBA3e4t2CAjSw
jmhdNcLSqNp8pYEBopd6DuZROp45mfDOIxAqzi5ywP/wHf8RjcnE5CiUQJICvWDHODIfR0WV8MH/
1u3gEoWEfuwI/mc+g+Mc7ZNaHQmu+Aj2ZUahnKXoigaPKdYo4qEBYqqp1CIHp1LbQZhkV0KiiaIO
ZeUhjbHIg6G1fIJvjYjYr9XAXpchXQB2DOd8XvMGWYKPzkvb0jz14sVKPMR/KE2AKb+rVyItFTns
6PTVMcl0qrgrQqLuB9Rr6md8s/Amkm7iBzmcOSO7+0rHgrlsaRnCq1ShVw0e1VNOiwUGjQvYxoOk
qAXg7BRAOWUShcMACsKTrDvDDRwP7vzM2G62KJam3iqgl3zaEwi5VYk2GPCNh4xYK/kQ93YE171q
CpDSt31nHf/OWQLpjk6Ju5FWwkQdCd3i6obFjANZr5z3SUxsAjaJGdpy1odFNEktRpvJvIyZvJxf
C6C7slzotJkmTi8wenb4ZG3dTxTkABXF+hhcSbck+BVVNxYE4+4jUFOhOgIbDHJZ+VI5bTlXinH+
9Zdv7pu+KitFIcISBB5rFQnkBg33ke8G7BPIpftM/Xy3mOYFr7HkZHmia61Qw6XhnwUIm6QN7Ee9
CamKpQpbOnAc5ifumQ5lngJ7wgwXBz9JWtiaAzt+J8rSSPA62EydnrGNyoppEUg8kNMYzpru5EyJ
PSZ0sfMvqojwn6pzeKk2KtCfmpP05bG0dT19uaz2T2JIx7eXFZPEvcqSILzzhg83pb6UWy25roxL
Y7dqqL2SSastLIOvAaiNBHX/ys6ewkSBQb60Z+4GvOfEcGz11J4nsEMFpzP3dfns2iWOI/ZeX74p
WXaYHBUZpeVA4/A5jd2xWvfPDi99ioD9BUjip7n8BcBhLxhlR4SagErJ2+ZRnHYQ/UMOrIO779Dj
6aPE065TMxLHxsg3MwfQTrNrgeEpZuSIjAcOQ2Ai5II+UpY0neb3hg+C/EAbPOTI6k7/FLZiZ6r2
c8+9b61d3bHPt97S6VRX8VN13RPuUxZEF1RlSlLnuUMPi7l9JlGoZnT1XF8uDmmijb4uZ8LlK8Up
OcmBJq1+XWPvu+djuKEVOq0l1rSEyYFFW8mp6CNfyZ0jAHeP8psBL1skogBzrcGJTVts31Hpk2GJ
KBtTiGTOfm2IMpBFueTLOKDTMsUyJh52wWMkcmQK8hpbGjBQ9UkirvTnXn1EjkJwMERQbgAfXoYv
9GH49HgLr8t+VRINZ0L3+JcaVcK6Bx4ypvt1af6AdMrsX8eetQ9zjScDLnH5GvXoJ/M1NIrDZoHo
45uRsH9fMlHWblR1tbEZQK1YgzH1T2SswLrySTXF55ZXPX6kkL6rwAXfMDsbPNJM7fepGWMmu8PG
yH8IZUE+TMVJgnjlpBc1JuWZkOLK7bsjQKwtbZL2aTfiuzWjLrynIODgxf/SKJstK+Rc7eAwcQCN
pg7yURAGZFc6802dGGcvud06+PE9+SajxqWHSRKJE84dRHwX6ztRk+/aLLzrzkpRbeI+aCN75smO
U1O5R/lvY3jpbjeitbPzrzy9cBt7WEAP3ukG5mG/CelMs3+X6338Nesq3QHZNVGLXhHS+PI+F8VP
Hyl7a6my22sohJUE4lQEbDKr6YfxMQpeu9txidYrUiW8KdsyzDGep8SBiu+Rl5oWBgQv+9O4RSKE
HGqDhmZZyY0yakxhhCvQUMzCeW1S+nSawM263dGMpJkoL9r/3MZJ22ssyTbZg6fH7Iz67BUfREux
N5BvdU79Cy4Z7CRH5X4FWVwoT0uEQkKq1iL83o/21n7PGDej81fD4550otHZygpskovus/EOZwIC
bpeGnSMDhkqcXTqX/s66UdyvkPK4ki52IoydcpeGQ3qGpLjfIaggDenKJtOcKq2xzOC8AEWwI9ix
AUvrfDnKWLTARTSF272DF6C/VhvloKnX3tOtFQH0ipxteRR/h9KlmU8bHOwEXnlGh1VFtrwp7bm0
p7za/NFYm1Sq/vsWFc5GDKS9ESjLuKsJywpAlWWNpOEjicFVMoPL0rMVPvm/kCgmSZNoAccKH5Oy
x4eFCbPqZbuwuvMBzWTyP7DMEso1hh2Dt5dn/rSh0ZdjV0nia7Q6WkfVI1WyE7wsNqI5FC3wy+0o
sHH6JTnU5ddIXVtAQoVP47XwZFsYIurjVsR865xxI+0LsVGWlJUKZezetEQlwKuaD7CVr1JOraEn
4iPve886HlEZJA5nwSKwBMnf4Fh09KhZq+tUWvt3k3dKDE5EF/hJGle8SpjGKHMMmfr669a1dwKN
T/xotDCbtQ33Ak1O1jybDaj4SKUWUlbzRQ3OD/LBYKta8KSmpQYGzEyrrwRFneNtqlnXu405DSOI
vbdp83MzCGYPxcjHdRCvdApEUoBryTkbOMHMnQGVUmD6NyM1P/vlgY9XfwqIO0xE56ZqsW+3FMNq
YWs8+EFWAZJErjbxba5TZxmfXUBX/bWcepzfAmilbhjQtPCpJ45ycME2P94rDNHmQj0Nwu+ApjfE
hBI1TKAxALVay7NTp4AgCZ2cBE36r0TqkpXZ1mL7iU5UiX0+0fMayA789jA3snXXdY3o1PiJJEGH
I9YiGzxCwP9ufRxJD/5pJ6zARW527ZToNu/z8KNdyFCXqhfGalneh6J5DEn+YPBLQx7rnkPvk9h6
zYJvn51XejwFVGvI9hTOu3QVWFyw2TRFvaXwWBeIFDsmjmLYlMIe/NOQTkKmx/O958+rcRAfUkA6
qWCV2ny/qqkfCQWAh4SJeU1oLTx01stdBXOZmRJLLtQd1UiGS5hYL68UFDBZ9YZx+3O9utEgq+Q8
nP5oGjw4ituecJM7IogHNdt/IQOlaHuK9Ss/ley6UJF4LJw8cvrUawP5lBfWTdLurEF82bF9VYIT
fcdnn6mCx6dsivF4xLgqQ5RrXn5plcbGPQHQvfYJ9ZosJBx3lwW280gSYEyjyCcJ6xX4PHVOGtpY
xJ66YfbftVwLpX0xk7OQPypLqL7tXyWC3zZuk5OOWfGTT6bBoEeLsJ0rjDuWVMCL2x43DYQr6Qsn
mgNpeck1wD2tKeJy8KLoiE33KKhi4oRJoNh4gsXO3jlFv8c6r3wA63Ns3QvvLRtGBon7VbmYeQ1J
Nu6thgNoM0a2YWP3WCbb+DKzHAc/j6f/+XnpTG0dVR9itEUV/OHV764DG4lfSgFHo8BgXpKmTYgy
TQ+JmgAwIn5Raz/4UkB0g9hlapM8DRIs6NO9SUcfBIt3fOfVQtfecXhEz0lWT5EnLqk/AbRs//kt
gY7quCjrsGAwpO+CxcmGS0XPRttB6v4R8CKFa8v2GuX3N5eyuGVx94u6t8NcwdARZ8TS5M+BJk7S
W0Bu5n/vdHdhbhEgIeGJd0YK2aBQuDWd89BhcGTHBF4QH3pC7U7sxl0IfL1nxw1id8hAOo3TtvqZ
cJPZfMdzzFWzWNW7st6cJnWUKXiE3Oara+7DmNLr7lCsNuBjSXvv2NkllJa14zxUVLszO3yRxmR9
mIQL1voWLrhnUXT2Eu/+m1DE5IAqMilymMinzEn9cjDKQ0q+Ce2f4awcHnlbz1t7XLBowdU9Dbii
33sx9YH6LIblhYTALKqunkhG4zsGRzV4onJsKqC5J54temmaIxNBftFnV8X93+1tZas6H7Utv+j2
+CypIDyjnpTXqhPTVObdmZPNT4ZlcbQ/eFBgPcU2XY4JoZxWWWxY5Wn77d9i2dSZswm1gzHej2Va
M9NERO077ziLFCOsknnKUV84fdMWnFEMBMFXIZRpMR0EpqMwqtM9K+xIO9RbaRq5c6UQo6JsMomQ
b5udn5W0+72LTndQF1HmXTYcaFbgbN7epEI6s/KR2V1Ep5nyLo3c9ypOWsh/ujy7kZaWepIcux2v
ydSYPYAn8WgEigZcx+zLnjvHVxzBr2tM8QWzJ1k8ud0dC9va7Q8VCFc3NNo0FkWNQ0oPt1ZJHIE+
dAlIVjd0C+/y0/N1WUWFB5XfggxZTzY7j0EKZIrb7VH6bY3Nb4Jnh6b+XdQn8YjMCEEF+g7POTrv
3AdeDprBjQ7/jjEf5U5Z0OgkUbkfyqIMP+51o8IITB8/HL7Musd5MHURgCT2HzDmT2xOXT6FlDIV
gcxCtEpiWZcIYs/KJG7b3wkWX2MjUWU/iMNzEieE8k30dWJAWr/c1ckrnzcQRtTpvA9ZkdYYwai8
1/q2IRcXvh5mz6z0DwZ/CSBgeU6QNWzrSm+mtIszTcMYj8KbuYal/0WSLvrj9fcplNqHa0wvg3dJ
h5jswz/bcrDLMw7PiQqVkHOh2FgwXWwwIClK71OHN9FjKPP/9diP7RaoWjgTEDzUjeelQOzS+BkH
BVPhuzi5s33RV5uweJRKrQ8sBWO9u1HR4bzhzR83J6UIrethgtGkSRQSVPJkaRvk+7W2WQ2jpxPI
JSw5pdnzT179CjpE8iivXg44EvEsLt8QKbETqu1jbCSvvm8pOmuF/QX/qcYo8IaFtbsuJfzVWYTU
QeaBvWP4+tnu2h9orXJajSNwCQKqv9qPOr7RFdRPVxPT/IcVcByEaGrKGgqYy5KeVIhnNU4RDc2b
0ls3hJfcch4chqx0dL0foiHvLWJ0QOSeIbpq8/3+w+4OelA0kU6LSzLTM3wirFa0bflGc2qX8VjD
lka4qUsD/El5tY+ACZrALjh/A20vDM4PYmJyTzpfxgkDTnzYOtBlo6Tk2lVhGCI2kjhfi+mtl8Pz
hS+KC7QwsdQKE/LN6PFIJPWfSwnlT7nx/o7BbHBZ86NgM3aRKqJJ7q/t9rP0Ee64Jg9pOp0pr5+L
46YRSmRDgLs3tayAIlj5F8oVqoEX967YIWpx98T5ZKNhNmvjxlNz1yJ/b4mIZt04cO0ZbjK98aVb
BONNd2rMYLWtSp8pUJNc/HTN2XI7G9JYTJB2CLVUX6Rvihf8Hr9I38yt06A0QZKRBTCQH2rgWWGH
4D9vpoORjrGBz5ks/RF9RZc2L/n5RH+OkfRn11WgY/36E80/c2qeGRgPnP/rzIj05kAYp/0Yp02O
QhfCejhE/wOtnR872ETUu67gVNnaY5cueJKJpvR8ztrobD7GL1vWx7wO8/allEpMzCyVowpQnof1
JYkoezSawkrqW0iQgpGtLD49Bg0UUomBrcuqXeZP67lWNUsnkscqHdwt9mmEMydOYhnnzpDj+czS
6ruogr7QZ0l5DASHm8tKJ6tN2XIu7uxAPqv27cui/BvlBZ0Rb9Gu670d/5WxN6M0O+4NQECvtv1p
IkV9/ddnCcaDCF4KwLSnWTRiB5BQtzVwBHVAJ+bOoP2mHGIzNFYqIkSuGOhR6dwWF+80GLLXlnDg
k2gDaKQjioSHjp7C6t5Fi2Yo0tbTQYVo5D64AX6bNksSKQutT/F8Qed3gmRW2JmbpbYoKNaQtHoq
KNiI2M1TCqfZcG/Tax6LQoky0QgPAeWYYQbNkb1uV7bQbpromGKMcDFv29q6cEO5eBBveL3ygw7T
SSEIsc/Ea7UG4V6yL+z5sD5NkIXoxk61jGJYhMfN5r4szTSuJN/B2Y3G9gc8frSw+LV15mvII6m7
PdcNhfsMOUr67AKKyyWQP62thjAQbMWJJFRdR+6iCKEagjlMcBbR6FdPI43vR9Nvwe/HtBIm18nw
AEW0IXDck2JHnwg4rIBVzR77+FsR9TixWgn4zEOsG5qJYzI5HcUjKvv7oPkidki/nUil59j1Stwv
SZeVLKoxzxyB3GaFksLc6AI0aAFeyrOgLtgDc+oA3tAtWEOgacu8/4o+/mYLg+5jCjcU8j2AhiB+
eQcpJ3M8iWKaq53jbp1JuRnXVuc28UokSdpt2eX/tz+cd1aYmC/5FVy2LI1b6d3k3gsNP5p9PFdd
Tp5eKozE5oQPCp77iq8Hwipp8deWN9g/1vm1UyV4ZH8BI5FSR26+I28LjkoDvFHJLHgRYnDhAN1k
lD4MyX8URhZyg8+/kAs8NN68m8/uM5XKcqH49AwFnmSr2+E40R7lGbnUNmKeLf5v7DMJ8ATRYTgS
gcVkMDVMVQHaaGcGW2+ytF45IvCbzmaisXdoee1MYIrl4+pt7pwt6X+vzjQZMyVbrIwW8WtI80PS
y1CPO+lBoQRuCMH+Nh3bQEuZVrBzRHJ0A7RNGz3vVXezCxbG8G3KyWsz0PifRswl3XuE2DV/sPh4
EzFcOZKLScMkw8eeA/rPUuCulPdHyRVX+I6UA00chc6l6EQBVzwFMpDRoLqh6EC0xPinngbb1yMV
giRM+G0WFowNxCjcgM+nUSgG3DNP+yzQ6nKNbywxb5VDaQJKyYDuV4cl37oqlF+ABWtPvNYMe4/v
gWE6GdO+KdSSc2VIb1pjuMimH6fQtD7vZMArrP5uhJXKWS1ClW6KUpFv+bANBPz6LZxP2E3/RfAP
8zrfd47Rk5cBZeHqEeUB2N4eVfGORIt0es4GxCBX0AR99Q3/BFb2Dk9BHlLsTPtLEcd3v2AZSc7Y
R3Sb5MZrfZWsZ9F/6gk/H4xpHWGF5Q9//fzDLExM87OvU6F1IqLai0O7CopQMChLvaTPQjNVdcfR
Sqp6mw1j0T+58Gtmrny0/r8ukvz6nvyPqupmRi4nn0iV8zAO84oWJs5qjWDyT1N+MgzcJg/U8Iej
omVEKRQ7KMiynlt+3RLo7Und7HXsC5NQoivxgLld/vVRZkrBx08Y7P6ur+zp/llCEFs4DPpC4oKD
XwtnJHH24JcbT2oFuAbnvitbj3h0jdGf1jlPF3hU5rkK1dTGInHLRuihzszq8nS6jWAifcs3HZ/C
yRwFdn1Jnq8eaO2eMXi9pTJg1iO9tbqbenoCFvwUm0wLnic2GgZq4siQ/7FStFI+UvuXdZEZxn+V
1mdeCkRO3HAAzwnXVi3Fx5THieoj6hGLx8EB+9B74BouzBTLaGtkz6TuMr/zGHzoog9EbmCjBIF6
WxinJzGKLX620ZtaRQFukkbGEOrF1B2OXKqhhmAsRaZsT0vWA2cpJQWmDTxTyoMRVDn+TInxwI6G
nxWDbWiXehiMSf4teus5xX6u3Gm24bnO+pB2xEbNupWsptjGKmvUFJ+qg1np0jw++QgJEKrdAWyi
yeOwdqTVZlsCoGMP1xJh5ldTy2cC3rA0V+g6UQnX2FGARdupF/2lnkShTT06Qx0d7lA5gtEluTqB
vlEKC3ipMoj1jihCzmlX3+AOhFvKB42B1QOZ8hM2ifEvOeVFRKCtgoPuyAXlyKDMB63XEGeQxo/N
FKOziT56N4H2RJOF7G789p//QFlyqLhZav5pxMjwXayY/yF9IjRhGozWcED2uzpEJA6XelSF1WfW
h6/hG6M4NrpxTPCnZpnaeDkWxhIzDyoK1wn3kiJmoSWtLnB4Z9blPMZ6m4FrcmCFcV7p5/vTnj+m
rxCV5OfbTnmwI5fI8rkPSopgrE3uAyr8yO1vuOYHXKaP66gkoNySIhnAtlEiU4GcXmTQ8dLf1Mhj
LVQWjbwI8WPHeCCVpF9jtSCslstVZYsK5njECiRnghaE+Jd/uHuzW9Imoz5nRgzDV7EUJmvY58q+
o3AP++IYo07SFcysZnPR9JLiQtX3EPPvEEq8kak/sPt9rRTtfmeJg4iE2R71pTIconC/N/+94qCy
5YJIAy4icWs/JP74D2pGIkbdeu2yQ/OV9ehipIHvrNCOknEJJMfIX74f+hyRV0xRULbvfx/Y5dZH
Wvg7danLSarowGJy1gFnLYXWYOme/+kHzrbVX9fjHxI2SAUq4rDBxqEOq4+WFb6nC+wF5SdQcltu
73+9a/bTDaM6shHY7t2aFBMiyl4GzDZrlIAJU8fbZwhdQmGL2jkqvT96SNLVBJjAbISiNLnXZ9Ki
wBaUOi2pHbP5S+s79vEtLJr9cGTcIb1n9C8Ml/ONFEKyIIRec4rqhWjLSgHPviqdQWmnh5WiGv4X
6QYBm76dzO6zik+DzZi1rejQW7xPGVSGs3ihnPGbP0jbx7l1OhOBTrJ0+JjRzeea/IMPbRWNj/WA
AdC6w3vNRBvkg4lCviTTdklE9eQbm+7xMJZ6o2A4owPSddabsfmUrgFIi0+HRlq1rfxi0ll6uRuS
Bi81/8KmlbD2bVqCutvjC1MI9plc8jv1dSMjDvrzXX/2RtY3jIt2MnvIWn9VKxvS8wnbAFUv377q
j/p6Bquma9Uo0aQzJu0bukmWA9o0ZI5dsp37rrT6NeNiQYMNi55V0R8cYn4wGmhyU+n6j6ZpHmyU
bA3YZ0VE6ZYbAu8HicTclC8cRNN6WbufPNeFVF5vGOHOZ0c6+lhbuoTyW5KMBS8WtSX2Gx1HtPNE
U/QHW78gs3EA0jwvLoccmXf9AcA+l3zfPFRDAh9MPkOQ18l/EzTIRRcxEnaItCdehm5v+ERMQ391
hDFk3nx4OSneyzwpogqP2sQOA4rOoIcX14PaTsbZaiPAZNpmUlTInUcGdaEX+3zUVhlvpXg6dm7X
d0bZlUX9DVRofTyUOMekBxt2QZlh2gmCewhefQ21zSWWo19dJEE2+4oSoDxbDZxpQgxrEB8T5XcJ
PByEJhIbj8GJx4kqRcDoME6IM45IjfaSOK3IoAtTbwhTbLv2Zawp1lOUPUcaltQH65kjHNWUKe+h
X16LHXPdnGSU7QPlaNlzUOk3/ljNkhoXp5q5THTc0igTBiv7GT/FI4cl9T0t/vhQQUknrpULChHS
Ke3QTuazmkGIbtBI594xQ+ZJQz4u59yam9gRlqndiaQod238DXnRJ/E4mqxFTj6Uj+msYCZImzVE
4HEllCvHlO3oNVK4Gog4gFElVmF9tbfMoQjn+ibtB2ain4nZfLLng8PR45KqEPdz7YAWFxiQ2I1q
pv3fLUDJ5lW0ajE72hDn7SB8Ms6aYCYUetxF+ezHfmeTVX0UGnCQbokqPo6T5OAeANzvaXiAjh53
MfkKy0DAG2soJfx9Ok/V4WDdOIT4EMitedtzWYxO61CzzFf+/mYcZsJIrYTH+vHYUp6p4I4HsaJ5
AsRt6Yar5fTk665W8EpXdup+HDGrSoi6c2jIVLYDNibBfu/OkRFLJoxS8LEj//AEuZo33vfQDZoN
5HnPXAnn3RgNZpoYLayUB96R7Q1uL9QyAdC3wLsAt4/sa9cHBPHbz2qAS4VNjbe3U2BIrs9+uhiq
kPWIRh30MQjs+tOKdkcSrPOKC2DDL2zt6+eOxop3V9kMoXO+Rl39UQPizx9nojm/h1ccN2Uy3KCN
PR99nxIhUsqiglOS5WWMr9Ekeudx6gqW/0DIexpR1UjasMX19uDehYNyiIoglHyDpN+03IMvKJaa
PD4oi9YB0xmS+Rg9eD2UfCiQSX7feZARheqy1acMZTd0lIRucKJ8tPoV0IN0gsbJdYIZzzXdoFPK
EEuAVP1IWcsUSS5A5xYl4cqc5OtqZPAEALNy+s/BkoE06SLi/JAzhbZ+VZDPdd+j0qwKXhJlCWCR
hDEuCWqBadEaRrqgBHmDLMfk3NNzJIQiEVfZ53CPLn8te9XU9iDf7aNCoFQQZlGg94eLMDAFBTMB
KWsFQrXy0In6HNLfDJUFVMMh1myp4DHBT7TuluewSkcE5LRAstwvKo0fMUX+WGPdtRYrB7MvUmTN
r1E6QKtaIV754BVSr45yIPCEpTqFdSkOJ9wmD6tzejmdYPeJ4P1V4Jww5id0tQidY7wueauXHz4P
NBIgY2JbhmrnzXdvVnXMqPgNRq5C2frZT4LHTEIoPw0NwKyPmsR2ic3uNA06Q2Q3wAg9AE1C4iO2
0Ol152jmuilIqdX3RArL0Zt95uH9Sqcc9l7Tf86DRSLPE4dguSlSSfiJYtnFG2pIn9v1evGM9M2N
lvAghaqS8GMHO8abjqttuyFg9Wbcep8PZvbBoRXyb81GBoI3yM0cww3gkS8tVdMKs8n1tLYCp3Co
K1eCtmdJDrU6x9QIgabBYNzh3M8C8mvhpy1PWCbNna+tbmeTtURjEHKKMwrpXbxqVaBwypNQzUlk
tqu68CLKoe6490HBsg6EhhmIGoo0caQ3WB3eilSSNH5v9zDZ5maVT6mHz8RW11UvO6A0tcwyjs8v
IyxqNAR3bY62/YH3W+63CxtwamZ2Ll0Y+GKfZHqObsWnwz59Ler5cx3GaYoUIBXA+WNPki6bseie
NRNA5TiV4Y+/7PQfomkiPJAPfpJ60UgYnYiIHm15oGHJ7+h116mwSFQQAXKwJMbv82sMQRM5wGBy
2I5cSKGRQDsEC3FAjO9OxOByzA7JhRVyZuzT2e2ByyWtELK4t/LgOJKAqbUu1mQTd5ZDtjHCdx9X
Xw7Xe2rxaw6oErGqZsK0NbRn9qLLvQXNP1mdgA0aIqMsiZ3u8vxrqnHZLP+o7ZCONuOG41C232LU
fayMfKgsIj8GLBJCQ9m5VvkAkVstYDEfiKs45kh8YybiceDNE2sTOGjlRrp4LnFQAqRi4idVSrgj
XrM5qYg0wLWsYGTZVebDPdMzXtdGmY3HqV81Ha+h7WIpSKk1pp/FE5/d2j2i4hnwJHsCD26iqXdG
9CKzgVwulycZMH5JcVxXpK7PqZXvtQc7uTtSGs2tRiIoNWjf/wAzWoU7hXPBLSWxHYrc6sqWCFHO
eXIeoQmvRves3d7yIpsjPYqb4g10juFdV0nBO5YRJAbmz0MdMucII5S/7alu4QBgHIUUZhMWpHkM
E6/o2lDuKsUMkOUecgU6arlQYMnPdpwPxApD13G7I8od3SvZM9RHdfuEG6Qae57mCpIgeVHW2/hu
nfjTVeN9mxVwTCwWxRGkqdA8oyFsmDHlZvW59uICFj8WGPNAIz5QH4PRn+F5DHkqlgAhCOgpxRPx
+r8QkmqGfsPR5FWtprfDhdEPefthOrH+ttjQXY9HsIi+T4OZ+EHMLX7lKBPP1TK5Thor1LElvVFO
zZ9u9ZtesXx6sYlgcRWGGOp/88WppEtwyGgBEYKFkkXWlgAr4P0OdMFYaz14y17QZeMsbeIOvE1/
MDDonp0xeF6BHKEyW5s7CVlpEmRB92p+zg9xhFXewi7LML0zQfWnAhDwvTN9jVxTrs5ks3qdw+qt
WOYoKp41YNaJtDPkSi++L7NvWOvowkmaMheSgku31qqrXXLSpJVlCI64LcKs21tkRTrQx/EI9OI0
PeETTkTKXw3wwC/sgfyHXy1BHBkq3V/s8wkr0DuMNFJdx0BjHri6jkcjCAJXI2AeoztFo52/yI5o
MjWh1jlEPbZRSLoCbIP/XsbTwasNg2Tsey3ip2YROHGhSd43cw9Kl5Rnof7SvAsPF+HnzgFFtDUK
Q4evbuaCLtMvnkgGEkMPcgkGuCrdOies2gGOr3aD/YJC5r/0Mt0d3vwk+tlV0kYztD2xR6vCV2wH
GDjJSAqQZjLmLVyHYZd8yCIN+gO97A9liaN7sqFWXGgh5xiZlOd0Jslrzz8N00RXXZSGHtIDd+ZS
da3qki+7prINIJJKZyk1jqqWkDOGvtlIUWyjnbjSLUgad8xZ5uDurmRWhglYojPd7efftvkBUbQY
fInBcmBBq8c3ldmUrrW1vJ8HtYenMO70S5QzkUjrWzz+CRWbWQwXeiD/yPqnD8iJ0dQqa9X7tA6v
Hu+vJja2ShxqPqPS/Lq+xylRLubd1iQrp3Gc2YMREoIL0Hrr9HpKbqtKhGzbnsqhKpg25B/PjKrg
MVg3nac6vxMv8jDKFXmahjqLCLlVTZNFeTwOK7c2KboLLKetkyPWimjkwH+zWzFWXv0BXim8tRL1
J/FQWT2JQKo6wjiEbqTuS522aa6xo69JufNYmwT+NPatc50dhVtW88BRaaX9CiFMvgUyvEYGzFOr
SqyMxojQHun/hxbKNGlOLEQvkjemfKMvFxaYiunlJewpvHU3SNtVkhjD99n5D+Emkd+027i9neas
kzSs2WhRk2luaYLXUpLP6vChWogYumGQxL2CFDRb4LovC1Jd+ZvSPr/RAN17+XWQxupK0kdy9buc
XpGzgZK31G77MRTuRIFBIwtdriKwEprfl/uhTnxSkzGECxO4s+aBkSz7Cjk5r6Gus3DmYW1qO+7v
URisB1GXJDGt1aSsRV9d1VdsrHkMGCN9ERLMffcp18xoIoK4Z0Jvcli7DD7ZQ1j0vzK0mY/q9xGC
5nno5ANr2QNrtBYd3A+9faoN8JRN5nRatN0i3Vi7qaycMUW+Q/GvkyAbSwwftzxXyh44DO1hhxD6
VLhZ2kqCG+r9LqBwl4g+JZNJ0Ivf0Tu9us6DjSoJyVsQ6MQr1RD3ygCrjXoNHjW7UiyrlEhbVngj
KJJi/2K71H0Xp7sokhlPH3socebbM/6/gOl338semXO5uR1VTcjw663v+aMfOlYQ3zd/EKEMkQNm
z2lcKrDVKL8OTwVevagvJUDhcj1FQGYgezQtwVXJi6ttoEm/6i8dxtG1pG46BVrg4IjIxrRsPY64
0ZtT1YpiPPVV84ZWvFRL/NNjkcJ7nmPckmRv3PY+lWQTgcOIwVS0sQGVfxZn0KzZBhg3fRaKhY59
84kMCdyTlh0fD80OFYgIvEgVWU2Y/KbRWvPydrT+iIpa/Vf7mrXcqIvCnComrYsLGG2XcRFrxufB
DvNTIPuQdxoFQ9K2OrDRykfr1R+4ZrTqRA7+WyurT87Sx6UdmxTJ4ztqhBRRm+OhtGCbD3adAn60
GvUAteymFmJfFzrmSUCY1ldyXkfJqgAzfJGhcguCVN3ssYj/EwwfaKr+6+HTAcO+O/g36VSfF8CB
sEr4EVB6cys5sJYCOeFMZx1hVWJqMuORKVjuypNMooJE2RG2gDs6TQ/DjE1VYnLHWbcKuJ96tkQi
IElhaVDSzjAq9871RY75B1kesP5GE6v7JUt+o3gpGmXqLSKPI/LtcDnt7GcF7PqtCT6jZ0/LtY42
aWIkbsxnf476gRE2XIIOdOAxraaG0BzXug9MlKv2PYIfTY/5KRVpjugp6vB+Kju3Tc01E5KO3F8x
sWUu6QUD5l8lqoILYWMzFie2NpZKCDnPtfiv5TwC056tL1EwkuTcSofmq8GJt8mxRwiPZf1p5H0L
ag3/DJINMaALdmznCvx3utGH/4sZuk2oC2lWHVAeWVCHfv0xwpLI1IFiTFhR8zdPRxGUmN2KHIhj
+rsxBiVpEcMpHTikQkvTqIkUeTNLqGh88Yoc3DRCi9XNtVPvTGCgNBd0jYYfeaG4MUnrBMWU5+UW
ttA/S/mTc7jxW74zXKNjsBJXFpMOjyUgKzjKNbqAlbiBjejuOuSls5roXu8yIfkMgMYwnWElr0jx
sECGaw4Y30jTAg/zQqZusX3KT+IafHm5eDMWAPNIYhcFccP3ewDeLzFWgUq43nggjU5adPj9kDJb
rXVGaRug073Z8Bmuiw36iDp2xBPlPhuB6dAY6Qam10rA9s3Putw2SEXnDUN7cw6mr5evcIyuzFzr
FNQEd/Z0Ip0WBMN3BlJYeh9nFWVjDGxGh2cfVzo6S2LoJHTQMPSXYtLzfEcpLVfL6mBARki2fV6a
gbig+SjQisgVfMB6nv6RUatiN548+bDl5NGf4X4MtIwxk+/Js38+QiFy5geu1slg7fWHJswh5wkW
O5G7n8m6i7RVpIZyHSI+t7p6fA64xVK3Awa9djyaPoFHxUAjeQUNbvuihUskRkAEzputZFQpsWIb
AUKEzZIYS8HP92LU8PpyYW1Z3K1GMv+WQy+tdl7F52kKWzXfirhp21WY4iycfYmHy83ijmV3dagM
O14hfUXRpeBk9pewST51BTvEnSoteztwBEczv9m6UmugEHbtDPlZVZR4t4Z287wSEUzPpMHlYzi3
/4UlltVq5fKm7ZNedr7/wFoUOmzBXNX7HjNIfqDBYw/HR27h4dyX0sYPhavx2I2Spzc/j5CEnHqP
6ySXJv2afLA3DhAVaCsj7Yxgj+YUKVTtKe8+SyxmfsMRqVd0Li3fohAegR3RevmiU8TIKOMFy/E/
Q9iX7508mVQOq7mg/XcJFibuxu8jQ5qwx9MT75YE3DmX1FY+LGx38BiTv5l9ZnohuXc4mU+Jl6WO
IQ87L38MuHsU75eNFgYhZhA3a3HMiRXjkxgzaajOGlNWSgcFnGYxhO0uT8HFewI/8upIOQ1Mf+5e
F2zO4FzfQT01ZPjExa75h/XWHEglU9Ha9QAdZvd06/MLKRj7VTVE5lzxJks+jmy70JY0fjlq3zpq
7cRR+8I8LuSso7nQb0ky1XlIS0A+InmIXmHVOCKHmGBojRVxtHD3XOG+OuqAne9OHgKto/Un2yPw
JJLwMdiOjbRLvU1Oez4lYsN+nOmRrDC2p1xIQ3KieA4WvHBUl3frqWvqVOszdwueztqB7Fh6S/1q
ZByZTwCVuFWJzxlMxGV1moob77yk5S1LqyNjfFvFnwLrBvqMmudDKYmHLvlpRs253/Dgp6H6DT7w
Tqiw1FzFWLjHYclqjnvY2IIh8qGuEngnWTJAsJV6HVoGHM5X2oaoenr3mLk26itKJqdff7Ts/MHv
n4lT7Yfretp1/Iy0qY7rum9ilw3qp+1U0OdKizkMnk7k1vGJ+clSpNJmuQqBVslwWmglYTNNR0wh
Iv2sOp6U7HG5wS+nyzinlknk3BH+SgydHK2awrsrlssgwk0fYEJMuYRRTajGx/IrLsw1XTpLXaXr
ah6Ejanx7TRaHHtsjmZ6FGoPG9E20DTvMwxAW2UHSJJCfXTivyvjziWAckNnuaFqG1o8xFWYD3ij
2YL5kpLtL2ILAuaKvR0vPvzD9//nq2jdc1NtC5Sn2jVG5RS/NrxZpJgDU9xl1+O7CXcn8S/uMiwy
kahGThIyl4ZXyQ6IjXdCVGQngrCneXihnJw0yBKAUndl5vEaIyu06FtGbh6bEMvgBQnPif9DcqSc
YdYAaEaDrU7STa6pKPnozgKVGQgueb2KIZFBgWTjsj449JkYcwrVlGiAw9AX2XGUg4J99ybEHSoj
xUZFLN7HZG4ZSDOoiTupQWwGmY6C7uaS0h6bwIE7muiJgBZLHxIyMs2GYQT6nnPVcWabnf+QOvEb
AIn+5l8rkqzYCZ9zuNgwr+p6SVJIskiRjjWaW8qPlUHBdT021VHEdaBWPQj64r6WZQNMkTpde/FH
8ItmBVlfQ33Ig9Dhue3uK10fR9aMDT0YHIaxtT2vzs9yZWKL10WfAGgadwU5Eb7jfxUwfeaBUDcz
pZSEtiDd/knXoUB7Ou7UoduUCCglC8OQUgywj6ATi4JhmIzrxncV44jHYPnWF4lvJnREWrIoQubv
pLvnxAgYuYc+dvf+val4ZgJJsMA4c74tvE7lwVU70MzFDSmuTlhhFOms8HRELX1bJ4XRr6O0Yhon
kOvI8kagzCh9+UJFnztF+vtZhHvFyh72x+PcSFY3L/lbxrOgD35F3JuXJjWwQs+18EZKtRjL5X1W
cWzchHoQkXUct9vNPS90Ki8xy7+IdGyA0qNl+iz9a6ILD9CYZcWrKP3Nz7F5gRGueH5lmkTSDwlm
QT8CCgMQeL/AWORb8rAIyijE4BOUCeFQM+k+cDMV1q7U8rTg+IQvBkwfKEiHYraWQHKnrnioPSHz
PuCw6pM1oM7QKwnLdACXw6hmIvaaz4T5svTliVTJjUOVZUR495+wc3Oj913s8mLqbPGXtoctfJqV
+iqhaMyc6kF9xRJ9prNPyIerlI6Dvn+//GyBcwVCqit5jeasMfpATKvSdkVl4zW4CekPadxu4yeo
07/xe77jWBdm79YtXMOGTFntbm4WxjTui6uH70gBXtHNq7yaAGXIJ2GMTFFkpohETCcZ9I/Jxxqt
Ga+IFI+rJpIuUQa6Wzc4Ro0v0h/f/jc0eq6aFZ3U+rJp0QNYxtdD7ismYTRXp0R0g8lhu8+bjPyA
6FMvqDd+j9nRx/A2vxhaPlpcZm7UiCPvS+X00TXO1gzENT1QtNiD9O92kUd3MCgjOiSEwNGDfoOb
T2ehDH0qV8FLbvHuXeGXhNHfQBHbLkDtf/xtyI5Gur9IL2kFDq90LNAzfhgsJXJ5EQbsbVfcoedP
bhmCzvK90oFnx7urZS+lSay9etO5WpOp4AkjFhRmv9e2vA6VlL7yQo+523CJ54X+UzmdQfafvrig
YVKcI/p2p5qm/sqLHpH6bhS5TUGcSrUFj2CKm2+fHNYJSAFemT16hA14xYWw+YOHLEpZJiaT4Tw6
xVVZ+SFBxT5ebami5Gc+gaJUNH0Q9PC0Svw/QgU4njJS7pNlI8flsM8OFRFp7UQ89ceSEnkz3V1r
rwMrohNI2zZV9yThXLRoBKGaEw7nbSjnFmm3k0N++42E1WZ17SAPPr++ANmEzQ42yGgsZnR+IuF8
SziF1z4JcOz9ikbY90WSvroGbDzcJCvIn6RvTOJB0WvOEkZg0gqc6FZ0wKjOTU279S6gytncwIc7
CusrvvxNDvJXAXqqZTDcpt+ZVe1K00wKDAzpmrkUmuGl201kfo6gmWcbfl3X59LLUEmfexSiJUCw
Ynk2cX9wBanUzhJ4EUzNLInbyBw1BA4OIw2TOsrmj9CUxFjL9WkycFgnItueOHGT256pd16288Tt
l6OrOxa+iLg4axRQu53INDH3MAyntc8vREGSrSf38PHVcHOjJWan4M1ELDJa54HIeeo72Gw9cmjs
NS6tGarMChR4k2s+nQagOtKNi7fuQL7YC5lksO9viL1wIdtwl4HOdYgrfVJEY5uvQ7hUtX9XiWoC
H9aRQghHsP7racoGKjEibsE6XX8rzqXnDa8+tjFqbxPemTe5Kax+8KdYY7ovic+6j77v1grK67qW
+bLdhSh88YQVPLbijMxAD2zKXhdS68bw+BBuHcbONNhO4ea6v6zhGxDsgmzKC6VjAqUKf7ZE0RG7
+FSYbP07AbYqBD1k/iigMxi2wksKW4VO66razvJdkD+ehr3Dnqz0l2dKv4dxyZzIjgT/NflhBYc0
kjcHrO6+SzPFszmQaW/zOB7TCjXmj9FMJd54fqFTnSzhUfITwiBsGCX2CL/JWPVz5R+rrG+dChM/
wyfaIJ5WT/2DaQnUvdJFNluobwqrkyPl0KfvRNtW8/Y/2vTyz5/3Bt0Y8AFL8FE2BIvEPS/vxZbT
92mNuxaU570CLeLB9YEA/vMrDfk/I5fZjzNUZWMwXDP/ohxHRVvhrXspWJ/a+qL16rc5DmWc0mvd
W5ZU3fB4zqWBbe3LgLqjmCHeL7MmX0RxzQOul7Wir2TMAZ9oSxSKzq+jh9xhL7RgDm5XrfssYREv
gaSVSIKfntoQv+e9HQtyWAkn2xRZ7h9nkKHjVgVKdn246M9mflsEi4V1UlfkEvQiTclOjgJsctLz
lWmfbq74jMv4FErWTZWTrgiH1Wwwxaasr7pWrMtAE96ZoftGXciDfjDmjEnRkDQnFn2LqzKpl18G
E4pIxp8s/XQsE2ue/sd31Z/7vTZm4+TZ/UdmNWJejLJO+IdyXhftB3eC+j2uMbQUmVcoAvwt9Tbj
uf160ABZ19u52bbHJrq0oW1LaG0W9iS3JvlvAgdtWfPize3osIlGq30TQ48+VfSW1Wd5UbV8L52K
VSLdfplILGCqbacXEhYbdNYCI0IPn9k71mb4uQL0hnYV1KuhRelU/fvmPO2M7/V5en7DkDsFbX6X
QzmOoKMfmihqS7gRDP4RcUw1PQs2ZMkdLj/Uhe4tq2wMninjgYuoZCX0PKOcjCf0uENvuFQgNLzz
YdnkeVKYgDaJd44g4MiJqX5ixY6F5m4hLST/zw92o900FWikR66zDn69urWMiJxdPCxvi3vNOGkp
PQN29ule9KGdJCCcGi4cYYoXp5wTipm1segK2ynGB2ey69LwZxmqpeOLoCEitwxYSDn0bj6RGPKv
nEztBZRqDOw1fxqySZs1u/lPtr26JRO/3mS4MHB61PHc5W3ZWxrDxsvfaMXa2p+/cvolHn0yGzFZ
Os6iEMeETW30skLliyM9FFRWW0AAa9itg93XPbY/dUSqMDEB3rrSlZGZcPYbOkMQt4HdaNrrP5u5
Zz3H06zJONVgzC6AqugVX6CIqm/IKQsdZGotCMvmbQusUqUXRLk1wZoFYhu1FvVu6/IxRb3nMXN2
jTt5Larw0643g/MsBta/LXpZiktaV5tMD+lm6U6joJlqe8btR5GdNUZts6GjfKkpj0AqAiDeP2M5
2XKUdOISWyiTc5xjIQE31lfx1MZXgsucwOLBH/QRejkZ3zNoDe5Qqqleicr7+fUa3dtNGeeHOBHV
2G0lLvMl0JM6cw2iubZzTuogr205J3AmzBSiteiR/I/VJ8GrXRpgR241wXZPfrCQ2BtBJV8fMcuO
8qGN3bjSj5SnJmrAW5YxlWakUypA5WH5miZfBBJ8hIoBGO1LCexpLyPKqwo6FjaCU4AkMt88kJWf
ODe+im3KovrZcokR1JNOh0V7C8OECwrtWTQKFqnUq+Y6//38tqHyotd/l/pvy/Y9Gp8LC6lKTdLH
j4/gOj9j9E9ykZsM3AnM6MXDWlXxSkj/YCea57/N0uvpsQAtKk0HWQQnNJaXKrCiEvR6jtlrfJDt
SssJm0ptsceta4nSXjfWi19rK7spnnOh4AnZI/50qgQcesij9cKy05hBFP3wML4afJ+JnN1zDVh+
iSSneA8blhR05y2w+uYeJaLmMVBNFtaOiZ7yxBKjpP6efqlWJXUxLGPD0Sjf2Z3CrJuVYT9+xsj5
At24hNO8XVsrrg2GJ2JYq9rOfreerHkmgtSrkOIN/KoSYs249ICjdKJHfrK1ZOtEulx6nZaLdu8E
PZ2mO7TWY6Lec5C0vUC/3Pb2lIYl2PwaYt463VKs+ixvDBzLYI2D29p7li+Zxy1SXbCqQQNbis4m
QZ5VM3MigOFi3nXkuF6TxITndGeBga6ErsxYOAN6sZoJp0vIhGMtOa/0VlIF0eEJLg/X4tn5ke3g
EI2DgQnWMl4z/Lno/D94kpESHFuBN/R4WMgIury38YzN5LLgwO1xWxiAIuO0jsj+a8sHhca2JtN9
TznFI5Res89XDA6VO5esnJJq7622BKE7gV0NGUHxx6QjRefFoiKVABw87WvsoIEqFQ+cXCo/EY9V
bsz7oALiKv0lQr8xVW4X0cPPzlV9h6Nx8Bd5ipKZHQK/si9/Ii29DqYeb/jvYNTpLhApKRuPdAty
7WO9jguER9z3P/PGCpXRIWLd1vKDXJ9vw+61mSFG+51iyW82zj+dFtRJSHPHRtggc0QPVl097HH4
ILVALS2czIMocoYUDJsjmTU10SkTdaR6v5mlFMx89sPymDF4aR++vScBfePe5ysk34/hNU67ZowW
9ELid8rJJp2rjsmmflxSxCa1GHCMH+Ln/PAH/bL3BvQLDXR3MRyy1pVDbM5/eK/RKEq2aF6ZkwmU
DBGTFTzTIOU1YXYXX8gbf2RLSDImVU0sgDKoNaeyeS0j3u6sZ1fBR23iyMXRV0zgTWxLb3BGc2c5
eD6zkVmpRq7HL6UR64ALCMaXeSlxyqA9qED/zQCrlRSBXO9ye3u5rB7LMU280yfH05WW1tQHR6rF
U9u0Hx74aQSAV4qmBM+rKmHKP+iMk6rczbNaaXO8CewCPH7HlaSf8xDuKKeZI+nJ7g05lv8ZQmKA
gMEQCvAyZCApk9ucHnbT26Vv++0SA+2JIJqOJToiMx8qEvgTjR8zB+cOlyy6dxavIxASUiGVKML3
9UXb7tDSEG97Thnjee9dgD8WT2L6ZnHLeVQlG7qeZN0JVA7C5EhlprGjfNkp7ojyiRPWUJJTZfXI
6qOm+pm+TWJeSCDmNW/ycRH5wrtIdmm4qFwpmV9Cl0FuUNN6TXnuOuF7BfCxMg9lBly+2VwMCFad
Xv3qNiGzOjhoHje877HpfPsifKrL/pWCkldykSVF45RH4Rq6sW1vBH2LK46TLpTfjqg9JDiAstyw
3cVU8rSdl3yfb42C6twdp8DtkJ14Zx1KMpX5nBkN6QYbz5RXjqlpTLzux28eG2QM/HpMgqvTk+bu
wM5R1LIBX6wl6BWSTvaNwfltlnewnnowyFpMl9lNM4bO5di23cUjUuKuchwgnq/E9GEtvI8E2Nki
PROIJTuTwX280BBX8k9Ft5jIK5/04b6Lqcd/Vb3Xmo0wqRWIulwnNXCyIhs7ut6km3y+aCqt7a/L
naCVJ/WqZeQg4sj+Y+iS18m8GsY/P+UcYSM5HH9bq7O/v93iCeJA8V3nfNBIrqdzY7A5a+UAfhaY
UhvtTNMRlvwX+T22EtvFVsQgpfh/SYe8VN2NDroauosO8Gj9FvnQnJZtUncI0KWTFHWteVreCrUg
kZ+0IDqvZ2mm2b5nLj16EcxP7f0K3lihGGiOV0KBwhFbmH6UapnBKhID2nKtZvP4d7yDwXGiU0nF
RtqPe5GwHerK9oS+Prc5v1AAClGDRffkMkKXol6MK27G0upZjBC77nl1ka2vV06Tk5OhdgDnPCiC
ozyI9VFZNBC/2F2LvPfG41G3AZb1Al1qKjnoszuaQWXZS5dfGAU2RTK4tbbiF3fCxWt5Pgel6c4r
2wt+c1573+Yef37Lai3JI0C7HNf9gWOXg9bKV6gzG5REJ8ia8TQxCMsOAeUgW5L6/0PmGA5wkNOk
PMsg2FsO+qCJnCdpyPttzqzyNP09awQbp8AZ5GHxN2wy6P8hC8wVhNQbKQL1KqECqomGv0IiJ5zT
VhKbkJDHRIWKdFYTgto17yg/DKYJDYLTJPgO727LhKl8msxZ51pJJcPOvhvdinUV2pPVDElmxbU6
qBZwAhywpufVUGmHrIqoeg4+ekt2AUfppFoXjPLI5WbxTmMS6mq7eEBOEQi0b4YX/LkiGKAqtGXJ
45plG+fALXeowWcTsRUtg17gI92jx5MFDF6IdBg/80ZsPl1r2ujE8eWWim15iJAd26bAcDGSQFDS
5TdZ77o4CIBvVzFgjrmdYuh5ifVXcrnFaxDlla+D+H0itpaRx5pM0DvJRGC5r6K+/0GjjGbD2oGh
rtJF5+22E090F62xaf7QG2GEwU6zfKUwGcWM+Nx0v+fIx+3f0H8A7c/Y/mcw2lmvRM3/xHbS+g2M
zlRNwDefqADpprURDW1N6P5Bi45YGqsmlYAvoNDIUwun9KbZekQkwXQJBrIXov8KeoQoAHrEdoNu
gNJSwxhPFm1XtSiU5CgKw23zbKaJDd89p0mxeTZ1dB0z5sKPZKvi4WKlpTgcqUVvLq3Z/Jb8HTMT
/o6EXrRo5mC7D36VHl9zUrHx091/GxgRAQgsXo0SL0WHRVRJZRbBnQIkFVvPjBQqwrnAwmnyDN91
Mt5+MfQKL9/prApmVvx7wKK/JlmIfU5YzCqZT5aE5bP8FQBqYKhb78yZ9aU5UcOLEnKBVyvcBGf9
ugkcbJiMzPnS1XiS3wwJ3VWjEjAOuh7HiH4YLSmVRbIEEDcZxU3YxdtAWjvhTAZW8kX0isPV3s7H
w2zBogF+zg3vpsjZeAiw4QVzFYSNaPIV2bzY2GecCNrIeVCZQFhLLdiunh6JPioiPpG8qk5GLwmN
tVwmA7cNV+PPcX4FJa/e0gO/IkBn6Jr1mMlMKnwK/xGhsl/lia5Q3cZJ2o3Hzizg8yiF94UVrXE1
pe50steXEdT/D26pmsAKzgxgJswEWUJWcdUhQSrArv2z7/AiNbKJA3TyTCAW/uyt9dCaYB/S7znr
waGBmpAHY7R5yen85L5qG+BymQvK+Uu/k0IktdA055BMtyHrWOVjebcOWpBgZw+HfqEeOaugBRGx
OGHiqkUwx6+kxXUuXhfOy3yL5SqWq1ryzu9jg4snf63J+nAPjoxDotLQhUGwHwGYi0Y3QoV9hDHA
L0M/do3vQUXpX9t1P2NqMxYJnKIfnHtIYTAwhg9sl4crWI4cs9xnYurnP1cc96LCKkOzCW8taijZ
NFbPDvxGgfBMu1kf+ZaKrMr7nZmHv4pg0z+Vx93sXoWD1HpGZzvJjEzJjNxMvLvMHFNVAo1qauM9
ipV5SCwvQAYreRO3LvW0qxY0+FDWwTjSO60rPzu3BsCT93q85/YEv8S1v9jL9deWmjLUNTy8bjwM
ZFGjXIaLZDvlVsuN8WNUbFU6NavtaXqfYuGvVtev+cW55Kz4VhT8etUNWKsu6uiUDEXrFZc8ymd/
C3yDZF5wmAHozlEqW1xPIbHXAwmoO+xHTRXYuONdfQ+QOkVJvG8Hbd39bU7XI8GAxafUuo4TRtC/
XZ1AB9BOe6XV8PvcyOy0OVwOd492Xs+k9LavvUxC224LX7fNsa5te4xdoafjCRQqLKJMG4h53cUU
NgP0uweU0+QxLLpcr38nNGZoVcql0mcSz+yVAQRbHSmwt8aEEbZgQktEDVUr9ebBzgActJ1izuEI
5kxcAWf1J2yT3vwuRvrA39RM31OernbNz+YrF2UP1HXpc35GqZ9K20fpaWpVQy9Dr4trQO/Tm44I
uUptUgqjSsJnCRFPGghAe/Z4CD+SdjM9rV55O4FgXHaPvU4We5IPxxVzgz045fCyidbRdqYeNIlh
FTnLI8M3q9Xvg/WNw6tpaHASM/lNLnCvUdYptsHEwuBDoc8LdTNEgzYd9CAZGvE4WeKPk3bIVJ3S
RQWVQG7alwzUHXiN14QATHSzXozp9TuCAUSFH0enlDm9Ubdxzga8vBRtaJo3S59mxETa6OoWQ8Au
YojD+ikgbM5OolO1At6BYgejAHT0onIve1cSkFTBMJNhAf0e6uXenp1+MO+X6rH2xh4bqr/HfB7q
IOLZ/UqQoeWHx8cdvRnD8FaCATJLF6E/R4sAXxRkar6AeUvaoh+bUUYDvbx3ud6BcueE0zBQ1ueI
6Vdu6V+jshqnt14nUTE7AHwJl2XfNiU+Rg5QOzCXGjeIP9I24TZCdElwtY7BvIqQ9OjgdahP5ysQ
2jBW7M1eWq981L8vY4WSTyD8HO6rVf8f7CBp9fUXYEljH014+i2CWGJc0JFx1A5w+2KK7IhUY1nq
hhveZXYJn5NZRaDhOCB2dlqqQcrdQsnZYrb0tcI+WSxEAgmP2w+w81DPY/DCmEaWrSk9SFFumKRt
QyY+hTBXwXQdlU4opfU5D3YZ134P98BGYhUk2Sm1kUWSowrIWu6yGNjH+2Al9ajFt+GCV9mSKjL0
6oF9dJftWzwy2h4GfXQv+6O5MQPQo026jETfmVIgzHVBJkuCIP498xWAYq+GjBqOFfM7XQPPr8xL
83U6EE+Hq6o1cZrPgrf1WF1xYpq+lv1GHGsDkBTsBPknLFgmfBRJ749Xq4Rva7TmEZAaPIOrRG3/
elJmT0Ty0MlK+oNyTSfUv8nUwoVqelmE5xFquQMTDIPOqE9of13qoYXlXVB6ML4AYPL2WBcFEZiH
j1sDK9fmS54abo/4+teTxP5KuTUExSg91zQ9in6ckw75l9Gce7NRhBYfHlTR7BeEmUb+PUnxv//m
2uKgbTnZ6aWRPaCqxKCOr17MJIVe5PgMznv29bALTUNZVaDzaHZW3yvnYMZKvEJH+nh/+6nCJyqi
uRVKS0EvvvisUxk9xgwqN1PcCii7AyrBzdrOUM0qVO0EBcrdMJtVR4nJB8Tx14KmvvNNRS2vslFs
EAuitvmCZkGnZ09s6h+U2rjp/qcZqTSyRIyW0B8hRh7tCFTiuAEd3DDJDozUq+HlcxNY1PtM7UWB
w/BHc8Fq9mLnSqRpeTMS3EmUErEYG5jYyDy/SIeLBp1jg0HxF/4ZByVjCEchEt0hysPWa9uoK1tn
Jpa0Dn4/TN+rNGO12CurwLeAYIY8JjMhFA30y65AXxPLPXtJZhPYA/c6U4M7xXyV8nalNmM8AhKS
X8H0GBaA3r9nqxzkuCLVxBUKefa808gFQVpKPyozAqK+u7tpJu6uQqZlRVIIjxZF3EuYP+733Uoy
fSqWfixnJYc35ymGjTp/bILsAOUdTlvlJaeC2rPHbg9cGEmcWH6jMoKAu364kDXFrN3dydzk8uw7
4I2D6Ugv3L0CFpgHHQSsR/6qB1WOUQAifEVMhy3tSRnurGcfBy4lRCGnZp8D0OyRGk55NcjEjS0E
9gaFB5bQYzdk1HwfpssIbdPD3suSDfhJOa2GxQ8vOkQ2dTjcN4bn/egUVvaW2kTrO1gtGkMgkHzP
LBpjwVC8kpQDu2gsvtLn/gYcf59AgsNw8+Np2/CS0WAWGTp3qJKCdm1gkaIvwFrNgjddYyYqvAsV
pwz1Cn/yJ77NUu+oJuQQfKygWuJa/WzlMY4tEGBsbQRYrkvzpLPGJs0dP8lI3Ec7PaO+1LkEOp6j
+JvjP0ohYgjZvEh6cSWTsnNyzlh5GAsmSWRlVzO6SHRf1rbw2285cNzX/Nz1Nkd+HYOJ7wXUKEBg
q+MBI3TPZE0++BXv/AAZ8pC+hqqRTebGHaBZ/tTvYfZmg4fnuvEvqysEs8ATPSiifGPeIv3v1Pyc
aL5Bj69LTdEaCrVfPP0QJ661ryAqD7lNhnUUsHFJSI1A5wnBKBIcG8piB11bal58MwgIyA9jiSTw
FWYC5/8VUWXE85FvDSDrAbDTlyvyG8RbMo5ql/yc8pPMjl9C2v9wlWp+jaK7wwdMh72Fc3OZKqPx
58d+gbaKca1o+Firi0u9r6smKhJ+Sv0RqoV9rW/A36/8b9iWat9LsrMo9hwQM7G5cKFScxfU7mte
LTMI2xk3d08Ae9gahoQJBsGFFi/AiuozSwIw6k62gSsuFE9B9RvCcHWoZ3b/NxQhaIKoXnNkJL6e
hoo+ozmYJhdXxzLYk0xCFFqFeb+C859lB3pePqaa8s14nLG/OWwmZrbx50RJRD1ywk5dXsDzrGJM
J4eQUyFWcTpRZt/2sdXj44zalIUgyzKJalpjFsQqZo+pcwC5Ed1ZQK8VQrXa+815vy42HH88vXU4
pBWdyo3EgZNLW5SNdeh8t33SgBVLY9yPrZBNerB29ESX+rdXMn9IIlKrcDrU8O5+wbW1YhxQ9XZI
WSxrBJSCv2zbYAeaLKriPuTLSNo5WpbfkaFmai7GsjPa1Rg4YKhFReiwJIQG8S2zKjxDO+xzSJMr
FkpJ2NVgAkcus0L5MjNDxfE9PtQhv6oS4v3UewAokFpGEUHm80PwY0OQN3VLyizCwnmZ/oF8mJ0J
m0KF50iMr+GNsgNgHhXzt3V8DvWj9puPCVnTvr8T5AksbX/8eDDLcEUshmrbRhi4PjqZIqjLqcxr
VXR7pASD87dP/7c5l28OHS0dyiR50u2jJAf8aRZilRygt11nqTFeg0darjHQHwtbC3Z3EVwcL+am
yQDXwiMMO3d7NwrKNmBitpPlxJjvWMxbNemfmaDU7E6/ZxUYlXZC+nSUbSZFZrU30S9PtxwBJQAm
D+BaQ6yPvMhfKpd0L7K6m7nk2xtLbpYbhl5WPyFeYJuo0F5A8ce8qaxod1YueiQH1e3zStrdwTDs
5qMsBOw9QgfAifEOoefaUmlpuO33YD5shIvlAiYK98AWWzicbbXcaYLzwDL8lxB6oAZV60mGNubX
RMHBOKXz+rMP1c1pj/pmg+ykJs76rmEUM+e975dm7h/1K23cLjB1tsxYnwvnDBiLlPNfPXUMaE2n
AzH4KycJ9gY/2aKUL/Biem8uhJD/CJJOr1OS3BKQSbBnCbKaheke7IALuRutZRvyvDceMHK+TOsn
i/ixxUG7I4W+aHdTDsptKILPXUSUJbrfiAntiWYxYw5/u2oknfJIP2TMmvbxJuOlAWbJiXawyMAi
lHFViiLGkuPYOShr6dewxBp78m7PkCY1J4sjQgWNpS7DcSddvT78ogkJyG3fQFXXhVFEAZIVxiyu
qJEq24K1/cthCpHi6kSaXf93Hrvoah2Ura3j/u+g360Xul7xGrIgC2IxNz33XTsiLz9ZAj1TmmjW
MKLiqEefFOT8xSUFzdrHlq0YOpel/NLyk84z0RX7EzJ32TZCxiwzUdCaQOtBk9p/WhEhe9CPaLH+
1CJN4L4tLYxnYUGxwp1h6YxISfnSprIqOn0xkXgb9FyZF+ax5fvMgm8iFkimj49N7tfVDvN96EP6
aSC1o4nqtx/OGJoiDGmU68gu3a2A8uYjLlvMt5kz77IpeBvpMx4KAqakjQgF9gqZ72lbGdjsVZzE
HgBWri1xyh5U1ppt5ramf9Sh+rDeohMmTMVOfEA1yexAKpzR3QepImU18r4IAmE0iE6oNBICh1az
bH7JD2bEyXEBBBCmqnijJLTGVAY224QXOHTyuMNFZC5YuRIPg9uqGE0j9KTfohttmQuO1qJ9l3iF
7lbBtTFL3huHH2ylpePCMpBWNQSr2Swncwh51gOcQGkO92q1E0iA2p3mVGBqktWMrRzJqG7vpXtE
hzAomOrSuBjy+8Suax8Ntw7ySMWdlc1YSndzNm8W9TKD1vXmzNHEgeHktg5pjy9kPqT8oSrks1aH
aIZ3wq6DbjGluMVDxXYssmIfaaS5x62ndlkDSvM5C/MOqKkLtd6bPk/18qQ1zt6CCJj5yhptjVLx
8RxwhtGY2ZVTwu4sV1DN7KyXJKwfNWWyxdH0dMCPCzaBL8As/jAsNRqR9DJooek8OhbjRxSuHRvN
YHGpfg6cKGQgtwm49U4dFbf+v+6N4G0WmFppu6JICjvR+s92s4JpL3qzV6iQrIaaQtgfWqG504Xt
G8Kz07uZYp2Uj8W0F6PtQ7dY8i6StZ7iUt6KuTT7mLRusy8tmLGhefA2x+HDus+5r6G3BBhuHPbJ
FlYkIin4LI0cRapwCpCzKT/DpxyxwZK9GfHHhpjQ3EBdblvtvBJ7Lp5k4/DgGy7xEk7pZ1MKZLtL
65ylNuRDSbWsHszI85VM7aGJ+vBDYxvj4tiN5L6VIKk61SH599R3q+8vzZZO4FlReMYvj5YBG7nk
BCM448kk3GHCKH25X1Zl8RoQdVqiB22fnVaAOQ9gVObgftH1T8ludlFLV4EoAg2gRVn8kT1LVpiN
XwEx2aDMJ0JjX0KNNWg/a50hYlJYfoj4I5QE35ED3cHxDlwTWWMxkwzzw+JWFfAbO4tUnI04ZttL
WLTv/yoHdac9VCfMRv7dJItTzZ/ybjQe/snvGIOBTgVVrpxn57ZK2RCVd3l26X4lHNDj/K1HmSD6
NSSjRyVK2HJ3yeUzDyE6jNropHFjIC5AdvI/j0LCjpRAZ7ZZsuADEvxmybdp9+3Bvg8oYhQxVygg
vUVCRh9QtBB4hi0mQehlfnRMQ0IvZDCqGRoKP2g/UcXT+Skpbsezzggvc5+Hsm59vzI3V/vcPacy
YveMEQDhsgVdkx2oIuuWUww0+XirsQpLxtaPxZKi7FJZbp52nzn2wLHolsyCmvy0MwYU9IGRnzv1
QLNNOUd5jeo9MFcnz8u/L7BvDBYq51/WIyrR+kkLyI9YVme1S4xmif7WHuYsZDAHL15qxXDnpdB/
PbdWlc5KCYrMV+Q0+MDsHZjnNo5DkGF99fF/5Lb3501NUcY8Om05gDpWJP/AQvpv0vkxULYtDChT
/Y5IP480Iaw/NwKveebw1sScGAtIyngErNtRRamS3CMCeccJejPA12Aa0bragtcsRPqzp3GwKmxt
6KwIe43pOonqATZlNbyphufj77pX68TyXQ2h8f0kwduI7wwjSooOJ+2O9vsqeJS6ZGF3zneMaCO0
ukGM28GInzJC4hfX6BAdjxYElE4L6JJfGVmbLXg5nZIrxAjdgZDxlSbKZbvX5/ROTrya82rUr89m
l7YQ79TiO3HQBTuX7TQDkiZrC88gC5sa7PLlWLv4Q5KlMPfFgQpCVeuLCvPr6rCNJLDsDjEUu/yQ
br0XBacXIiCmJneTZIwGxa2yBTGnhbFrnn3ZjTpqsaL2abo5MYIVKXjRc7WoeGvlT7o4gXTr2jDj
xxRX6WZ57o7RCm98cAzYdvTTIkbLSxizCSay5+qpbVs6NeMSdaourVE0MyBWWaaG1wfSCgDHrzqi
wFs7rAXKqx0tRbbVnpn2eu8wk5hUKEAWkTXHFelpqE1BozSiZyOsLIZkHq/brRKwLVwwTiy+eqCi
BOuxVHbYInM4qrEMv/E2Wcylm9vvoxrltZpiHzBZhNGm6B8MQyPYyaVonIzFHFeRyd7++hQBTWff
sJH85By4y7IVnHtWX5HYIvoQ6ftsGy15l+d/WTlgPzgpl9BYmVeGp8DAEIzFMGfmPfNf28SXMmpI
/9cMLXUlOP8ben/qcFg3SnBQLs7SL/4We+LOdzH6M9mwKi47g2M8awru3BQ0LIYlKEjWtj4v1HCn
5NfVEKfDXNX0eFL+M8s7+teXQU/LCJcSxOEeJMu2PBcu0uKaQJwRz4vy7O7vlljiDf9X1zFsS8I9
6K8Yn4cuxgeGOs9ocyNGtvzIZ3t85F9P3jLkrXYNIWvwtx2473D/6e3XakwvV/8LR8+QnNiFxv0q
Reh+Sgf6A6YRtTA4qxDccHQxqwvDn/4MeIrAPTpGpvYJXbKSc/2YIGsMSCab7NTY4LQvNNGiIjH/
BaSvBFmuL5xYdoa+9NxIHtr21MlNAeVV6ZWjMEDUBG3ngTI7VZa+nZ4CCoxSSx9KeAtpgeknZ7S6
rcolfmLuz8ciQTjW7cvt6wHCLc0yYvrsJllPxklhyuQeHWizMF9LOV6A3Juu40a4q7JEQQDlaQaM
3Ab64YuHIypylj73udjhEz2/8x1q2M3n3EkJ194hkuKEJEfj7hKboQODqDXbk5/2v+hnmkRQw9SF
UkuxFK2aNtZvmA4mgf8rx+W4BInHNNIL6KFDhB27B1mBg286dM+BaBPf2i9RgswS/pKwNu7OuTUz
SfXNnSbLe1DSn5RjngHgioxp+VDB0BwgicAsxsBO0iDkV1dULROPli0cGPc7Uf17PvP554Tx9sTq
oxqwarJ0HN/utl/hWQWMYHI/QWDpRB5Wi7xA/ISuF7utb0d+zzUx9cNLtIOLSoF2quvgjR6U2vXS
S72LAT1cyso+72k5D8fSVYV6VsJ2sdxUIxyffFxjoQr5FLb/BfyN02dx3u3H/59XWja1lG2i71ar
FdN4gQoJlA8MN+lHxu0KSMtbrq3cNDuGIH++YXACYRa1A3Scnq5E9yc8FQbQfsQB7qBYzhK6bVDz
lVeCozet1mkaT/R2rhISNGRnU/L2uK9DlhJkxQ/+OBAjeyo/B+V7IqUkHnb/L1aVwAcQGyk2BbtS
ZVUwoSyhGMzcd5E6OyAmbUUBFzFNfgunCURmeyW2MPomBSsYeVB8wA6PTJLcAEoXBADurHZNPNk8
9bUqO3QfRdt6mVnar6nK9tiELaSzcl1+KtOIMpQiFbmz56sup6y0FG/LwCPvxXPtKYxmvUZlK+Je
LCzHUJmYY/4UnXz1zvCLMGbZyE6h6oPlSUodKUBunHS0T+0+Dp9Fqn0OFf4u0ZM5/M1VapBqS9fX
HgMVLYPCnY7z+g0nY1gHsmG/3oyWFUsu0lufvopgiRlCG6GjF1gbAac9GE6hgvuuNWc6qlHMgYzH
IMcYhNjQn2ilCmeMZyUPy8A3Loid4A1GBQGlIUyG7HGXIBLgexRdikCiYzmdkfzxDecX0ArDdycB
yA9TuJbH7o/FUZEJLSjoG8QCLfdWh1soLzjvUyEBfjpeH9tWzdC/1BuTJert7DqYqhN/KtOFkamZ
8VHsOTj4vymndBjwP59Cy7xgclMAzQhkRqmbqKkW3by8gOQvv0bXy/n8Gtlo5fsT3M4anmi3ShUT
GbSnzGPI5OCbtMptst3YPI3wYt46jlUuXlMcbMGqX7b+Eh7IW+/fKzpdsX8Qo5Qs/N9yypqt+S4X
d4AXk/WCRcJY3CcnUOn73sq1HbWgQke5uM2gBS5niBjwfdHowN5Elcvo4ieNaV6/ylDaiqrUdu7J
OXvWWnYsMD8UrvnSDLydO316fHjSEeDbFQfhyxr5ahgk11H7fYIOe8pl26MPeBOE+385l6JMXYk3
EzKDBdM7Radjg6DEjjoGMHwQSdJBt+52Li/Z34oq83vrnh5Jl3Pd5Hp9ij8BhlARmgrSQ9oqTXlj
eI5W5oCYXuI0Xx8ksers7s4yfxycvcC6dhyHSM8erWuauROB2V2MXZVUIkIPxIShGEnVKTR14fnd
C+wrWUVQrFLQeP18vJIy8RJIvSoCY1MXtQnnlwARgTm56NomIvjHUDtCxt8KHmXZ/zJgPdtQehoL
67JOSrBtrEjAmoqQ46oBUTx1ZaF/NqLTLS2AObhj7SnJfzLA39pRV4L0aYyGezZ7oQFSEFvzyGWO
l8ku6fwGRWeigQqpLEriY8fD6VzIun0ntEP8Gzmu2vDajxrMUnGmIV3AjczTxj4yUbLvAkzWqyh9
3HHMvSVBZoWtfauoRKABr3hvLdf4dQdsiX2CJGnalC4xCvEQpgRKA1NdChJ7QGrV1RxDUAcEg3PS
YB79DjecYG33QOV8BREA6Mukw68QJbdTtY1dDcahioC88BkEywy11jfpPF6qruZ81xxAdRRVYWAt
VaDDATSzUYU6w0nrIVsR1yW3fF4eEHayg5MxYwvNT9gKcH0YsZ+9RUtXIKL4+SjmWP+OaNgZ/R7f
dDfQn1uQcgGNHVSacFxN+kTsy8qQR5WtCbyc5pGkXIG233T88iRNMmX5mVwD4pH+mCigZkJiThr+
kx/aShadzoxjuYg+c2VScH8X58KYE5I1alDvQJ4K8u5Fg77VzTPezXPPzsTauDyGjuJCqeMzi0H/
PnreQRdQp+i/GfPBD4vkjs4e1Tj1+J3g4jicT14zXBqToXwxTyEUFxxM/3juM8O5Gcdv5TronkTj
YizliybwNd4Gkk/Ohe5n5vh1GtLJ915IEBAs2FhQXrQhfiwptfwaAzf5mEMyr+QRVdvXDj/uEXKE
eJoLSi26TgkeuoZU8ImoDj7f0v4ZnRF2zp4NuoyqE8Qk71+xxRvSt9fOiqzn2oEcr6x56G3JLecT
wAW57ChjBT9rNgtm51DVVMN4J1WiYMc/3ySwbi/ohO0j08jvg///BqfAzzDzbN9/Nvy+mLc+24X4
AX+eszQNyX+ZmfIYS5LSoGPH7WvuboErPvqRcekXCGX+4mGBNuhwsDOpO9eREI9HGPzqB9BPYI90
qhI5lYrwjjV96ZuIVgb4wx2yBqHS6HbVCp1ObZsbuXnmFwaSMLCbX6SvXNtiIMzBq58bOzHAHQfA
HAyRjI23m1/xBoSo8m55v3jv2sngYFU+eadfG2lx1aJ7/3DBoVrnq/DV+qVLGj2+ZTpPkNAh8gym
yCIYC8x5yk9/8XivvTOZgnXmMfkK3FBI3d9vEeSJuqQ0MXU94XAYX719KIPlgbWg0Vhx46RIHeBK
9ATbo5ZaNE17z3fk9ybw1xxG7LeLuHc4nxo2630o38KemuwJASK7IZXyM5Alik1XyQi7DqcbVC1s
tTYRAblkWiaRZz2CFIYFHorDGnNuYPKwYdLcrl1xtRWcQuFoNf3VhNhKCFPMS2FwU8wlQkwIR0mH
GvPi2Ls9udm+TX8Y9RXrl69IlB2sBp2V6kbxu+vjwieJeMd+7u5XrOtiIS8933VwE2KFHDTlAPi5
q+yJ44X0iGAkx8Z9G2L2NH5+n4k+OPt00+M7DAS5f5DF5T14Cks2P6Y5niN1UbKZfLhPpDF2hRIQ
SaorejnoDp9ziokb77YiPQWOrMEMNf4P23nkluCFT9BPgSdXw5Gpz45AURwUSfLZfgf7CUPRViC9
jfu+ZZ7txaC5q+H+Qd31AfhgyglVFEcBotJVsNoDnZGOyebzMLMM24PA0/RKdHHwMCUxcAcNUrue
UryD3np8pneQS8Fiz/nFvsgq+cZXaNNbvrHtzHqyPsTEq1WEZL3I7rBZKG4cLpxoOTEvoEemSI0W
U+ZXsk7OZXcVWou/NBTpc4j60I1r3duAjAoyrYdFxEmqcI6PvAeNMFcve9gSdI1J0mBcYRt2pOFW
otDx4KI+/odXq5ynhjXLndZiwHs1KjBA7pNDG2CBJjNKTwhtq7TBGyYo+ETj3ZP+Ke+fB5IRfyAM
2HSEVBDX//e9CcuKku8KKNnJvGdZV0eoJkDExFk9g8O2j/dn7Bjgem/ycn8OZJn20mz8JifHA+p+
1BYg+NIJcZE9gqLi5kHVebrRIpZxWrWZ+yTvTsRRcUr6ad/9ECDJ7l0dMgiyu3UEFf/HtYTOK6Qr
iA5zK1RgKzOlnxb+yx4b6P7ibHkWM5NV/Xl+DIb73fE7yWP+9ujmqSRAExjKX36RmuxCa1fVcjHn
+V7fRcUYYTQ+81W4RoYCSSoXh5qkyClQz4/cr6SG4V4UHB4uhNxe7FXMkBmq8HBoPUrxQf3wj39i
mnWxifvwaJcQrBIQBMtBfNHyLjWnppGtfC6vTYQPtsNJ8/3ohnqgVmFMRB2AtxJcvVzJZ5P9VimE
GqW7Wl702h53is47+OxKLvFO31igmj3MpYOZkIV6KRAtBHOJJOpODrSgLuQISab/9XbEiryfDuBF
kZrS0OZtwE0/4k/Yoq8XxVA7dTDxX6RT1HuiKUaJDrwAKTsqiQmDed/Ua0NOVhrO4Zqlh+mMvf2g
4Bh9UMYIA21F1jCf7xsQRd+4lyasS7t+j8AxaHE2rIQZdh6Wb75hDN4iaRhzyZaPXtr1t+qZYp/g
6BKHKR2Tu0Y4J7F8AyBShoEsqvX51/ERb3OYtQizTwj4jEOoL4UZA2G484p8EpN3Ecquq1b//Z4w
hiNXg+ApZZxwBlLkfDvAruI/J4itoqir99UzArcuGfmg1IEUeM/ZazlYxWKvoL8U1ovRovrYftMw
sJZElEGi95PREN8XXpdZdg5NFXZYF/g+A615W6AmyjI7w9NBnvXED0JKdveVMJZIz90gfmq1F+HM
Kk/xTmWAsJ+J4YHab/1cVnx5bqLt0K7cCVgy1SbF7htU5FcVaD3Ny89/LIhJOdk354YemS6WmAds
LZPIosMrua/HLLvSt9xJ1lbq1Y4CnCFgjzZ4dR7+FXnZPY6YtG9mBIGuQqbBJ3SERXDEufFlSLyb
gvv5LKK4yRj3hB3yxHmZBcal97ldSfF7U3wtFBQwlFII43EFuEqeN5t5fnl/g3qE06r5JUm05Khl
+sWnUP4/O2Nb3/1UEYLiVvvJLOPwqOeWDikQ+PJ88cj84zO1dKCwl8fXa8H61PXX6R44EsBwPqJK
UGj8IWzMMw3jwRXnWdXv48vbavlWCErCsETVgZZGHSfFo/c3vjhbdBLNrjzKvxfm1f1E7289Xh19
5bzLXF1DiAJHM+c+1wo1j+PQ5bVPu3yKl0CxrB4fpdCanQD6nBYrbiBohdynnzKGEeUETJzLfUPW
4x0rzJE07BId1VIK7Y0yjirtIBgw0YC08X8sPvdjAjcucYWwpVgfMIrwBrYRd5Ta+XRXnXeG+HPd
9y7k8ClGlNaXV0CSDtLBt1XK1PMzTqxU7RCFr4nlzPgDTh/PEe3J2nxL0geBUZtQqIcmxRdj7rPc
T2NYhwcuAjQqauqc4YMbSwZ82UA0gcFhDSKWwJgUJfsbgjiUVdDYL+QUt9y5h7+8sZ9aMkyyyJEy
GW5Hq2SYqPKQyD0KTNBJRSwY/KeSM74RasbkqI6tGETMWBvyD3pM3YvxKp2KXI43FbwO3nJ1U1Zg
aVd0bU1KhyepOXX3tOd6RQmiQdxrdMrjnGCZm5ZaDMXicceN7JP6lQOTmNaYCSAMVLzehe3d3RuX
DAHAwLgcoFKH41EqJqloMWBY4JAqDyaw4Bfv8WGHGsXFYJ7DTdlSp5pGFl1g6LeH3MfEJkPrYzjO
AGodzfJsBIcHTYeMaTAU/afpwjx/TEwwuT1CKXAGx6fqYGGI/5BZ24fYiy0kjCq2rd1dKTbDH3hb
7mYNQVq5rxauszyLcJ/7HzTMPCQ4Ch2C/G9CNkEi9Lo+eLGOr0YclV35sQa78RKr3QUj0PTqIsNZ
70IBcwHqjS9ytR5I6o3X4/JT4FxT+ePpM+d+WdChmZXL59yRLzUG97zTZCLv7M6SxCBF271GyW3R
fblT45zC3yolh9QQygqa9Jy9gnE+FCCVpPhYW3FpDSpqz4jZI0hLeqjV68OnGldjq7yMd1uTEiMW
fOgU1Ha5l0IznnHIEuzBQdSTCHVfvrx3smiz0jFlsP53ucEunLjocC2oyelCwgCMSf/pxIMpTt11
LgUyic2fpDO/7vkDlD4w5OxpRJH1/MiQK2jbooqZnKv2XHDvGO0YU4vCHjq0skInXquzdyW/jIXF
vT8DVZKSv4VsteddwFu/kktM2wEzF/WNiO0Rslt54YGqB8jUjoqw4lzXkfSDqwnAFUd7HZkiRuN3
gbi0XrKpXxipM/WzWPJyJH8OVE134SLLQSjBVZhbwLfDMmddJI/BqeyVnZV88Qcn77K0sUvPn8dc
EwQ6JQSXFtkJ2uVQnCabnSt1vfcBRpmmQFgWa2YoqqK6lli2MneXhnfzFbNa8CAR5O4fFylhoC8H
NmSfEu4mQDuTr/A0uaA1JFDoEaLp510FLu0Ur30MT9GDCYn2MWrwTr4uj6/Ux4ZEPlAhWM2Nsy7L
/uHk3u4wUhHUd1ljt4SCZ42FuyLjNG3AjMdajRGNIq3He/+7x8WKRXTmz2AQaqilODz+2tB2e5ax
5gj/SQp03atzZiYZx5Tw04MWB+xMObiH5j1hNTr5DCyL9xyEGDe96cydifZEAlFFwEnQqrZjcPH6
ky4sM0b4ruqZpy+O8H4rYhuxZk0qLPsfzrT+gHmW12+dDda+gSk27npUso7iYgdT7/cdN0r3bKAZ
LcRppS7XwaYuZ3vRaDPLENEZHUZzXdHdVo7q2CNDD+N4LiTLcjSQRW5p5x5ibjENZhul8TsMq6+q
D3Y3JNPEWlTUhfFURU0NsUrrGqkPZzrvC0U+eMQYo2GfA4Lkvqek0wWF5bhZjKvtKOH+nfFBRTCY
4/s4wfnFo4JbNAG4+mP0A2hVgR0pc0gN5Jkxj6Dm+YNcU01s8XArl0nzViKpf84CxECzpy+ucN+z
aC/t3Ez1a7PxHWTPHjZG4rX068vNxgyQ+QF/oxncuOcTigGG74YRbK6bvQl+XzcTN1/yxRfp/WMe
6KIRq7cXRwGxsdGPiJCvjirBfkBD+XX6UsE0xzdA4rNk+CSIm0rx1Vj4V+zzXSelkiBTDTO6nzMx
HOD5a9wbubEvjz35FJUz7qwmn+wnlKY3IGC7tCA9iVb7aK2jRmH4/OTR1vFxVcw0SbCQz9ZBv1f0
wYiueoWlpEJGp33akPF9DaeU+XvYMxZ4LPSKnOSm4kca7amps2RJw5qcwAF8HYRuN0VrOnly3VSF
8U9KIFKYZ5K+RwXqkbSKjXlE+B0vOaTpMJPWOxZEML2AD67W6QtMT3k/4ILOadYvy/hIa2dO2abV
CsFHLEVoUt8yMAZOZcxKvBR0BVc1nUAR9jHXNxVcUWndG8UN5AuPYDW9PNh9yPOXYI+CLSfLJxNf
b0L2EK7lNnwFAxzLsCeGjJCkut+lEbUSKtMCBufodkzzxf1YzkoNP5t3fbMaFtCnf2bg6uddiI5n
H0nlugHFoftuWF+5oIM79f/RR+Qobz9/iUqF9SU1XKMI82RoPv5T+e+gZlag/tTapyDNYZVvtLlo
kxQs0NR3QOdsG8IWEpfFuG0ogyn8LgCOAlXbLpI8IUmX71sHwq0sSvfpHcm3CraXtGcAzdLG3NK2
2LR1PMn8D/O9+bwKM1/jYeWp7/OFb8DxvJvdQj3wEymrCz/rcm60WZgM+7aMrpVTCseiPwVROLSg
kU/G9CiAL3yxYHRgNiP0EeNbi+3It6wFnWzmC8yzQVRT26A5YiKCvHUJFbaMTA/znNJnnBQo/Wlp
ZCPZ1QE7aCZIXCGJUp97Q/L4Xwn00HHxq6DuT6XbR2SRN+XLkyBhXt0uh+VdYRFLOxE/XOWFchTj
i82GNFfC9wEKiLIde2YD9NFtAz753jprhl7GdXH2Zgwj7tvGmcq5ITNvI11P9z/MJGLT8zeWeIrF
OQxm9cD7yzV3s6GPgvXr0iW7HUbDd/jdYV+IMPdGgzsq+X25j7dNUvGz6Br/HYPW9Jtkbv/cYkfy
CEhaZTHGDaTEfCMh786T0PsJveU+sXXAhbpOufjJORW4KtzJkijPrDB3xHAC0YJM+MP4dA+/StOb
uksJ5fg8jBQwGqajHaMuoKCxbPdDwG/X9IoAtm76Gt2j+38q1XQ967KHsXo7Ngay6vhMrDRnRjnU
u0NbHSW71RsD/uTptu82NrVPT2W5DcosfCJrPdoC7t/L0Xue2A5SqI5IIPnijgbW6xKPF1m1uJ9O
yIglbmNdN5zvOWgMW1EkXCyyNmKvl5GzoJ1KyTKibZ+6x+DbHOlst1aUEiwtRte4p3IZSbamDim4
VjobP0WYfCmAPUg8WsG+KpfDsJwq/KlVkVJs0Yc0Y9rnyqa2fBw+VrVjdex/gP1J6Ya6vkzACJ5i
Xm+uMDK8Tz/HLryC+GQYQvVrDjjH7kDDrRZmS8Ts5fwh2RFgt8a6FSIQY14H2S5RjyCcy2O6f92i
N3IHzmr6bElo78rNZBeEC9KnE81nRfRY/c1AH2/4TyPJ66gMIFmI2PzG95ReHAfYEbfvO8d+fWZT
DmYzpq+1TQhQrdA75aC8FI1dNvoz7dC+qh3nRJp3u8Acih15dxO9egvrZfYu5VVIuX/eS+Thr8Oi
dyJXVf5vvQ1aHuga5BWB0bJnGEpaknmgrqjE/gkieijs9baqOMy9mj6LqBIf3TTs7nuAc+7TPvBc
IZns+bYgMcjfFLj+78cnN/SGrqjvXvz7KG/T26/5EXPoxBgCyFH+YFmBf04pTcdzASUojdhbEfK4
rF77BcdDEJ5yLgkaqdKyNiltQCNOPPqgYvoFTyboa54qTY3Q8lwS4W9vrWv9vykHs9kLIc/9Yv2o
PurNDLNpQeqmOyx2hzldkksd0ITrDGWfKgjV1+yYDFJexktIwTDEOUNF0OOpYemN3GyPNK05zZLb
HeU8/d7XUe31Fipg+3ReCuOuxXJvz58dcnQcmbBeHu4+Az26e6rSVPeomwt7fU4cvpxaLUxKteA9
enuvtITIywA2a/iM+U9JrhbNYnTVSARWf6n3e/DxhH4e71ehm/Kh97+4hiALoaYoaFmZkqh/e0jM
/G4ePnbQtggtI9TlLranTZ64/Cz5jFA10nLNTwwJ7jJrYPHp9Ncln9nxvVtm96DxzaobGtk3iWt0
kswyDtppjLIgJwuspHZbYvAKojv8gFuurKg/fVkHta/Ay9fryVJBoyv/24Fh9zDvQoT8cLLYAbDd
WxltRvCCPOly52caN3inP3JViOmRJv0Qtk0PDif5og2/JvDYsouoUAOfncLvgIcGf9Lte/aNxUyh
pxVlxrZQRlEmTe3wLfBS+R89SaSDucDo4AzZOeWPf9OJ5lzL0S6KFo/0vhBRdEVvb0UReAMJyLLY
SEIdThoMFC2s7juevW9o54bj1PaeJvPSITDj85CM14Ji/+NtbxFN2LBM2rcUQpXIRGYqgQ6AuNTG
Mj8RqNfNqT4/PeelK/hOSgCHcTwJzNsw5hkrKveZA6KqJTHaCb7+VHWQbWKHvz0J2kvt6J4i0U+a
yLZCijXmHFDypftZYSCiMSN1EEmrv/Qz3t3a5MM2kVVbYot7YzoTPkoE6ut77V8HiGKh3McGuarU
uFBJK7cQS2u51zXI4Qoqwb7Ua5fQYpIAXVy6IEgYxCV/qe8Ni61Ub8mQftH/Kwozg00LDBf8z151
pbftaZxj7T/0vj+JXfAfOk9o/8mZ4iUIBJPoGvtJ8tgbuKshHBHKq7pyhmjvAbxUlhCz7W3H+AMB
EutqF3JgQKOnA6uvrtjWTaqI+GiYRBU7yOV/7OMBnEfAF+uFGhcxQv1OgJuN/PQYj5spFZ/h/8BD
3vPyYSShyfBVxvqYSLIRVZPdXGr0rCRLMQFJkiSGmwPE8emPuKcvIk+0cn5LDqmkHZ2/kuHmvcoW
1LTJuV7hVkUlBSdh9RCazJB8K9Yp7ewg5X66/+K45qrXxL2gTQWfSmrugcs+TyrgS6VNuqCW5uxA
RxxIvBbbld3+P6uNCQE73y7r3DN2XfJQMucxO2wo0Zi2O4ShkNKcy115LnMe2X1VF1zACkrpUqj0
K5GolkrHOnU262B5C3Y7fKzbe4wpfpeyYS3pp3NpEV2XLvjxpqU5OIprU0lJ33GQssJ7KidelMVL
c8VdrnJROJn4ApKF1abQjkgWj7sbrlA4WCsSyNDInTCUfISiYdgk/9YaZ71tDMMLqsRenO3CcHAp
YIHPxLHkU15pipbeXqGuzLoTQdWFwYsxzDpUAJMi0AJM6107Tb0m3jSoMGceaRgaVB1qoJ78hJPw
eM1CnOtUpyrU8I8qSNMKmpCjCn67eDhMkZdtgOZPuSM65/yq9G3pzcInK9i7IIYC2DGKvBq/bFwY
ahcFv/6JK1i6iVsCfhg7y0y6ZtwBSpd8JEaex47NwmNKTyp21xL1yM0JA6jivK5JY80jGF/+Lhgb
R29Dm3/wcrMCWRG8bcRJuQT0bLGxYLmYO4hevmeF1w8DkNExwFCpR3/EynIdsbN1B7b6tbfiSy86
8LFXw8csmPwIvyjwYpfPzMKYaijyFZI6ybYTve/gT1YtvUyLorZo9T2mHG+lH82ysSiDd1EO0vIA
sN3GH9+Bzn8PhOOi73xMHeI7bJM10nSh9hsY2sESOgqsM9muiLa0A1RWBuVWGynS3jrKqCauAX1U
fU7jXwsa0int4heI9clMsW0utSQxv9SAMi1Kwsio3PfdLu3T/CohBaXUgqaMpDM3YCmu6Cm18ka1
sApl0OJmuCa7EoWB74tdPxuxocYC42SqbwiLE7fOfmihZOFSsZeGTzAvAefMfTU8Mh+SRbbM+jgG
88lvv6gy1eNyRZDDdUQ90GJ/0ZrxNWfjeUZAR7ZMkEYUE7boMpgMEiL9AvX6kSPYs0dtbif3ecFG
TBDez83apyj2eSGTDvdPESWVjisfNLT5wrob3b8x715rgPWzjwpMd1lwgmG1PfDCMp/iYrOdTngD
Tn3ySxqJbgAxpgBATrRqTH1lPHW0jsGiFteKtmJuhaWtr+pK11QmN39joRdy1y2iGdB+jwPYp8qD
6UwQTNvaJgAGieQyl6zy9M1CQnAzKDtoYjbr9YNUkCYoz6Rp2MgYFDO5HdjowEBv5QwSULGsRxaA
J1A6rmbWdJSmlxU2hCgPbY6qYuFTcBTbzNxAKT9YJ9Hblb+ZlcdThMV/X5Wh7FphFEvAXyQndFfj
SO1xzd777k9/Tu4dsXKlr2/JfiXy8V3ZXBTdH9aVfSIXJ3vIXTrelyMz+7+lpCyTuamK4rZCB9bg
5QUpUiz8m9elAg/2q/RS+dcDOqQp8XIJCbsnk8O26AOlp21QKR7AqWoMHY8KH67B4ClERD84SNA0
ax3KS+tKnMyN4PVriS7uTp6Si9RXBep9v+eOqRTx/K4SoZhn2Ll8w5JzzC6kGI1T0ppC9/7tpEkA
mOk91MQ+F3VfaKvKCv4Tp0Ei5WAlUoWLSDalk7x9hAkanA8z/vVun4jbqRIiTv6m/U/Z46emUrKL
wz58+078NGu5jf8/ikMY5Npnaq4AnMO1fj03TOvab/4iLAK36QDVDmHLu0OXBuAKNZRUDsYk0Zbi
GRomTYsOCqKu2QlFFd3hx2A0LfL+mAk7Y+FmJKTN0TzQBVxK52ft3kpEdR3//kZZgSY7AecOXfKP
Jj2fFKsaDFRrOiVYgz6YjZHCnB9TQV5Db70Thba5fZn68YDorfvvASLkrO45WbnPZEtINwV6D83M
GftE5KapG0x5xgSt8k35LqAEgn9Wpy+v27Oo03q/3vBTREUmWhDVPIcU97/0gSQd4y2eaQEBx67O
/EbyjblclJXNwF81MV4KeNydgmXhO06DmOZIMehU+DoBD/w5kU/e+a/Kr2FyfU47z6wfByMX1Ws8
w9xGlUts/Mmnk2b8/o8JyUnq1TDEWmyYoeCqTqSfLHRS3pgpXJCHg3HspFTaGUCFWCKhTjxwf0sl
F/JSb1cXarWIoDyepNKvxZz5pNfYhYC+IklvgW+57PPwPJ1LteP2BL8RabRxS8GwF3f8/IPN12KX
R5QPup6iPjmuoBwRc/kYfUphWwG1vG/jIlheHFJWe3uq9GkC4A8qM6spFxBmc3tTlb2luUwbb2uI
+KDu8DaP1gEV5l1bWb1T9mNt0sq1xMSA/Bw3MKHkEFSaoip378QBBjMDBrl07/4GKdlv1UC14HXx
pEGpohhNS5yHgLY72FKA3IgLP8JvTryy24Psu7659jCs9/OT5nPoMaO4VWWDqLPlZSFVkW3dJQjM
Ru73vXMYsq8R0/0nzD9v2QBtNV/cyJM9VqPC6xaVhO0C/ryC3YK/e00Cg5i3BS80oSyg/oaGvihZ
bmrF10nzVfqaxGWqTUKAoAPSnfYWHRNR3JsZVBcDdlcV7w1f1MTjBqfdcjCIY48j+VZn7WLkIong
2HKZt8ju4hVkukLGMExzV5cwi6L39Ayw9fVLnLfYGbxupNB8o3dsObPXEVPFm7Vq/4r+rvoX6mSn
3t+RDSCGU5aRFi9PMUW1oMx9bBEQafDqTwy+MHofH+4vDoBptT8G0s3mHzqkc9QmxABMvgz6fzka
tUlAFULv+LBSeRHN2yteAK4j2Bn8TTZCfUxrKsC2evMMvELPUz8BDjFt1SLpgUEMQHyOcAp+PEAN
bBYmbfsHmxQtJHla52pYMQmJMIFrdqnGiPXtwb8J2/ExApqipeWnqT3F9perJsfTCCeMg7FZUGd/
t+KdPUGtwaKedHOpbbq76wwnhTbGJzNSR5ADtzIpfXvJV9us7fI40dtpt63u4WL2vF07UWZfbv45
fJTn7w8XaXz8GodCka/AEBGqFSHOYz6bOOpslFl6elyT0qS6gOpb04Gh84pYV1zwPFf1KlueCzls
QbYyv6g6lFc9PG5WqOCcRzEbNdwYcb6OxaapGqf/X3z4hVwBB5oIDwvfTQ/X2CEb4hsJhZjErHzX
NrWesI+R/OgYN55rAtVsuuljeGi3UI2AKniHKCe5Y4c9R92taxQgvCBIXhv2HrkF4ZAM62MLTCeq
HrED98hGEE1n4GwAZE1c+HkUTUvLin5g0f0s4tduJC8kXszsE1eCYLjSvVK0O/55pICZgCCVKV0v
WThS1hTvcuLxV+SQ9uuHf/vCaUrwBXP6jUlG2js3t9lHLm2BjszMCvIcPWxIvxv0R8Vm/hU00M5j
w+gbHzlmcghAiT8SNM56VsVH02oCoIUYoObBgy2d6RJ1bY7vdiWUtjryGuvf9yzzGW6OqvNPOOd1
7ZjDbH3Bb74kuJArEDE9j+6yy0+eQeiP5219kGd8ARn0QFvKc0xUJjdGOQU+QVEdxqJbRzykWTOT
Zs73NY2W9WOMHIraFb5vBd7zfqD+xGb02/NuL8a/SGreuJvBuekmJWQZnJAW2eh2euecEIiNm16h
2A8Ejdw9COcm8k1DqKyO6b+ijeUfrW+UvO48aCLwjYf73Bk8XktHpJHDaIBhvlNDV809SFcBC/XD
pyX6NT3V6WQtNkYZKPYakZA5rZNIiwIpSF2jxotRUcnheoHRRcjOUnb561fR0bQurQ06smdtdYah
siZ3cZU+qxp3bK4qjRjlm/h1QhFNy+0kCFEVSFeoUgkAzO5MLOfyownWN2dL/FV5F7RDNaNldi9Z
d6zxKdxQClS1bQzW1vLBFZsWNOd3qzBN8xz0PNZokdUUKrOyY89w3tup/gUuky3WttjDYNwMAB3Q
TNl51ye92XAP+GyfwuQDOY8St87+5wmqE/+o2kMSoizCi1bTwCS+TbXs/F6EoK4sm+pD9rlpxaZ9
XAc0ZoD0Brj2fkRbAMunrSpRumHAkmjTvof7OOQbpEbFIguui5Fy0/vy0Exhx3Kl4EjnX1uKRlk6
P0L7DGjKn5EHfukAOs49KffVy6dAEPA9YAmPHl3J0e9jeLPSv0bw4sNNtb1iNO09stXS/2m+DgM0
6v1e1jRi5lS2RBJ4QfoArNE0ykgFQ7W884m2dUAR4WlgyTBmadsw8XKfBfvaLnm1cojsVJgnbG3M
5DhQvSKWLuZoQUycKwIYSBn+bFb9ZCisQAMRuqMqZocXnImptk2D6I1LTSLqtA3B3FqbIgXwEqh8
5Oq285Me1etdALpZkxHrUKARhAomdRcGKCK7KVfl0RvDfhU6zHFkOBPoFlEaxStjCzDW38/xPDy3
XNga3LW6zF/7J6Psl6xPhytyZp9BcpF1tC/MI+FrWIpZ2R4/oOrE1ud4C8E5ufypMusg0tifWqX0
FFW0uqN/dGuM7uk4tPmgZ0xQnqte8TJhRqbIK7IJAC78a9if39kOh8jJf8POf627O2Nos1YsnZIj
7PFsGze7iCwGPTvOd3ZSxRCkH3p/ZJolbsaGJtmzi0hjVFIpxSZE3J7S2kumfe59W6MtwlDNVYON
8EXoTZbZ2TD7ZXSeD8D7IW9JSSSdgJDFJJnVhhv7JWiKTF5mAwjmtjxXE9UQMuNqH1D6ktwurKzH
Zd96KBbr4WL6xyouA/yrBL+0wUH3VdysFAFCBxb/EB3js5wOnRNB3lp3Tnoh/OMFi435PbOMY2PH
8zbvhq0Ua0KWr93OarLxZ5X59qiDMwcWId4QHZ9QIrp7uak03hG29gydK3YpcU1SCI5ZFFz3chbg
OUxpthis4rOCaXwAJRAH9ClkelDs2k6TNsfQzgcB6/OdBaPQ07AYFijeezyF5QJTTZU3tDlkqmbo
gPkKnPUNmCpNVQn9H/s1JSe9u7LI1gJ/lYmh5Y26G0I8omIHr/LwppXIZ1Mnn6SqNf3WAyqkkGHc
Yc3mio7C802tb7IquP/uL9ZtlMfn8qikNZMtoTB4UagTlg8mpZjrX8bAcTGG+lTX1YKoTWJN8g5M
YbEWIfhEF/YuU4sGSdb0yJ+qHSvTkICE4fFOeZiS7iAMHF7O0kmDo2IKsFBJhgNsvwZORZ65KGx+
5gArEep8gXqSWbY5AGC+dV/tUuK2dI3oMSGqCEw56+zRi432jPOfsGlvGRxzp4RfAuVRVCvv+scg
znUw5pPdlMjLNzAQWlMiPiEo3v28DOQgp3WuH+6MpBocIoAp8LTv0PeqEWn/lZ7g6c793UAycyfh
wd7+1fMtb8WKLL8IBJkLokB9Q9auszbRR1ak5rZygFs54wOV7CEpy41pR8R3v5NIey6AFN8i6mz9
4yMW08mBxMJT28UX0OYSr9oTfGg2Lz3MAY3RDzadtf72HSSuWWVggwg/t4HVhDx1DSx8v0u34AkZ
/AGUCMIchgG+SGofKnObS95da386tjgo9fA8lBGO2mhg0yBI5kQeZIbae7z6qflr3QSIwHv4z2fd
/jwV+EENeWjLtBXrU6EW47EI0Lsx9wSM4+GNrtgRidJc4y94v8Ivw7vnbkHlornxxVpv89PeXnaV
8RIML+tZw7OJcZ3Zs05vfUP1NJhDqbiguv7ImLBTNQDVcSYrMoQovDsmFgRv+OhBUF6h23bf3Drm
Op6OyiU5nHcuLzscu2wA4lYQep4o11Rlwu5gL4MjVEzRyqR1zkaj76L6gSQXjWPS/MIKofYJciC5
5tE4GZHSikbF+hbjBfzUxXY2eAfyCqUYg/CqFRTKVSt48IOINfxFT0c8/ndaNIbBbHwztAeMj42E
gb6oturUxp5jUztDRER8CiP1JOnR5JtwR60FMKg7aLE1vQ5KZH11UY0lPqJI/QTgLcEsvs1mLHac
4y/vLckge8WCMja8MuKw/Mn/YerV5dLSi2A40sWwdYqiknxoAHZIYJnQtJpyNxuhMFocC1P70A09
9semBuEyJ01ocd/uneBm7pvXZzGUtMk0VwenCo0lNUOalr1wcmYmwUDb7GA0zs97KDD5UhoZMbeR
Hz+vxFMxuO8SdOnkZPNuimGHSJsjqt3SATtuaFwxE2z8/adBliYOyJYU3GErbSUtXg8Iq4qLEOfb
OVHRZpbOo5vKkME6p8VUmyeiefLZWYzCKcPuCAFp3o/aLDpZmRQW4lmyn0CA5ANYnCL3jy8Zr6bK
LKXIQiaIGXl4ttrZi6dqcmlw+E+4sU4O2BYV7EKCUASRLSQi+Jsw1CksefGpXBnp/dFXi+3wp6i6
Ulkfi7DZqX7l6iAHbxyEFbv8ee3SglMi/ER0x/z1urt58TnLsq1CYQ1dZLZBcdP8Q+WF1HVIz0oP
3cD6TMPDp9Jnw3aQwRX0xqEw2IdBCHWbtFdu4+T+6ZqLEyTHlT+xH8ZnPCeAJXcR6w4VM5yHPJF9
vaLz2uYga2qv8Cp3heRgCS8HmoKfCAoEJvLF9qfXwLhryquM2PydYbTAb5TDqtMDdNf5dZ2AptE3
qKkg39uSPTdPP63NKGMqdbv5wJRwmA53tHo3c+YpS0eOL32AfePkT70Oq8LexsZGdWxH3d1GxwZZ
WGfKq3qkrb9tSp49GZxNgi6la9ulraJUP8YQiqAuwJBa6/l6KioFz3bkKhaKO8jCg9cBvdXuiOqi
noy+EeSrXVFtr+d7CDJUmJr0H/I+ZZQ8+xU64H9iRhDrRL5w/FUrK4trIIRmEUq7JGDXJ3krWk4/
Oa4AYiTmoJBMqgcqcipys78Ba/OnXV6xNYnxM96+DHcb7v5m1bLawXUyw9ZMx8zrVKfeM8DaHwZf
LDYaPRCWWBFyGA+k0559cdgHw9pNmZjkoqwtu6XfSlrQITVn0bV1640lyTEeJvmlaPDTh97iAPT1
4gFjlXPnCK7cyAPifkcuImNxq+XnUj49prLfWnB/0MoDAGPZpKEO1wl3NZOhMyEZHIN/h/QcBFH5
m8ZapZpZ1P2zol/A1TaOj3w87BXO/9MKZ85YhtRFYKglWjPdSn7Dj8DO6Bh/kOivrcIfrcF9nYBJ
Matqn6U/b1xcm7dRxERRVZ68iwKyLZnNRVduD7PUdr6bUqVNkCtYAlgh4OhgJIXLd5e1KpnEo1TJ
krzX6PhoAjjX586Fb0g059nnpupcNFN6l9xpUTIcJYe6UKknY2Y2WibLZyR9jNye4GTV8gJCHdF6
VgWjaozZ9cwcboDw8F2EPgEe7nNM7cM2t2TgT6NlIt20gLkUTQxs0Mh+7eVIivUDW+6P3s+RoJJh
T5jtCGP15sm25P6/BAx/2M4vHHvy6YmhwqFRuUH9en53Tgz5iZolCis74R6mtpIj5A4qH7hs9pDZ
6eqpWjKCL3PtUpUubzK87NRaqF1DwDd/pS3/o0h9kpNfQKPQ1FuIcTbPPrZpgnFD22Z5b786JBfi
lRb0TKn+RhFI58NlbPVVKRI9dDrkiQHl4UvOacDV3P/bXwRZIHgD5xfGAE6iJKD8Jx42RHIHMlau
6znwxlZVMnKX/MXF87UvJ2ll2TvJ8xb9+UkxqJ9ysO4kPh2NsRzIOGYtU0ppees6zIM1RjeN2buo
kjsY7DCsbTctYyTOX/2Y34pjvabS1xanAWtKR0BvqIzDlsk0Kn+zBWRu7ZNhet2pfo9Pz3uSbuEb
vwK4TEjxbatZhEXqYoxGF3+hUr+HzQXqP+CNEUIG2Qf1wcHWPqq06sOAX0rNPCWUpxFiuDP6HPoW
z92/tG+x1ou1SvpkrbLhCQLfzQQUgHHuIeZiKkEle7iWwNcDiKlXGf11QEXhkIjUDGZDeL2WLFYc
t9ipH3UPzfZh0U1GkxSgt5A4vYnj/3jCzgSYpIKLt7gQLZd5ho90VzYw1jiqcLjQoFat8DKKENz9
jkVJue0i+Ko3jOz8R4kYBxjquQoU9h7Fq1ictj0h/LySJgfqgZNo+5K/fwcYvPleiM4IhtT+4wAw
Wg8Wp2uz5zb7mNG1RIj4N0+bTJhLxjNltbTU2WMQEkC7t0+mIzuRgijgHYTjWN/U3zb5aORDTP0O
kIU/0IhMQbCQMG3fsnMXMjOGpzS/LvnEK3/0QmeooFOv73HMAlAl/gXk07pKBFi/5FJjrbDFmYkk
NwalMgIA+RETM+JiKkHBGKnclZ4xgHNbuXRCmHBfS8QWWsVKz+byJDSsszmwL2oetUVG2TQtwtKV
+bCX59w+qaF3OwCfiSyyOgJ2v1hogOzM6gKiUM7kOXsF9U070Bexkt5uF1nz2MuKCDD915Ws4ONI
ICZnbVmbSHkK9sPcZY10TtLv9LZhOM0kHMTNdkLitPXanhLcHovLUg5AIaC9Mp5V9jIRhBFn5e+d
Tpa3dL5RfoF1tnDTIk9YupPYwQAeoaf89plt3zUYlylHVSjhNF7WYga3DT0YJXzfxVTdGqzLeBTi
JdUvYX6OVhnBLaTkW9SSqwYZKexcOWMo5NsLvairwSlJhbY92yCTB2pMAiOuyLZQnwiWTL1wP19Q
6eXUQvYK65YJvktXZq0ALSQYpnpDqLaqgqU2MfHa2Tc+l41vhuaaTXFcOv333QsdueKWPOVVyRNc
vzzpL7iOTCn4MyqUaAgA8NzvWXKj6o8bmJ+ihBX1ee2c50U1bcVSiGm5VL4Qzhr66m9Gd+Iov3Pn
Wq1ab0oPdBo1nsV8m4Nj+tXkUOE1Kob0bhAtA0mjtrw/1VGidabTMdx8yF8I9x8Wi8ijsN90I2eA
xCgU/FP3DHcTREUhCxUP+XKxAWt28/KNESVHN+enFr4spUtFtvCFVyyZ4MuydBEXU/FnWshGkumf
uc/6f3qACmPtU5mqkS8i/R1L6faK+RFLOVyS8hhulA+PXiEZmsxGakpe+cS1N9G3h4fseLg9elQv
0EIHZi2d1Vl6oRAI+6DaqpLds4eGYbmWUVk7+0xnzgq01lzoZutrAXM+XoPhArB+7cx2/SKtb8KZ
wD3iu7Olpi8Pt58VUz5W6Azy7JNwU6ZSopQNGme6Hypu0grGg8cBz08ShRA/FYs/FFcdn5UXPCwB
ooFb0/bnV/hR3NFbF7B3hVtz5r6LTzXnTl3M7cj3yGJKkqh6Z9z/1UY4xVkTLWnBGRTWdOu1aPMa
/lmThEDTqKU52b9V8q23cBZTJUcjsFyLNVOxL/luBC8KPr54WrLUv9o1dbgccZfqzRgvCxgy91Cm
WCbwTVRzivvAl9qs1XjAFk904L57HkWvahIauacnFTO3gOJo87t1AxayW8Htjlusu5s4ddr/udMn
eMG8sRprlNFNE14sWY+8beUvP6xQCRYeC+ufXq1nAWULXOStWdHs5oP7eBpVaMPw92+7LhCJ04XA
za80YPuA0/1rQd9byKvrZFXrDbRMgX/pbk+B8HNMJ1+OCJAd2ks+jjA/Opqjkvg8UP/C1kVuPh7z
Q5S0euOchdO+ay4oU9U7a+aLtaDupusR3SAil2hnRFS8WqhCrCyixmVW6H0FSyhWY9d45HFSGuI+
OhOIMQCwW+SnokQ80tAF61oW3T3nxH5O6jx185zr2XXrNaKoMgzrGa+5UCpYtDlFlEYjglSHjWkb
YhSTa4RIH2oOYFd5uBkFrhf5ANc59e6FzllO9rGEI83h5quSXh3qUXRGy82lstZHFmBLhRkroKyd
JbjeFUsJ5xLVVP5niDZf9rbVI2lkmPidi0sHbyXu2oNEQFV4Rm/ZA/dFk9MZGYsjS7xIATuHDm2Y
dbBECLdZt2NQvfsaC0XH57PoVCrRb9SF6QmWZ2aIlE0OSNGaS+ou0yGUlM+KH/Txv1kajkubnysS
zA2jp7MjgvGu5UqsMsDZu8kHeFVG84yY1auLiLbE0vVukBFR8IE23AbhLNbk0waaIN4KnyAtJ3Ij
eRhYDfoXRrdPmR/kpkS9+XS5IIvY9Mnmq883y5XIQt2uoVk6ps03a2Is5CF2XZz+ApY6zCqSO+br
EW5OC+VDHI2u0rhPcDWTyMf2G9sGvIuvSBnZDIJP7Dc882BV8csHnmBP+vwV2qpIixos5Mo1Us7x
tRpgkSM5Gx9L8zjvP/5gw2KEwrikdG95pZxWlVI4wa3Z9BnycP56CHFt9ewbxKz06ucONtpq+kWU
kKyLtrssHIVZxChF2hToEHgMaRH4I9C5RvqsEbEMRzPTmhEQTL6eJdBzNZn2AeY+3po+47GA6kDG
8BRuPeqn1qKLvm4YSoemEVLjv/ksYXMzKMEklKuAQiAp3O7TYOa1oBPZIlBT0whyXJHpEsy3IaN1
bA4pqgGR2mE8luzkRr+AMExnnbf56/IFEosrb4DJJQza8ok9fr7wuTL14oc2sXKwlXtAVNlGLEMg
R/6zxqSpy2GfIxYtdAOMd6Hw5gU/N1EXKyqNDqp1ZnEhY3JH/sTAJoYaU3g5E8sCtkJUs1Ft9dov
ts8uMHnP+aLU28u5llgfYzeA5p76H3eZm5+63hDzvtGsmM+AMQrcZrfj0tjjeP6+mTIwv8ziLvzL
SASLCjxW+73qWTb1XMIVs8ntGrw7IcLKyzjzbEnrug6VIltuZcs8MNu5NfmFCHKuhhsfzoo9gxtk
T+/gkkdZShPXa+OGJewjJdTgh5jP0jR41e55wb2diTSts5MlTRupN9t7xk8UOSypKrTYP0nM2XPl
px4yrPrppDOZsQHOfsp1g1N5C2CA39g8IbyQuyXrhX8IQJiUmehhggMtQW6dy/f0C8/1goIetz+V
GbpHQvIsyyLIySlYeOBRK9DFx9/qbmIxGcvVu/P6XkkTcrsOlOd3MXCe4QURbFlcz7w1NdAtPLJW
WsKqD6/rbpe6HprX4Sjg8QXd+2Wq4u4PMVnjKSU/0Qov7R6E0JUNBRflOxkWyZIUERFH2BbGyRzZ
w5cZgaXPIU1VknvDuBTOO8C01bY0Q2M7Rs8BS/g8Li38t1wNWkY39+KXKeaXRU1PigFCFtrZ+0ag
rmf+8wa5C+M/etwVlWrUIu6m1ZgfeSR5Yrs29k3xE4/zBvnilY2x/MeWL5Srjh0uO5DxAqw7X1Qi
0XFnOI+R7rUFeDnQAZXyNypkBPGMyDjvEKM695gz5D6vWQMPGJ6g/4vDplCXFguASeOwI73d11th
/An+FxjqMDFJ3s9kZMt6Z3xpLaqzpa9AwkIuJeworlaPzU3suVezJGvJqklN4+Hm/SaVSXL7gbZF
Li0bu5hIZ6mzSPWnJD5KCyPJc00GfmO2bY+CA68/ob833RWrqS4oM52GT4q2xYLf/ujTW0I9iajt
/UUbiNnXVgoZXkF2p6EY/4aKN9cSHUrm5+NdERbaSeGemlrRaZzbCwBw81Wxj7jjo8M7wkj4sM9s
CWhWPRiDGGZTsJ9+W3np0jaK6GbwKACcTqk0uyM8W5i9krn4KpiJB8sJVobAC2h1fXCxwRzUNd1Y
ZqprWXfOV9yNAOlI5TDwRYnm1PBB8POfvnWX6c9JtGO1EPChMRq+f7mn5YRHwE9uKC+SGC+amXXm
5DEGJKPx8Hgfby3XE+W+AABkvtC+HjMbw646bHbMbl3r1Qo+BvDkJ2c3s8rdbYWgLp6/jhLjGtAb
bxSTfO5Pws4X7DZFaCezB3sF4tv6pb0GnsqHiJ2lIlPyiGCJgW/Zj5x2tc4zdnSOSep3RlpS/l7Z
dXgksPYzRV/xVoJg3JtYIhrvI/ifsylfFv02mIAuiQT9zQyPMK/IkzJkyEethZ15M8Zp0Eq1N33M
uL+bdJDZI9SGLgFwwIDg6LXhyLUcchvvWqGGNWf9itep0W2PaEedrqdIG5Utqe3cRkrqw4Ufuz6b
DtmE1IeiRaNUwBGeonW1pY/MgBwbW0fitqIJHPI3HJETFrHPzb0MuP6FeCaNuAFaZ5K6qHYcccZc
lIyppuMFr9j/r16BmphPVt/Z7bn1CZg9sQsbl0SoX0hDrtQ4mDWhmY63PAMtjSznh+E0+Rd+uHjV
PbRmxUSzEe5W6dCrEdxfLyGyfIimiGhxOwtf8zpyAK+rpQKzUk43bWDY5zBpjNRlDmzSYh6YS32p
BQKQYZ6rETgG+QHoqciSUq7lM7EG2G5nuzuPwKmCjTgv1ZhqaidmbxMAOUBN9l7MgcPw3mzOp2FY
mvxnuPpL1xlBaQKm+sFuJiAItv8yOLtjKe/sNWLpCEJK/CwYOoMJu0A0MNA4ElgyFSVJIEd+j0TS
xFrUniWzq3h8E0QeyGxb+IUsOaPY+qkcsMFP4pwRzO1MlJf3WZPlSgXlwH9K1vtfFxdUSbivGaQH
cT0FRuHvLBpp1zS9N1hbnslG8VPNJjwmqJPw6EFfJuyS7aKHkoK3NGN1IVQkuDTgony5aa9QA2Qw
d0NHUyrkLZecpRHa3YAwbDRkzSqz7CpQm6KOoHHHkPmzpMEbW8OoXjvWH1GOovzh3bjNK24o2avb
nnc3SkKm6rHoc6YP148dZ/yhg9J01G7CP0ixUp3fWCI8Ken+eFx03I5bYHntxTYCplLwLexuUHku
RDd8U9MibfeaVM9T9q6svmOT5QoB5fHmI9U1JDNVPg8a2wobb7VV9WvMdRXpFCklnv1IPwGEVYbf
surLX44bHGdt/ofB+D6P5CsVeP8CB2g2SO45Sw9WgzmvdC+yd06gDdlINMvTe60w0NyyTFI+UTHB
dxU9QgUHVtEykrXz8LzShtwquqyR4WghWEJD6O2Quq91QGKiTjbamymqUgtTmoH0QoeyL8qA4vmC
CAAc0u+GJvSNPlZdzgWgcWb2qE2l6GoRnYt7xKGtqLEgRVdxN40PzKOXNLvNvgXIKwm+uJo891Dq
CZs0g/4zVpoSlz35L2on17LpttTDyVF0Jp5H0NgkpSZu14jYBftKm/x/e2mJKnzJEBMYFU53LTmt
fMM/QwX3Pmyyf4iy66kku9WXEyCy3uoTWm6K+mL+kXesR/vZ4MHsiSWcvpyzfTqimeIgcs1RrlLr
ADm0qNn7qEX6HMGrCsf0aGxTm7oKuuv4bZ6QcvGWQsyyZIYzTNd5OmM+2JHBl4FkxwpF3dE+Fuwj
G95LtvMsZo/ZcK6VkamMCksUqbJrfxx+zRDrs/1kcOYHjJvX0n1jaPvncc4QJPnuH8PLjQ0KDTC8
zbHPLPB3oYYDZ+RkwhM0COW6KiHnyiDphMcdtnRk6cWTV0E1flhNQVVHmM3JV4cNDXZnUNge+Q1Y
dW3xCG3RL2niq2MfiBZzqZu6/E0gfy0cm5R9aX3aKQThOzwR0+alVGCUV4ELOzc/envVp0dXanyf
4RRsBnTQi4BJJkq3b3nN8opEe8MAvh8NkalU2abTPnvzYLFRZRhXLVj3Cm33cpfOD/fdhrcJ7ymr
djh+ks1O9YBglHUBYOJNrwTnS0PfDJFUdO7XTI0TfRatm5BAbJkwjoe6kMckJuWJcpLyeeBT5zol
NazDnvBh4V0MYs//vkRRJjpfsaKm1YtOT4IIvh4Ur9KTt7eaGgRkE55PmkrITctgGjXTibKyfBte
jn62Y1Ywzecz0wFmD+JEzMEpscNGuOtl5l5wG67pJbD662q9iSd8x1JBkXbI52uiSMJB7vUZIugc
dGhmNRQx2aOeA3Z93kRP71TGjMsBpcpkFFhBvJgk7KamQP2QXLHSdhwuO1YfWErlcWOq1ZpkQpVK
bDFHMri69DPwK2iF/ZE2OWcCNcieAEVL5gd4dsUOnq+UbsaYD1NdSC/vuKrEAb5eszXdjRHkBJGm
SDTo4QArO6Y8SoFLw6KyU227oDPRip9W7UUeaDDtpAxaZBUdo7hZfSeVvC3NEhtlrHDZAL6Px9eM
8udJ7FRQk59yBLgs9bDEsnVLTgOp7PWa+ah/g42+fGIxjDQ+hZbvr4jROPh60mNoXTEhOIwMxdPB
qhRnQCcNtd87Q5WrU5FOL/s5xuZ//GP6Xe+fSiaTEDm0KEFXvOO1i3CH57aPXJn0KtVbgn6KVgL9
lh3sKDEgSldM2KTy49HClfOhjnTYBLqy1Mf4/G1ynkSsx0jyYuTyDmrxarZgOXfI76fFmPUORORB
MobQbcoJkyaYSb0AD4U9CETHw9+VZBYPM3I6ubP0Xqxdumoz1Rj9iM08ryyreZRKiAn4eb8pirrt
p3bhqBX6wbgs9TOmz3qsA9Rk8xF7bzAlB+97S5tqA7rm2YGg0ie3hkyf//+T9yPgPGDs6tOC/BAE
dz0qvK7Wz8rS12X/AZ1zvHKrTxG2oJK8J9x/pcEn6bn+H/eiMSL6QiHk1GwEhdbr5VkmWIKRgmiM
Iq2JBBgQ3gxS6mn/cfWpbIUEFHpZY+7din5kYYJw+iwOOTgsWCG08BsUn+nk08SEInv4aSE71npv
caARmoeRj1d3nMJ6dpCfWDiyNTim58efLRSKtBkB29O/oppIpNKLP6qsvMlvoFP+qxBcgn0zqHZD
oFdJWWDyMK702/T7jA2hYpBFHnxShewVYxOy6uFHFbCxujHOlEAvhwogmtIRGHW4reVP3R0kBOOu
OhAk1bL89N1hIBECVdqDrj4LWfyzpSvld6PvQ3kUkJmOby+0dXu9iL1VDCGkg+b9W7UQoeWfK4kJ
M8rYHA45vvwAr0ihq1SISCPQvKmF0O8HUWGsgz/dgP4D3kG2CbUhlFziRl8YqIwGOoK1H2+zt17M
qS0Srx3yi8LWbMEdNkO8wfbFhw6NeibbRUqkvIJPCQscE/4oh1Dq/mk6dSuw8vySK4tKmnpg07su
sK3QlU9OiMxx3oJ0KimxzO0YO+sXajZlpJBNjIcYhb+DBjxIdJ54C9KlM0l6/+RSoAdd4KXgruDx
6T7PFpgJAMfzIsD5BrlXfSRKh1zk8tdvXqjRvsYmwTFIWKfrqzfQx5PMqoKIhBjgbTdE72wXj4Ol
bkC6FKcFEvnlEPnCEBHkDQ6IIXDvlxk2+prrzyNy6pmc8pWFPFZbyb5uJMYDzmoWmqUr0GUDcrWD
rWL+0dA6ls5AZap0WReWtu4MM4sUFvvkjcExqnH3+VHIEaqG7fTYgnVU2VKrW7HmgIv4bB8bUk3v
UGdMmjXuIZ6kJjwJpfm6fJBYUDkE4ac4eSxF6ZSrlWenDAxsEkUgNnDvCO28eUbieRQjyOC1SegW
UYhAdxwLWE6TDGqXCe0aYiTgPywloEzl5fnLl+9BEREvtrY8OFVuauaeNwd9T0OkDlLPyuaPhAWK
j1QE4USjMYn00MAxWh0cYYjSqUQLimFNDsDu1aP1Hnq4zVwByENDU/OiYU9VUr39T/d0El+RH9xG
8XZYH+5h8dZcCjS+Ijv2+pNR649AXQtsrHX97P15E03cRBnbI0yOl4q3DSFiT4oo3xy8AKX8YKGz
eogcDW3JLgKdwoCskTu/sSMOQJzYFs3dNhyp/JNKWg+9xlcwsZ1GEGgPm69sOdbkR0BN/n2CUUW7
iorpZICuToHN7hwULYu+aPzm+uOFFihIEVyyF+/4mxQhgfhNMKozmR7DZ4hiO/q5G9C8oAdzPizS
mLYltG87bTw3SpSCcPk/XK0Ri9A8vR7aFalcxUkVil59XP4BZWAVPsVyFrGnz9djJFXq4JUZNaw2
zMbHZYlsQZYxETcQUYX1xhLtdo9aNv01D5P+mw1Q7ptS/E9XPQBEr8SyqKPNjaD/PaO3U7RYt7iv
anPg+TfKruTkLd6JpOzMBYTpc4ZhlNqk0CgEPtpzRr89WI7825pLOvzRoY9snnoTxdSNJEGADmgb
PGe6qo+u4BjxwqvJb1slZRUgMtehTiYVL/JcFKZnZcLnjAPksJ+A9uFsKH32jfKnODTz4c6kdg6q
lWALRrm3tqJWJzfzZlTC+l4tSJznR/FP7mkTCFS/wmA8Bl4RuQYcJn+VRy7SCm4G42g0LxK5CUSb
K7uzGuikWbP/UGCJOEOvP2n4I4JRYWw2ZCgH9b041JiV38NVauFuFNvDxLE3SGrYhW0SOtdqhAbE
HAxCz8sgMU4Fn/ECU+ifIETmrgsxWP2pOXRjqVxDIUSh6nHL4odckD19dVTSDETyu6bN5muxXgCs
5pJHnDgQvkqnailaXV9yJVRxKzbb8kINTifs1xpNXgSJQLJD5Do73qq/Kh376N0u7d4SbgSkjTot
O8ChNyLZ2IYq8YIM/UzQlrn7HDjduXNYml5j8ILsQkxFR8itD6/3IaNs8id/1UTIqd84MUu+HjGA
NYjlyh2Z4VJQ4UukEQ7gaDBeSzjvdWt7DtknXvxiw6kCfAyjXQ0U1CdmakDuj9k8WoXJ+PQGlKO5
4Y3F+veiE/trpLToeq3oRLoOtZPaY3pQ0qTLYIYq5zXKcbsbjW852KNquG2l3B1EDDzlFcxt5gB6
CaPgOT/aOiPmny+9otMhoigKhYm9M5X+Im6JeyYf6f/EyYtO9h3ffVN0E1y0MsfhnUYbBUOS+Khb
TQ6CR0vYGejrBLMYR2RJ0Lm4ZZdNEh5vca01rEuDxe4QKQq61pPRn5qMGkhewNEfItbWU4PIeWRQ
Zsu3sJeClHWYQopnpyW108pBBce5HGOu+3+NNC6Lr5RI3Jj1GTPA79XwQSc8Gi2RIzeeUO5VqJbZ
6k8fGsl0oduAL5hvv9qsMt9cO5CIQ6mUA7EvSfY9SZEGMTvEqk20uX8zGf85QP3fnwPg4LGb0ZNM
etykwb4WG9mriys5CygTDhsjcqwz+GHK0eVg6mS4RALHoff0TL/x4HcX7/QdF6VrkirTfC0zkhfR
LtsfPXF8gw4UETl2sJUYgh1mTDG7VAB2Z81vl3magJpxDKBrILjREJkzxqNgAA+P16bTCJoG4DFy
M4C+N9wD6lZyjfOXCpiZiajXBfcM19UNAumLlIdXuJSzfkuFHgebgXiZkeNYn5ABxcYrpoocV3zm
7tzAuIWqEZZKccrSHb3s8yqO8kNQO4Wgt8LCQS+/v8K2sD7yYdotWSdnzQWLVgXPbtEa7GnFGA5c
JuvwWkTYnshrIYZ3EoyGm29fMTfTAw+Gz9s9foGTu/QX7B/c8a99yrdNKXS/QIWLfF6Ym4c8XyAB
mutjl4dz5jfIWlZCdsnaksfARpeN4gba/E4p0KwmmsQqWlWHcdvowb/7LL0HBKmSWugSr1RwN0z2
wPDn1XlGBZUXU3ceNpj8/1iCSZzSYckziNTG3AehFTQ9jhYhjxX7oGQVhjCHygRHTUS+4uCl/883
VNYfGyBKxSgg2KjYVQwoFk1VHKMmHs3iaB9Wg4X7HENwn2VSg6miXNTFPc7/LwSqJdsK/qNPZW2A
GWM3qV639x2YwybV8Rn8oYcqwhWM2MbcLxjMXMf7mcllK0+YjtIy8aOc8uTrS8uvkqAal6J4UBI2
DPO95Ybthh4eor9pK6pvr2p/eWMw1i2nD0FjFFW5xNw/34qAwP+N0DnjCelGv/OFOgj3dtgPU3fG
SUQTwS4utucXTpG9NH419xdN7KDdrd5Kh5HDHovFbqE3LKRHVsH6ZCIEnRVkICE7AS51+pdsyX/f
4aBDGYiHhIhbdNODg7m+4uW6B8fAqD4IPqm0HCINP4PBFySPtR2iR/fyqTO9UbAfeQ8f7zBIrgXS
Cyr3owf4mfIs7v3dot+Z+BmREaTggQi7Tof3BXwgDsZU6n5vd67LBuvB1Ku5/ZW3sKabyallroFq
IXZdTdV1TC0fbLD5SVchijxRJE5u5lwLDIlVgRMFT/j/3CENZd9bNjMLXYqivhy4ozoZFftla1AG
wG6SUdNVM4erVEuBavcf7Lz9hT//ENqQwVYd9edPyUUF9DP+X6mfpLrYQs1xWhRevWMEHXWNii21
2SUVg4A1e39uDPaYlSzce8aj3FhdNzNJW7yQjt3VCCeflXgzNKrZz3dBdGIgpxoo+i4f9OHlRZmj
B9lG7HFCaSRpamLiLUaESVZsyE2/uuNuUAGneergsIMzciVVLdaFDrvx76lXxrzxz3kygwumcA4z
EgZfGSEEk3m44P5NBsSxzv7TW/8OFJam4arIazfygfQTgcavm+7ERtH3U/U6friK99d4fwv6xK3r
1Gn4gyYbTvkqCC3tp49j6VcvJM9ap/Nzy4vgJRIYzBIrY3qFbromMNXIZVWYHNYXHExGz23UK2cc
oNYjQq5CNcekZniLEbHzIBsWSMqK0ZXI2DVfDH0emg+3dxHxdJNh7d1ydPianACb5xZl3LMoFWOH
hNpmwKqomrCZjkM6y8XLRja04haCGHhaD7TES1jcJqhPXUkIh+TRXEg7TvPpftjZP6sEfBTN7YXn
XK/aZ4i6Lr8HeMJmHhzRt6jEjenXBQGdx7ffREOgdSSn6w9SHO1wDfP3riPkuUZ+MOsMXR2ovleQ
fxbhgjB9bkeoBcjaDeuKwE2brmXbh+Otz0kAOz/x7b1vVaP3PoQ0S1QmM0p3X3EvY9v9I5cwoR1A
f3tkQD+Y1wzJKO2QbUQgE1HiQ4bCNYuWXACNkY1W0K9PaQB5Uv1lzfk3axk/qmzNtwzXUV/JTwNJ
YFdFp72wvAc4a1VifAu90gOKqDl9tBcr44g2qjXNoHGHPiaIcAhH4VZlm2dvi3+gS1bYb7evXiXv
Ml6p316hOlxPOtI0hMn+aE5h6xklJ/fUuhED32yWRLX+vJm/uTsrvbxtLRmwkld74t+1MJu5iGaU
Kfdy351n+jTQYp6My/n4DMG8kXCBHbhQZHj1wSzQ5la5vVD1sIlhkTEYwaHo1E83g1adsGxEyWIW
DcUlkefRvR/6QJ2GHAFE7g7eSsWGKWJOevqtiYx9aC9GesvDDvFdSLKgUH9eqEhATrDrDeSZdsSP
u5ZaAYS88ZG9E5DwQgwI0otDyTSPm8q75hbUUoZnlJQrnCeEG5kOoC4NL8/5dt+TZ98T6/+oRs/p
Yngodo99iy6w5wGOJx27Ocjrq1s3Y/fr+lCYXfmvK94ZW9xd5GM6azt3Clskqq+DWff+DFfjpJEf
5C7cNMCibuy+OrvKnsrAX/PR2a9dTnjD1V52C1WZCbfc+NIpCluNrWH5p7kta60SInbsd3uf2GbR
q7+Je1cqntk3sr8LtcrG7UTdacfyQUQc5uQ7ni+J5gLLvDl5Xm2NpycV1pnV4Tdfkw0aezl0PLLE
i6qqwVY23ubUSP4txBQFKHHI0BtSbnc/T07+51IKWkbRE1KYje6RPS8/AYKIvmBNndUfWsDA9dTy
v9difmf+0BebJKfN41WDa9t+9ysTVJjwtOvIy++t+Fj7tEXcYsEaZ1fo3RI6Dl60VGDNB8MVtQ3Z
pAKe2poZzcqB355Hf8El0KGkXZ+nWwAVGW3+paQQAQiqBwQKHotmw1yN4Q2kZnfh56ingR2IGjKq
fNMk2q5kIeswXkwRgG62rgag57UIDlAnkiU9F+vvNMKEN/ZLtbdbV+H+pM4GxE88rBgTQ5baOSPK
tqYqWR/u3Pa0B/kkyCQHz5EJ/hcMYlqdIqgxAYtjKUNLDJKSncKRLP/8CArFHRCTFst9KCTYgmdH
S9mZlauTW7+3QkbB/JpK7VlAElFm+v/VHSL0yTLi82jku0KavuZFzRoXq3XmCn7xOMsedj3fSrwr
jNjiPA288fhYn8TH3nFrJp3Lslbid6J/pgFDHHA8qg1D2jXXtjdZdCkvDFysdOZH5vH/y/AfKFP8
0ekNC2QdnaAOXEnktO9w3JVQu8JoSdnmvnW4umjwuMmXLXlLQqJqK+gAfMzbEeHovAn1DE6IwE3Y
QzSCuTysUVR4/qDaCA0w07e8B5+X2R0MY+DjfbaeilbK5saG1aaxYa5UG/kkZGxp+EOvQUQ2oTXr
14wtsK7XtSJxHWI7z1Z49MxhHmcRu2K9vO1GKNQNaJfDqrVUN/KJ7rz3c0zUH2keJNI0P/zgmhiC
ud7GJFQgni17Syop25t8qroFCEWPRofuMM8V1553hjW6htbbB+koV7vlFFZ0l0UT9av8zqhSqmuD
lNDOotp/fPC0qsTBxbnjzkYTLzhSk6lUCzWxoZe4xZVCUwpBoJd213vw2RVaxB69yr9YWb2bLaZU
/zpjokIIJZSNwTZ/nTWVDK53OBQzMSlibK/v0JpoO61mPEuMy5+AIIgWqpSC943KaHc5tOshlNBq
Brk35xHRnPW1GhVa9lKZIX9YYN7r8h1Uc/aEHcFRfKOcCoMyt3z7ignCvLCPQdVVQ+XpaujWPA4i
ECJSVZulhlrXyhjP2JgOcOV5oLUExAaxr9Vhg0HWlR0eKcJNpiasVTTx3fl+msvqk19sIQdVQVcP
YbfXrFt9kDYMN/6uIEERHXlyV/wz/kcGNedZ+3Okbi4zvYoMAChlMhlHFHmjqH8QeWKX6XcGfzct
4EDgg+4g3LYiAy0ln8z1gjl2rnSqF31tXjiYVU2aPdhvJfbpweGOaGT8wXdAgav0Ob/Ly5/rjhek
9fok0dFSEJKROijB5mS2BChcxrJ6MPFH/pWiIUcir1SwrRaUR1fotg6aDCu3UDbBOMMgf6a5oi7j
PR/PzhJNKfJoGUY6JzNNdM0QU/qVjurTk2OdFDAaK6p4H34TECgYwfjR8AXjHhD/WdfSAaMQNRhN
pxf95pYT+RCgxT5DgCIW6IEF76DFHLdnzxUcw1OS7ayXVlGi4O0BMUJrKVf07CcA7eLULxVsHeHX
Nhc+ys53q5E1tmSzSLDTGzoQZE0iuNOQ04bOaz+9DwTHFJS3FFJ5FgZ0Vt9voEBub8IinORAu8gu
ovsHyns0k+q8lGh8jCwI6hvWHqQWwGrOb4sm/sBJOfFxF/c6iMIuKHFSJSsv1MYoxOOipstVAyNJ
S92Z2CX2Z1xZCf7rHzeVb2bjJ2E1ge6pHzim/w3IwIE8zyxaeDxOCpmta/FrirV9bro7h6FcTC0I
H2sgrINljGQiIV6t6VupktUpuVcWiiFY5++RrnCZcNDyVsbPA1i54evLBIp4Q8KqkWwjZaB2LKKY
IW9PiHgpfgU2xhNWNWhAqQk75QQzFrK0dNMN3iquWUU90R8tGYv5S4DuGrRVEOzu6c7pnYwADDe8
Ur9BwChaSYDXhngNUXio/AVzdugkDqclkUVqZ4GZ/X8kdUosAGsW9DKIrlqRSMe1zkMAvXItVwxH
SWLVw8a8wS49mqIzZ7Lt+JgQk7xXwqchtryA2yVfq/2rl99dY/z34TpSxtNkZz2lNF1bn1dAFS53
If7g3EJuE74eBFbwZtPzlTeCT8nmnmTMq5snivsS0D/5psn3SrbFRa2ISkCU5G1+45ZZueWHgPS2
MKt7F6i1+bWeU0nUuIwDXFgH4MUaqLqNNbOepcdKpgFd6tMpe8J6V3CI7Iluw74/BmVxrAp0TTbm
oyFbSD6KboyJ1EP0DEaNR4UnsnU2MZraom4dXj+SVxlOhpI/sjuECpTndnpQP1B0Sh6MvFMvz51p
bIYJB5Tqj/VHceajBVVVk+1QXp2Y5kw9s0WopUXzGjvUHTUDc0F8iOYzInZRszMa6zGsYLwtwfFH
Ndd+b4zpuOsdu0TzYKBzFxUNNYcTa03JOq1bpZS+RW86mkqRfhGMlj4HXa2I0KCno+ShMOi+VSd6
PiNw45P7faebL7dRm03uLL8BkVqG29Xn0Ni/gc2QM7anFflMoROJRO51Byan0+/70WpdhOpWIgVi
drpuAGLav0WUMlZbsi4fUBwIEIYc9jKHg1jJuIQIGUof7TquCUf5g1tHCIkFA/824I/Ay+hDZJ+z
SappOqGYLK9sk3O27bZxrRtSbV+WoErc7JTpNBKXNaxPm1rM/tjojwH7vnvKFLa7xG94yMlXm+wD
UrzmMBbkHbstDW8INXcgOW56g/tvfWhOZlVMTbqz45UbV2VtKHviCRiT0OxFKP1whb/X3vYUIL2F
vDrR7Yhp+AneblVkqNehETb6FyH4ZAlt9drRpIhR5YASNzAJ8wvCra2MKzhLWMaHQaeU6rEnK5ds
GaDj70vyGgRL+4ckrNxD2Pxx/FeqP8UNoQ9nVoUut3nFIFgoDRMQWAxXFA3pEcV4pDDqxc0+m0Gu
E6giSFO79eUb6BCsAU7nOVuRG3k6xrvbIBheozZqpxsPslhzpHY67RdBw9VwPSye2JPlN5bdJUK4
sYckBmNz58IyNWrRuYydwO84vGDQeAFUHvSFXBOFcI8/WPZ8OaS7ZqN2XejGEoUlh/2M3b2xlbkq
ENVobV66pWzorQg2DoIB9l6UBrfPULFZ5RFZmNowkoQRyFgtHeYAThowjWK6+gyh3HPUypP+IwmB
CQGFue6+2je+9crUrZ5Ggqg5iF6393boZeEvkkm5LvdTlGz0ktbhIttSaig84rxWUF69akwvEcJf
a49TJTa5T3sjympOsutmsTPIzbyvhU8jPuKlI8glxZANEoxELYw9671z+9nHuIDcU6L39U2Nz0PD
xkqzxyuXKK4iAWR393nnQS47RFKwgSHB7S/ZGF/IfTDQFlU0sbB7ofqw/OQ4kwwLni0b1POOTZah
OXXDkWw6H9lkFxERcrzUdguCNuab+NeQJ9+iPfP+AA+vIzXwyh0eKFloPGyiOUlcP9wVk/qmDR//
1SAS1xj1OQap7sDARSijZOiEnslFj2Ziw98nb66N1sYM+wl2czdrMGNqNJjc5dcBJegFjFd34eWA
SpB+5bHd0DfOu7MQFUJoBAclN+ezDMCVOcaYCfDaEWlEGn7NipHKW0i6biqovU0BRq8oDvy6n3S9
4OApmsRZ0U3WYEhp5rkbXPKB6xi9OYMTn3Po9bj3JeXzkMZVYN+hl+67QfReuVotoV2DKG6OB57I
FlGfkBd+vkS/9Z2HxpNPGM1Y0CLAGVZHzPnPZZyTvMK0IJYzNea8kF8EhCUwR3SvMcPG70XCGIO0
G/8FpMbOpQRSMbZ+PYPWsI+tRIzFXUKu2QkYnFQZHN0YJloVlt/f/aHowl4+Tvwt1fk9SzD8rNSV
egu8Rw6JJqV685ETNZH45/wiX+a6qwKVw8+hyyyBh/1SEr6d9PX3zpPQ99uuAS+95qpV4JRe6UQ+
GtkphrCGq7Vv+cKVHW/8dV2P5ixlG3FgwzYGHeauBdn0TFBB7cLmKvCjvlOjru77zh2v/D7chJvl
T9ZtlUU5QW52VjIvb+6n1MvH7L+1P5Ttw17Ndb23Ug23apYHWzS6KtwWUK3PbCKmiJ/BGpc2Joi/
AkdCsHZhXDp57P92pS/TmItAy1j5jk9GqitmBslRu0nAxxnatJ8oaxDKHpQ3DJ+fBeH3Qps9EmT+
uq6+x/ykKsn38wddQKTY7nLAy/QIDoAtR2SSlRxdgb887aa2BsQF9jC7NWLo6az41+i1C7mb/v+Q
OcbsWgJUOxmJuKWJiTHESitndR08G2CHpM2L0kMYhgzzb5WmOXxwesy9l9zH/P+o3bxvZ7dDCPq4
ytFCWyYWAf4aqzTtz42mwCXAkU4/4eSL2JTXrnYoi3wMnQE+BYn2goBQLevnLUxpaYdI9tK2I3i+
btWM6bFOwr6m7jnFE04/Dv5ck2Qk48JgKg/1uJoC3Zv/xbH6GuYek8PN1l9bB8PhpWMwQRe6HVid
YzxZxVhlU1bxBEe4+3E/EfuTfp0yvFaf1Uh2xMVUoGvixIxNQ6kgN5Q0WPqLjI2aYfi0RttF/5y3
W1kVtp+a0vnPq+6nRqKKUtxFPep+lWKJD8gjMBCHRWWVFeWhDpgw6VF93dhOqcHnxc/JRpjW0h6v
tANp4kpMZ63RfA+NCPtwXVm59XhlYH0yHNRUutZYutQ975YKSKoAY61LgsvlGLBReURGyaXeW0r0
G0iQMxRibzZTAF0cieJ6HBpkXWrsYJ3AOF/zIdYQWJccgWiQqoZDnBBc7HRavuOfah8W+NcpmMKS
UK133g+eihViEzUTh9BqqGVlEYAK2nf8SPqQrbiL3uyj/woU8Vfsu6P8MmUNFu/Ck72KPeTc83nz
AStd+EvBau17kFkfwsOPf8uabhmDPjqciULDqAg678Wn2KQ8owsy/9qxdxVj7AeHzwoUT9otedtS
/FmP6FPD/JtF/C2FvOqYEjTGziZBvBB/oCtRhqOqNFoiQqBqyBFaUZh9CZFQLrc6YgsaiG56iYEW
mSKiaoaOalHceVh3z9yL+Q4RbanhMA2UMMN23elSiKYAX2SayegpSJpXJGKLDFKbkNoSWh/PriRL
3jYDdAcsKrEybXFwrRSonI9x/KJPKohZOOMBAWRjgpPgKOG1oWaIywhfn7lfCTj8MmMaH9Za+lvn
ub/KuxV9Nu/8iBOJRVPGs2tZBR3383UTLanp7jkXRAmJIysCzCIFUv9e3eZ80hnc8QSLI5ADrs5F
EESUi7XtGix/nWmRocOuRwFfhyDfMFC4zuAAUWFzF1PGnYWKq+8VUnqo5UZZ3Kgyn0Pr3C0kpGbk
GlQqKL76WYyYyzu/PdYsQLq3n8T2MbJQCfRSKGxR1QWBzhoSsn38mVmayijyEalhnwDc1z0JYuHc
FlE01/06MmQbQoO8tDVlE+sdsdBxn5B9/eWrdOQw47qgV64ysKrj9O+h5JnqejjPnho2wtl9XFwg
7xMtreIgBUynCE4+9GMPAQ0+4uYXsB+t/zBeIZSxGIdsw+gKl6o+LW3dqmcrKfKDAP8/ocQ5cjmf
zreaZVo2OxZawFFjZexWsJ8woRJ8WQrMmULg6TSorOmDthQKa1/XNX3UscXexF4cMLWJ9eQvV2Lo
O1RkZToIH0nkr7ueajM9IccjfIIaKFxcyYzOp1lM1+DK8dRiOIAdYovAF2KA229GJXa5MeRXy4SP
9gO6IpcWWjeSd2oNJbxlN0wqDvIemx4ePFvOUCUouqpl9ytVChFoyycoxtn1fukcUvnD9WDKqG6G
rD9jMqIRnbk6rALmlU4Yq5ZIB/kQBSnuf7xdQzQsQ+F/FV3E+xX6PeYLUiNSbaD8v04xxQMCHroh
a/GpMejx/0W705I1PR2s5tWcdz3I/WnWZ0WXBKeaQbFffSBQkLuSuC5/oottwOcntKbPg2Sy0E+J
HOKAyQr87/RQAlvaisnIDXtYmkpzoZE/oH3zk16D9BEFHT2zP24mWKHIUFzCD8dxU9a4BjbWbTlN
34aG/50Etx6FIvtRgjb418kiOStjj7NoyqZHP+WpvFolzR6lSCbZKOrVDT/IP4/g2ta3kuESyXkk
m/zB/oFe8Jk3ip1j7bgLOEGb52oCdDsYyneIY3lVIEHXV/7gca61xKlLHa1hxJ+iBAjYee2SLpAt
V5o1YYcnAgdoxgSkMhIqKBmLmPPkv8EEwwXlRkvcSCjxYJC9JOIW48604j95nKelShoJtVAQ1E9w
uGVGtco+0+MpwHImeYitLjvFqAXudLSIt+zZtGzr1gtz9PGLn0GkSxG7skAjrhfxF/p6mVdcTyZ/
pz+cWJdsyG211uXE9cWxgK/1TXpz/a4ejN9UwPzV0wVLWZdlu07P0PbqqqAH0mF5gtofP2UAUTWc
idtlRPwM4rBCWdgJW33Gdi5/2tZuvmSBJkfKNoYo31tCrSzmPMrmXFYLubYm/AcCIj6jq/K2JVgE
K1xf1tcp4+4fnzvT866F66D7WD5vfyGaZLZI/7Z2y8fWhCbDEMbK0+mSyM1QMn+18/CUm3lMTW99
JQiEuNGvsfIoxORarn/OscyvxGF2xuOfWYs6BgV8bfcXUzHNQXx195DeGa+Q34dJeHymJpS0eP71
2F941iPXKpM0rOhT1n/Lurl0BPNyvYfH20/a8URMHXoX1+71VhqFlQt+FOl/1UpLfJ/RU44x7/3U
VpgSpS02vSldMQe79dWSMqG/oalQC62G3o7vEpPXrnWZRNQXxDmm5W/JWlCrsLQK3CLJKvi1KHYc
KjLPuvJuJvwh6hQsJI7Jvq5eqOw+1CP2uIzEpU7Y0xoTKXs8wfnYdNzIcq8Kbnnp4Z/lGs1bt/Q3
yaHCprDUNk+QWJRtce1kmuye/5X5CF/FknQ/EwwYt8j+73kqahzPzumvcn8Sn3wogoqqDUuvXD1z
Glsn6bxU/ZY7px0X37zrZhwC9x0BPPHAVnnQxQq9MTofeOun2sscBNPU3KrJq301hdHGOYhu2pNk
6NBoeW6+JtaUJZIHrQfuI7h8kNsQHqaDESFT+MaDFUznjA9IGvgoUzCA9mqwG2dgwsvI7qp4JBXs
O4CHkJmmLtyRpV0vxqgJTODvcXT/f8qNQEvZinjkrQSHmle1ZhFp2+GV4fV8E7Eofu+1cP1gx5lU
TU+dgQu0/XQQEJH8QOgyP3kO0nFcDU3PAmCe4sT90FVuUkf/MbNwmwz788GDrg7WFpsD7E52OxQm
95N7h3PdDpVOd33eKHIu2xm/voR5dNb0apTyKcVcLfk7plkuC1u3rtvoFVk8Z/9voOwFrPawF2IQ
U0zHNzx5dH6LWpUfwNGS23R+L0Elk3edATAapMF3uDvztqd6Ytn7Nb9uOzhG9WJsz073IDw5PFG5
CC+JU5HO+6V8hMU7PWWxqqtK93tUelpM94UJGm6tlpBuzvZT9zoVQJ3yRAuO+wAC4ONrZEPpDYr0
8+3kXmKSIYZlLoTnGyZFkkoA5amfnUY1EQAUcahWT0dKBWTUJS2lFjiEWKHD53zle79oz0cPrW8t
XdwzQXbolriRvJ743xSIjYv+11Ulgh+UnSd1efDl/1JjFcT09avgNVdb3o8qv9+rhyDiM62IaRAw
B7Qe0otq/aoVOfgGB3kbsb3Cu11XPWgM3BMXz77spCgSd3Li3lenJTnO7sKrd6pkcBI2e2ajFsMp
P6K1FUOnEOb+qHlkWoi6MA81UpQHbwMERqiU0R1bJN81PPCAWVpHXUlSkyqAP+UDH+tatFUN0ZV3
V3yUTusKzBOAJSDcjs6v7/y1ZixlWYCgnIwGqOUn2wLrRro+zE8aP9PGdVlWavmye2nux+SlJYK5
FXFAi5Df4JKCAawDqw/fHLcNpm886+B6fNBfdLMArDhq/8/nSmz7xTZOl2fnO80CSiteZUboqOKX
hxXrGu8sC4w+xT3576zjT/YSvjyyrabjluaEpmWXLlITv010KiYUcb9TNdZJYyab1sC1a3XrB8h+
yTfsp+EK5ogCo+ldoTQ3W21Em5k+At29Pnjmqi40pDieC5yPWQCoghS/YIFCEmMj8UbSA3Vs/vIn
B5d86UJYyVuUgaBYoG3NhZri/oy8Gris+ZTFHdsjsoQfwZqRolmCv/Lx4AIFD8J/33iv1JyvurDH
gZXbnTXSYjoEWTsMAacfyclIsdRu/2ppDM9VjJNaAE/QAVHGTF6SVFC6Cj38vGhR1G2hpQu/h+A6
xvNJ/z46Za4tAUEnDfVsIqkNJbLD7I4ojI0kp3CVz/qYL81zbCIJhVuvSR6esgWBrJzVBtzrFU0V
Ifn+AsxjjxggrIjbrUKxenh1As0OuGg2tQbMQTtsf6R0Bj9jKWRCGUvwsQjvzNHCHJokkvB3E2v/
2pTeHRIDx3GfHfkD54ozhvqX8dQdARghXLczGI9cv7x6AkGhm40sWR4YnALvUBLLU6En2luTgAbA
s6Wza1/jCcgwBdFI/fYnSUzhpXwhmBHGvZoLiBX0SSmeADiJmBTkwbUNpZlvNF4lWlravEcd+DZ6
fIos4xzWOZbCuj4IH+peDNlifPJ5B+WJqzYFn4XNHIBnDkVqQFc7nJbRl1IkElmLh4l1L7welBvp
LipOAPL+ZEywg1HS80pvqrwxZ1mge/WGC1HcsymiKfDBgOJn5NLyxFD9nRTUTpgoN4xH2dC4Va9e
qiE21oLH1YKR9C9xEAVLJFnftVmO38gkn30TrotIlbZfymjgIi7jlEDU5mP9edmq5PiuBo8sXtL4
sFSe6CTDqUMVsqiufEDumg2seUAQDEeQ7iBSZxDTqbaI6a5XmwmNqheN4gxjdaUaL5b7fXoWHdqk
1gWLNlLeLNH57wio61FoHxpUQCsUr8G1awVEXV/ef1VECpccn91qe+HPni0ujY2XstsgTxwK1fgt
xo+uF9OMpyMmsI+O40Z0fM+b/59O7J7LIGcTRLjFB+e0r8KYDms8BMgsbNcNzABtL6QCb1EbQVNW
c+jNTwy/tEIdJLNfmSm7PYNX/BgmQj2p/R+QyBpbKNEZ6/hF4GR9GvD51CIm7Yal1wi/s2ytgpd/
mWnXVz30Z9V7jGtJz1X+CyVSEDHjpI99KC/gFDPzhE1SPcEZKKcgFJ3K0Y7hjzwZUNKH3rAll+Zx
Ts8FjNyfQpnigXsllGp6V+L9CUn+TEteIS7NCImTtoNMz6LeJwbflz635lGF4U1EOf3sRh3wyPJo
fUGs1D1a/C5mswKq6VVv+xp0CKNbVWx8nqXM+Q6neT7/aE3pBg5bFPCK4QQ+C4AdQeNc0W7OzNkC
jcp8tx/eGDWyoNHmIRcIc/eVqkXK/2QO5mXkicCX3ZowIjQc7ApNfuo57juuOg+Ap5vYnkcqxl9k
edwji3mwGU3TUcaOztJ53LTKyMu+UfASp8VLp8OEhqJAINMkVIQviZwZdVzp9T0omz5vmfhyg1Yb
+iIhRG0g9x8R5m6iG/IZwO9WAzGZ+8YyOmkb44JIHVjYEN4Mw+hh5T1ZE094v+vqvsiO7nIE6+Nf
/9gffBmI+A4e+S8duVba3nVTUq6IuOf3ztFEaMGWKKoPtkYlf2Q2ODo9mr59n+Hw3qhlAJZtuP2x
mR7zeXLTUUJG4Ttb5o233ZDjxOZgNmSiTZ8ya7kFLwDUhujpqw3vMBYfvj86NDU5o+wIOOKlsHNw
X9o8cGwPM2Rt/0mc9t4vaIJGkZAaKTXMbLkZJrrPAGCSh8sLsb7OqYIHa49N3vlULQNquTVm/bZL
7Cl7migJB7qn9Kry2O1NDRSHDPrXlWIaDn/xIEx2qwCwk0ZfReEVvECb69KJzyvNEa5lAleJ2zbo
WDvQ9Y1QjwPhSkXoikWFV9bzoatMfcLeVzBQWvigssFfrjiNLxykPKFScjCeb2t3Uo6JzupkHO4Q
l2He8b02Zz4HPlKEeO+1r6Q0j17HxG/yvcuOe197ReYKhck5Cb0lT5ZB6o5tKk9aD8Kw373A9HkI
mcYqOdUKMtPMjqfMSACGMmzG7k+VVR14DunFHGjNS5/1GtZ8qMwP7w7FoPzEW4H8Yxy8c34F6hH8
Fk8mFF57R42izqbpefE2HfgiBG8DD3LPUd8LizlFVY2b/ViApEEQ/3mC3ll3AY2sx7vM2qgwuY3/
LQCYF0zPXAu6JBogWUhvjawKfhzr3TD9aGX8tqi6dhdw+7ZUnhs8PbsmUSyL6keOv78wSJkeF6Ej
DJmz6b9miYYexu1c5rT9kG2oXc8VTEQyHWjEguuhd8laUIIud1HAbWj6oQrabPOa29XL3zzTXbVY
2sy3fyzCGmSn7/z5hMm62ATkWp3h0CmjqULY0eLFYODsYgMiRdlvFYSyn5lnmQTqabH1eWqIXQbn
LWUwQGV/xKJyoPCF7K9K97sVa0vMNzJ+xWQqRG0iMXq+3U2E4It0yPvaEpWDZNKNLeTNAtvm8YuW
tH6qVa9dpr9H5hHRJDkfPko8V77BLb3wRtN+ABcTFLWLL/Q8nMcZPzPzgHDT6chiB8qDg2bUNqXT
rAozo3mXyBFHWic8lfufbhyeLrk5WD0afu9DAB9eQTzHnCa43rMhk8MtwtsYk2aB+b2KYYvR3DYb
VeWuOvOV/BATy16PSZc8Or/tfsT0C9n+9Cc2mSAos86t4VeN2Sbw/a3wL9pb1l8xp2r+FY6Qlgky
xjSbcWMZH0FTMulgF21CAzGMbAbDo8V/5pEdGy0SxeDsGAzbJwVH+mdRhBslN1kewR9x9GgFZ5NF
1vZxWr5+UiiJAYtVWr7tjLQ/nChpP+0Tmcdi1GcCUWeoPSe9en+JobLVWPFf7DHf9gZ6uKMlL0OP
AQRuwDKEvrcNZiLpepDHpPi2/a0hvZDhXE3NU7LO8NgkZAhXFLrP6AiyvTTN8LCAQg9NGAHrCiDA
7QCAndJj83lzosvzfCB+3tDs9fHQO4RPUj84QlC8hlzuN+6cKVJyxoIMaxl/eXiq2suhK62NxYsw
w1T7reSeJSgS0nKFOcf9KOLGt2tc0p144jg2FvLvvKWU5Kz96HCw0nNCbxs9IFvH8afAkfS6GUj6
d1/RcNa+nOsvH62xQukJXJC8bvHD8h83khaOGBLCkm+CYqwMu4myZ+avtFW9dIp0AWfKi3duJrEl
fod/XXYiuEYWcm55b1zrYoLxXYjXY5/yfRLGs3zviOux64X/y01LEtaQQCsXKLSgI4+T7/sGr/gU
2VejcLDev02RalxOa2RJCvrkyRMFMzlwAHT7wTBntWzNn5dt+LyD0ZYH8pESi7Tt8ai7W2DK1uiL
jGDE3AvwNJquxkbxc5sTZaFseHksL3oEqA98iEYJaIgZZ5eURXRVn08dpF9xyLRZjtaDaXvw1jdL
Hxbs9pwPPryRHEhWOvHKjOfTgW/aJ0LmhzM2fypLFuhbWneiGJkK67+TRgQBYyRJZtXl0k0KC7Gu
TUda4Df6Lk+q7BrDLNDkwMjkUG2G0e7BTJ+HjexuPAeDnHXcj7BVPNe2O4QZR8sTob0gjxSpyE71
cRyiPOHRddAdi7tSemmuZCJbsTWQt7jf5ctjW9qdESM/sNGk+JpH1GGZEa3U0h6PIMdnzSeWz6Bx
eSM/dqsdx1zDXOW6hRV1q8ALLP49uBS3GvUm3d1G4VXD5xjypiqENA5eZKt2q6R7NdKVxnf/hQbM
HkKZfSUP6l88HyrDKNyQin2AD5Kzk5VXO/0SADAP/NcgkkGT0bum0ctaPenPaj+YsHCtPFljzDl2
y+LB3IDdWawBJqcNhkHbHuPCkE6QMbBEs9RCOLD/+2Pg7Cg6qJaEbltL4xys0Y9ytc6K3lUe6c6i
4g25xPreR7hsNc0i3q9Gh6C8C7RJPPtWNzgK3wRGVRgdfIvVboRy479RL4/M7zg3OJ2f8no0gP7n
Crqomn2gxTxuqkoeHwR9cFnIjP3E/ZES3j1QAulXcbpQ0hxJthFZ8KIahtlT31Szvt07SvDYnj7F
Yt2qI78NOzbd+3UBfUtqDFmWrTZdAAPdXRZom60hrGDaCCGert4iRSmwhv7xid3pleneh0DRG+AX
Bs15yMkMdRF4ty0EkgGBgN9GfDaN4E1r+0ayn+wyN7kaPHgQeJ3/BQiswBigIhHeZd5NWHd2ClCw
REi2O4NPSFWNQzLhOFFJjGu+hiNL28AcmvDlTGBwlroBN556KxXZW3Hfe9WG48lab70GXBoOPCkq
dRm1BFmpzEcTWDhJ8p+/2jij4c5blKvXVsV4GhCtjAWvWyc3Jo1KETBsbDgBN1KNbCOwlccMQMyG
uz0WN1woq2v71x37GomEtKWAuaTlFoE4EwElWjlnTlOIMPRh5o6x13bV30do14P84ux5cYpnB3kq
fSuD0xFvaYj4oA4Itcq9CImZwhXoHWwLajdYzwJaNcWkAyW9sZVyr/bKDpTeEK6U5Jj/rspPwjbX
xiXKW23Z/m7QwRhHMtpO5OXMOr+s+5a3gNsud/qkyRCLaEc/xHZF2S8Kt8MtXahvSXOwL9OgLfgw
wNbldh59GCPslJ/CASZYcx9yXAsiLK4jwTKxUtE4KcaOMu5sXpd5fZHmnlsLXOlnhrSTs5WL2e64
oycLSz8trI0rDitjcySJuA7V03EHIlMbFOpbH7mqZssON+jN8VhPE3rv8503MhPPixei4Tq7KHcA
Gc6ZmHsj3ncmTMytLPsJqNDMRL1uxYGralShOwtCR2WZn50CNgBegBUBgzXFsjRvjter5i3w5t0Q
9nORnR+p6d2HbbezPwYX4aBUG3ljyLWzUy8QH/UyFMekGCJQmCgFtt5f0LzhpyhrpOWTRRN2bwDP
0zdFJMTTOZx+FiX9JyDTIyiVncF4hgUK955zn2bQPmFeu1iP64MfVajX7yQMbNNRHxdMU/qN8i6V
WOCrkQx4FiMoq4/9274AFTNFa5tTchSKISUHfFXjZhi/YTgDHB00UUwtlmu3l0bs+6Ij+hO+En0C
JMyQg+FyCYECWi52tP3HWYA/fjRDn42JRxfs01KXt43lDyW2IQLhc+6jvCf8FxsAxqQfb7Noe0a4
dIF+4JLkWiLBEO4dyNuk8AmIROMfB+pDgkWUW3mgg8rXnNlm6ltYD9OApOK4/ueuHbpGtq3FOuNs
XW4uBR70xIBXl6MJI0jvfzHOmv2hWecAmA1GvKNX3UXvzfmHl37qm6jXVeS3+prbqqsOHC3nlceW
7DDiKs3ogFURA4OMJpDrGcjjzSnCuyW0uejt5HEr0dzxykj7NujPMOrdJP6olQmcVzHCpHBfF3tR
wnZ8/Rvv1b6dBcxStqehz1w1SjNwxl2pheRmfi85gi6d4XKJQth0YAcQ6IVtw6XANwlqqf/63CzG
xRQUqoA84XlcSMXDRF5TPXRtYbvdKaF4Od3br2Vq8Khurzns0EsTEbFiGGIZEqZSsSQ9KtBbna4x
1FvVB0rWoCgw5cKibW/mL21+RxcR/LpUyzEZOiPMjnDFm36g8Br8Q0sdvpJee8Y5NxpnKdLPfAs5
qzmd9AA933r13OsLFaXagRR0H2f+yXy7P9OJ09TkA1gIFTp2uRHuToDFGzAoVpnKB9OiA6IXzqyp
F5LSoTZHmwBRI90vEozCehXP7e4Xs/svkd/Gth/hRqQ0zPCK7Yo1Qw0PxHKn4oiseFvl8jIO1O75
pRGq+IuAEu55rPZcX+6yxMGjOAWkJS/6V6UvvXWL1p4xtEYGXKDAOjFl7WAQBzl/e9Qz2WW5f3yK
TzNOyiIF7C7hQSJE+tuH0Cfy4jZjJ9Sl6rXnnzg6cR3AD/jnSaf6rFOYcCP4jYgPux3U1xMjlk6q
cR8FkhflQ9UCJRlSR4a7GlYjbtsMzEGdn9WxMU/yhxqFOrIm++pvOEx7ZIzJatnPwHZMn8etFQxN
uWHIDj45luxOTX2KIc8l5cCpz6seiRwv8XSu5gtmqC0ye/VRidh0MndFkMSp9oNP+DDUJCP6ACug
dyboeHl7jIXIpsLxtrFpdh+iTfFQ7pRiu9ajtRPP335A1pYbsDe//cY6AlROZDVS76J7lZS6Pbvb
8758Ap+PcHq5tTncaa+1IMgdtLNUa1xccBf8MU4cy/i+FtS3b/MsLX25txnofYeQDawkdY1vIT2+
IVTRNzMIV2964w8wURAb2YZ71pDvzS0HUHV7/tnFlAmqvIKq9dYXBPIndXGuHMAOK/zzV8jbj7ge
CHpQy3mbNQQY6/LTD9WqLiSFDNMDSX3v3ljZyCS2LRcyQfTeQrjh49jx3oVUcE8iZO/A2WNWbknZ
kM3TEfaf/zzUn7L5Vn1ceyx/LMc70Hh8D+PeA4b/x1RTkOfg9H1BzRCQeKdaPgY2vwjq1vYwcb4R
8YWYNSFlt7RQ33OaKQJ8XJXS1McyOzTL7QYfIxX9RTNZS3uWMgK5MonV2wab8eUU5RS7p3aOA4iH
cD9nV64N91vIe4Ddh8dxzu9pjpiBPLzpNGFfdIyg3+Ufk2N95I5mMpVJX9o3wcOIC2tR4T/G//ru
UQKXE5M3tThif/UfjjbdLMexNGVNB1mldsP9Kphcyuya6Vv/C+gepm1rzrY2Tdf59vFCuYIRwvKU
aqB9Q2gtSaKlBLHY76IW7EkdJ8tRdPwMXDYX2SOWpi1h4Bv6Rp/bBkcaJP7sYKLIuz4TiMH1UeXp
FAXX8hV0aw7FEo/WKwlTAJ8PDLLaghrkKArUZ/bQzzpKIgVuoBFLbniAKI3KGNG7x04Fv/4QTyXc
Ueci/9Rnk5eL7NAKyEvQnahrIu8KF1XX7gFn9QibRu/yLmcWdmJ7MT46ympUEq6ADJXzMXJ/6U7g
K8lclKM2xu4Q7PJoeITV1kz/FzmCdbUGCBpZU9AQ3sE/1vtnbNgrF2d+WnOWpj9PzWZUeQEC/W/5
iOz3oxCWdxEefKb3JsHgyiy2e6VFd5wE0J579JPekxNNZ+pPNs6YkiXz1235vrTUBO8xkLQjG4yt
dHpIcIpaPC61fkUOs84Jfh04qZOgXLy5rJzy+xPGYRz+6D/ZjZWPYaFPKHAPqM2Ntse8PLsi8/CV
RvfiuNQcayFsgoXB1gfVsUOyHxVbW7gwHJHN5WMJFOW6kC5Tw55d4MqhEyZffzMq7H/mVumc9SSw
KDmn35zkE1eBNbcQz0ZOc/ntg3wDF6a0F10OlWTUq5qBV9u9jVSBwXyuTscsql/31UwXrqJ34CSI
tjbMKbHd8eRIsYOwGo9gb0xkDV+FJDdzSgL89EKWbt8rEJY88jOL5W3DlpDxh/vOb30HI1Mve6fJ
ZBOTjSPKhwb23ikp6yaU6X7GbrU76xgjTnbZo9sQBcbjSMzO/qwLiWUo96Zk0M8jGQiMEEHJoHrg
TvkuLVYY42ljm3c2O6aJPmy4unl3L770S2sCdf8pGFVOvIuPQ1sp7L38pNzfpY3lOfYiOnZO/qZL
FPZr5kgYhZ78aB4dBTBvGwwpPrXbeskzbzz0faf5P3dt9S+MXz3FwFf1BTnc2p29Pqq3aqirphXn
icsbfT5r5fpHOLJWWSoqxiB1Z22/O7rzqoviiP2CpFtAzn9iNlfDSW2k9e7oXwCX22n3ZXVRuKOe
gBBF54GBAFLpspngOe79U04OFCXKjQnTalUgjrwn68wfruKOc3wlKhP9lT6Mfkl7NFCzhEYJ1P6c
TsZI8qAOGKpxFsiGItjnv3YYuKT/xCG0JRtJa6OVhTKwUDHFWFmWKMHt7NBSKssdCqpGkDvRNS/H
KwrpIeCagCKoMCTwdOFfaaU2mDbI+R1oMQZHbCb8yMqPKiwzukMX5FqUg2DXMhaFuodv3Q1TtPoT
EyyuP+Fvj7ul3KxCYVBUXcoZlK3LTnik3OalwHbR///JiE5gR829Ycy+FwCsZ24HJ934gZ8Pep/M
8Bia1upbjUXW2mQluBVW8TzA8IEqEaQgQP/6HkMqq4+zxjlkHp7svwEgkpGmEDidbMxqE+YFbl+7
qIt0fqFQF8mZGIrTpxVgatyg4Cyeby6Vic3YGthPU6Dp/c4p1Pnw/W30hx0gObT+EvBnQ0T7lvtC
nXznHcPRlX6rA5XkfCxKBxVP32uvyYfrqtuU2a+dhS4paw9ZiHwedQqSYJi9fPEMuOD80Mp/MsRi
quyeZ6I4u+G15d2jVkti/kIioz80hPj2NhtQbBslYWNDIHWqrg6HDo03SKZIan43uWvyS9o88xm7
KxD+8dm4qO41UBEKQ1WgR1GY9LCCX3e1TY2LtTpXUaRS93WjooL8+wJU7AWbYnzmoqJj8DL8ELZG
Mc8hY3MoxEsgndw1G7S+yNE1GUDY1/eNnewPJbbc5f/U3xHB9SVods7N3xbWMJTUx5C/ltXe/RZN
+yXRfTpcrYxjYithFzbkXcCA53QYGJl9wUP4y/udNs6CVfdXUpxxX6IrG4lQXr80LPe/BWclXsUt
mwhT0au23QSlfDnR5qUdHl7tT584istJviOpIlw0NNIl4yduxHcjR79gUpPCtll2Z9OdJaMPxcrQ
4QdgCyFHhOVP8o+/d5JpmVi6lWkTCxBRCRHd4JHs84OaE8n64ju2/Q3lk2mruu9k885+uvYKn0xo
p7V04xsaN7ld2oZNNnHNHrp/zMSeHjOw+uqS3+OW6CEWy+n7dZQrnZzw3SQZ/Hh93OemfO6RCD78
OtqLItXxaGxU/nXN4bAOZ/UXjqny68gj2zi7pUvaVQZLW2xpSry1UoSZDsU7fkQAk5AUhR34qm+F
4s3pRQgUFlFCOwLrMw5n0XNSQRZyW0epw2MnqpNIwYUa4Rs7lUBH7z6lhXzd2fKzMQFK7hUOf91T
cFeRgOjOjDEoCia/fyGEfz4n/UyTacxdKEynYT1fLSB5Bfrmc9grsWaNZTq5s5VO6IhH3L7mnUfa
7hq3TuRR7YtN+OLABd+m3vO+nvoIcFGG4yb0soxqt2PfMxAfTjG/cxLVzfFIXEHLWKjmZ8ja3MAC
31lOIxs5RrUVneiQVRgPyRJx/o3jxxvB4I3Vy7J+uu/KntMM2spAvXpxV0CJ2LpSV4etdyj7nWqa
lA5EYGiOPT0LGThgqunJc+B7wvK+w127mmXsIiXgzuNZoY6dQgT4WAsz5G/YObzAjHzsizYY2ven
8KSM6P1MvodeyFT+oqFnE0nU6Pvw3dgoCt67pOqFNzsuY2uuuLMJ0Lq/q7GXGRstklQladXmNuCc
P7g9lJ1VOy96Db4ACVO3Du531zCWnWCqCxxz6I4SZafNJoQzVQXs8YrPDhrhRhEhTIJaYJ5AVEoj
JtGMRsPp8YOz0WgYYDxUyLsUvkSkmE7PcqX9I/+gUUi536aVgcgaRy8j3F9Uw11mIUK03c3Y6Pd5
ohmeNSY1QLg1v8BhWN2fRfuxtH6uI4NN+hXvpAjaoJ8m5vKiv8rrVUUAdI1B8IhyblRjfnSlajCH
hvQYmWGd109f08SMnL9ytZtdXNxylPfq8HnFlZWmHdz5hhdlXHFZX6TiY/pUOVPhAtsYq78PLX50
SJyAZN5XSLa8a85dm+qS00AIjzvMEoNK5tq0aB5mDL24g4nMdIsbBCHxblCYlcIaCKpqC95dBaZX
sQIoFe0ROFx8kajCq4pn/xyWtkjlixrzRZyKCAjPk+y6o4jodaONTvV10AbtMuZjsV1F1ZsAHuEA
pI3H5O0c9U1YsdiPxEXzcpcBS72+uFIcsW1MOk8PM410WKAcuCVlrUv5p9uK3QL07IyW/D7c1KtI
pUOET5DwUfvnmOXYz6oY7FePXH/Lny3numkcfJU5n/xRN/pr5BuDiizNpxVUyAJkxBdbkE91nQ1E
h77OjZ+JWYFOYGYyd2TxJG/PhYKNIdpkWOtQZAGFzvUa7hu0Oc93GXTJ+cEtQXx7gFAiTP26T5yF
M7HXJWFsyt4x2LUzPF1S9JBaK7sRmbkKl3AzA5t1W2NeFTnHYuT+HOCViDYtaoEKPEX5rwzepuyv
ilsOLhoYJC0uB0jp8n4U7o5pZAVxPGjcyyfCvhJuU8ERPWOR8Nxd9vukGd0h4owBCVFOGJ+vmbGO
CDRN6YxrVmfGKwzQvNj/4zgM0teeMdOz3L5bQdg5mcbV5QHB2AwSsJRtFyiJY1pzLMffDQZl+xkw
Y5dZUGDbI4NoJLYPeDufOoqTvGSIC8UhgPkDv+lTNfNwXurOXknhEQ4vPC/eKYapT+DbtwDv0B+a
228DpBGqclF1IBvIHNi4H1t5xpwQR2jmTpgJsGOnWhvPhPi4i/NdH/fHqY3SaYD4f64agcaKZofj
2BZ10vNHJUZwVmKWegIOM+JlAEG3l7v/PB6F1kyPoW2vHqrJSl+WFwpF/dT5zgyZHBedzRzNdVGy
TFYA1P0sdAwcozu6tadMgO5TIU9mp2leVRxST4MknqqGsl5EiYt0az02cI+HGN728dc2PanmCVyA
9oqXBfgSU6sQJUXdvS0LlgvQMxSu6HSCEgMX6ulsAPqpI1mVcAUd3BSd5d/a6Xn/QiiZeTluIqPI
eBNHJejhbraL9tFcK9l73+jcEd/JT0W4MM+aPXad0yHQNb0mGY2k3YonFT6BhO5T6D739v+0k1r0
ZOf7u7OwG6nyZi8VUdxSM3J1S/zq06pl2QVdhztdY9Di5QCoUArszBR6T70JtT9UVVo+fzy6osZq
iMShHIxlY/bI8XNqKcczVzAEyl5qZBwRj5k8L8qipgBM7It8Qvrqq0/ow4Sb05oEPSJTnTOx7klE
XEwddhhPoJtm05sEyHWtLAL5OiA/QtETUSlAGwlbh0RPl2VQI8uCiVLw3dC5O69FcLDt3s8FgFHU
e/Kx1UWnF7TMh3Z71fC/GQxr8RTADhB2hJAonHAOcFTbw4cKhSaV9SR9O1W6naq0zAs+3Si6yk5p
BQ5WchAXWvjOyOK8XNApDY/EW8H1MTPM9FKS1A1FJZ1DpvWSxfwLZ+aSlTspg7K2GJE3Et7zO3C5
BFQSCCRgzlSAOvBCHi311Iv6GdtEif4MlKf/99l/4p6BrViBnQn6YlBJSDdBVeUFE3jgngoXZwsN
rYEf0zFY0Yf+m6iJ8TUF7mc8FUs9L4WrZ49ERAuSEILL5+weSBalJwDtTbJTit6hTKE3e09wGvrC
mfcXTVm4wuBqq2S22zCLfSNlnScnpNy+U6BzRpkrgzpGB/fv4f6ZTYDfVA1GJakF19gTC9XmYubD
0GS79rKQmQJMmvnpghEJkkqY5YTqJ26eH+FG79AdmgZcM0SMmHBIHuxp0AXs1RlfHtoMkxlqzhwX
kS2kDrhjD9gNZBznbW0gOUvvyDI6RMEw1rRvDsu9/+46Xwg8NmnvmfMlESlKfYe6mG5kPmpIHrs6
10ZNHt6L6ywULkKkCZVPp57W6Gg7dllCBsSBWXzfVPfZ6DmZRtoHVDnXW1gdflxOtW84wecx989N
Lve0PHW+JXL9w/dlCniUmjt66hThoyoD1BPzqZ8rYrdGrl93hZRIRJsReqKrJtqVAXGuoF86VumD
x74xkwadnOcW9cHZghFsdJh0818PBXEUmj4rzyMKzp3q1XoaCxAPCfGR9XNLKam5esZGDRKvX7oQ
U/G0krdbKx1cbzEWPT+G7ZJZJR5cVqSqHR9ZD29R6vh2tpjL7mgMhbwOZsGWynvNgGDNRQWgNelZ
WPW1aNCxGzI3aRo9o68ZfIjoa91u8x1WJKUMmhzRv2KVZUOVph8guf1/zYzUT312KdhzlUJIHKyi
F8vdffLIqOlQa6qLCTeIGPXlwVjzGmYtBmeR37U3ijdWEMguTjGtdzeikobhHtSHxaAARLmBexIm
1w6ZBPHLhkyH6PqHMMAfxMy/r+Scn0wuojQlBG0zBRBOXtip1kthAMaNTcAQEQ6ZdtxfBUWYQThh
XCWfkeTf7CfAY8ORyJ++GQY13gJ1DB7VgkSiEzg2XsfNiFAoOSO9j5LXpfa13Xu+NGQSROeO1WUy
U84TssEiVbDaZiIEtk/pOsDZIezuR1fm+HnipmFsX1VR82gJB4IAn246bhpDHTlDMKfQ+rG5MMf4
LhX5XyUqVd849n0FStGBH625oAmUB7PJB60RSI1tzdZdw+rNYUGsJpBcgkZ2cJNWSv0BflNqXBWV
Tnq4EjHq5g7xadXFrWxnovJXpbznwxs51b0vx/aWQwm1O+09TLXNS4jyqRYv1TznItAdU5FGlf7t
XbFy5yO7d9mu72AWZcc/3/HS+CTKQYJWwxd8a/vWNeL/23xI8Nh3zYDpOJlHmEKThZjLJv4pafym
gJ9yXzuwtMBWXuMECQEibWcZsPxqaf2rs5PvJMXaU6WxnPtFi6wTyP6t4EjOFKVPdl0D4ZOH+H8N
CbeCwxc1Uo37K69ODRmiblqDbd0FU9Tb1ZX6uZD1wYVuAE4Ic20ypAMv29IKRVk0QIhBYgWiK4PT
/vCK0M339YreGGfJHdXpDOoKAO5DivTJd3+9ZNAwI15pwqI9StcQnm4/gz5MP6Ba7kmStDgmhzh0
BhbUsrbCIAOkpBngQHxo0JND3VLNVkspj5q80n8a4enLuQNIcnzQhSPnoMvOIl7XfXqo/scGdfAi
Q4r95mGYsITY34c9Oy48jiGVzdzWGntS2ql+WjZFTM4MY+6/zqe992emlMw1PDpSnzfHGukGbkm+
YWzVjV1ZXw0y+AsIuQdY32taYj68d6snrMMGzwCfnkRFQXboAla5FU950aGzEFf2hvVmN+/HxT6Z
eVAfm+ytvWQPHLo8zVPO2PscXjiNegWN9HbGNBz+dIe8FqDJPizmNiD4g0U7Hm7216+NiMno7xGH
KTL2f/BFhLvj4NRbRD06Xbi2bkTVd45eIs3eNRmCeRRV3Ej8KYS8a8FX+iBJkfI4vQSTuknkmTZy
ZYk0raRW3SNH9vegCOcNXtK55NplUpWwtDLlO7Y3mtksgaq63na6AE4bOKMTlM1Q90SgBvyhrw9y
sM0wbV9O9kiblVwPmBuLEywRGCUpEi2da/sj3tD0/ondMD/qptCECwR1fMW41VtAxhajiKbr1g7f
QyUJQ47hA3qyG/6Vho39lynSx8hx/Gg0AQZkJudwssG+O/iPHfhxZOPHdbD3VdXI9H0yOXSk2Oog
pRA7k8HMbGhSx70RaC/Wo96JDSifbHnp6J17qc2Bpf80ITC+utGqda/n1AROyEuV8Hp0JswJva5+
USPrikO9c4wS0oVyrJtyalEF74Py46mQJjlrU3qT43GfPBKpop4j2COz5SGiPx2HfvQ+snlcDMXm
+5+2lbMHwKgWtjMyLBD/AwsZ1UY3i/GH3FWUQW5hL5BRRBUt3lyYIvGAwHSg/vFT95rEpXlRTnph
xMNtfOg9SsfWMCZcot44tUEnJubtCVP4ia3eeSS88wY1lGznHH5kcON85EX3d58bnzZthiXy3BqH
sx4Wkj4vVZLeU4T+xbE4qyFxLyt9+xIiRZLnpk+fRxMz5gxvN9IiDqihW6vXX45gc/5O3mh+Av5B
kcbKmWN14XspuQwnsXfG/JJxmgDNKKzMM8dYxatsPb4Yhska5vjT9PsVhmg+AXmo1v0rpfkCuz1t
3KA0v5IU/VoWR4bKLmMZ4N7szNBJU9UqMWRWzbiPCLmkkdKhDP5k9hOrMzv7RNNbFbkdyJ6y3loG
NSDSbBI7D2c4m9ChKaFsvLz3r6KSeW5yBidD34VGztMquGHSEHkkHwuSCrr5mZn8guaxty0wZF4P
YMN4lI6pRUdYxMISDmUkNRkmZZ2nLM4sgVH3xVRhwkSX7owQk8Rf76f+XAI4ip2rgfRNu/Ans0V9
D9lCaTkpXwFPSzSRSENdI5pezLogtYGbWWa7+LrNPFk8vOzEfF4Q2RZtZImy0v4bScLBVY1NASAt
6H1AjgNDVOwa7XRXW718OmPkdh45QowdMKxL7xrdxu7M46AuumuwkizEfJ6Le5Jgjk6sYlpN68NM
2derHPYueUyPYfRsAVep9ZJrJaq0IJpggUrcMm6pJ43YoiFmqE9+djtcca5av8UI0vEqmvbF+cRa
lguAwCgmL7IsqqWDdT8+1wfO44dN9kiyF59KiRrgOI2VkKecswnl4TMmryBbtmfdvt9z3G2EeBQG
qMeoUKgvZR8n1mzkRAN7xTV9bPUIIvTvfX3WYYGpkabMldJz4b6ce7RSqI2z0InxIAXVwonOLN59
QGnqP5dWkeTfGjEAspkpyApYS/8m6jS/WdSwb5vpud6n8WuzUfGwwbVf9Et8+6cnFoG9VA/OFDU+
naeqeAHOWE4E4qtpywaDidKBW5NjDO1xdK6V6ng4SfQzztQhs5MRLb2h9Egw53FiNHdJveIkUYwt
2pjMfa+oj2z09EItOEnB2/Wqd5YQz/QEJLXy40h4SWOMF8xXpRfM0RKJle8enQN28sBB9F3v7aVL
SZvXPJ7PB0l27rH86h9o9Z2P7Nkm9USF/V+CVYmGUoqijUlQi8CNSlL/7qY6bgSxDuKkG15lpOPK
YgD0uQjgPv2/OxIEtW7SwOIUtc+iLnVlakxlLO93ETKNKgH657wGG1enMto4m5qy0EG0gXpmzlBZ
HHbi09oqOjJxcL+NSXaC9m5OGGytzQF3ic5UosT8HZz+tUq6Q2iAp3SbHYNez1sILodW/5NvHwHi
oXcrpMZuLqhPMKQPQ0RTaziuV6/vTsuMhdpadDkp/XCmR9wLcv5Sv7Cr7YfMfq4R3ga3Hf9uM+di
SCCF6hwFoAfuaUxJNMxu8ZQvnpucV69QqVGNPlZFlGoBJH9FSpeW3vICUmLd3IK7NALSyJCJy7OV
LXsG+D7P4rQrdJH7GOi/XaLeDC6JtHKB2CfSO3X0lTNfkoUiGvnSvw7w0Fch4seuQrQ0w+uGHf9L
v8neXMEoRt5CPYTaCM0AokzRL995uha79SSsGWpCQAaf64nZwdKOYpoqiZysPIjBD4QNi3ElPrib
TJ2Gd3I+n+PR7NHy4g/hIebcjQ82LI4gouHdgK7/VTnb6wG2vJGF4XKa59xe+B4VSmG6XUGKwBTZ
MOhV4Kt5mTVubxpKblMR8t8pl9CR7nQmwofoQCgwvlHOzBTlh+NSA/7CzRKuAXI+l57XkrqmcG2z
YcH103dFavxRXGKMxVKWvpJUgP4D5ydLMU9lNMFvgxsTTPQTS5NplrsbKNT2YuHczzP1JkJeQHGB
mjuXwwTy/rBVjAwMpUDLplxJhr78odltv6RNJ1KMlTpKHpVPTHlxUo089JYxNEcEbspJ3p8yJhGC
fdRGUZfQe6ikp5tJ3Wp/T6CAQGRkd2zdqcNc3mQtzWv7dPiPIQwUgUKNAx832BQMGiBBNoGjjqBW
3LwI8hHVTb+vcE3dFJlDXO4hxFlB+Za9tJx6hucLezq/xBPAci2WKMvyK588E962E2Wd5iBmyl1G
bptIvDYQiHvQtFGYknCLuADLUvtdSBIC02snnALImGzUeXkrc+vawn8q1TbYGDQvZVhcWxhpFYiF
J6XBKAHLMmgjFDJPPwhOCY/nvvhARINHl1V6rx7gvDriV6fw7V8D0o2EP77XjYvlE3UX/T9h9Zax
zRA10PHyejhja3s+/nbtJHK4pBoHn7E05NzMPhHy3V3MEuwem/rIaW5ewP+b3891Zc+TCLwoh5H2
UONlyNfUMQz//lxvQt8Jrf9SvDvbT59miUMaZbIDJU+6RY7mAyA7p+VMQSV8QFmHzKbdN/kbfLHd
9ItbTHFl4nwWsM1hURxh4E5WJMYMP5NCk5GeyEjBfNxUQECQHLgXNc8o0OzGTq4wcdXWK4tvA4pe
DsRZ1X66swXV9B45Fj9paxhFLm6e9GVfjQyfkjlTNwl221TYDfJeW0bFg4shrxDPBHqLn3Bk1XHJ
/QiEA3EH2TFy3lJuH/yv2cCOaA6i4kD1EpYjD0yKq+0UhzP1VJd1qy3Z6FD1vhSXLNQXAmiOYms+
xSWQ9PRYdnKeDY8OKHYkqkBNWNIGKcMTpFsid6JQHDF9lkHHdM8hU7xeG+I01n5eQ4Ds3tmaG35b
0vHtv4dPkJa+fg9rbWljy0mh8K9waKU0XGV/p9j+l0EsOxixen17rf9rMHpKFiKwgR+sGFdd3EKF
6+QdCN2ZUsZ+nS1Oect3c2Cg78Xcv1irbHXtg8n6SYVXXsJZaWHygLu2BpvrLnsHP0ds7dsYODFp
eIzpcKnFpu1O6jKlEGM4jGCv+LC3elmgTUBUHalfPRJOZenFAQrQg3mBWVZPj71ViDrWSQP1UET+
6lMXTW4URXNHBRKLJRZEmWKhKnYAuaiukUz6Zolv3xAw+1bOfW+MYa/ItEvG0dc0kjy54xQcIPlK
M0c6Hc2T+3iFcVtUZW3wK6tdXquRA73XE//zghrKxU+5RfTPKU9Bee4FUfc1MygegAcFXIcP1VHe
mICTV35DRtTzGH68msh8xscpB86IOGt6Y5/ogkxfin3YvEo8VeEiuZHpVSslQGSYp6gDeANWR7BV
Ojd9ye9+u81ASYJAZ1DmecJPPKxlbfwWHH+tS3Co1so10P54if+nhSS/vzqv0pnvYlrqezLrMZ5f
lvlYm8Zw7aHukloLY99azlYgfsW44QOK8aw+93yemsT3xsLmNHDHMxwzj0YMfe5MN5P3wrrizqJW
G1GEX+RZDx/lwvQ81opM+xUB/8M4uSEsbsZtN0gTz2OsL3/cO0owgD+csANmz7tdSCc1zErwfhYt
Y+WfgOBvTWAFapL4YXr6Qs31JDOBafCA+ACMoM/8l7mlfEVVKKumlBtE+dCH+PlPUlZVvG+gl1/z
ugjDRSCBBztST/wOX3U6FSWPDHdGW9Dr8v7oYb0gHd5/JbWYk7+hJkkodNhUnuwS6wg+y53ufmpk
U11Dsh0zpXrTRH9IB41R3M+9GvBrH+CGvCIenhLtiq2sOqvl/n8aJyRDlElghRzujrYVzp0Avo1N
XXII8uQLI6vaqTCm+iX5xzCh9Schr1ZByKmI3hc3AlqVGAdvGXEYKaLBdrN+O+4TlbbMDzfVK8Ed
w9avZXthfdodOY15gwZdjcCumYvXmaXtgv+HQi36OaDigXaShPAAzOvECMjL6uWjpBhqCySnmQpw
gqMOJrVJ7u+/C/pEBazpHkKweN+hmJarM4GRzuB34TWQ82zDjCvX7tSYha4lRqGAGfp/h/lFKqen
/YGociQGrHjpuQ0o2+iDve0He0U/SEAewMukfHj7bw44bdLUeIExS2UNp7EG63eOxIAGsEDGaNh4
F8P+BDAsxOmvk+pbB0f/pw4v+/qLZPWjp4/9prz9s42v3x6ZJ9ZJmQv5kxLaowMkQ8p5oqHzvUrV
fIRYn5bESHrdQlzp4vPFGiC+pjyab4c3QLmUYImo2YkRU9dxWHPAHUr6SOCiyrNxU2uqvKRhzhZm
sjkIyf7ONmFPjczsPS0xcdCwrSek1q46Pv7eZiUOlelLMTEgLg2VsX6Qcsg2nMkzB6aR0XLEDDUG
sjGugBnAYFwObQGJFboz52SAB6Ce9h1REoF2ujGiCrLkywV1qY6gtntf2Ymb+1lAzjo8lBYoqOV3
zmtuZ6S0DtrC7WavDBCoxH/ICj36QaKjexn0cEbXgrGBcvbOUeWzIfrICYoOJQZMDv1QE2KLpLhH
X64r+0oiuAru8bYO9YEBNZTZLEFpXxRZw6xZNRGsZoHJuS6MD2w7jiEVytJCoLOJatzBvyVA7UOU
b298tqjM5/zy0m5IG4464kLRicXBkHteR5X2iCzFe11C6ssiZ92IL3++3J63+1mBqsPmAQ53LC1y
EpLdfwDXiGjt1SdCg77gonpk3He78q15UzV5BiGg9VSjVYWeFUcaEgRsjE8zLoh9LgmmfhiUaPqY
2OgtlZAtdWJqxT23Z9Tv66WjNUx+dT5j8Q1D8Mzg7GoTQgIVcaVabGiWXbqfSit+D1BFcalFpXNb
qlaX32TpMDbCeySRg28l3bAQ2bJ3tlQh7iyS9tLtD32/eCeGnrXNc7HGSllBBX0woU3A/Eh3fdWD
xR5IQ3wKm+2Qy9hatKEJxlmxEq0Wo8+K2N2V4RkTQBgVk+eusSQD2xGEV6GwDyLve9y/lZFntlrN
ZaPJTCMzH6azzzo93z7vUFqq1fQalQgjYARryrj7hLNweSiIwP0DH4PdGDR2Nxgy0C8pWW3tAyqD
Xbc+DR/aPTINL/rohLtgF8EXaupwp8QwQEh1MU1gEydp4QrCwP8TRXYqnxgMyqsq4fWaQKl6wPXd
89WBuWGF9aXFl1HfBA13tlMllkmBWfkkZf9cVQvG1/KmGSVBl47HuVHYvCjrX8GRaBZNWMj2htgV
nbUsUOZ0nR545ePdPFyIaGXL5rwBvpfBdZ3JgBdiGC+DiSm7GtG5RxjTciNUosCXAamlVum3ZEtQ
oVTDk9k2NWISfbXCvBM+tu3lWgN7xPjMp0zsmiEBHdq1IF7dTTtUtBMA7phF3MeBgeJODGBsgmFm
V58JULXbf91y+XIa6tjp9JeTnZ152ju92MYiFzcClBiFtIXmvvD17BErMgLBky+NDFydYDaKuqGY
DK/dDPcjIYha/jdwgyLO2ExT7lyNai0fHZCplvFIGlo0R3EvvhNMneRYYlPpj4pwkSj2Z+2ECiuv
bViFcAnjENOnkGSp39By0owszHYe5Xa12I4C8hMVUkd4f9MrQysntXINcLfoLw1it0qaSkKL/MFd
d2lyA02nWA3Q9yPXGTY47LY8ma8hasQG/hXShzaHepOLgAGVOAkgYx75v8jxD6BtCXCdo0JXibkK
6edTAKuHq/yqfppHQmJpcGrp2o7rDs8w0W/gh1yDwy84m7lxNzup1SIw+SnT06Yz6SnDjSIFo9cE
t3oW9Kuzl46GDfncrcxIuPO7LAd2W726o56pq1aZbtZuxEae5Fr4f270ZCCVv02KchqSTjH/ZpGE
wTmmp7YthB3WWS1z3owtNR+clYKS26ZQUPmnFmUkdZ4HOVvjKssoNX3tXW7e1LmvKUtPcAenP7RX
abiTlsPdjjqsLDM9ngVa5Jfs3shOwKrC22qkoT3Ey/pYRgLGidWrH0IdFZCAtSIDHp/E9YaRnser
Zbd+ieRPAvn99puqVTySHPa1tl7rZCv6hu8q7fGvR9/yIOr4N3yABpnv5QLEgDgssECr88ij5uw3
T3Thi7SZvnNaSr0d+KsHe6/QAb2ByNg6+4NQxZdg3dFZzLNONofjuxqdjcF+kWCXTdyqM0uJJ4qq
eTceIR1qwHAECT/qQidtcm8QCaIsEhMmjtgRqD28epzlXVIdCVxsylZ/wKWsq9xi/G+R8Oxd91WC
IxiVPMigyRnXMP6Q/npwNq99AxaUMKiyd7mKDPqI2LM3m6ZS9rc+zL+v/fxneWHoBWcv5vlNqcWD
vj0atxkqgjL8hL95Q4q1b/uTeZGVDonj3u35Ta7h6eWwr5GQvV1Neg7BIkSMPz4edmUAll2XEHUX
9DuRttPp0e2qDipRlHQfVCij2tBZLiXwc3mYS7/c1ykIy+fGRMHpMIUj+iWs53NTmE6X11unvJDV
62+c9NYmCbHsLoSkQa3vcMPjVofkVU5B0ACoH3xNM8cf8qs7HM8//gCXKfOxVFrkxjI/pIGMn9kb
h3PDCCGnNgBlUf/DQVaUfjlSc6c51ZZbqvgh+evxIp6dfm9yCxaTZ2RX+w/bkgSpvxXsbbTJPj5A
VF5IwRx/BiNzQoL9PhDnUZPk3RehJg63yOvHlrmhI6KP1Oo5ukPIusNl9FtcXc/we7vSCnEMrOTF
PYWMWghKBcjVALSR+FEHwg/pBUdTC+lTbL46yXSmm1vd8zs9Y2vmJwGRif+4SITt3NagSnZCzDk8
2Qtxi+lI2n33q/aWDbVa9Zg+pp7dGVDa5NI3raJUTlPAqk9qSQQh+tm0RELxcwBMbGuwhoBh5OBC
GaabSBU+XBePk0ZQczvVHZfKP1BJcmCwB3ameyvu1Ed5tc03bdyauv5P2DjvX68jXTDOnajCFFkz
u6L5/PfhH0+yWyDwF8UzjCB7BawXNUsdGMR9YhhcBygmn8qJZ3wgZVEYQ/rG62GRq7j2Awo2hcmo
33WA2TgH1sD7bwvqLmJfWwmc36DoefqBSFHg/DZKOelNWJJXpDN9RlA5BnuPpoKs3zsYvNKvo8Zk
nqGd9VZepRBhZIpzEtisWEsLwWgGaO4+Gc/n/pB6Ojln4uZLIHf9LPNyHiCpKKk09ChspuBz4vxO
AAGTMoiFODr8f5e2N1ChAksmb9c1KOVapA5ou5PNtk/H5bSNIrfdVyPTRZXzQ9VgGml6fmo6E0V8
5Ps3XnwdNitztSoPk/R8QO007UsKx4j+cIrTRmyFf/kW46S/OD8R0IBRAnnGmDQat5kpGmKRIq1m
1X1xqOaACNzzMWqQ6XGF55yuGExrNTKSOOcoFXtjadqOPk8z0l8ip0lwmysJ5tAGZBMjJ78iVGNA
IX+/5hFIFDM/xAUcJ/vkaBxSQznYJ7hoFOMKeUN0wbJ/xdszPTQwPeJQrVKSgmL822RMhPaxt3kS
BRaPSzAr28pvz8deMivjXFNw4k87ilru12K+R/t1+qJj08fI0dK8hoEqwkFZ/j74BbJSTjPDk1YI
eSFKypgJ7i1q3kBpj1qItWTeLozm5b/u3oeBpTwYS67K3rxI2iIUuspyUfN3UE03nl9zIswT7pGN
ZZUm0Ac1lQP3lN36vh6N10KUIzQAGr0W41dfQPJCHimjrfFUCPC9KpseOw4vx75WorFg7kr+ldAF
ootl6bqAUHn0TiDsDElBnH/t/ccKIpjIelrxbyHh4Z/rT7sHxrf0ToJ3CxOsB6ePdlPfWYfECG97
DtjbjyB63PkrZyaur7m4P3etCOF4Z1hWhUQEh6q3f94KbNuLmX/c8WfVgBU1wRzZ7uK3vQ+oDTUR
EMjVTXrbhYzykecxMQSx/jnIiJ1z6m3sjUGhXjRJ3ha3+HxLqW12XrGKSvXIY8NVxxehXWSOV9fd
yHpHcM9RENwL0T6Mo+cU4nLmEb3qCfhnztseIg/lRZlwEtALcXDge3bNmi9Un3JDSmsf0p/Wt3gL
1AqEtVSDpDTgoCfLM1ACQcPN89d0u6rxSFa9cx+boYlrs+IiLKCUeB/0nxxf1YwHbUJ0kk6AjEoG
ubsEIjiL2otF6buTl3BgAixqcBvtMATqiuZy/VPStCvxxvPhG6RDZ9r2f5Hu1clbpr8EYom8M3Ch
jT5oA5Qz/mqUVDDxpIeT6Z1CV5RMGATenekmK3TsL0vzONgtGXMOtgA6BsyGdQ5wwha5L6bqQT/g
DFq7J7+FJ9tKeK18kS72RrOGcGkotOMQ2rtnsiGXF1Z4GNDoCyG19nBNj+7veZ9OAPGU66Bo01Qr
K7Sk31l1tzjcwnp6JvcipIfpxKKECwC0tfYv8kw6elDf4sLXP40WIyDS3heWKFN5YQbaTsHb7XDP
8746zOy6gAfAe7KoMo5LMKU8jvXDHFSDFnknw1H0+1zIYCxzMWRXrFwzOHare+ujdVS1CefJJBGl
cQAFCkcqmbK56JiKRyp+mf20S3clnPsOVNUW/SAoDsdjEiLLuX9arYA6SayX6CqGz/PXJj5TVxZx
OcfVYLImmk+/HKGloq6Aa0lt8AF5SuzVFOJ27qoDjQFt3ltiug8sF9HE6EqJpjE4ST6Zz4WyxMjy
mLiQ7xURUKIUaHiImPCL8oueZX3HtFp8i8xssqa4vt1nczsfZiQNg1IsU+sJCHOaiD2U8jCayHba
Lhs09cRswkcOGYGzWHHw1/Y10ISc0U4AJS9TriSNZzMBh6TescDXVAbcXJq54vEkQTW+98cD1ofv
opyaT63jrGV+0ynD7pFTOmpJHkWNDLsW9gA8tqfV0x1ex82n0Q7rnATjJBrz231fOHnw1nDwQfpV
eFUhxSXaZE+w8L95qCjqCAhSoMfViz8jHAElZObx0bs+znColQDUkmNg0EeATYTpVkf0qJbdjBwx
SWOqOh/A3bNA3Icenak/jR5AqxpSL7bcSnvtpyHk9HTBSUhQNB/yqknNegh9DzQjFwaZamSz7iJl
kFDkDxQOLUHHDpuJYW/OGsm5yqL/N1F17SXQc+9lkq7PBBI7q9aN1G/EY9TGAbdUpFLvhN9DHiMa
JT366j+QtsTy1uXcmF4kzTnBHZ3w9xftW1YgECjYXMV/bEFrtcwxK0Upl5E/LOTMGvtMVpyM6Qzw
GqTAo2/9WDIRmgftVBnmRs8y8YM5pbCGt+DjBNNIbVeJ026w4GqcXoX6SPYbgbF96qupDzYnxRtT
bqo9XXTrjQRKjsOue6KdNj09ZykcJKL0E13coeQujCefSWb25AHejXNmdMTML11V4xAPQLAKUrcG
1Rg9wIhXlSfPo31+HS5TK5SpXPAFqyb/Dq/wNgXuKFc1ocMPR7dFb10Ja72FzkM2vq3WncqXRXuO
Zk59jELwz/B2wA0Jo7mnawhC8QH1obeMHTfOy6ki3FeYPrglRt578aYePYxe6cau51eI4WgJQo32
esVve9DDfSN8+YMUgkZSOC2OTSAnL0mdsABBankZQDx3SO7MtaDMqh/VwWJ9V4CfWc9lqMdHBTTN
gCxVGEpaHzM7f4OreBYpbI5pt5znl2nOlykKzn2D+7FgNjC767zJr+Y+i/l91bvY8mdIjl9wySXv
Uh63xsHgcq7KobBnb3ybrnJ7TRmGjIQX/fdV9ft7NeolSx8iG+DK6ZeAfKdDnqNbzk2n8HJnKvd4
kWTWXaXhX/GEvG3pYmxDSNKFj97au+nvxAe7d+A70BcjsH7OUlL3bqp9K9vJ4oMInYJ2xm1NNAJo
wAdKAOFWNPEy+MKTr0w3zcdCQIrPX/ioS2lpFgtVf4oEBi+SpzOULwo32aAfXmG98vnbhdEM41/5
uva5iGb7YVhz23HIudfnttNmLUvt04nhUMGgEMKyYBjY47V3hBE36VTBHOlrirZWuJQGnsRUScO3
kybNrk4AxOBG3yaIckUIekaY/LESUOjp67emLx3V/2JPi3KHgTMffgNKt+zrtbg+xYgdRGMKQzd8
Gfwa/7acv8x1zPszSRLYSlbhuUa7D/IFKdDmQYJ6sPPszIgHOiTCN+oc+QbA2mr6U1N3wJUUMlTu
IRagXF+vjwYgW8LGpKyU/BDTKovQ5D1za2QLtWeg9wq4nbBkMiaiMvBUFTXzjNUjtEQYJ6krBsvm
ATHjooJN5H2767Un572jGdxFnBnzrhlOUAQ6yqJvDkcPNPqc/+af6VnIXyKN1gkoIA1UacRIREjS
p07Ma1jUmBNr3lVZrXLoQuCYQQjX5pA9TgqnO10Ygupv3+7mfVeA6YOCpBbCNQzK6LNaMtkLgwB+
mxGURoXL/vd2D3RNMo63h+OIZ+6n0ZgEqWBDMyCH7JzsKw2jPoXurJ3CwRNjc4xNT9/IjLuckA87
RtdDXiLtS6axbWGVW90ZRo2fbNqvgaZx0FnhISYvxz6VVMqfRlz6xUvTTFEj+Lkot8rv1T5F+K7j
5pJTQq/JVvwDh9v9QAOHUvoiBOyERwm+M/zp5Ww1Kt2xMQq4HG7boVBBegHeYJDOHrU2lxQE/sFo
/s5wA/URH8PWuvxnEdKwB8jirC/bieEmxJNyc9QxJ3wgQIeZDU2fqijwdWHtZgqI60uFiNpGTSHw
OZNGzgPzGRInMFnYfS8Cq4WZ9gphBeULGbrWJgpbZl8UNI+yOjIEjFLqbO/E3AGMrwmZWS7yZZW4
vX/BLeiIsVtjTnsK65ZVYjm4DsNiHZdDAzQhGj5cxqX6SV7WSgY+LqFWWicftvm7Lg6zgF9OTIoc
MRVFxRz7AYUBAX4kIGqmgYOnkPbsveLKCYlECwMfuSgeS7AURF8HwE7KadFrVmDYMjREC0xne/re
6nlBhIPWBLOgqfAWIWpDX3lNeuP55d+a1rUKIoK5CuYUhKAIpCUj3kpV7ygaCGG+nNIGF06BuQS7
kPR5f/YK0BRJeHMJw3Ti+MxkJ5vngGax/Hb5IR0zslopAZJ9K1LTesWlWHdXrcFcRjgeu0j+WTo3
z97Kha2XC4CG8Pm0Dnk9aQsPd5Qi7dE7vYH4oyo8k+cc/1Pd7fA+hUWSZrnbuAACILzpIs9E2dpX
YIkjkxC/mucsvKS1xPokju1ZMI3utNOfPJkheuqnQ8Q6fCGzJTN+j564Bc2PpoFliLh4VPcOA1He
5Xu/K+lJx+Ma0G7NZXAHA7sHV9+5jPP9gp+w02f5Uk0hOlrIwhCB5SYui3G19dlDyrANUMJUq35n
hVgOhkUmckDxAMmP76ki1flvKA/5r9+3XKovCPuJtG8xY6cpO0De22RxkkonwTl1rPmUDLGu7oYb
1iY2UcQ+YIO4Wf1sP+CsJbzjIHgh60EFTAY42U0gnDOSI6SRDHcsoLzjMWLC1MCHcne+ZXUEf7eS
e5HW+de0qIeqPvlHu1oD6GoZmyZt8VuTCGxOjS8+Q1+afxQfsgcscdtR6YSx93f4Ad0dfhtfDem/
XUSqqPK+EIr82ydbCV23M3fNE7rJo+A7JVeBJBImEuuEsg/pe7j8kiaTQ9Sk29BkJBC5bjRLYkos
3O1seUifYVSgOIU9PEam4PxCPBAKArkfBBhzWjF183wcp476v62M0JpDyUn1Hev6+a5Z0JvZE5vE
H9bPh5xeEDvaNWGUE6B+Fuq1pwnDdsV/WjWUpX4X6PPEt7edc4d1JpMUS+C4v2MfCV7nXNfIJi13
7MeP+rwJuvLE/04YonRo6AXrGjzy2v4oC5UeT4Gwrkj1GI1VJFrMIYAl9hRxLCh1NT0yPtmz8VtG
uHm0ifPg0aTyvLkXU7KK+A3UWFnjT1nHIiOl35nMT6fKamCvjutvk2i5yZ49tShagfVWTjniaDPq
yRFj/gpbaAytWrjneEnkEGSW1wcEgdtpOc5QKRsvpUWTUu3iop4IRLvjbm5rjNCrSs9sJDQNbicE
ggC2oD59jE6eKGTyF3MC8pY+OhzwyC52Fy1cDPTelSwFRodAbFCPKEAxt6spKATcukjRUst9tFpk
grS0SMed4VVea0ZtW42NR2tAb6L1VDgXFy1KkHtlHl449u3xgXeRKv1jYQCpCiSw8tcojyR6U06n
m8XeuErD4vp7rXcAzMU4MQdRUgCcKGpSc0S79Rxgz5VVQo5xv3K6UXvV0VxG8KHAotf7ydlk0EYw
mGYXSSLIYV4R91ip94BXDdLuQLhhziVfrFO63mEC+CApQ3sQIvVRzOfJomgQO1lc5O6dJeYINNOT
XlL2RfoLSFeQdQ1phwRr+R4kE1Q/ajMMiz1Vh7Nv3Bsg2TVEBAnz4GnH1btafUv80fTSRIQyTWKJ
rH6N7DGWSBYwbKytlXvZQhEhLJF2XXLsfxWCdTHeVai0vhk+bSKmlRs4Dx1D652T99jrqE5rJOJD
+pL3VsBWv3gCnNrtnMMxb6eq+2nvD8rTKXJRBBfyREdCH8LBeQ/ET8NTgesDoUOC097KVX745pKr
Af20XiBinaYDmTF3b2qUpjGAe6u56MbMTcSbde5X4IGeisedrEBrJoElBIEG1U947P5nIjOozRQF
WoOV7vWIXe/di4rH8vfPGu/51+5dGUl81SCCCr7GWiNhplSf1TMqudrkteK2DSM4Kx55ltKGMT3k
dZDBgydJqxpJ5YCelQeZ5bY0nr9+JObvkOZB4i1EFWFbA0rO/siX51l3XO7TNNIglGKQwXnCVhws
fqIgB9ElOhuQRoiD5k65oCbVxf0zKhc1vj6MfmvtW46OByZLtOK/kxZIN+LjDNOgDFKMiYkh1vet
eBc6HQpADPUibsWIzZq+3Ql2YCaWrUIiIv5lWfwSDhuQzZLEXBmc6Ywoqf1BBVyslU4DxT8wTDlv
fJSeVXWE7qFvWE5f2+noF396//s1QIuLzbb2AstioQ76xDNlJeLhPSHO7G0kClUiySJZwqHlChGJ
fZzcjQtbthU1BHthHdbTwPwZgXX6KdrC/vPEttgqAjAFD/XdU3ZjRZF0+JBmxtpK7nL57EAyonkM
Fz5IpHrRfVygalSh+wsevgc34tr0OsiouzNapNmZ8J7ZVYBTqs/ZXldAdT16uV7C7/BAEqqAlSLH
k/EFYq4/IKJNjrFcgqquzpOb54852WB9+9aseZ9Vl50s2Ke4/3qNvHY+JofAIHECTj/LWoriqOL9
Rha6WAcT4yE+cNY9S9KR/a7mr9ic8pwLWqsIbP5/0YEWzQ5rKaIcbYMTruDMrZJ+/usBc9aOTWvd
WtNSf3Ju6Orh4b4MKzSxdK6t+uDHmro/tJ4uWcsds0gj0K/gWsD7rTEUpvqhde1u+WlX5kTDPPa+
/bULgHH9iRKumqAb3Xdus0hEJ4I21EZlG1C/mcOcXiZ7ihKP37vEia2OAtA5DtcrhhF/vlzH5SZH
bdGXEb7nTgcX9PbPuqNQ7UOuf1KgqdRu/4v6Gxt2zybL9S0Rk182RC1n1Xm32sCsqZwrDmqrheqH
6O/Eipin2ut+HqLoWdE9wFaNEvEw30ke7W55DegRHbSM859aSFi2tJ8sqUerFfUXD0aj9UUEzEYI
agkKHMNPk3iFNepm4PI98uLrnyWQilUwquGl5ReXoq3GN/YhTuy9tJyD5IePNpzBE83iAjvoXmVN
iiSvN/46Bia0kXo7dtRpz4W2bFhLetdLXinRg3ArsQPAV8qm62yqCVpP8dPUvP4XG+RU5cTRuoF0
MLjHw6/SlEhWA9BPWtWP4uCg2fh+qSjC0G1id7trF840RKHhwQO7/t46twm2w1W5zPnxFmDJ0GZm
+tbWw0NqtSYRgs1GUgNUJ64Csjfrfz1yEBYDThxxK0Bn5dBH5UtDn4K5LFhi6nVlB+cQ3p/ckjDV
3ByCVI1GE+4yxV93Ym+wLHBJjqxPP+huNhf4h2iiHg+M7Nrzdi8QmmGHHV+OrcsMTOv/bKrHELLS
Y25gjxklRdLKeY2GHgSzsXzxBY6Zxa4IMS2TBNwEwyKb6BIyovwnK6qYd+ydq6nKUVyQFbq/pxzi
klDl6DmNckO03h4Qu/LCQ7UF+DABR05jN9FAbp7Vxcnshtg2DIQKJUrFKwOKt+DNXCzoUXWZwOQd
1wOhLI3WxfYa6kmQTy65XAKxV4Q1xhgySDLOAAJSYx6YD6gkwoURThqg/G6uykJh5VzI4I4c/S81
TOfEQWAi97/scBfTpUBQjWL6CkaVVbPawJU/v4Q2ZAtT62uet7JeNP5OeuM4WM+oVEutph/auOIi
aDbGHBJlQIwHERnbmFVdPp16LNd7zU4snn8ecQfTc/iMdZVsghKmQ5orhDanht4sPW1IfvFmmZwI
6FZZQv0p6yJ/4RB5QefZxWKp8MWS5RCPaYz16HxGYO/IDx2zc9IYM7MkTlAygXMMPo4FO/z5nKfK
Kg8j0QOcz6cPYCpObASZVObybwUo1hbs+gCmCpr4nKnwYiGFQ/D92fhbW5NyWoA7QuOMzsRa7qg2
r866ZVKn0gzJ1nS4XlEY2A+rJOXMCyoDeN8PTYIN7rQYiQVFKmWxv7lQzhTAsSKYywB5B65YQnd+
7ylKXRaxml7xas+bCE6ux4eu1H79qW80jE2yaWNN8SsEMalTZeNmIu9KZk7Loa2en3tT0WM97Hjn
6/iTtWqmicX2+CHMHVy4tRaKvbaqokPg3Xww/gj4IYe42DQa2LVGvlrhigzpOwUQozwNPguw8Rue
5xkuB4Z+jDvey5QaFXTZYSx2C3jJpMJRm3e5xp40sIFIZuO1G3x+RY4alIgUa/gF5pYwwCKOjABk
aPXWBX4rf1eanTht2JWdYJlL1MU+jAq4iLI5bg4iAVfsKeoVPoDvpxeW7NKZYUqEL9O6gqU/u+1u
FSihwccHaE1AMR5rT9bMQZ3mYeoH+J9jxb+Ky0CJFO3puIRpJImRF2LGrsSbEby7JiQ7Uyy2HxJY
QCo9zteaY63hAlInHFWaMmlu4PoWQxlcwj7iSRW4TEZH+ctFBQ2ZRaLRKLk03kXtbiuC5mdH3pVR
IYHzgDMwgoqU7u963JbL3JfMPMXOnAFsxgPNwLZ+80a5dWi7fP0f+pa/HwasjxePR6IXuuEGGMvN
myZDDcsVtKj24Wjq0WnOaWbvBMfx/KZ3Hh1JT7O2cJRMytJCOaeb0/RW0i8E8uOmJ5EaQ+msJ6RI
nVUmIcXAU8iYvnwqTUDA0ucSnUDqQ/ulukoQudqwd9gs6bTB9NluFGfi/T7cKqzMcvj6lnA7b8zN
bpC3ExBuMTDTcQcdCkhhC+V4bBEXI9mfz7kGWWWzSwB5L7Y+05st2ZMkcGWfcVCqLUqisSD/jMUu
mIQvcmP9x3QrvhMfDaB52W/EEWbx7vEUb3YwAy2n4LB0JbGi0IsxOpHyKsJDQUUXuOCReEdgOSR0
/7TsXiZMTByqFfcfXtqc/upVhr133vHOKkRZcA9ouLdAVz6xQs1d1QDyvEt1ZOcLzeTl9Do58rvl
7UWkIoTnnTKe/wMQMXgUefOyXB3Jqgb1/T3KelHonb1Vb5OF+s+rcghrawyfe48EsZYPi/UpNf4r
bG2GNiy8q4yTe78/1Z2Hg8/ZWCsJPS/7016W7/bxLmhirIf89QPtcsZ6c5BcQgLlFDwmOYE/fHCL
EpkkbJRlpqHQRaIBaN8owAMjNuhYDmMkMhQX7tN+9ltfX2hpOXRiUHvlkd65mDVjpZZ9A/eQ2cZv
OgqKpJ221SHdB2ThI7NDQsKz1anokxTaNACeW2qU+Gwge/2TpXgopzM+8NjXpwHI85/ipph7Zs5V
1dXKf+DlEbll1fmlD4GflxP29jWdo0ZNSmedkVKll1eNvzjVQhPW9zyRhtProCBZ6u+MxL1i0Mw+
65BG6xzwb83/ekqRBYbPdyOiuwT6SXsCp9vKLQQe6yVfcAxxM+qMbLDlLlsBdegDYrraOGOF7a9+
MvIp2DewK8Km91RX7deY2m7h08XQqs8BmoFXRf2JGd0SHg4Vaa/yAUBHv5L4Fi2rfyCbRONfBIaE
CjJGccdQ122lLx1TIWdHn3Aj9vsYv9r8y411VGcrk7J3dJ0PfsXJzFWj/ajEGH+35l+x/WCcixic
BtayAOYEJGxvjPYvkMppy8pC/wfu/OESlKHPMhR5/zpbz+Jm3XvGjL91rYQsB+daM2tp9oPOugXN
SQDr7/XfDK3U6BjNuvyAQ07sTq17gBEW/CDgQLAFMdQCAN6JGA698mem3qEAcIi3GQd6VFwiC9/2
ED5L3wYN7I/qVpskRy26AmJi5MG5XvVISRrmIXmDV7xPXFL6/NjMy3GJ6I2HLoz16TLk++rBqQOr
zlDgmVGMB978OMTB6TQzO8xnOZswz2c7CtqUxA2IAd93fdpnX+d3l/+NecXegCXf9JT1gYFxlpt0
NOAreu8W72P+h+C8lcs6Vsq3dENI+b/7v8TFid9aBmluHE7u9Mk4latggd5/vLTVfA5Pkqpqa46u
PSDAvxKS5X+DhiCPhoTeBBq58Kp12V4vrUV89ShoTKOp1ElE399o+HnaK2usmu1wP1DcZxuZqsWP
N0wtHy124LYhCTt9Wp4ookmtYT3s1fTuz9HVCXQ7+dpfhsa9bJuAU2eQuw/UrIjV0arV5pZJxpPy
obMMtGu3LmHO08sNM0mKOa3VvcvUQfv8bD2k6aigDL9cjAmQxwikU7EcupwVYwwnfu1HQMxCQ+d5
+D0nsmnVS4ew4y7zLH98bThi2w1bTsvlzMPQtMCgLZotYt72Jmh8E9wHOFdsCgCMFt/M0QxegIqZ
t+OkEBQIMPZmuCowEfkSCiQq6LvIPl3M7cynpr8qm3gFl6B5iuhsTJifclVrF5T8hPZfc0k3BDnp
8B1KlbQ2IU8wQoNsJIdI4BQLWXczml8fyZRaRdWcpQ1s2lnw+DJNHA39sd+rV+tMGMvs2LlhxI+6
0o8VRQOg1/xM0O/9P5VuJzrkKAoV9pPck9haw8Mr8pmrq82iSvj23QnsFaDUTvEQFZMR8juN/8mU
IyexjoZCEHhDoWj5cf6Acub6hcGVwbIIINBVczJx4wu8PHQddg/itD7IrL/0jexQgtjyxDMkGIoK
jUKwE7CcuLIvEohik5SmcJKcWngdjOuJy3wJXfdW/mD3pEwkqhbFWFEMicRNKmhpYpdx0GiyORS4
iNrisv+xuZXn3VOXCmJjXN8/NUvziPvyTrsj6Jj33q6fsJo7ZJKRwWXfauQ+d+NUpUkHuT70KLoI
EqqEtwje+w+hhM9220v/XSg/lL79501qGwmNjxi6edSXjzrPdlPxaPGbEJxC+NYzY680El+btAcn
gPTAdo/KvUlS+SlCTLv5smNe8+FvszPS+BKWt2oKrdgGH6B9MhtFoQCMRP8OjQgsSStJbxzpQejI
YkSJGLOpRt+uhRi7FPCNWwU5FLUqvN/XlKm6p6dY6IkbBU3Us0DIIeOVqIyVcXem5INhu8T9e5hL
nqflwrR6r2QYGtVTL3kX6QtCL4n5gsYZB7hbl9WTGP+xKgdZBGH8DecnfHHHtGxDuM5RgFvVw09g
sDxTRTBRVR8SjTUd6akK1GEG21fBqjjJeaKDz0Fx76COiAYxNTQXxqaeAaNHam+niyso6RGKpXZT
ZtCTdZTSV9XVvcl61PL/M2DpE2pjvjAptT7AdDsE2M4DvP1UTT+IPRXqcvGRpM2CT1mSaVwpJ6ax
c1ULwUfg6iY+IMnX09xIFgGj1Xsy7lOS/NRkn0othyZVsMWRnsl3q3lvmMGElbOActxVWnTPzFY9
nYwPePl4c/23hE3L7nxTal/5pvHf5l7q/+EHrnDUDn0dZOmZjDzmBsr3ZAxXZbml66NFupeYe1KS
bb7jJt8XZdBLJdFgZZJ/O0PDjb0/c/WwIvL/Ky+/VLzjrZrcCpBSyOMGHAatSk3aymJ/heeB0vrP
2jrDDxXmkjqlWLnWU5ijH/QIoPlQLMImqf3hfdKQQ/JJRliMidcHdZFMul+0Jlz3wIjHc/FeghQd
5l5cYuiR97CxFAY9OuHuv8FySsUjs7EECwD+TZNXRgm7cbcfTjo34L2ZsGO8ZojhcZLDcFyz+jYt
JZ/Epbn8W90AusoL+iPlhB3JZLSj3ooQ8okwdhDGNBHgCrARzOkoueb4MfstGL2DKwzQ+Ix3iSiz
07xJiRuRzKfVtdaqYgqUjs+Y7WscvvMyZ6wJEIlUv0iVcIUBNS7kkvc7NLkXyTYQZiaaGS3qOal5
RQG1gWU7FahXIwkNs1HQ2XIISnE1U8BR1KDCC4uUQ5uFQnL57Wc4WaIBiqAZ1+ZNLqM8BSScedH3
0BXxCB72GH1V/v6XdvW8AbE+Ar2UQHZlVwnsEOJlhZdAsak1YBWnbnqpacEddYwyB33ojqznJKPR
3sFG8i2e/SZ8uaxxSdvYc87Xa43jpUGzHz+FDj2c0yhciUtVQDgOn2zvnZ4dw7VXLP9jggwSekmh
3J4h7uDusRudfM1k0tnBpufeNxPvDQkwR+3w0BHVB6lxAPb2V3A0lMIoPoBq85ur5wuoVmVFqIrm
xYOeaEP+jeV7u2aOqmI1UJR678NQnyWuU7NL8cOuCwa9kUEfy0EIWRUVgHUcsZrsKOGRJQwq/SYr
AKZONBR09SDweq9NKMvHt47MUyYK2JZeAF66LTvD3MqeZiqrmEl5MXVNT/FD2Ain+mxsQzRcFpqC
0YOgG8pKaKdUT4pFm3oNPv0g6eA6/kSmy34iRmCE5pAHTlznCuyHb91iKpnAwfT9nWjQgEXIRJ16
FFO1G73iwvxU/mdJwXwrx1RbcUwwiUcM+UtW1wJG2YJc2fVdr9cyan3sSxjPh9to6CjApNphAfuJ
fDN/BL3lTRLaYqlebGcx9APCLLUrNe3/eEiiPJXwjjapIjkdvkYZPp468JhPeqWLDCgiHxpjhv9R
z71eUzYdHefyYat582J5PtgAxq7SVLa9J40St6Oes5lrbRkl0q82RdP8hbwW95Jq0DRClJPMhuER
zUQ7UVuun8GBUBAya06qgJbLBXqawqIRUiXNTGHR3PCN6fZusWxOwNiCW03Q75+kHrjfNgBwPXS6
2vb+3ocr3VKM7YlhTw9xXwENmKhWy2XILC88tooR7R0dISrkPHoiZjW0XT6I7aK42GgMoEXoX36W
vWYfrMC/YGZ9vLGOEoRcqOqlh4XT2gcpX+y+zGQOU9LBqddsMxHnhmx4y+wVlnAWZuPCtO9Qbm35
/l3mlp5lCzCIeHQaXmeMmM+XHYEK1yPs7ciWifMZr0Ciz5WaIpssCXBpLLFgTiEH3IdO8bxdkq6F
ZJ/0sIDf31DgJxczmu49sSlrqtS5nHXPRMR6n/TtnfnuZT+lHqWhIxU/PNYQdR9YGuCZbFIeldvF
JlfT3tX6EFD794H6uoEgCMGHgCm2wgoeuNCaT+ftPzn/q4s7yeLfHlOfcXEjzGJGiHiXcOGgvJmk
NinTL+VGS+f/vS82WL3XsC15EtOKLj6jVUSguA7IMR7GItffR5zNmXdFQtc1+zsrQ00mXGEISP6N
tHwQxcz9FOYQO9xOF51nhguf7751jwgu9BA0SJbxhgP1uiH0YZe31Yyv4ryeZdmB23yqOIAPAscT
89g68ynUvfM2YfB7Z0cL1wo/dkB05yelglqhw0BQ8/R1f0oC7HrvVFxHKGAPVlHQcq/M2rkk1hT3
k0Knp+CB1t3aSxCiUT/8f8LdwhesQL6iqNv02v5hVuZYIIbWuV0PWsp6Nvz09wfxdyG98HlnutjT
CGtIh4FM78gLhVpARGjGW3U4jexl/pTPpuZrHpxmBie4GZkoZ7KBXZX8sspjccn/AnPEb5O7CaXl
tARp8nR1WQpJKFF/CS69sfpDwjLuTkhsOZRjKaYqkUdKJiwZsT71dq0FszLpNyoA4W15PvI+ANlI
QTzEzjLkWe+sOrS0rP26f/wRedoUNWaq52QtfmRzMt+tCsWoikogomfkLZB6+2C6aKeSy/6qJlN2
p/xaqAK7weNPwR8o8lNWazOQqKFopR+bKODmIGdgMWORlyKX/1pL9Kuhv1PIGBiM9+vmn3aZWSGs
WtQ9Fc5oKHoy3Y50rAboemqbyJqOMetiSKRXQ8JGLiUHwqQebPrPk4NIxkg7jroizlP49PmpiO3h
BGET1oFH+NPtrow2E4kVpgJizaASUc080G1LS8bKpFMeNCDIL/9KzYah6Y/tHjCE5m8ZlNPMAkPw
6ZyPyhAki0A3zdkhPduh0LskwNpA3mqp19lyb2jcFLo7kwjB1wQ+F4kF0OhkHiYlebdVFwEz+z64
p7dvnFOvFwOqYc8VqiMl5w+gAaWdvxWDr2N4vHRcBsfrRcdqCPSe+yB2fH1/vPf46nxXFZVg3ofn
i42EPlUA5pbwIRlmc2UNKIV0TiMjIJkBkly37QcIbHpT1RmvlTfDsggTV48E06nijQwWBl1LlWUe
qV2DTHwSum1MlUgdYikaEoJjYO0FjhUgLd+Ebr3+vIPB3mmcK/JdVkLuFE4n1s77E1QWhf8t2KNQ
WKbFuWEZRhghUvlvUq1xaN5U7OyrduGliE1AaoV0aqQFzanCUOuqtRsB/vGM8tP9pmeMb42/2JmG
f1BOh4NnDz5YxT6EZgpYmpj8l7bV4/dPYMyBo4Mf+z9pdjaSgu0F9gWjEgKgVRXqADy2dztv83ws
RFaU+2KCxPdKnBZWeWXftUq3xP47BWKT2rRepklq16qmbJdnV6XDVKj8r+qtKQTFThUZJqcAFWX7
3K3fvYFM9ydyPpwcpSrfPmiiWs0kz5qa1KQ8d0H0y4+eD/id+hH298yiH7sfGE+NX4pJ3ZtW6Dnz
49o/DbjjArC5ijl4DjBJcptUQj683K5gyCTbaAx1y9j/boxCmpm5+vQ64Cn/Xy9aSWH2RusWk32X
nLrdWfInH8k/Ie+H8tAYd+kbMdgcMoYHChDNCU1Brhdx0PG8F/rt4B77N1f5trx5p78j9iun2dJY
qTwbArSxa2odsHqHspwWup+iJga9cGBbPZMuYmKExVi1Y3EYIJ6WseTTzC3FAA/Nas1oumboCBm9
aU10NbdKjMlMJxHAf/ZYmTCLtB1xcbW8LFTIPuo2dTSJmc39NlwFA/MflfIVYbx9FLfADygsWIBI
tpRuhO5EyJ3MuxCdSknuLL07cLVRPehl0nBflKiLedo14wJ8uvg5j68dqCK6W9ekKdYeWXiFGlIa
wULWqftoaaC0TUBaUJF8SdtNf9j92Kptqk41l7Qejj9bQaaAv2YSCppjeTWXxVENCkV+KYR+f+wX
bDra3YrlrIcffYN4l15PI0ApzopHQ4nLFgHRkGuZKdniWzIK0VUf0BhQoIk02tXw2/yWTCPvw8ml
QjQDJTXzYBWmlUV3GYj0d5/E1T1oHGoij1W6Fk5erK1lb82xiG19BDMA6veqLG4prlil25tipE7l
ZTfL03dWSPOL2ESpXx7xFlAbATwyjBT09NBKOjw8HxTRh353rZ/svGcvHJ5x8t/PwbjfYeWf3ury
R2PAZslECdWMjfNS+ATBlW4GfTukheN9QcLOW8SSLjaBF1CnKVFlxv3hOKVk5OZeSDZOvRmLPqPD
s24ka8pQwTKGnwEKeEVSHsvLmu5LxKPrlzozNCJArBiR218kKdmLTlE0E4h1qDC3HCG/Aa+crTSc
ZTTX6uxkpOCbMF5U/tzhIzJ9uXfOciQ3C3vPDXqCJlkUwY3nyGFaFxS9339rfv+ujcsb8nHOHm2l
v+QHKnCFWemHZTyIj842T4fotTeONPdr/rt4qhs52w7iJD5ylvd4qMnr37CYNxfr41eKyfEkR/wH
fFswFJBEfIqbNhGRySXwwXPirLMM1tEWyC9ukBTn+NMuGGYnDq26r+USbxupkAHvCrK7f35r9L98
gHF0EqgkwF4+6FnkEBXT0CbJzISfYDBIv92Wzoky5HtpzPx7uMshmsTYxqsimHJeOFzV/gK3cjl9
KZC2CLVEut8F0C6wn8+n0wfwXIp5DhwFoiHWHzPFmxqdwbCi3MQo+Pje5CxxA3osX/Hov/8Jb0PT
sqX8zCL3qQ+Kv/oOSBzy0DBd5kqENNHy41CAYJdYdwFqUgSXvcU5eHP6JB8gvwWAT2WJsscfsM+8
CDY6ifZn9jx78/1tm9c+k+4z4+R/O3YzdFjjuja6Gji7y2i4zXq0OmNaMIRaqQw7lSWtUlr/kXYt
u8hqttfw5W54R5OiKWmPpVPgtYIVbbSqg4bTckO5iMArxzfJ3E3EVyZ/GcsZ1t4zrLvUZTq1DBAY
FEpMeN7bEENGh+6x0MSLaqLV07cychN342RQfFFi8NynI4N9a0YlWG0NDFvX1G57QM0AtcuvragV
840/k01Ub/ZYjhQIn+TWNDMV3AIWiubyGNPlkiQ1bYvR1pJOg4t+89l9LbHj/ZLFiNQhO+jLjjMb
SNYXK0NIT/QuSy8APAzU4hURFycxRx7I5+xbZ2APce0V0opmZZy+Za0xPitIxqWSBd5aX4Fx4A1l
Q5TcWzPElg7Yq3CnayZp2519jIqHyttv7uUY3ZGC8JO415SRuCGqOb9x3Hen2LKphgQotowt4RWH
ZSwbDYVqvnUkb76iWKgqOTgnzXZxylhgZRN1UDoWzM5iXj9VNec7ClSM7E/YV5hp6fz1wiT7XyVV
AE45Za8Kks5zDbZKIh+1nfIrtkDH3gU2Xt3Tzb3tznfvVZpFN4mdBW0FijPGNj4hEB4bMDaaptba
m0OzLThM5hjhbIzxjjL6kRFBtq8sE6GiWNPYIjiFhc6ZqrRcjr9fHmp+etGqe9BJvlDjrwp9kdmQ
6we3VarhfFIpAHDY+Q9i6HPMM+C0DXKOdMR94Ld0Opgd1AZx5EE6qn0IXrAQcyAMKdPZt9fcw9E8
/3jKmfUDGNQZgK+kh1yy+jtyHuerrbNINshmXd39j8fo/CdEEiAudsg1kx/BV6dlT8tnPeAAG0SX
VcS7hN1GWO+VaKfVjVVjKn9i22p8I00G4PPADnvnrHPhyP7DjTClm/j2PU57VSHcPMoclOHerpgE
ObsMj1yT9t+iJodJ2MNCplUAxrFmilkZKacbNIZFdaC91UU5n9DNKcRVd5BXRRj+tdljJkGf5RyZ
EMLFspIr8Y5pbnBjLzoUu+NgGTCvxVWfapIA/LFGyi+wBIBLyVO571Q8MpeNhRcHL3apUFHeP+2M
dkaDek9JdsI0ukHGfSR+0PiT4lJoLjZS01qwZtJzb+a1mI2L/cq5XS1KvsDBughDpdc/+x6SlwiD
Hpaf2kjk5IvtkO3afDA+hez2xRL/RpI7WaHe4noBfAzjE3ByuawXHl44kVXTMkHf862ct94d/X3R
hvzLksXz0EgNEjeQK3H+smuVvbjQm4NWtDXBPQFF8vo8ZYt4Vb7rCajoUmt5P0nBDAsWZTybKhpt
+gn3gplmG59RIhvpPx/sW+ZEA0JBnZHos++f4acjihCpgg2q1kKwVl3g1fEVJqQy7IYaLPxt3d/v
Tjk2RHQqghBg43z89uZYSJwWQB0rI19MnQdcKF+Hgvt0wk8UCoZiOpwsADf2VRE02/SZ0D76qtJ6
43PsBoMhbfdjV9AHSdLu275uoYOFkHCP+Dmji9f35JgafhSsBrH1SbdszkQW8q9Ga1TSZ5cD3yKk
nneoG7WNlFd4SUHe0dCyrDg22SYpNACxqwjgX6QFxw/o0EMVhsw7qTlpfnxW79XwmimOGIAAsLWW
o8savhpr6bUiO7/Ywdhzw+9jUL4eaNXe40twmJa+cDiOiHT05CusMeEfnoioectYA60wSKFwD6xX
FbJrbJ+9rowW/oQBorPjftqN7RcIaGuZ2ljLv8Fv+tbQFMe7u9lXB2fWAgjs7DxjQwGRvW+twiw1
sHcUsaunqlDLCkyk/GpyqzgneJpF4w75r/991kWIx925dFPKuV3iO94SOrDnbdhLa1PRC5SRQVBf
IV3mI4wbwHeG1riFiZZbAEP8YS+uvkPfhC3828RS5FqmAb5D1C8RpAAbOQqdkienFMLunzBjnhH4
K39vH+P/BymE3VtSASRzGQliKpG7zwYm8VLfloGNLp+ihO84jm5ZPRBU0TSPhCKyk7u5fgFyjc+8
2y2RS6zxgDejLCDQgJVkK84+Mh83r2GlcR8sdLmKTmDIJdXIIRlmguLKv3D7CmackI+4jMk9mj2V
PHAnKhRfNgDI8L4/sjmLNJWHr0V73wd0tcwUFZPxY13MyOuAYndiYv0DKX708Ae7QhKhyK8iKK/5
yJyjUPWRGKXy9FAs2CkUJKlYRqGTkofLGTiucdAmT6ukJpDtu3dhpp+X2d9ypFH5ccF93vmu4Uto
fBmDH1i+MfYpyErQBVU9j260BYp1KsRHUJziEZVzrCOvRQUdb1chBhNxgTv5kO2DWJcsJZ0Tmixu
zayOZAi4pJlNK8J29NyNDiQuYXbZ9R6TKVNX0DU1AmYaLLHyIpCT2do+HspkaPzopSoyE/POTPUl
pp/Rpu7XwFAkEW84qiNFcaWg1c6JvRkSaTX1ZL74/De5GbyoYzVX0qgWQaI4AJ/2zfUri4HZKPQ6
zD1oHcaz6ZeYA7zMI84afnC4MEe+FXCRwF0f48iKIfsheNk4wphBtf178yvHLNwV7zLn+oeLt5tp
Rhmp/njGI1HcjIPTgHgr3v8v65bNfqnICTeb3HTHROUkoRwafJAqJPBah5E7SK/FSfilg+eokLZG
0j6Qji+2np7Tc8x0h8JDipwV7WmUbnQxDI+MtXSTNyqOjbHHOVHDaIvjrM3gu0QQJIsNSxZgh7Bx
TfDlyz1jFK6NZffnRNx+IpH6iGoWEd+e8WwgiIBBig6IX2bHexUS9OPMmb+tP7jU7veAy5mJBbTw
4iLG9u7YQ0MNwW0D/JS8jPPh1p3A4PxDf2iuK2/cmdHQTDULO7mvdR0Pi8AnuXWU1+6085cGb+fV
RyJcHXl1PmmhbdpxwQ5P+fUwvdlCm4w3F00cIxA94X/GQW0Qfq2LUEx6UxEU6VaAqTqcq3q2npzO
S4UgQgYo4yDtcNydJWjYJlT8zvQmJZFPLlJBXU+2UgH5R7mAv7fsIOr3dU+aYfczO//Dz5fgwRDQ
AS6/JWGFb78qe/ff7z/iJCXm2pM8lv0VD/69PhU3aesF4Qn9UhjFzP5Qi8O9L83SEGas0N3ONLTV
EYzjdYW5wpL7VT2SL7f855EIP1gDPerwG4uxEmXLHUVm49Ye+TnNJlniapPl1DwkE6i208vvk/xl
zYvNcDpnvJfZgf1aZl9gStU6aS9HPozL1YXe8JAmlkp/O++sfzrP2iPFUfSH3k4CHWH7Iw5BWRh4
1F+xVqCMoQhnDX/e/ej2n8tdLJiqknboiRZdeaCpMOZjaXp6RcMLrTb7nDsLXiGgn3IZ9o7GKLY1
U3e3KWnsr/O1z1cRDCDEp5nN674audnWd4ifuDDdUbJM80wK7XaYAXz0EAnL0D6UWj3qq0/4xPgn
jJpaRWG5tzuqfKo12VuUDe/4ZfdXoRcF51JjUB0kDzMqxyWJ8fTktjeNcbBG8UlVk/9eYWNx8ILs
xq+3XCVvoAP5e1V5v2R7F9SJqq+U0IMYRxoRPong3TGJWoiAFLVbyVGGCmOTFc6ysH/XKCAYUJsm
oZtP1pJ3k/c21/+1w1JGiVGYcen1xVb6eoW9vk80FgrCeUOcCKABuCRqm6FXqUZ+Q6QEQ10tOAaL
7i08oNUFTWxO4I57lH6eiqEZtzzHGxa980UQA5Gk6PP2NmhZYRLtTVEavaJOgADFzwAebiTwZNtb
S8VXODGgtS3pwQJysorIYYIwt8sWZ2g9ACNjDCtnitXBCv+CpSK0MiSGWBdFSY9iE4f6DHGI/AZH
rnzhu5NrAiSqhzz9bXK3yrnvpQOX5+kuq+8ED8y9ZfEwANOS18jPwdztYZrT/cGj3JP2dp5YqrnF
bv65jqUYuMtf229GNmThQuIF3gLroB9H+9vq1K9wzzW+TVH/p2lKdWljO1Z5+qbFiq7D60Qwt23R
B3ImpBW5IGziQqXMNLw4+SBqHucKtJz5f0M0ftInjMwoJv4twJj5T2mFVSA9j+ds/MQgQmWxh6Qk
csOdlLsdc6aohzoQ91tx/0OHVG97/Urzqz7M7kKt1fMBJ/5U+8h4QgKJmzjG/hfeY13RwV1bIMqD
2D4Iv95XtS9FqdS5ylMFvqj2S+OLayaeMJZzsVw1450+YSOoiC+7DojwWN3a9sB+72o5o0PkRmsf
Li91J7mIdr80BvGhYx9jlqYefCAzw0SLrMlWBwKohNn0jm8f6D680m027Od4RRmNEuP3K+vuxp+3
9QEUZTeq0fwy/z63rQEHoZUsXdwP9wPdB6Y++PMZc0rPqVPLhZcbEcE2L6J9t/j4urxqBt9uPuBH
+OmS34wI+7P9aFN5UD/2hVAjRtq/V3vKQMUFqKgRilO/fK3rh9axVc0rIrrM1uu/Ui+eZOHAwHbZ
odIZZuV1EtXRCrdZe0WaFni3XTE4bJ20i10dcZMuO44slRfM3KyMW4txLN+96TnYOnMSS7ohf3tq
Jsop/0w8vv9zj9nE4DdfouBsZjGw7xifA6lm32pyxc4tRMqCCIHdlO+9IvQ4rZQtPgcjE6glYJ7e
XaAmFzrkdlwPwABwwYFdDHPiZ+R0xcNhYVGOq66SIrAUlxtru7BZBDmZg5PFlsEDT8V0hfedO6tq
6kDegzadoetj8TXdCJNqs85r/5guxFAAvM6/D/MFxBPaqRGBv6sVklUkDm1z8rHaR9dMVOEIPVC2
cAsyEXPTJX1NGcCGQUo6xIi+abKCLELKPn7L7GhLGgl8SCV+lWF9+ooGFgrx7jg5ONc94+2MoYQt
XDMR2SaddswnHMNNLySkn+k5AlTo80BPsDaivM9jEE5LrYKPxhFmMxcZG2mOJotsf7Jr3QzBL89+
9m1LKBjo+0aafIE1c17RBbj6zudBz+7mmXrWnJua+4nCjFLflGgnAy/9wrzhhoogMjApMLG7Mjlq
EQ/LU5nDAdizJdBr5O7zWovu7/3XDf0gkZfM8K2eeeDUSXcIksaOanhsuID0vFwTPsQu+gibfSQQ
70JnZDMK0fVYnbMNoH5xnKyQId43AvJ4d/M1ei8l9T1zhSZQ0UU+veTHPg/zQMGceCjJAoLkjqWS
1PW63y17xxXl7DQ2fjdcCw6PQn479EMwYJIxk6s9jHpmv0Y0WYdkkskzAKblE7is8ShmCwVHXEYR
kfG4s3G8o9F+FkUjGABD0z4idSHNWNMZ5MQJ1HAyr8DbZYP38T1a27a0YzQDvbDK/KY1m9DJVqiz
bIune7UtmBP/GYtl67ujF1El7CR4kmxaCN+8Sz20RBBUvyzptejwtQ42c/KZ0PTA59kLh2/LYL8M
/y4QxsyE9ySqpuWRk2x0D+4IM3zAvcCnxRLB3xNp2gGxK4o7k5b0sIbwmTk4J2eUJjyBd5t6E7xW
DFfSQZwgC4kGsPCu2BDaN9TBVA0JC8tDvwSw6QlksVA+/iBhmkToyueCmKIfLajMDuAdkgzZQC5D
fOMBHim2MBtXrEDhBcasfuSnKcn5npcWOEeBvzdxHF//2uJxmGATIqtuv+toJtAz5FAeTImhhEuq
PkHA10845CV3QODjGB9fqS6hcSJaNmMvP8GK90Mq5djhQtTmOZqCPZDSlpLlOrxYxxChsGgUID3A
swEb8vr2fmC2xcK0o/Xl5FJdbn3JXDt0/m/vV7+5CNDvSJujQY54wE2zUjQ2Afb1Ae2g1ex8219V
mBcYMWvfn1zZTrX7CUvZBlM91U2+qE/WVK2ZnHqQYWXws+IcUtv8r8Hn66TIn+hngLkSwaAvOQtS
3dOKCyoyMb9wVSiC2GS9hUKvE49jg3ELhyBhTtyeLg473CXmA0M+ZqdJ/4NLkY+yLn0gAsf4MRv9
1FVQuwyzmwVhcC3wrubaOd/FtTQGO6ZYpFe87sMDY20l9IowQo5IsjuLO6ZU6wkycVZzRvPwVkaU
jS4oVlhBKNAiGxP4baYtuq20hxXpONz/R4PTNle+Zj/huny5HsNjIoTGtA0aW+pas+aQSl2XCvTb
T+I7jweErCvaeFQkm2t3pc/J8K4AGtKiwwcANbFFPNxMle15M3SOCG8RXNwkCum6JR1aNWUbn1QN
aYdjlLvd3GZP3YfqFle9q2LqoiHql9UOXQ6VFVhxPjuRsJWyxxl/jxMGAIgWlPizZ+wtXJQH7EU2
MqaTjTALx5pKoJNhu7uAJCVkBz0LGxC8h8kbFCCSRWoTaesHO6CErKtO/5t2dIrz3xt0r7ddtFWa
UygRBjINsEyWTnoWjHO7OXGJcFj/2EL0NsKhxfwXe1Q5Gi0RL/PP0bK3SsMlaEEzkeMee9Lg6BgD
1J1Me788XAU68eAJXf8/Pkab0IynbrR8HA/YGXbHEBl0XrcudqsbhFtYmTY342doMbhohNc8cwHr
DnTNAShTm1zK1vtJkt10QaVXKiPp+teb/PqBrC5Z/4n44Ihhh42ACaKcBSgLM1cjGdF61oiD4K+R
im97S/9ReVeah6Y+BLep2zcY+e41ioy1a64ODDfB8A5UNqPaBQmCVQGYl0P9/KK8CvVHiKMmVFF3
sSlQ9A6aXK/MfKnhv2oG+5aQAWyqjIT3z/GG6Osj/pm5JHpLvlAYadhaDEt+BTI+fEtr9miXBTLx
wMthmHy0lgqM3FXcMNtiyWaUhw7szW6w0NjP4IK/Hfy/lNsl4l51IVqMwI54q6csovXcBRhfFWC3
h36XrEHm+ut5vZnclSy2cBhdSMfOcBP1C2YJEuDSqklPqDAnwEC6fwFrmiGSa1GMFeK2hCAXDbpb
inqsnoMdfPfLpDEqnE2CgabyYyt8ujvH0AYXknUg/L1jSMjyn8dh5GIiY9Y0hdqO+Dq072XwyjE1
LHMngrKQXD9BXS76YJnE7EYE3BWmEFq2ZS+vTxTAu2YDNESD5Yuj7s1kK0kWz74qYGtAUwVayNus
P0/uu7wS6VYYZ1WF2YQ5MbA+/RSIT45CfNpa6Mbx2pfCkpvR77JEZWW0nKSI3X/FKhHQCRmNqJsj
GzB9uWN0OnVWbcXAYY45gqDT2J6GdceUL69LWAlUf683h1frxufgZSOXW3+cWY7hQu6FhIa4zo57
TBWOBIPg03x107NMDaHcNu3J59nC0XW2wemoUCgbZK1U3iEbyjkzLiqlNMAdsdhL3IcrrALX2jsT
/i/pNeFCaMKCgdlUfSN2zT2pPaTKi1k3FIf+GewF6AN8UuU1Sawx/1IrHGR7Vb8pO3WK66hgWbxS
mjcjSyBRJm+EBnO6MKW8W0TP2P1U1Wq5l44WQdA4yyd8vmEliXRmPsB6R9PPSxoVssypkKuM1DxI
6FQEEomgr85E9zc40JZ8ve8hRwFBBO7xNV1y+rKDGhDEfGFvuM/fDgiwysiJ2vh+BJnFW8t5qtIK
6+4zakGxSPvLgGmotTNiMmQ5ICBpNN5IuGAZIPVIdiT1aGyP0j7htu8ayr8rOAjZnBkbEcDc3YYa
bmD3YOFm1sAdRR2p1owf0QEKfKQnyc0ViBwtkz86/IFtDVuhwTdc9XsSR/qHvC6epfS0EMwE+O3d
5KqoX+oCg10v4yDHmpaXxaRlVZrXeczM+73OyX+av25gyYxvQiEVeXkEx8lrn39FoiQ1klhMyWL9
jZ7yYVOMj1JtspRNcA1gl4aqDwQAtZwstqeD3f4o7YP8lBO6lGNXUSFCwXFHb/x3UFahf8IBruel
XkQjdOfAHJ9f2Q+7yR9vBmT9kDuJX8AzsFeKvJ2pYr1w8Y6BOthKiwnS77ABdN2nh33ZTg8mFEUW
ZIjKkwk8I3kQUZWiqRvDDaSxoJfsV9GnHPQETay2l983P9bOUXNA59dWmoP8Do38dUYUkihHFA92
U84X0lqE9we3SUQ9jdef3sCMN80QzWNUZWa+TBLWSnjBwuElF1Zwo8nakRPnuJKleuAtn6kvsGT5
ZBxtJMaHKM1VQugjvYhKCot4FiDRed6NqtZmKkFVZfEUajgN5jtdrR1c1lF5fHs98KvwEPCED6G7
SOSdUh4erpi6+gzV2cAf126QCuorAMpUgB3ZEWbiaov4yoZPuz/tiDIkfFOJg7Q6khSePFBkh2oX
OoVUZxXen4ee1GNmKBcV/SBybo6LQxzWk5kfPyDdEGF8F0M0gyWgVv39edgJnwoTSPFLyVUxnxYZ
rHOa2xGf48ZSAB1+SJ3FsawWxxCPDdv9eXjk2QENoK84xHFMBrmNz1/4SDngHo1j2a+RrlvKVHE2
OONfl7LM0Cus9f5cGfqpCgxGvtZWV3M9CffBuwpLmJx9mBh1C/EJtz5zTbvRG6NTxhBdzgSU8x0V
kkdry4bcy3EdFzwy+VXhr4lqVKiN1gHSV5fnaegc3jUk6XTAYqtjhBaukzkEVRtlI3U6yD3m7gT/
Vrdv3VYUXQRAPYArZutAJQSFsg4fN/qmcpTrkY8DE/TEVc1N3VVzzS4LkBHaRDGGRa7+J+9fizGN
MoLpTprnIdB+A1CCEL1xwb/x3lWiZYEkgIx9h/7EflnGxXgcOo3NteUdumqdnP39FKjn3IdLB38s
KY+9knyoWl60iOPcUVMGlfwpzyWj5Z/68t6NJryEUUDwuV8vv+5VsnUOxMB82Rlg8oKUTTQaklij
4J7dqP42RyV2jy50rlEdJhPp2X6GPPnB4gPXmKj1nZ0wxkJ/64vXWKRlk5gLPr5fqH5iyvDn5+Kd
lbdOzkFxoY8zQD3MGgRfHiyTqM5vbXkkgKZcNuMY/PJ9CQCHJK7/+qDTOsHH0lug9YnvUIusoIcr
3sAkFT2uyvEe9Y/o3mqTqqPG8NChGaIAfBwZR+HLeP1n0Su73wW7k4M/rDfdBe56hYE3ytZAqFt0
LNltk8tFK+1M94sP1do3H+O6VdEMv+Ec1/AUCDn705R2dVTQgJ3YCcqnXfRIGCdE698yGL+2oPRT
6B8Baev32jBQ3kgwl6lKJ6hqxuLgYIl9xAuN2qLnDYExgFQ+thlYU1Xa3cXqT8NJrROKegVMnYLh
LCI3cuW5+xhlEHpMGlEbt+2KP0gNfUtsp92VsuvU2A/qtAOQKCNMyFzvcGGREj9iD35hoUIxueuP
61AQdIMKlbfl071HLGHP+cvUECNgiWqk95cPczCnbLRqZvmiU1It2c29+cQSigkKwq6GCtoTJpDA
lZpGBMx3cPwZ6bPesKmeEjxja8kgu7TklBqlFc2YsSEZwfj7yXlJR/9Rd+8pPtFf2lxcc6YkX30x
mcjuA39n6smF7UqPlzT8WS0o+/PuRP2xpyLGJ/8YB/L0EVU6oHgTN089mPiu9xRl0w8yGMc0a974
biccWHlsStSqw91pJEFfJYjTQnOMENXBxSOaxN0ByvRr/Fe5DP1MjYoViiZWogh/syTQJ1/+MpXM
S1m2n+xKozE+u4Ao2Omqf8fpIn4/AIEwvCL4euzVNS78+/5rliZJ009lc/5ZH2rKC5b6Q+T/0vr4
3I3EiwIX+hKlQNvWXkt6/YT2GQXr9fFByN+UQnaGSSCKk07sRVPJADec8QXMfrv20gXPchA4zS9G
LPE4T0zmHu5KEn1WK7nGkLie+KAAsGG/uHHS/P/hEN7xHxboeJ1t3IEb6nitCIVf2NprTs8NKDfc
d8nV+pG6gv1izR3yfHtncKsRC9k9Sv9PZvWGukVPphbg6DbXq27S7Mn1/v+ACoHnACuTsmvUJzEc
hR5WpbNwUqN26FH4PrGyYnV8IyIq/08I342e6C7uVsxEkiuWOqRHO7qht0jba9q8IUWVtfqIUVmJ
0nLs0KavcGBhydR5f/3oGBgeua5oodE1xgvyYO4Q4WDBURTiji7kvv8GS9jv68JDzdfo2lu8LwY0
qyCV8t/ls8MvCfSFnriQqgiZ5NkyCFathSiJY8OMCuWuEhefr77RHOYp9CwXdGQZxihkIZbpm72g
PEkeGtZZOo9ulJr4+w0gx9WCuoReItypDxPNw7gXx4xUUruKgDvDkDank2ufXqclld7w3SdRBM1u
V2y8VFTttPxfqwFkwXAj5Hr4gxrgQKFrnTbYZAi0Ykv09RsRev0Bk7bDxkwPv2cF4H0XIlYrn8fr
S85cqJdy30PTi8hRNTfENCNgT/69eK323ucVBfV4cs9d+dd7WP/r4IH+4CyuD3CynDmL+uXFBOMV
pQQf3VJH3HyhHOd3lK4coIzjTg5uMlM/vy5C3kSKfR5n62unKI5xj+R2+MaNivCi20Z94dfXMuHi
As06mRtSMByTRkXvqEKk5omSv7jff+Wbn2HTOdByzknB9LDbi5+Pmh1NLxLf+lHiZO2Guwh68X64
qWjegb1V26jG6yqwTX2qrpX61JJDxD7HUYhX5TSxK2onHbke2RRpEmmA8rVglyWTVONxhGubrwHR
XnzMdqo2cAYr0W4PkIUktrVcJvSFivyTm1S5PjYw6j5UsMtXos+kZe6bPhSaKVIBNDzHc8lEhhzY
i+fhL/rQ4kKWZUm7HtqbPZzg4CgcOpZglF2HNR5favPYyWEs3J6UzZRqcD9L5mvTSSFZAEi+3BZx
M9ZfEfjz0y4aBGEs7NtnH+fbXhBEPVffecTJKYEXiB/zpl4K6mm+OuvuY7VZnd5PjxfMLuMQ/8Wr
Ua9g6o5dvWPzT+HYqVds8jWIK7haDid8xz3mIZSnxLnJN3qqtlOcck8lZaeQkU/aeY6Cvgmqo6Aq
/SrL4UTh90oGIWW23Ue4zUfh8oWjUc+O4HLaG8t/lFKkcEV+Ghhdus6P3cJvkZpcXQiI1+FV05CM
urdhWsEg5flc2P6GOD9+g2sodC/PPqaJadbG/YpUjfIq8hG5UNDqSB7IEF7HTItphcolLiTtLSi0
EZq3G2Dsq6dBxnCs2CEiINsHxwA7gwlbXzLbY0F47iOh+csLXNW80uB7u391C8zwfq78/NZ4+4zf
253jDQt9ORK0OCV7F1ezEvQ3HyL4R2ZHCpdrs7gMtwNzt1G4XRTphX04GJrtZZLybg3Ab+/yVH/P
ZdxMFVNjFb1C9HVDM3mc+NLtDoT4DIlpPQUWKYzgvgosZu+jdOcQf4F+sTToXWr8fhbgz9mRaiq5
YXqT+5HWDgCELnRFUcM5LivQCt3OIaimGP9UWra1pb5Usw+OnTeR0of33ukfuKj2aN/z0fKguZn8
itKn8fR58f5YY3N4ubGM5jiVFJ/L3iDI27Zc9iKJyIMtvZ6NSAInvPZl8ADItzJLeHCSZ7FOYCEx
jE8kjq8y7m39fOxNbOskuOnj1ciaMcxq2BYyHdtVcAVZFpyspsFG0KoRzbKfV5tiC5xn9pmDm30W
3pba1wT0MVceSnzcS+ZGVS7+j5DMMjd1Hjd1ds5a1iU3MluENkffAIKMJGSTXFw9/DG/0nHc8ED9
HpTytUBBekD2rnEUvpxiHR98/L1HXeYEmgJ871At3y8d7xjQvpPzH9Q6Babk94sbbP64YKDMfGo3
DLg6fJm2/uNx3fn4in76ZIyVZy+h3Wzs24DX1F0NyVemoU4agIdjXELO3cFdN1LGAkS7WKx4tpQB
gT5VrbkaazBR+LQtzjI9rqtUnqNS+UGnMrlT6x0WcKWxByvnoU0jOP1H8NB9eJ+gbJEV3jXRYu+U
4pFjWLqcjsPC2pvDUWJQVYFhZlEar7VUMvI2bt7Uqdmgvm9d6aLMbkQHncmhw2hLlkkqC0sROoLq
f+UgXsRTg7XR5cJee4qmJkUj9LbMsnFGKa4q2Iy0kFTEjr4m1IQXDrpwCwZHlMxR1f9t6GUVxnWm
98cez0RO9oN+KJDNu0hgOELvaocY5ExuFDc00LSlinxmbWNqaPoweCkH2++pz4NT4ZQTwQYAqPhz
xgx7Rfe/oESRWfERQrwrrlwliLniipfmx5dEwo02F0IP/hepe/dzEFlNaH+C+oMSopq9tIJVKIxJ
wfg47+US/7nqZWw2a0ugKQCYJim7xZA7NctBUf5brOcv8mypmxAxLzwZy1vlAttwThfmFdYvL66c
xYdx0asVVU4zFk5wzowNW41zDYm8+72MesyOoiaeEq8sb17jYMrT/+ECOJM1E9XK2fLrH5rKc4KI
qOP4UWkplE9JvMl12utwweZUnjJaNE4Ka6fh3+3ujP9ugs+onamnNHUKXiPehXEeuvl/q8yd73oj
PtOQCPbSaSQxRyb0UpEq9i3rnn1OZlv8kvBz1wwklQAwS1DGNy1nC6i6h3BfRGVotCXOsvn64O02
YRV2FJCPVJiHy0LxwiT+MatUy+OtbYbpeS25uLksD+ejKFVwCImEI5hi2hnDtuhMK9WNnZMBeRnF
4UEkyNE67L7zhJRBvB3Ybd5bKQhCu9CABmKcAGFtL7kENZ/zdnExVSEFvzqz/9eGCbKKYjiTr4Wx
XifImrqLL6wSd4WVxXQvPZqGlHNUXURusn71NzZVhdwA67b8Aj5RRhQHEFHQSIitQi2LnvS0cLK3
b8FyGWAky0bar+/ikqn0WNdiblzKPfUGcjILNAqzRMZZwMo27FcGg7GrhXqbE6N4J/W+NfavAZYm
Kbsln389KBsD22FKQWhycMyOfT+52sQvV1CEJO7XqPZK1fim1mTX4FDQNbPi0eC9i4RZ5rIxOe4j
joImCE4oEaf9B4QKB99lH8+Lms8wbrhvUiJ/K23tbjIfHCeKHZy9eErcrDwKgy+9Cha3wVg52xyg
kO0lbVgDE/8XeGcSKKeDSzBjHKCjVCQ2c+7KL7sl0K12flRcH51CRhpzFMSKLT+Sg8/HC+EEZHPU
VvaSz+86zf+pLOzpE1ov3inXfStaSrAKgtH1mrVqG3s4PcPV4T3ymeer1dNMLiz+jHq5iBNuFyhA
uXtShvOVclEz3TOdgRORmgInBpnrTIvpOFSJyRUHJTU0B9dEJuhDMq5p5WYynVtlrWYvn/oJiJvY
fF9GA6Kta+RXo8Slfc9+urYaQPuMfWL3FEXCTY7nMAbd+brFt4Qn+X9T1r4X2EDYFqOhyMfFdREp
JCbiPLibA3IF+bdQeAhDlQLTgpauSuH8U+gimhG63+yzrmXWCUVEG9mzF3al3+WF0PdcsBXsMDp1
gd3+bwmSfo75AtBf+16f4/AvSanw5u6D3xtRSReaIVcLP+c8GrLfQrwp5sMLBjV2G91mSpyeN1u9
u8nbiIuaGSfvzrXzvk2fVEQSGo85gt+Qe1Sh2AKkBBeSGLDvxgEGvfnt15IhaOQCrjM8TiKtkQ5D
ZuPqCK/yZixLEnb8vHbEL95+ZziLeb6+AoDKe/PJ0TkCOlHgA6lZGwZLyo4NnGcozyXaTmSuoZKT
T4+ucOggBpfgOGkd8hwCsq0RSPzHjgDgtwVf9D2ORRx7+CeR7zUk9MhpHbKmklnHY8dQUD19/WXA
DN4ubGp9Xo/KQocUfxDKQjxeAJKyh3edS8W5LzA5KA3Z48TWxiAMkM53CBrwddNT8OFZAGopYtFb
45i1cbMPIQKYCp+3pxamsaDu1OvEqEQ88BHqKFTpqLpdmQeaBJCeFdrTSNNBhchK03Xlc8Eu+LAo
BCN4XOHQMpN+Mu+1fzYbfMKhts58TB4Q0da6DXGd1tzRhDbbtRDtC4VIcuLDGYJLr5QUeD8EXkBt
Wlo5GjgNky+n+MUIEK5QPdlW0B6bQyJ0ygI6eJftSYk8iiJGt2XPaZGctewlFwOsvJl1bUIm3OKS
UeN2ZksqQcIwoH873HDCU/lpPVOxOk/TD9ZzO+uancuMMc8HRuMVtWnqL6MEqTQ+fG96hLHwmgNF
t3KqsdMGuxGOL/a8DZFITYckTLwzJXYr4FB+VXmp/JQP5p+jHFw+XJ3pyHqCizRfOxRCA+NK54bx
+r3nEQkQsgnwTo0iltgJeDaeV/ECuMqquoz4EdWfEzAxRYpaAvY8dq53IwRjGzTUTBSO+I3wDX/5
9pfx7ENTDiCoWZq9SBr65sqw7grU90tJva9OuUOBHljFV5xDbL9LoenRjQXKQahf8INmmMu5U3PL
YPq3uTEEYImGUjoaYl+B8zbzuxLBiWVyLoAcWNqKpgcoI3Qak34Er8APc6oJGCglDz0jdIFGNL8P
CE0J8g4ezeessmTZQ63m3YxK7wjrIG3yg0NmoE8MMYQUsyRbxjij/mJs4pjKmEqd3NFQXYaOf7Xf
vbw3LEzGQA7HJzLSf9cFBV9X+0hX58sICuVqyA8POXeQPjLmt3W4So167jepx51VpeaFQi4QecyT
EssX/OVRIRe2KV/1/XUGihClEO+z+IxwM46I3XgZ2S/xMnEblJl9OhfUh0tyb2acpiAHVZuxZV5B
wA2zqPj6DRNc1PB/5HkXQnaggbXQQnkl8Pcq0Glr1+CfYyPqVKrN28bhaP3ZYdJt0A5UfefNVAUp
M8jtlwi+ypejIjRSwZdEObHo+rHq0/GcFrhcb8HoCWnuqOATDH9kqhHAqfIX1t8Y6Ai4T0/dWKOK
IYrSrGJwpkGvD3hmJ9+dPMWyL36z6xzx9n10YZ55PIo9dmpIK6dOzb/6YcAXMnR68ANcj2z+T4wR
tyMZeg1sJFIRj6SppGnVtohCtx8FvP4Sm0YECjEFTNtw/j55HkcuDvOAfvOU7gjBjnzfNKMi5HRB
Gmbxhiiy1SP1bShFhi+24VG3Zck6oUt3WHzlKkwXRtLMTnXpHxawvSvHDckrGAJcka03hyP2iG/O
N7IzfePDqjDlNRYCk085VVfV6Ei5DmnJSbPb2/WPg5kAok54DPdmmWn0JlEGjh0A6pCdWTEKJRIA
gFurde5RaNPBk0enpjNIoEQtH9kOpr+gi6S/gFwym5sa2TIDOxmVxIMvA/YPsYYwsV3lTNNjFiIM
b8+r3axSJrETt+aEaNFQ/UFtUzaHRVHYpOO7EQHpvShgSiosyAaAB+3MOBGwBrX1ff285R7M5ofC
+xsKlFLVprwFqWjEeGQjZ0f1WYS2K7znH3SpmaXUu25bDf4ZuEJjuoyIeUHM4eoFdFeCKNqK1/GG
xAaJJetuPIaFFNL/suBFnKZODJZf6py4V4HWYt9jeWCQVWkIBJMIccpjigZ446ppXuYCD8L3XqNI
h0sSIgoeOPj3n+h5Gbq/G/7h4m7Q5rmt0ZVqZtgtXpCUVUy7Eor0TSpQ3NdzEBL980AdXxYWPwBk
Ho7OCbG1RHeLNiG64JYhQlyqduFDcGYNRPvmRKy/XnzvaVl3I5tO/UUiAIGajjaeSXOYZoTqFNl0
NNwXuZuYkxGRXShz/X/5M0MTuLA7LauwCl6Q10/gu/ZqbW4+FkmGL1daNTdyZvqvxhQM2YSZAfIm
Gx8ZEEzczdBgc0YyPTAQ9hVPP3cXUrE/PP5kKS7vLMqy2Hq28D1MMjqR5Bud4Y+aai/re5lfUwwA
RRNquPSsYN5HPrEEc+u2zkdV+ZuiVdpHc0dGgVWsiwAC6Gg0fkHPww5LpZG5K4B7iLYO5FbrYMlt
iEWRNf3SK8U/4W/SrMAzafajq2YnF8YHO18l6PCP404bkrXLhQLTHQf3+yXnkjGJ8jGF62HeMTVD
IyR5bD7CsWI2OIDYK6Po3nk0vYvTnyZE35pv2Yxy9ntmoopSXuXDtgD9wqkgSWYJI6GIqF88o8cW
ptKEwUeDdgIH40PEQMeKhpLOXJS/utOTO/RnUDkPhfvU3wfMoSaKCfxBfwjp3XwuyDoP09r3igmz
MowZCrzGiZxYtTEpPYh4AbqjJzYXtRPjHMaF7LoUV07fNYvyeqVuc6VCUELeqzgTTLD1OvYtVe5a
VWzUVpkOC2DhtySx7ujBa2i3JUqH8WfdHpTnUPnrM87UVLrrf8+xqJPpX4sKUQv3uG2/z8+1XcMT
cRmyFFxewBDybDcMlYoJIewL5HBnQ1Tsj/SRDnZDQ/GFu/sKtWcs/mivvruiqsMthtAlmMFv2oP5
5Kba6FjQ1JMXIC6Cz+kWnR4L+iOuqjg4Vi7E5Qv23cATAhBr11WaHN1VQ32TEs8jg0cfzrtgal8+
zGU6Nq+ZZO5ICDh5LKrUWxmWws0rpVYqH/Su3SA3l1oN4ChhSAH0+dJbwH8DOaZPjIHBcGgo0psi
0ueoQ+n4QLrLKL3/w5EevRyCGrvJNV8XsDnYP1wKOu4ZNC/mdMzeH4CHTLnGFSVTRVRJ5c3PM11H
IjfnV84T9vK8TpWFNYJDMMt/VbyNsRASQWyZ/GAIPTIaOTOWEorKvRLBX477bFZn3i2nLo79lPYG
my/CcBK3ERKV2SG66Q/g/HvazL0BbFJlJUU4DlPuUXaNzjtK9M1FtIEId0CHkOH2ud7IxJinj1Pv
6VfyV1T9l/GHseMihR1XjbwzP/ivji+PgVd4ji4rAQPc76FCSk74LS8zmuDFzZl9qeg9F8MFtD78
614Na+VTKnd/Ofm7W3aonaA0RdB4vYBJ7j6GifCfChzKRGD+Rc9PlBFNG2intcfi8ITkdaDrjOs7
WVtAlQnjAatc210XKj3lmzvYMJjPUbHgNOwW++C0Ooc6UN6Y6TqVf4U/t6xUrv9+tHZX8I1wF7LC
XAmsXAa/OPNtS8MyaE3stNBL/pNYYPXubd530U7bGpBXKX9dhQBy7u/S1bGzgoy7oNia+gaKiKOo
F3O8gMSYennqvDpn3yeXaiNlKNKrDPucbyCEHNjbLjWG8UrygHMhs8GngeYNRVr9v9t585yAWXSH
+RGQBhfAB8Dnsj1tag5BPzed0Qw+sCoyI+UzAjnDSWQL6mU/NSgL4A/9BWN/SteqeIh6p3Tt1U8i
8vzb2r8kgeYu6Bv49XRvAmTlC5ANfBtPds2LPgGYmLjwJ7O4K+KSEI8ICT7DXJ/eMcMAOZHIerOu
BhSSQypTu99cS8H3u6du3U3URUY/YamV4U5ZBo8Wh5LazPkOS5yhUAswms6l29UECxCHLbHU6jxY
xH5aqNwRJNvzMFhhovlfUwP5f3Zg3HXGWD3LqAhfW25J4SBnTQoKaqttu3cGtqn3DFV7FuvAvIBy
eKzapNbS/OwtCmPXmvp77T2yvFfOoO1mNOB5YSXSJUYkIdEcIuRasErh6SA6a/GlKQkEs4fUp4VL
GsdA/BTH0oirWRI3ft4RGZyZXwtymAFhOz3gkNDvWSpWwFA4VfysY0zXhB5b9KZKTpZ3UDWriYIx
7wDG9rVHwiAXViavHO14OR6o07bZtaZtUkE4bdisp0r0y5InUkAcCAJgYbOJkgw3NQX+16MOwVuQ
0lT7HAZvX0pGC5HIsWEtonXSBlk/jJIhAmOtX8g9fID3/UCx9jqpFMYUCUXwvTzp6LsNR4TDTEJ6
8QB+V9B7ILf/nCAAub2oob5z08Vc+mdXx5dcTZm24coMQqMZSaoP6AKlzbc+S8P0/cIgkLg6W/fn
Ks7S+pTgrsE7poE0KyhwTJzew+HzXZCKj1Q93SauN2YqcxPgoKX64sqeg0nQ0NeICRqxK/neThZT
4nvMpLmuaREnia9W+WaJXVDRZBWsYU4DVBF4ndZswkyOW4Ubpe8Bn39LNN1SsmoPkmU4A+2Vz4wr
J12FSs4CzoXRyVd986K2u2iNHXd76gw0K9yg3GEzGZPv/rGkF6I4DwWKl77Wz4JHsnJKJTge8ojS
T+V/5V/EZid1JhIPrueOUegm/bhtAlsszcNbpYw+NltZLvzW7Le6aqSaEDtNhOWjg6qiWtBJ7iQQ
IR4RSID0FqmP998lRnh6tR8ne4zItwO8t5mJxj0RvYA/BTidAz7akc7k86owNLZ8at1JiLHa97h3
I0EGVfOpt7CHyj+TrUn2JmJE9wd36TWx48yu4L+VKsExBs8uyXTHYuCRaJ0cANQiyzJwxzX/EcQt
ibQ+sRE1MKN1snW+eEZf3w5/VZMHiLqlxl0glnG0FyQVlF3s6C/L4ZXiBqhGyutyXdPAtbA9JVZs
9W8o0vvf+siuV9zAviinvgV/Tv3293wbeCGS7zbR3EADt5KfA5cLY+Qf4amA+IFAKMGS7MA8PnAj
DnicjesoP4oa/BXaKaIgvCuSTKO0oo0aPXtJ14uI0P7NQI9zofR/rA7tcnLtJXjrLVPUB+Um41Cf
sHHksQP2eLFudOqkeJYVJD83wijpdb4xFqTYAZQTfCWEGutPZ+Xz43mLG0/7/rGl/SMXEznq1umU
uTyltotOSHfZ7OGSSVL3HrwOiehsAF9KxKbm+LLjx/8GvKxuVj9YeesmFIRqRgTeObxq2awv9Evy
W4X2JFTdxlv0qa4rbX6diRbccZiOOKkx27Lms7+BhReq60Bs+ComHheX8YoNQ7anD2aEr/cwLVWn
mnSLQt1zsjp4eTnVBtp9kTzMQKHMbf5xXiQSKt6P8uI8fL5FXp+qMhBOheekVu+hi17zxw50vEKk
Yrvq7qRf9kmEmFg45AbOlFKlkC9Xs4SIj/L6w1tGEHRjxm5M5eiUIzq6R2f+cEN224s20w2/zhUH
CgsrNvbGlM+9+SGLflLiqWinX75lSrW4u9LfIWpDUTTmaDVFft3TIkqtx7piPX9SFsIdITSv5O/H
0Mz96WjpMuG8So5q915lkJzDXhl3O78TDDR6rtiDdWPwEAqvLfx/O09DWQXrWgNtVhSzkj6Sq4Ec
ZB3juK0uezFMr4HdEyQo8tCZyQQQC5+q2h+2q+Jsfc9WM6PvvXid39lRLQjf8yG6rNnKxBdhG39I
J/6eqnbGvKCkQVciY7O0CIfK4kv9JJMtvQ9/Q9rz5niwyRe4OeeUgfPpBiaBzx6k7LNN3yQX36Tq
iLJynzkbMVyU6+osNqVgiNhF6RO8mCOXyTDZxZRxQ25p/NXfClhuyriiaAzaEmOs9Zldw4D6y/IC
IB3x0M3llIXvejt29ACnMlkeEyStkdPnHDFnlehc2ZvmA0GjoQvaztZko9j3gfQfY9HiEJRtTOzH
YBQcOAa+8NBC3UE5ay/uVKQjs3DuOAzlXPij4Y90kygtgohRCKhXQBuUCmwO9/mpIzpm36sP3diI
iA4ZBb7XXExAnQhVh0j55m+9DfPLJRvjAvi6FR2picSSURkrHtxxcAukNF/HMp+dakC9gf/FoJXg
oNSPh49rC9XcbfsabwWzZXFRp+kz25jHULmkQAz7P77emRXpCtMYfY8PJ4M1+SJRa4tTa56NWgT8
j6jYnZCKkehzPgGtLkdIfwpjb5nvMo80KfhHIQ1AtNQppscg8+wAMToOrpeBJOK8pcM6TYInWyQn
EvjV6y1zcxyh5o75VNV/EOdIInHQdGVyu+6jCPI+TOjPrD0lGH9aRpxqdempe7ltNzZd/oDXSog8
eSju0da8Xm6oDm1B+5D4JnLoqngc5sCBhMRQYVu9q+4Z9J7Nk98730s9QKVVe0B2KaLkgKMx/zpl
jVEN1FlHMjGxf6yHwm6xkO9ywpp4ERiCHQGY2vs1ddcNwx6kDWGDJ+ALM9UyXGACN9k33ZFh6L2N
ZCsTkWfw0cugqUtE93fBKh5efltgRVSb1EeDJr+X8GfhETEqM+YWfUleDO8D6tehNoO8cp0cevw5
K1j0GVqcMS2SDkJcwwbmNRNcE3nPiz7YX30axYl1DCawYaXiNL2xC5Fb0biPChXapIMWSWoa7QCL
gCQZiTAO8TCpaJ/AWSuZPhw0b5nosJyn4eBxif8v4xvCsc5j4N9mmve1kpsm5YOQsiuDw9unowUB
8Lag6sE5FipPqCveO/KgolPX01qKiliBwl+lW4U3ZscVTzPVHhq+yQG18aPiXyteL7dOVHgL4aOn
owCA8oiC4+FOlfZ1rPOyfn9CeaH8c2RJkbQj2ebr9krAEbW+HSxCMlJmizjDjrtweEp/guDko6SO
sXij7cl6FhxPkt4nFQ5w/RF5ChsuO5vwahRqhhbNzmXaxKcyf96cr8jeqRGZZWqewm/uEhKkrkdx
3dqxx65qPD3Eo6LWKZ2titSJgP7LYFfeVrZqpySXqMwfVdBFy6jqGhghOkxsbLOApff1VHUlJMG+
JQWlIrjUEFtzIvvdqSKP6M0yJe7icruWFo6+JzsRae/UNqnk+NRwQzqSLAOSEg3I6OGfh5McIG0R
B6+eNmFaHpL/71WXVmZ0q0gnSQQadO7yQ/udqYThcwTUhZZR4SDypo+g5DRnooVTdaNTe73q+c5e
D1u7C7gOgNtziTIQuwfJRgjKgNE80O7NQ3XAZMbf2hDz4kSP7gUGgSrORz0ik2WzN9vDjpR1pzla
IgWAWgoZ9K6u6LEe5paPK1UlYJERBtm2hfb+VNZZKuK8hdYPdUf9adP6sKGddIpFXdqlpUIWQryj
mRe8MO1dmi3fuP3rQVHCGxr73sHWkE0FkSI2emufPTvlVJZnKQWCaizWWPJlUmEKE7AMZ7siGrze
AJTb/LfRB1RnM0uaxxrR4YpzXGlfYqCjfr/D85UMEcAENH6oyax8h7mVhvxItBe3Lt3cr17jFK+M
WhaWRedBXd/3Po1PTamBDAjCVoB1ED/0pIfUIuPhDWovhip8KCaptt4OaqNIMdGEdzTlewybzq8N
lnmKexj0LtV+ZCHjKgla9ZOLKFh64nX1c/+8+voOTsY610UxxdsT7CfM7FiywSnXEwciBTJ3xpQs
NX8swiT/pt2PxP6t5SiIoJ7tKp0RkcrOKL7b5CZGxXT60voE/14Z442PSNTfHpno0MgiTYZJwIsY
Ng7n0XroWpikXanhqTYVwFGg51gNLEC1GsHVdXVvPAs6GsuesJfCYURlYDqPDursVPQA715YFd3W
dL/bSRtFsIM0yghTFx31cX/wnf4qO2tJkwuUdbTBUSnR31M0nazyIz02jYuU7EFcuCWLo+BasZgm
fPzgM5Gi5vvhEONlu/0qFHBW+Unz2APkqOAUqooMKGNFbn5GIglIqzj4rgjinwRRghawSgNC/Y0q
VjVOi2+TeGIqc7T2WtD5uUgijKI4eYLCvdRVsQoyE36dAiV1zfc7hFg239M6BN+byu9wgfURVnMN
WmdX5RiHNtQ7SQLzSUcNvS5SBGERkQSJHo1Wd69pa79K09L5S1aLzgCqhjXCF2Dtq58CL/IGAunH
uCuLTpgeB7pIC+8qHwR37Zr7z0BQDBbpNp0OMp6o75kMqnOEV3QalzppIISbR6sbk4DMD5ae/a0z
Qgd9TTFdXS6GHLvIFHliy5/gqNAYCbGY5GsO3LaGQrfMEa/nf5cKVR6Ph0M295qsx6Bswuj68Zf/
l3xF4UYwNxprGSD3+BfNTykW5cpoZCxgCC3culeSAfTECD4QeBPWiGtiOgYBUyvUTQQulohjrN4x
iu2JQWs129IPQctQtMPlatDxs95KcbGB0g/ruOQNmRBcOcGAhKz5zGYE0E5aeuvjDY5igU3es85U
dHriRlVaTsk1ywHb8er4r1235SyfjZ95YE0riyfJH4Ku7aHhCeBaNZbaPkqX2uSvz639KtXvreSJ
SJuUoTUdK74llt+YBqcx+gwFgYo1ih2DcvyrJJoO0E3Uw7mZuKbcgnGRNqiEFYusqT9RZGA3Jf8A
Let4YTL1CGy2QzCrsbhQbTv3S70o9bGh0zzdNt5SS1eLBWcXovvL7jKft/fORa26fA6HFfcRUOxu
IIKPqJIRfhFQ6jmmrO1shq3GE/PJAvSqH6zUWqaxFeHqIxiTe3dazJzR/Fo4gUO5WmvpmUfc3oJV
3uJsnzcPhSvm4ihZ8N7YgVGYVyRnDHQBlIv3u62rnrXTy68W6G0Gq4Ck3FxOabipZZ0f/IMXFTpZ
/hLS0hiqbf4PwWotlklQ2/dk4JqX6gWxEe41tMSBcP5AR1K/2bZeppkfG7UGpqhnXW1iM5/aysfx
szwpmuhol7yxktEaHaYNzR8K4Cmtyq+IEmVVfq27XFGX7bPatoJai/+kBlwcoD1RI5sDoBORo4zi
CHlRzKx9lnfgd0onsmuHzZjgYZQLhqkPGD8ffuBa3uQPiMiO6Gsk+akIn9HqNodKarkxY1cJwq+I
RrKfYdUOhMWthyVqDn8Zcu5EjX/+fZh1eHwfhXgO4HrmCke6twMrXP6moy/figZLbQrVmmGMxqh7
1iLhPLA2D1a/OPpTvhKSShOTYFhxPjKbIkKuQr96p08pG5whEIWHfc7YCl4UkVScqlQ8e8kaxEAs
wj7pixhPwpFhi4l9Yn4tZnNz67ab2xGqcI5R12xbjMuenT/wXz11LoMXzcPmhGKxBGw3Zck/Vky+
43wXPo+sSZkOjayvBTEa1ftgSLEkg8MgAubgHG3+iHA9edtbcRTpBD8fbQ0mhCPijKcuGGr0lWfJ
TzOVYj3QSNjG9qLpSN9nt1IMt1kCW7ARJAIjQO84hxkOASc+iXI/4nAPI8H3KbOTMj7ss0ALdKXA
8Za7gLBmkSmJ26Y6Ia5n1whWN+3eK6+ZzeIqMpskCLGKqWf5+pXjyPXBs/mCBxTD4fkvPCWK+uN9
2OCLSfriRgTQhEard/yZuGxLW6LBFo5254n3iFqX5cafrbKrpldkEdlVs+ZAv/bf3xFyAuJc92YC
MOs/5tlx9rbsQRkJU+qj0s2xTa8rvBeh9xlSkEwei7beSIQxLlDdxM4F/ButfL6X2YqI50Y8z3+L
d5ErmWk3v15MqpRNn/DeH2lzBbmzG35VPotYVKEpyojX63Vxlemxy6MGTsvXlMcWACgmSeet/tah
MlwMoNfpC/sYAgEBpynQq9KpFzGv65cmYuxApnncqh0SLJWuPjvz71ecJJWIjJGGaDiFEZ/obhRC
Jk8OVIHGkXcWJnimkq9dVVTlfHKW44FfADZTFXSfl0p1NyHdJ9QAN4+uuMc06uylcMWEp1BiLQ/l
6zmiC8ilRdIOiGJToAjZ/WMM+hBvRvX9RWsKkHTO5sTyUyqohrKNfEzqcr+EfrVuHINo+PIdGc8Z
3lWRQIfZ0D275hbwkSBEee9XecIrg19ZtqAFxJuWjoe3t4CRmCgpcJibs53U8UCQKIgy1SNOzOm+
uZvJX29Sz/w45SUAyuWUhCmAeo/Opxv1AZkjakLQAm+sFd/f1OKGkttXVa6EnztLc2n+fDcoxUpc
sdAzftPo4XIX+kkceeRfPk7EWsCVrp5fASH/deuVwdk0DmfF+zAAQpaJJue+JB8ACNjyuTyZgPyB
DXj5ir9yO7WvWBMlBCMp+IwMi81X2OGM/9oJshcee5fj0krZOwBijTM6iiPyxaGLSS9SE5Xyd8Os
60PvP1ap3TE1Gsgc6fVZH+2ZjnLGLoSBnbN8OJHuo7ve9pZkEr4a4Qh12IztNTZVEAnLNjguPVZ7
8B1OfynZCmis9Cc+HhLQC71p6x+V0mGFL4cWjhmxRqOzmBRJm1EAVyEClRPanV/RzPyhFAMlSVMi
UuEfs7ey+0XDQ3h77S+ScfxWPeVtkyKZgmpFzlBWuixcw6JvdVJf5NTy1LjyCj9+MrQh5IQkgnMQ
8xNksHJHiADrXZMsB8gAJ7D29gjGJoJloicPb98NQxCPXiFRE6F0eIvW4GNcdiXlqb59L2+rSOjj
vS0EBGErhTBQPUUJ0iMYrKtvtvS7GqsCMGfDdAB9R7kaHt5SvAWBoB2+melqxtQed5E0YhfZYTaX
Ogx5M4XdjqE5Cl6fbtuPfrfsI94Jc5WlbQCMAtB5+naDeuJMmUIF9cPFun/5FW2VKKUazYUc81o1
EK0nx0OebWX453qkshQWupW9ivwFajXYAg9RD15vC7FiyUz0x7zdeejYFO1J5vcARoIi1KkOiD6B
I6grHmIGQ7xWALnMeopMOWSH+dtepvX2do3I8qHAXUIAVSb50mOFFD8D7wy4f40frZECDD1ZnZGj
qMosUcYVPQNdG5VaJuzHXp4Ci2TkSXWI6oFu7Mb2IOMGobfDF5luiPN0OW581TP7JHjHrRTnWqux
pSpMoQtyr64wkZgxzWX+fKW9YRNa/dR0J3+ZX8yeOxDuc2OOY15ZlSlygGAWw28kAksmskMBSQHG
UziiPoFcLhbHaX8pNLtDkB6by/re2zkfV3bZt8WuE4QUq6821TZ8wZ2WOR9cXUvZBqKKXipcmYWj
Yotq2KzOQCmq6xtfdKz327A0iV1HE1SlyJstfcfiZIrpHGZT2ZhIXGJ2Q+4ALQDPMiDootHa8/J/
5nQwCVprqZ+Jy13tOU6uo/0M8iJH2CKgUTgDmMhvPIIFxclskQjS5e3pUAVJ4Mlvm69wxDs+ggUS
oYymQv0/Wl5TVVSrTbjC+ucnjWnXPE1L6wRz4H67eLMqERdykolbGsQu+9Ir4nsNSGxc1Qo/98BJ
1Kr282h+rFLYuLGHZHE0uwQkixk44S6Ho2tL2UlCvcZi85ZzjpptVU6tJOoioqfUOU53rCioM/oK
vacYGeL4J5p1mddWdhNj2i7RquafjoCzZvTkgNuiyHJr8BbE9qQfq53bqw6lnnXm0tNd1WQeDxea
jTLu+FVkZ+XEJVxsINVeQKjwg2BaWlZUmhE1ddetFLuLVXb+ODt1gHudSlUe8e6x5gy7DCBOI327
sBLCp4fBkp3xMnM4glGvMFK4/q1NYeWGXnhTAR8gY71UR6eWQw6cceCYTN0Zvnp6U4gj60mSh5TW
o3DRYv0zCZ187GR889nrtCRaoa+pTf6gC9OJOZtElQsNplZ3FkmEW9swAwkBdEHcVLU31C0p6eF1
k+LlpLyxU/eHPtbGUV5Ww0XlNMkIo3BKscEY+1rp48JyHIK+w4vOPdlUt2SjDnLDyTeZcdko8ACG
uZY1vpxuz/aR6NbHwlv9j9jUrjzBTgiWGsGgvatuRsOsf3+EEgII3EAGMl/dOpBQEVmxreuSu6im
48uKI/FVW17EX9WEEo8ih0NK9zcGvLPX2ps9y1NFisMKBuv0gI9N33D2gl9qKw8NvJVieMkR0mIB
Fb3aYzC5uv7T3uwYx96U9ductTPfUxd6qXkIiVsSeHVP/ebmLdDUntCI4CUPbj4JI9lA59jRTave
xKYZ+ppK11ZLR1NvwauQ9LYMT8bwHl8SyWvIF7MPdwCfV6+oG7ROgSTNuFpTwtWZ0gn1hVn7CHfi
j30eoZWfOwdjWZHdQPv9xauQ/Bu9DqF+g3GI9PcEbA84JdxC6TsdWZzzNKwic0UC8wFOqKIjAQMR
HyxdtW9QR1aH1iw965sdHdobeWjjE+NpExZJRwU2O9GrFNf4SvwIXt0UuS2QUduGSGZeKc0yf8P6
Ip0Wa39+Y9HYz4gCvZvIY4GSLqhQCJskY5J3j+pEFLh6J9oK+Ag3PjSO9M1BC7FOLCHGPIPO9eYN
/QEbFJiP20ev3Xc12ag71ymWnTw/PwyB5z5fb3l45tJHi75BsweHHyERW89heOI+doQoH3NRboKJ
XUqOsVudevgMcqUz3nCXSeUwVCZKC+XSNQy5CP7PxpPok7bFUiXeLYVFJKPVlZHib/21usGrFtOF
upJ7OMg6yhzefrmYEyBAc6ztoVoCLTeC1k+j1fwr5xSoyWWsNhVPviNld6muREKNEq22QKpdSTif
/xxJ0vpPy7M4D3xJX/tmsxM+PFHDwWw9cgRCJYNM37ifQ76og5Nctc2Z1R+tZxrHJpQfSr8Y+7Tm
+ZgLF0JzLzz/WYiq3lOVSiZQx3bPBfbLexr928Oe+O+mFFrDoHIp8sIn+yjvLZXTD/hkL/Dwx4c+
taMhG4SNSxwAiwq8kUoMR87Ahz/O+vFV8BZO+HriOWHb7iUHh2F+pArfyC4YklptMQO8PuXzWKjZ
y+o0vckNWmZW91tWQC1cHPS/o0LAWl2LSMv73l2ha8mCI6iXdfFYiAkOeclS9Dl5AgUbngsrmv52
N0sQuHwlNJgamvGxgVRqfmkq7l5PNTOMClqWM14yHPPmvKHUH0N9FjkCBwYj9kUQafjtL4JBSSp+
eCxqeyQhFH+tcaZF/UtBiVsoHj295oS5QPMvrQ0L2bvJXemApXbbo00jjPJtjfEqU7AhMfhf4b9q
ulgLibJAX9g71yFImNPfLJ8srK0FETWXXa0oSbA8zj6d6baieVTppJ1wJR4SmhykxnnUFe/LvITE
Ck4NyV8K9EoVsJnB+zYYYxDOxmrgeB4/njHp3aHUB96r9c5PMU5CxuvASiBS94Ob1FXmUlWxoqEP
Tg9R8IguA5+xJ+lIJ1Fdva2H2c/7N5LvuAPON44Dky2llmJO4qqsAg72DCk9MFt/tR2MUkzeaScb
P9+be7L6UrTtc7LjwiOpDmAXdpcbac3Hdj6zdqMXJwno8xy3mKEW3ego0d/qlfX8sN3FGUnrce3i
iLlcksAIpfFeVNhNlUmiUv7XrXrCLS+8zrEjz72Y2wwGIW3uCFsHZTghsZJkCfbXfRsyaEcR62Ij
5g7oec6A5/ldVWU12HMAGGf2pnYPYYVzaeKvVjEDtKMf3LIZmeBsGOoxoqyx/VFPE9nxLBK1xnyo
DPcXzYbJXSY7yeOKog6BJdxa5GsDHQ60DOUIfYyCG5MR4hA5il4pRmGM5oUaeI06Wzyk0+JhQ/el
/0nzU58oTsvxa47MDMENDer1alpoHuv3jd/cSD1mssXzm3boNTEz0O5UFP9OiEDtgTsbqCzro1JJ
v/vABeNWzTJvivGsgYYKAnXLUbNxvIViEl51V8xWKmHxKRZFXqxnRI1Ib3apwGmXrbauEgrhV7MT
D1O7Otn60loL3jRZqJ2tId5T9+l4kW8IKH6bObDTsfvXyznQ99YAAX1n1Q8aBc3jg1hitBX5HxMD
4C3QjaTtumdKaWUOP8V/5oASDE+sMdjCrFTVOgc8NLHoJbttNKc6wBn6JvTD2ukPgMrpj8OeZFXr
w+NMQuarJRQXldBpeKRH+BkmQYe1E4DLCvVnXaO/0raj9e137aktU83A//NZEIpSGZwRiiyHvAEA
kWnbrpxlnnEb+u0gck0Yh6T0ha7A6e8xjPCNzIS7gpVgWi5Ygxs1lkQFCNc0VjhxG3gsMoop5ozP
v2WdJR/CjrWldYVeMbfQKbN5PhxqmUc+Q8d16B88pWBuotXowh/3UfMvh3A4rbRRiw3vN75N1dqb
3M3wEsy7j6wYNrPLouGmB/atMogZ5DRB43AOwhQgq3bj7EhgNuNp8Tkx47WfkWa8ngCKK9zLIFEG
njiVBmNx2awFEncM2N/rLAzMTROlW2kRxwjrZ43qaCPvl2UGzuPHuF/b5IW8BlMLsOj2qGVlR7bk
ErXW/H7tkM1y+CylG972zvBmkHUpEtVV6QXTgd2zdJIXKUU4TOraCSzwivtzVh1qMz45ihqCGHzX
CDPQ05ybfmSzID99of3UiT0XXDgtB5hW1F6me5DSci5UBnNKQaXP2HF+kaSZHyFGcQT3dWvxw2me
AI94UwDup5SjMQTuqeHJsdLzmTcxInlyRssXeZ/UGW8on+pzNyz0FTq0KY3OjmhTT9B8sx4FG6az
B9YVHx46PBxPe1eJac3xJY5HE8JcGLZAcNiDqCddfXwjX88kMSZYdpFqYHm6aLR0lwGaYDuvhfoF
h9BksXZGLWcrhrVlBd1g/l6IPO34n+sXzPveXXpRkWCezParNOqNNb2dH8QtoiQzddf77QEHcZ5S
mVcFS889nm+7Sc18mad/3wQUbXcgSohJZ5npHSWNB1b74k/BSG69hXrQyLQfSzVLzI5A1NJEmFxm
ArJPJvDECCVER1NTOJVFIqITA0nxpqi+kRu4TyXf9qQ79xVAWrqutE1rFeie+ABX2whjhoi/nHND
IoNBY+VtZlAZUqVmLZwH+SqQ7lDhXr3frXpDe9Wb7PYT04z8S6pmAz2lTzw3gQbgdFjs7u/gpaES
l6/TzR7C18eb41y+iOAju9D0/vrRVsqCe1/4jZewe7VcosRYq2ThouNwcZx3NBPY0hWWuOCE37c6
nzH6ckOyfnxQBHf4a7CUA5Le0WffDCMpIPTBRfLQ0ZmckPNRmpdjfAqY9Dobm5sbWPEQP4Bg7vFK
rIlvR61PRurgXun/9aynm2SvT7FwTb4Q309FH9kRSKPT5u9xT27aR62KoIO87sBiWoNQvyU0OHuE
8FtF6enax0FivexeneAdQramjg30GQfQo4HCx1eo5L8P9KnPU+EaoTgQlOvPGsJLlriIRQ6ZfNlk
6T4Jimu+gTLZCvkV3JNUepk+fIqtWo+j8lVVqZ37MN6k82Xo1OMK7s4G0LZgkyhZ/Mfdc8PtMWRz
ulTR4HhhJLF+9wiKPUw7PtOgBJeevLA/S3NrKF8d1qAp4VfMyct9WsWDuuDiVqRXjEeahM73lsO8
yQx3p6kHXvpqX5ZwPaWdJRim8E6ysPkbit1xwjMBq7r1HpJPkn67IxuxPj/lnFrFasLpeaUG5i93
lOj2tMdJALPRo29uWV5a5q5HcPKiE9b5dDDJ8LnMaieCKQ/oOYU5tzzttLP14aWn3JnsQtz5myBA
RnPeav5c3XNrPUTfTxS5uUGUpLsMMMfaLmNCN6bDM5A07ebEgBrCV9oXh/PI3q1MTpCSv3oNQtNg
s/yid9jNQEbXYAg7zqSN/eS8K7CDJfNy6yZae7j3GYgJOIDaJyIp2s4EWhF5CdjAokzJcB7tFV5a
hGmzQsmltiaJp3GBL3QCYujU9z+y4ukwqbUkKrP7w5WqM0x3RxFKi2xw2lmYIHQHhHvbDcjE+rTi
gwTj0g/xa9H+2M2m1VKqdWAEgqCDq5QgrPVgLbJ0i/54WXmtqkRfVVychnXMc6ErvYxNox9uoQIq
/H5Ikh+CJL/z9T3MgedkLvTIIGFyWEQpwdrVn/xvr2j5YWO8pFz1zvpQYuXtWyxhpAaEroiDaN0i
UhPULyTi2bJgV0lJydRZbfF4uraJp89UfjABdqZusy+tgeCxxNwGYjuh85T229gQB8x6nl9F5vM1
JnbQuS87DaUD4aaeKd5B+6IoIFU3bO9Vjt3nn23QVpUGlcxxZ1qWZZdpVmS9yqksBnUiw+UsEeER
dwkBBNzkW8cIPQ93cKMcce8okW+fAbfeiV2127Vq8lepUrZDUGKiUm2Is8aP8GEQ4yKeij0R3gn2
Bn9swL4D4XATOrWE6Gi4YY/WUwmjKt+joZjBE4F4auvlMQq2DTASIwFIgEroT0rrYl/MNqbJXyrP
oV9OkxQzsWC6y+iWqp62G0tHbovqDBJsLVImuV5mxnYSLWKyUqvxQx+/zDq0lOOHDK55svx46wxq
7HUR2yAQLn0gIfddnhhmCNL59S3FhvDglvI/zea0asBsxmF/KBDd42Vc4iwZAbYVc2OodEEYKgPZ
TQgvs6cjyuUhypiFtFl6whMHax+kaxywVRR/H+oUqCET9fy4lr8xeGAB3E1AYP2or81zvtr0XYHC
jhmC51IaKMbsYAbkzTA8vryaKS2zEMCB8ktxZCyrtAwi4ymE4UA0JDCRbd6KXmSgUZ+2FQrjD60Y
TH0C9bDySopsHsQfNOC3amAaGUdBuWEGk9M1xd1MfF+AjdPqs+yDNwoCuy0GCoA7g64iUE5p9h/8
VtjGIqrr0A5aa9k/PENbY02A5RVINrgtg8FNW5CXHnW23gsYWc4GzQrIHXLpazrDaUbxL4tDCn5e
WPck0i7D8RENg3LSpkytTvoKPWFaA8OccOexuCzRwuH/8MBXHuk8wSZ68W9s9Wp4XV6b4x/DO2EU
aE5zTX8PinFEX7v/WJqgJ99yD2VSEw17MewVFNF9BIqJwsP9Nx2w6lP1YEOZW+cHobQzq8FZNS+Q
u3UvCVoFwP1kE/M9FXqZ7eQL98TRDBr2oHmVlCeSprKPnwR/dM0vVp0RkAu6dC2N/pFh7sQgvC7j
FKDd3F/q7YG7HjNjmACGPrhTW+KWGwmhCVV+Zs/HMJCCf8T07W5v/IKTUVjxqdDvx53lPQ3s6s4T
6b2KYQEU/2XRoBHOAI+jkamSUvQrP06/9EOZ0WaUO74pYsmFMR5nVk0vmk7nW4BiI8WUDhpcoLmj
bxIhCSGh9StJ0y2K4eJzaVCT4/7y+CyiJH1Sus38N4Vo8JexXErm5yQo8PTx+JEpDGP1owGJmxG+
OQfPWdAIbYl0s6YYahZojj6qAnIYzyM25MisFrrq+lUT9SxYw+DAl29V906N9f524kYDc9f4KfcB
Wxho6tlhtvKmdyIvL+vhpCyvXAg6FotnoTjUQfXICK+uY9A+L885D621j6iNlemjCWJIWlOB7Aga
bmDmDTnMywqbs7DlK0chIadi3B+wGOgT9zFT5wPrC7vFdkb3hI+xkaY7RwXmsU0YQkrabole2vAI
Ks5/2Ng79AlTIw0b7jpmxXJ1R1G2uOwY+I03OXAu9r51sm0lUuJCA/MYqEJnUTvv56VjodOh7vSt
D+E7Kx9WlhRpQRWNZrk8xUCCiXZX/o1fxQsIE8ac8ePB+Eh7ZPe13lk6U5928+qkZHOKeNve3C0M
YlaGbX1JDrwsOtvEBGSKV6VheH9nH54XS9ZrVxxIyoQsygWp/epa3zvWDnwWnWvt9gJiCBq7QGc1
NqtLdjZzFuXI+4UZ/u1qA7fMCMW1xRLURHMpoErRGrYNFwbjfiwVgOeyKeZ/aXQcb2t6/JHw77UE
TqOv3H8MZTxk3eDiv2bhP2HwkGVINF7s7nVUf7WFzSLkvktr0/260zRd6hX7CWApKOvO6xApzGhQ
pnebiR6k0dxC4y6+hCTs7zBjMxIrHfkBbhhgoPL1gUaLjvwXQ2E2mHJzWxXYDaYR4swyg0nZ8/p2
4DNjCv6rZAYk3su7CHr76JJ3wK/LFVvo66tugI8iuqPogPz0EWPbHreS6AUuJ6y3PuMqgDPhXpkU
Ol9X1lFw3+h4XBDREAz2Y+AxXwZY8FXovQYsz9IzBcF9n1c++F4DGDPCKA13oEK/zqVgGV8rGx6/
TCSu/J69mYSWUZfV8+5NhNymhEzmA5d6LcqyD9aA7C0OcmigGEE+RV3exS8ENto40I/4PWqDIeLn
azbsNmYSPbKaJPYGMZf4+CK/IM9qNVJllipM6S6b7pMhvg/PKZhxz3ZeKViYkQ3+v3Lk5qLyQG6J
FdR9nt2xEDVMqLiuYdp5sKAmHZsM2WhgTRw7Wt+8R/gkraQlt0uyzs7eoFgdPmQkN/z5TFEGQ7pK
L3Xp7pWWERTFObe/E/ODFjJHEZ9tHUlEw9sJINP0FM4K8IXINM7xNDOrsTBxSEmqcD2Y3mWqtb6n
hzfKPPTphHhOEiXKNxLDL3LeOfBi3XS64A0dwg6/DMcasGVai2MLx7TFV8SypswunoxjNiKGtgr2
z5Y1pifQ7fCY/LGv6m3dbhstLJEhjzS07bm3/hkFID2ZzzFDOKy53o2DooSKF/dxR/0Nn97sRv2F
1hHoqgPiepogTtrvDGog+Rof8lkOHha8QxLky67EVVEzXxhv/i2CwcbEVm1sDMGV5jKkxCqIS36i
XErT9J46QH682/Q1EclRDrTxQDhMd6sAJBbIk6VN8OqExYANAQY2j5wI/LrsA/zf346P0e84570X
5GBM0/IZcoGR6hPaKy6plBEFFe7WjuS6XmgcrZI4vo5vhsH//Eagc4e5GGfEToh1pOLKx4lwbxlz
kEVCySTV0XjEfnowCEDM0GRoSyzv9AhNPTs/eseon/QNc+jWm6eZPaoGbT1LLbbwj1b0xb7A/znS
XPnzVKabh9Pu1pEtLmV7LUulpOo32TrWWvf1/BDGRo15pzLeKBVI0PXXJmz1QA0ESeh4KYXBMJe0
xo0Fn+crAdU5j45U5ytlLM7sh2Treyg/OaFEePyIV/baHuPL/NmsdZyY+6y2OEf/B8bFh/nYI2Wd
/J51fnnS6YwfxwXhfkoCFUMUWkAbXqD/QhZYLs3U98aUnjinlvm/Jl/FnlK0cwDWU99e/ZtjM5JJ
ZRdO6VV50Iqdpo9XAdNnNd51I192s7tbEosIlzkwEF9LqBzd2lmAY1B5/nEcvLHVEl37FzE+ofk6
QhDDGJQG1ZXUwJCa8ZiHZlIWVhiRpx6yqIlOB1+JKAvuDD5uYaMLu3EBjuQT/6mmc/eJZoCgAtlb
2s5Gd+JyMu7sUUascPfEE7fAEWiKzNF8kNdzIpvNa00t2ah+aQS7Z3J/AHkgMpXzUB1fWDC5kiVQ
KyzKcqDwxOl6vNOOxVJsuV06Cco9iDXyRSWyFqvU054cjEYoD5zGRX/ZkDExotnLdN9KGJJhZ+wY
KOhFlG7x3P683VNOfJCqxpK9mAXS2KJ10Y+s+FGm4Rr0YuwU1c5ChfiAM6NRb7pWItWK19CccdhY
9Rv7Lov9l4rYmDpBbNGnNQ5gKDxjBATxsPIV4IUzu3q2h2lb7ZXdqKHMZtYBnpwFIzPfM2E7ISd9
ENA298GJEblDeZgihV302F1oUdbZX27nfu0po98+ktIs9xGf8L7t/M3YZ+NSmB48aaem6cZl9NT4
K2xMWmrl1d2heE0ofJBuW5Mn9ccJgpIhn8ip+TSIt5sRyjk3/eatA9feGKG7k0MVi58ppcaATqSM
kSbPu634t2EImdHpbql6D8L+Cy+Rz3QxJcwJNlWanzfmpuBT+9PmdUL6G/AQxdhSyc76zJF8HxEZ
/r2Tz72iXBr3MmRRPvNjtuhmU2Qt840pg+JH0J9iJYComAiZLhP9MMRaC/Vxubd3cEzZzZodNaxC
AYWsSSgdGjpL/EjwlFTYquLdyNudnUEx9e3Stpb/LZBZSGwDFXrUHVUZ+GPGR/Yapi/bBzhyKMRG
v226hnyhFbwKM/rE9+ZJBIKCWISRQjmU9gCKN4GxP4NEn3cS8TZzzIS92z2sAgG62U0C+b+eG94X
YoLVMHBOtEgp5ArzULUZpcoG2lAg7bxp6rU0+cG5SYA9hBv6wA/wGn2Q3T/EjvctYTbu91pvet5t
MFkQIzx9N6EHjj5OBPkIOBJy9BFXuaZofZRYs1KSMm0WV5MkBou7ASySjA9JXjp3it0xdIAgwloN
GOmzlenMHkQYcEDOnhPTF2DD5iD87/M11fz3l4Fg1363oCKpql491UdmUJND0OU25oCYJhrucdEq
tK6X4noUe3CR+JtnkMKkADtD/DCQGENQg8eWgjOq6ztXuyVMrthqRCncXqUgyo+WkQN550F9Xu8q
WpzuiMF+EWUNFIKtu8Dp/IHdiUFXCru33K9VYTGRKwD7knhH/W+uGJP0q/FVBmxvkd7nL+xv8b4D
lgBZ+VLP7jfmK4FFgSrwJL7dXx4YC/g/MbL2AQ6pL7IbV0bZOf1omxq+qpPZTCHLYb8oglwd/zTF
nraoZIktxmfkADtBXYaFh1qTaqRq5FTBm7GMMjCUm6dbMOPFp21JNOAbdSxuUmByg3jGOj5UagbH
TAcVpgCRZKhVDgEeFljKinx/5QqVTqWYPcvYhUdH3Nh1uGdKlcotLhjZe3IqL9B54ZJxwn53Q6wW
+IKgJbAK1yibGssTEElxppre92sMUPjkdIXvF7+Ip+i1E6pYp+t/oz26fnrRvJDX/chsZTE9czMV
/QU8gp9DpqShd7wXgsRopijPX1E+nLZed6vbZo4USMY0WTU0MRKe0cDABZwiEDXOvOtRnIG5gBxi
gvWVtep5L9egEuBrgM59K0IlBLQ+PaDoJliUJYEGAhE37ey4kfF0N2npsju8Fgcy3KQ5LSbU7QCD
JyYlwiSUt8FtOY6H78Zq1ma2+pKblbKXhRo652nlR16SG3Cq9Nbp2SqAcU42RT7HKV7302wIUGM+
T+e4BpLaRJuP57MFqPC1eK3dLABa72GofUXsJsTLHYTw/OkoUwkVu4wmFNEU2J+/8XIxTQ7CTL8e
rdxnxVnw8upEYCS81k80sRmP4/+tJDkKsim7GjgWBywB85G9OiAi73BGwC5dGVHn/LPCBZjOHfr/
kkdQAOWVQUZ9ObBp9MPJqIQuPLu8JP/esR3eJFQI8CAIQybVNy2Fyy20QjXuZPSkbX3nPQRYDru/
ARim0zJzp6siv0IbjUnBq+a28SvVAxYnhzs5go2V6A5U4uEHqSl0TPVJGyWV9WqIQicPV9P56mcI
qtezPQr7VvTHtdaKr4UKJbMfxigvPsf4OmXGsoGNpaTmOLuQWJTxiNCMxcjqRKZdkgaroSicfw+6
jY4FaOAz/aTpd5cPZ/t0oreMsism3QVa8oMOKYWf6dhtiebGqZQn9LrelAsKVFPMDGhJZ0a1mnWs
CPzjue8Z1XYdZ4FARrGki7RMXPK5gM+5JEE89NHpPTJ9qN0IY2h/MJ4rCp3Fo6jzOAvtURe//rYr
RTJnWZLvlrDBH2MJiGsl0a/pDNbg2UdMzRmdxjhGtXEv5+3YPFx3XH2k2Ok7LEF3IkDKU7DWFrll
mBdLVrLLeBrug2oWVYnP5J5VVd4M9I+4iuKzhZkPqZqB2WZKQvyDNXS0WNvMEt740rYadNnbmP2S
4mOP5BZffDHXqAig0FCqATLBn82MEm6mONUXWTz4ZdGfZNuJR97aCRicsuz/gn3Mgjju6HxvL9mN
1taOID/tUGd/Nr1FDp8+WjhB5+tsGXE1wZ6avNSorAtOwFQ1qZPxaU+d3BAnqawyxKLRjf1T9i7k
JHrNf6uBVWmGtnE1sxov73LyQCY8f+3poZtGfyJrowRH3ekfC18NFJqR4UxoCUBGQu1wu1GQPkK1
EBbi1b5l3Rokd22M2ny/EvKF1tTa6T0br0Nsp4meFBiRSFd3oetE7pDVKox5QuB357WUvVpQQSAR
+jc39VRXVexTpAHEWNVSizf6VRquIxGtmAJkiREbTm3kibSpASjvZ24lg3qhBPTQVnJaRs+mExPL
LVIDn5YiqPawi6QmovoDtMCGhlADOByAgxy8V2ZnJYH0GlZA5ommJqJNG12vpjcfd7QwTCjV/Id7
lmOzvAy1V+qGz6lhF+f9wUB5gy51hNuI0cc6k1zT+5kz+a5Ra08gg/q4SGVD12yfvI8HMVQPnfQH
ICBFi6WKHgGhckJfsK6HuHhqGk3qXwxcDEVSmXXbyzPpBnSu1K1QFfNsO4jWWmLeKIkmwdfirPM2
OX51WRBMS1ROSmK506SLSjnSnvu5kWf91me+WyHkWeMbO6TgHwddC5Bwl7KNJfK0zPI+Gzap96SS
w+zHniTwf7TGXdSEA9KbzjHqBOLYkDbXBImDVgQOoFiECgryz+llylm4L1GdEOjeUUxx8t4TrztT
Zdph6PT1RUSEzvzlu09/7Z32K8nRsu9S2qv1w5y1Y+XlKG6R+UnCDcAftE9uka+GbMOuSrECG5Z5
GLhwaQnVZVq+jKMw7W2anXMB0+Ni3Be7h3GB25BnevgL1hYLz+4IS5NFitLvnYnVE2/J7DjLG9Xi
GLfetJt/bF6TtIjuptgLx4OZmuL/KUBt1MGE7ESZYbETV3Z2419UtT9Ivtv2O6X0PE8pfy+lVVga
RjjBMn+qjZW8NsgrY3RiIamA++jEycIdybT1WMSj3qalp4PS0Wm+tY30uqDerXTczwn0Tj21rlt9
bmk8dbHay6NpyQmPlV4tBlpkt0JXcE89IUUo9VWMSrqGCx/KE6Iyw6nBXzFcWv6I+369MUM+2K7z
oFnqs4E7U4LWSiGkkO43mc51iCtzH8jvsyNexOz3uqkUqwfk+xBqZD8iZ/gSozsfpYbE1dn5OYK7
ZGzrlZ0IlT7aYtMeVvwcxRwZe0WtFU6ILbPKfk9YdYHow2mpfYCJojbEBPqM4qewE7jzhPdJmvOn
64hP343Cop2f70CnQ7wWjxLJP7TnCMwz/aATxrOOqzFxvoPNyyZEcwm2+3Yy/TOFwujDkL3SephT
7TRxEOSVA9zOJs/oaW2gPLnDQQNxE4E6f+MM+1/FX4TzOEsA1BwbMstkhuvdP1XRw9neOs2/vxDw
P5hZn2zjvRMoiFeGKzPYoTthIyOYSCFWzkEY0rSMCQu1SZq9i82f7kfcVzXgSyjMAIcfaede5DzO
NartPh8PCqC4G96nRjfucFwJwqo7vsnUnA4+S7vNX/eecwxo5SKZxiV5MBVTI1QEDwwqDQDjitol
AZ99f6l0focWetT10BogZQOBnJrsSX78dsSsL1wDTO/y+TQ3wjMPuMbGpplIRPzB4284jjr28Q0T
1b/n8QpYU7qquMR0ssBB2Yl34zOI+a8Z1M0LOE9KFCMBYexsFh9qzniEuGndmb09mAKCA/KrN7UM
envSkaATA6cLCT6p6ud62qlE8dwp4xKUPw/skNwqfe4FZvxC4uN/Oe9vDZoeICgKhy8zSnLlxbPE
wpnrTObQJwDjCKFgxq5B9SwcX90H1srb0ThzkAgrKyaMcMezL46PWHjUQ232+nefOQzBfeIPKui6
cu58P/0SGasFiz2/JO1Xb7ftbd7PqbjOaWEqdpNQcf9W2+5V3AKzFi2fie0gt/Eawebh6yzS+u0O
DIIER/cSWfxHdmaj6S0RI2niTXIxkiccuQqoBQGFrfGAdiizYAA14yf7QYuJXgDAHPoV8VPTcTGM
T8Mdsdf3zBCoejhfT2JbIpvj5iQCBymsihmDvzg5SlAA9W2dRVQLTw/18ylEfN+0yMFFvN4Ai+Lp
QOYn0WHW+MYuy5za8riy/Ymkwr14KYT3ZtQDp0IvRK1TFnvo6ynFysEy7VSjEqfmcFm46mXoZT5v
QMn0yjN2ogZk5ZAE00s5nRdy28S2VALj+3hupXqJmRuRKfG4TPYQzTxDzBDybH0G3KLY+ArbyBGY
/gon3Uvto4jaE6CW+CJnMVJDzMZViGSO0XXTPWTGx+TTd0KNzT9WsC1x4n7W6hvkp0Las+MD70nX
Yl+AqtepvikjqeJTtzEf1bI3Q+SkbJQp218M6tXW4CrPdtntxJZQ7WgNI5Q8SGE9cKxaJvIi0gWA
eGcRw7swvDkbS5yXOYwuH1yiGrCuOouBi1vxNQzz7wTHHoR13YoQ9vMnid1e8KdiNJvonRNVoA0M
FpeyUZtJcMaHjOLaTxqPfV1LE3bO1EFUJNsOU6FhbemHth6qwQZuMT0VmwdayP1rh8sXW2XbdPUX
x6L/FZbJVIrbfHyJTTDhdSsGSRJNX0tbwA6Ngir+NQjCj0bY01kbdsZKNC9XJWsidcHT9FyHqjVh
GuupMlCnLKprCgi2+WqwoA72YtT6rpbxWBxzFa24oKp88CFXJGmAYf+v7qsyq8g0dRqdrWcUnbeu
kBraYrIYvRrLp6Q17aVkojH3GV4gWLnL4IePXgCvJuv85CDoR67uuOu+czsldXSdskI1PeFmynVh
LXw+fAGrJwhgJeEOrU7a1FtyLbnaJNxCWcpBSgCbJt4fdWM/6oyQYpcZdlJ2TdFGzmSG1IRpgmKz
t91X/uEdBjgZf3/veXkZbwUx0mnraqhKQJGhy0BBX9458MMvR7gAewrVlyvSVUo0SA6EdE8r3SA4
dJT9oYP3bdb053A/Jr5npcoh3KEUk94rEE7tpCCg9CT251OWzMLA6Hj4lpdGpgbbAPJYd3WeKRC/
ae819/4Tsk3B3Fe/izynWC+tx9riFNRxbez4RR1Dk61UOSKK4hZvZ1hnsqMuDnTtfGUOezoh2ZSK
Sp1S6PlRfhHwQEQyt4cKPdihn5xvQU4Exa0BhnxrtoM7SCKmXEv/QL9SVwl0HX+MASV9E87kJ+mN
n8zKFujppR/Mpdi9DKRWGUQmPe5uhx9jYPzrc/LLEKgnG+GfggNqONTiYkJOX+pEA4GD1OcZtUb1
HtCO2IfpPIn/34hfwbBt2j+hFRe5fPWiRq6bg07Mde+QbdrIIDI6X2eQPYQVJ2weLqmvcjTxj6e1
PU858UGcJEYTRxCs4F4G4qf1lcvvrHO6nyijTOvgg1/iRGvpevrM7DD08n9klI0XCLG3RPyhliWs
DGtTMgkBpcZ6cgBe9I1XYgDI0adY2ZoNm2QuvRzEsfvU6oXF1bzaLGPX/KNZfL2Gmq4FwJgx+bhb
ZYEObRXjBSGdXJ9U1p0lLNajDRb1nS5mxQEQaMyw3+jl30gN5fGOmKR6RQlS/iUG6T25LphSXbVk
CN4t8iHnRIfIDjiCAgFhDYFiZhh5b4gGDyT5SHFgUR5wCjJqR9YIM6ArY4F61XcYzMNzCPeOPw+4
/1zs+WHKgRzWBjawmpchICMS5I7TjC9PRBIJebRzqyWw61vnCvMN+g9JIeHqhnAQ4cmyODE+lrUX
FnaB70BIKm9Qo+Vkg9QUowqIhiHMNeVeVsrSRv2RUtzsdEnsHCDnS42b/YD4o9dAx97bsl/bz8Nc
wRkYpvZXg7iHs5JuG3HaaGBx/Pin7/6tVXfsKjePut8hS4IJOWEbUNrgERfDNMtom8xe57/rWe98
h0J1xI9VHkn8uM7IU67UTdo3UCjb6yNsxz+2r/RDTw6FhuKjfbEJ0cYOWCV5gZQ+kYxIEBBkJRH5
oltGekDsnoTWCvXdW16kzsi8ksKT18phu3T2ixvRNsAkZRAvjZOYcv9Jv5Upi0wgu4q9qDOqhif3
TJabjBk3VbwBNWdN/xSfO2O+HMQbkTBVMHUmgOG0dYxt44YZzAJyFBX/xXvk2Yb01L2XFBQej8Cn
c1Q40rAhJC9XSz+j3jhMS2sv5fFpimNudiye2uJyzViuNKPshsvEGrwoHPQA1h+RZxTrWVRugyzH
bpvHbfTcLbN3U26khMiT5VMghCViaP3mV4R8Qd0Ke/894w9ZQsm0yNPYlvOSmUqLHnxNk0O3Lmz4
G6plAIaBcpwUlsko8BM7vGtie4s2Lm4u1kQAOS8WxuNv5IIpBXQu8wlZjJqWTG/JA9UN+cFoUy6O
1MiqlMMCQJXApqD7cpRDcaUKgC998yeEmGIBGcMYrADbXMjJW8TVVjpiDrziDWE5BK9V0AnGM4Nz
5hJsC/N0WI6HebV/ZVEVjhpeRCNOQWZ/lmT2Ra/s3PsvN+5RIJjFGKzrjgwJdTN+OiMsg3a92Y9K
8wrZzt/nTlsDF/rcvFMAS5IcX+Fzn14nPOqVrD/jh2enclcvNLZheRNzWAjDQAaXBtoM6DfRYwul
TseupGq14uk3KTE+gpsoVCVX1Ujm7kuyhS7T69/ginpwiYVBg7WmeynbhiIM4GfacUC8cYnZaLJu
alZ9V/q/br+OHrc3tCphldYbMWUm/lkQyk/hsVI9trKbNtK5D/pjBFTj4CT3JCMvF7LJg5UexC3K
pL+9paS3lgaM+XwsI/hJtDlGw031vMx59SrIqr0+IQGIeMx23Tlo7YbnK5l4ZBV6D85MNpkXhf+p
uxOkSUCwi4M78p4kv/rEcS7icyAHbIIbdScLpTtQTIPvBEUtcDH/175zjqKkiWILvKu7xsEV9Ayo
unagVTxiqfzwLJ8q31aAnv6LZyYY4DBpwv2ukQH4biyi0hZpyS88+QN+xW0yL4lQ+JcwHb5vEsk4
tGIQFJ0Ie2dcs00AkpHM+R4eRlXnOi9nivRou40tYBuZcStvltwYHn9Ty6xMWgJVVQcNbAlw+ApR
GFsLYnQgPN45+7J3wx8NqYs5XD1h/7IIervasNzDO7wg83CsNAuj9gA9XBmWNwyLlMdfpxbzmRsy
5G5yhizoDP3nKoyvKtduk+g1c2vd4ueY7rvw5ghFjpdwFKLYisAx0VhSYCPGWEZssAzd6c7tCudw
aGWwtyuXbY6Ph9ZQIihu453L9wobmbHzdgQa3tpQ+7lK+8scfXwijUP3KavCktjn34lTcRVoosCM
a1v+KZq4TqS9GziD+j4k7GFmq4cpdaojMKJ6bYjTPtFsGdDBd0FZvzpaCAAWaLYV+IJ06/sf1AV7
mvB6xIjVnvP9OXzOw+3ZwFt2YSlBvnXcPoYjaghCEpI8yr1VMB2JLhOiz7+KKhD+DaNtT8dehN6A
sR+KtHoD6C8Br07sWQb8eMh1uZE1LmacBlMQGE2NnFw6vnM+DUxx1vs6orn8aiPBut3ZY6nOMt07
hFSzIapEza9kXGzwQ4NjSB9ftXH7W15qW60yS3FmKHPcYH8DhInjYe3a46C7QE+CdzNtpHrRg5O4
qy3ncgPgVnV/Nih3NwL5CUmUDIiJy2SudE6osUxAyKVz/95DvmkgDEkz0Lj2U9KnwOEbBJaFeUzf
6kagiDcXkBvzhPja0HWIZv0Amvbi7MV/jAIZ5jNWZL38aemcm0zmcsb52wUhJXbPAm6BlIwdqiFY
6FvIk6FYDiABdAC8DvdRpHEPrzH/DLQZLOULtXxh+X+qm5AU/mZ7jWGhSIxkYcB1gaj1Klv2esYY
SzlSZXEIrd3jDBoz5VRoEUWNXlqsnnieizqXE8f5xG9F8IgPoDAudchmSZiuf0HB4w7lOxyod9SM
PY2LRt2rgnf05nL1JSg3wqykGTLcBY2kQIIu71pprEFftQtcYdYhAWd/ZWAAlGNJbut3dz+EMc9V
QDBj1/lj/xWUombMOeABCQ+aeGj3FgJsdYYVhV55w0woI9RrChNGgI8zyUTupBAt18HhfxCjJNVA
VBDDhhGwDXs/w8UsNeHhS2Kl80QFAZQ7+VxOZ/UOQjnNWyks/zAZQg519/bihJ2R48n/z78eDaju
ftKTDoAwZ98SFqPYFZyn/5mKEY8LV16mnLk0gK4G6CJelKfzTqm9W6rWHUESXKMkS1p9JYG45dGj
mYWt9VPBaw9lBUllJQxtbxneCzbWP2GLyO8pqz5t/CwjJKE0CgjujJHhEncNMTm1hObWTw73zKOM
2D4LDB9/yZ8Jp7JtLaz61Q+/yyQYNupFV8lFMlJFEBmT4JLOHo36X7CDmsnthhil1iPYSgBXWYsf
GjNf0Gdpn277DNtJ2TOyuhx16Ttj33PZrkrSbdS7jKU7UlwSkDwoBYQNQLOWjItnNeprWdJp+/IP
cVO3LwsiMtrf0EvEl4SK/Td8x4MFiMvqUtV1LFFsUzh7D6glRji5+OWLsPg6NlMNtwpbI6qYVktk
lsU7QW4pENY+hdB/1P7UZQRKqvg4n0TIZz8wvrBqGNOoYM7vZYHd5ZHWpWmExMAIySvjsmouVZGf
1eCu/Yr2xW6gjtFR3GBVaYR/W4mTMnGA14uX4NmlP6KHzZ8U2kr7e3v0pPVP1z37RIyovHv5hbp9
EESn9ddFaZgVneJGBYfe/jxkgC37TIABjZ6EE4lH3GJSnDH+DozfrNJB4+c46fc1NSGH9kd+LQeu
pX4y38ZVfgHcJKmI4ncpCX/aKiXKE9GFg8T2od2rlIyJmHnnTG/WmT19O9firDaytTxTtoFQAe43
J7jc0iuzxYCuXyMoQZKvn1CYn4C1PNPbCTXKc3tQ5flWL35mQS+1VlFhQZvfHQqTz+dsT1bEWoce
/nfpnDH+2mOdZIWhuVBnEP2u/jIShslyvkYpI/RmpjW8jzoe0/7Tckh0yA+qX3L1E3IFcZG4Spzb
JEGbueZTgu8547L7aQ+CwG7e0CdLqc1n7cEWCp4LPuxG5GlQZP0l11dffx8jtlW8BkJGYlPLNBcZ
wUPLlo/j1hziIfYkgkT/encWNDklwMIEkjs5y5+Wdwix/cG/+XHl5eWCqfWzcuviengQMZlUALIV
HBh/D4yyN54iCfyHuhXyvNEVrv4mgIdkm43UFVLJMOqjUS9V+r5ztV6ZAT4D2+x+BAAYq3VkRs6R
LIhOyHuXgxlvzqQjB4VyeJiomPn2oMQlcLH5mhMIDiUFUwpO74YPsD19IKOYfHBKsQ7jI3df7CWs
/swEEUHYYpyyU3drL4Sn0DefoFBHR0T9JE6lZ/0Z/55Tc9nkJVE2bu5t8IlrBPK5YyEkaFW4K+Vt
uGlnPyIg9Za6YCxKfs0kNZnOdMJhFA5M1xsUy09hAXGei/xkZCQiB4pe7YLwCqvGBvvn0WUqaSYW
WeJUJkhvky1TZaRm7DFdiI/01VFw1P6iRpg1DQoGAq5lU8mglqlk7u5KTWKI/ZdZjkKXJ8mg/093
vfaNQ4oDNMobnCaI8GyNjG+gA/zUP4UZX6lKJ97sNVYovyjA35iRBE3JhlgRPHmnuHtntDUWykij
tG1F077n8w9nqnC1IBkSX7lKBHqvMn4lBUDZBpDLLatu79iuOIgRzOoT0jds0WZbIy4BxESs1YuE
kT17yPZHehF8gbEBpUGdZRvvZ6RZ8kAwlVvAAP7JT6Q9fql5BOk+M+SxbMHw4bAYRRdPCaKwL+qs
FAA7jFlmH4Vw1xuBr2iChlYd6OtVlhds5kAaW+MpnY9sCtW2ILiRDlWCGb2vQCW2ZQMizAbDnmrN
kxB8546qNccE7A7bLx9TmKiEGBC5BoCZjeVYY4b2qExMu2unrfC9C3zaTOXkfi8X23ewo5W5azkp
0DiJv1ynNIa0FtGxstnI678PypkAkTmbu334VVCE5F+NsK19YCFCNh0zCiEaDGiip+RkWHHlI28a
OInI0xW4p8fTrWALz3b0sQLRooUUxTGEuAUQSsQrm0s35yeYzorkArpQEp4NFoj/EXN632KG4e6x
epBEXSDM6w+y/NrgWVWZJ21ir4HvklS+FDz68EH7cS8yIQ9GVNuSvIJZXke5PwtX85aoFhXKqxtn
6qo9fkPdp4K2yvIinjEafbKdwlRE9zJcsK/f92A+7SlHlCfN/PHOUrD5tgXxkyhhrEk6t1cNqbw7
178y8Wvlx8GcQpVdAH9Fhh9OjyJVNE206W11VJn3b6kZbJqgmLpS6iT8Mfz5DBTZ6FT2adfayD4K
SOsySYea3FENHgcMI2jtW93cVGcRVRHKOYAKXohv2ELpcVPXv8L6vdSQzafT18Biav7QJpQePmU9
6tFoc6VM+0bWaXVm4XPnkdA/LEafLe4A62OKqMto7G5Dd8ta/Qdw2Kzhc8vd9nZ+zAMPupyLdrVf
tmn9VHQvOG/h9o9KlDRSxuY/hQQn/oVDObjlx/4C2UYS8dEfZ8L/mmCwIhTlDWtzrM5ouecp+2y9
9KFa4Qga7/+fYxtd+WvO5rWIY/wdRF6ICfz/NfC2hDAxUDfSMZx5xopDetbVjC+Qo71RK2ajT/9E
bGvzbxJV68z/o9QddyXyGMAmQwv1qBRrqEusTeQw1M6HPqewxqRvd577X16HtkoE0eDKcNlKCdjn
OyAKbla8yYSL9uJOBvcC6pF2Nnkxhc39t2nxG6+cdmASuYubX6x9G4b3joRh8MG6WpnNAz8DJfXM
ChGXJF4WkjwUUXRljq9tuWi1FuU55Z30ntfUKR/2wernITJHux7h6j3k5qgNan2XHwEeWSxVyd1R
Y8k6FcZeJ5GDSR7v8oiJ65yfjnGPuZWzSJCF8giZi7y6EX2wD+URcETKdbMfThHc9vduyT4bqqHP
ac0XG6yhX5LWdhB5lepWiMYbKbNKV8RCNrkEYfMWEoMZnUgOfD2+M+ThF+5eNSpun1Sfq8f1Hd8T
wNqI9ksMDFdFbpl6Xif67P6WPswrvSG8s1KAtErtvFb9qvRp1xClZWwWZWMD1+L/lf4746O0LElW
JBUTlV/56zGUhgofkoI8TchhjVnCmf35rG8gIaKet6R55i2DPrly2Pliym8b0y2HiAwwvx0pB1XA
vwgTmRWgY3QfNBH34LswLKUzGpGeKLlvMt6J8LTixoHHVZrpLGtCpboJdvHy/k4ABLReAtNkifY5
ThcxYGIialhMCt8InLwbNbOZDvhXOmnS8+/uJCNv6zqjTcXlKus8v4/y5Rg+jovfhA+HwTHDPrnH
FHFB5ejUPZNZIAG/fjiE8D7qnnGEyy4VZJdLKdc2L91ZdEmBaqpO61GthwY0R4ZdhJ8wfO/P85Xn
YAONnpJAGM0h0TGbakhTTJCQ/1fKsB7xWoO4Wte54KCYJeHL/ScBJrzZkZBGyrujJ4+Aet31apMg
KVKguTjBq0pt+8LiM1nXs0MymmyiONN+rD02RjEKec3NLuLX3IUtokQB7As3kx7ttjATgNAQdRuj
eEVc9EjZ/dqAHwX/SUp1OKpPT03tzJ7qvL3rRQD+qH1JakeiztVZqW7GWMgy90jCYnM3Op1zOKFU
+dOJapHKqmzPqTlTHPY6rfwzwwopkBA7G+SSUcL58Iu0/nEsKbRylvUfwa8wDKpo8d/kLJUbJzO6
eQ/KAv7eqb18Ydsbee7zuRv6iI0XovrUszs8eqKt0QIvx4f7O4pL7ZapAsUbN//bJcxgYyXpHuiV
34FKtMioN1RFxBT62Q2euvzWZlk5/drLZCCgetoNNxoHqvdwFv9M3rB1s+qHVdJ7a3nr/4bEmaSM
zPdJGM9r/Z4Q7zhR/axMWfpCNZpa0dpGGM8dabKz0JBf9rp7Whp+xpl/II8d+23nYWUqNY9dM9yR
lORSM8uRvomWkItvyd61uxTo51PziA7Xz+gy/nX961sz6I2TQZN6pCddivY/ujqS6rB/7WcN+z/b
aHepAqrzYqf7S+CT6t8spMJizIdRCfySCGLAcylxihRfAjU4tfG+rZZJXMChsgMJpHhR1BE2eCtY
y5UKgh8x7RaKAqNobGR1tQ8iUKo8pkzFkiIa+CUSIh6etlZfQT6BJBQQp5c5BOI3HhD8NpwrRNI+
lDw7ha2fU6QKoJj9jRf5DhJnp7N/wBCTxSc89LU7n9n2C9VzMYniGPfxzLUjGwZwtQkN+TZ7bMpy
RgQ08Ni+abvXS1jwBfKT8qcz2ZYwEgywRIZPB1KJqUyfBX5i0YQW+qatsmZUsRKrc2Nq3UEjoAeF
HnX2oBfHSXGCM10IqFrkKOgRAYTnR8GdyPTGkb8fsP6Y3pl+rueSifTHNoVcNjZD6QCB4i/hNjLp
OkbdzAQKVR0rbNOmuBH4vMS1MBKcwxZaG/vDeskLNo2NVGpkMKfveEG7C0/GV705WJuvlxpadmaI
GbxnTn0HqXHN1+YOM04laUdr8G59SwJkQbgIIgqX4b55s5aXt6Gg+C3kgqzNU9sje1sN+yCF79Kd
god9L/Y5qZ8rvE37zkaicJ6EDrp6tn0JT3MezvjeAxQW8BOpbw5dzdRwFH6jO0mjBGY42rmGeNFX
DMFirx/UWeAoU3R3DX6C+L/p0MApDHlZmta51iiUsDCDKaJMYaN3//zFLCpPUKbRluvcLj5VSVQq
dlm9Ku88CuGIkiWxMGncFSlTKWtjuneag7gUVlP1/WNgHMcAoNx1PyaHsFIGouaX/hz6jzMQlQC/
NWusPNeTgv6FxirjW1T4yuDgNhOxZ8f8jolIfdTxZld5EWVbC0QOx4Oj8l8TZojbfNeMFDsJfb+N
X7sKb2TZZsG4xsnGtI1H8RFdmqyLbtj+0kTR6b21VeUgvuncgTntjI2NmWkbwWo7MEotPgk4eeBa
ohyFa/Wk8RoqOsE+NbLFh3tUDwBmomtPD5vIwdUpBtHpiC7QaGMN+0/vbf9NwuVNFHGJhTF2dd0B
AI8dHV2Q+srf4sOsiPlHPP45M7QE8IH3d6DKj+RXAYp2TViRbZJls5C3abBn71/4TgpoEz3wig+d
GIIDHhtOxXBxpw9kS4F65iVZQIPzmnZf17OsEjNDgtzSpSk4ji1iaK9b129bxjlXzAvQzO4Exkle
5+sguT2Iuzu34rDWMKCn2pG0cWPDOR7ruRo9IF925vJ0hjtGLmOI6YBvPC6yaBZRqSV+cRdXM6Qw
G1ec1f/e9sClabykH9NtorWowLi5VSQwFoUwl3THOibgJKDI+fwik5qb4VdJSDhBh1eN36kpHKXe
JHL1HR8ZatT6dmUZQ86tf+wUfL2grj2DmoI2Le/C8mFxm2ALMZMYe9ft43aRkOMHoc3auoGKIMED
dY0xOXcOb/rj44/MJQXXnPH3LwOH5g5nWQ/qdnT/9eZZVXizaJ1zhQQ0dawi7rAv3EVG1a7XnDJo
exSeT0D61Mwaa4m43oMsZqBA7PHSVxb6FJPMQQV1emVqGwM9a4GDOLEIU/n+XKEv29bU9AOyqyZy
aKF7Av7kfPsuP6GOuiuD9NDLsSPl1TJAh/tFdWixgvK6tl+rWxSGxzOgSCg+p2esSU4l3ka9QuOT
R67ZOsriXPTTakckFfDJfJhtn4L5MVqJEynuv+FFa/fqOwHLtNogwD4U5UgUj1ozi8o4D8iPP6PG
iIjeinTnsY0di3T/ZSUSQcPtTtDdnScpy0wZw1+M9wQnEXPy9ewS6y3L+rYoeSpbkBzvypq+d0oD
hkgndk9ay/HYsdd0e6/PVdFg95Qe+zD7RN0XIW5nFYpImDhVVcTbhU7ULAGBPX8f8yufOFmqojVq
lMXk1zSgvWu5iDo7GT3xH7awKqRE1QO3sst9DS4Sry3jGHBHS5BGRLsJTr1hhKPQE9x0vaMHVhQL
mJYH72CqHHPNEOM7RAJSIv+fENcWUvvwPhdUqHF9njAZ3Zua4Lxms2a9HnwPWlL2ObLP8dYCF7eH
usmE9OP20F6U5MPvIK+qxF2PSeU10X4mCd4ixsuIFWapy6wmWuv3BHv5k9Bwg4ze5A+yrYe8Z8cY
yDa68+5t8VehtfAEMIWEEYArNrSlGwXk23PwH3AAriAP8TPmfQrsKj4EBU7z9r3ulV+C3OCNdV41
ovT8hA9/bbnfH7nE1lAIO2MtF7Jx2sAPRAbVQNw0sMcfO31+8RSUEUuSgT0qLhVSU0qV/FIGOt70
T1CbSHv9E95BlWTXJBBtHKbijOZOuE+iagpXn+gVXtdSizoAki61s2yC0T6rWQDdwtXbq4lMU5L2
PI0NWuM4ldoXb6nAIX3irVIBPiv42VYn0zFLmTy3ncyIN8Ln1NphDkkIdnwoGWnqaNShDe0DVksx
kH7p6c2ndBkRfRWW0h9Mh0VCIYCnvBycoQnYwl67NLmepnTY63m8Jn6gfGRlUwd0bYR4N+077A17
zIfTOS0ei6J+1MnDst9qvwTvVHr/PosX7b9FoAGiffYC8Is5nPhjxnNJMaGTocoPgcc9ihB5qP/y
Lbg0QNR+TsW9nU5LAKyjGaxj3A3v2tgl+Fw+2ITpkw5yx386pHg7TtKFJ9R+tYRu7cKOmLoMu7x3
0TqL6FmdV7Kve0K4Rr1XzeHWc0KusQ2jrGQgffPaVvEtcdObQJhFcc3xU6VKxYsTL4pdxd4QLjMK
J8ClJUBvWo/KGw3HxNQ9Yi8hPi6ye7tPElHEweC+yrYZfEnuhrkQ/8R+IOWXF/mplNoNkkOarv8y
TjGikFijHcUNxNdjGWYCamVZdyq/QewfaxZ4XVpAFiQvM7Un6+QsHH02T3x32SxHvkgBcPPsMvdy
uB7nrp8o8r2VBTtFXV1MPgVEMIrczhKlhOTjwFTMMhcsLZs3ACgf2OY6u/iVcqPMsJhKF46tCVrP
uHphpzOEvtgy4e2lWIhg8w5RsJdYVFgyrMM47VbxEt9jekaXK7Z2kjsDpzHChzFbCl/qOsKtud8O
agxkBkltnfSZU7QnjNDNq3rziDQt54zuVuxHogb8POvDee98q/tmCwK9dDuuao2Z1OEL5WDD1EWM
NsSW6oSzxpflVPciljMhqNwgYa0x+CZs94kgFRfy9ws5MaZ5sb3dD7CkDO5xbAhDqQHdJywrEAWd
LQmDdiXgYygKdvdmYFxXRiNAjDwvo7M5kGuaC6VIcdGPsE4II94EpFsLYRVNqVkLdOVF/d/xArxo
DYNcGh7igx8f6gf9bW0NrtNFo+2aQHqdh03EzGSuE0+XP4UyOpWzS8EaVYDtbqTA/NhiGntEa0jH
Je67Cpcl51CmediZ6EG9sBqAdTm3IeFxh4d1GqRk29i/78g0YnC9cBKuU+9LvkQVdDaBoxw7gr7Q
qvofHAjzvAnw5eCKYOhJ2tCZ3sMNorjZoKKuMNoA5G/b7gbo2IUzu0SAQZhbGYzR9e+J5CjpHqvP
h77JaN6SSqn6+GXMYl/F03rl2zRBoNYlIIyboiUgHvlA2M+Z14GX9AJlHibLPuCL7GgTYJ7nF7QE
+L1cu/n8Svshtw4tlOeYeQKsVwP3uSmw15anNZEZbxldNdxNBKndmoYvX5R6aRsvQlcita5MLprL
8Q1273O8O6BpR4jQb1HU1aN5OuJ9uZnvVMqCFNTkYtF3SW9HgFZCwWrRGEOzCetoH2MHiHsJvYM3
QOjZcHI4VKidIkjTKtJrdD7A3lVvZ2MAej11sXPRg1A4ycJ4E1mIjToZZOLTT9VFNyD6eWk+FuGY
qlM7XbOQB56vC7+EWiMchlAp07aPxBuAgdakuiuTTDidbpmy0d5V/sMK8UPLIqqvUEqtGVCzfwbp
x0c1BsJxlywQTjCEeYbR2aybgkI7cPJUDZ5IwDmplG4/h3IheFtoa+DHGBKUBAhI4W9s6Wfi+mv6
JaUruS5aU/PTAKjeCpFBASNBALSHWwDiJvaEmfhzSDSUruMCub2+DVUl0W4eYhY1vS/ATs+ggzfF
aui/m/LUTFDqj8Rb6kmZJWBuqBxITFJLeKXOGravNtkM+blDjDLUNkRsRrF28AV/vgYQ7b4KiSlH
gemb/Y6Owf80uqcYtEzyrOWqJQLdxVsk3u+OJJWELiTrowdGRrgSBc8c1IyQoBpUTQ5fO+T6NjPK
T15iOAo7B1jq99OtXIrqjd2Fv5IJuaX3W71gh5sF3TzLEIKwBuzZ6utIUg14EvQhUnhrNn7oSHDz
7HtIpBdwd3vJNheetDRnYUtRpmhLjbtljivfkx/IQOuLHwp8V39xv/6JOQiC+qzBIkenTyoH5DeH
7BHW4iBBrsDGlppB3eXN6uvPX+/FLCaOhls7BjUahg6zBguj3bUtfL62lOPhHpQYnmpqnJURABzn
7cjyGTJ62dRf+IU+7HeNm3+CqkNJPMBIdoUSBIvW+VQO5Gt3Waf+GN0ElONz/pkzUD9pA6hNcCQM
o4Jj7PDA1m3nkbvVPmYAU1y03AaR/KH3aCQcrKq/PHgQboC/I5yeTilZG2+5hbBQvLsIEyYvj3f6
Vo0zsiryTH0DrVyhQG8GxayDO6a3TRiFJBIIbqluZv/MDigkSQPlNM9BIaO7hMAazwiQb4ULlhRE
NgMXScR4SBF01+IhmZSj9q9lXYIY/9IOTJyejeyhfS+WtSAz8OgPvaLcgqaLvbBqIdb4peC2+gWM
6AhvpbQyRMqfzXSWg4PXHSzuDn+u6ctxvypW2P+PsgZPEU6VfSbwre371MkAzYGehwV3ZnVLOhrY
bc1CrkcISKXbu23S/9QY7WR17t1tACCxqklGl0vG1uoW7FoaKJufnfq5DMV/D5QYQwtX9yPHKf/k
eXKj7JUSPcnpcF/dBI68MDQTPvxgCFLDjH3kcV6Puag3xo45/aUpw45q/gMDVq9pL6/vJhvuBdmS
xEHgrwRKzwnodaJN8bSRiynsc6puz0sfOz0/xYaUMBRcCqj5yZE92wpdFHC5IaGJS8HKU+Md2Th+
voeizbsspRvEntKQLbePWsBNPKm2+DKb9Pd1FyhagiXBAO1V94u0JO1yjjamAvND+k9AIFqnk9oG
QtSodxfNBDh5JCzBd62fVGqR1T4hosHluNdZqwCMS2YfMYEbAc7eIOeZ8HSegyRVuNnsKi6Er6Dr
Jnlxqxu4WYyaCQQbTuJDzRR8cum1/CiWuVdg63azOM/+HvCiI5HH6iRPhMxcVRrjh+xdq0GURqpW
K0vSjhnrEv4Rjq0sxnzHDdh6yECy8cZo4BDloC2y7HPBNUEbHuMbnSabDxzj7jGiuKYtrqqEnepb
S+OYX+/x6JcH0IJNZzbIAdemAzYSdV04zI+0cr0u+VZfA/FKKx9d/FUvsf8Srb5lF0UeaJvRcuZ7
So191+cnwZksauSpEVALousfGzpSvCMH0S7/CNt6C/r1ybaGu3ix8ILLHxPGxBV2c2Mkf1fqBI4y
RF74jbkRyxhQf6tFoh5nBoLxttU7CGsWWdydcvwA7wB229lZpsg95T2XXVukTDDzJllKEPIfWrCb
erFq6P2nIuRsM0sm0vceN1mzRtDffRISQ0DK5pu3lwjTp1Q86YIdJVm2ho1yzYI+efthNq/uN2sR
wOrJWBfWRZQsbyyLj/J+RSq4UmrOS7g4EShTiHQktwRar89T7QjlQQ1/hro1ekNiylshQRhBJQuE
Fdcw0QQGJvZD2wcwQz0Cc6aMGsRc5iKtsyWTNnKv5qmFIA07u4hu62n8Y8EIl3KtsZdTQL7S6w9g
xn9M/z5NiTTbEvKD8wZA03pK8NbKJuwCIfDEyW1BoObn7rJnTBVG2JYHU/KjixraeSRQ3h9L5wMA
+cf85BOm9jZvq3rT6LAjqJ8TOHXEUsMUV8ayVMOUsytdav/YJVfVrpLi4uU9rUZpJFs/5YbEv1ES
duL5F0pHO76tsDr2K5PFMm44lKwYhGdohyx35dolyBbAp/spru5P+XIhwnsBKJuvvuEZvLEtqm0A
9/3/VjVG6jbxxegxBp/bDBEHUaZNQxwGW45azDrTELFhX8pAQREOLENCzC5ffxCo9TT9OFjOmyXK
iNx8Vp55CnbS3PXfBKU3WVlQdIRFUOhR8JGJejzb1nrUjVFNHRfO9CSlqHbe6mfvoY21PQcWuGH8
WrUp8wh7S7CTL1j3vMBcBsnqjsQjCG59y71ox8oujDhxMkXplrnBn+r97BsFgmNljUAdDjhqLCKG
QCGimZu21HJ+uhd+KNhPf/U+PZlRwTLkPUnXyV0lMGegxVb5oBjpTFw41EkmY9UTr6+cHKHwTr5k
4+lIDtSJLYZTbagdl+ofBaLU9FSW7/kqjepV7YrHuhlnU5+E/8au8iR4CH1hrxHsmP4WXah1OHqq
k2HCWEo4ONlUVmfND22jK3f3JMKht3hxM4EWpKqkAUAk0q3FslxaHhiAs6vmxQqMYC2E/Dd0UPpB
yLqvh76zgF0CBE7i4IHBJYHJ6zjOiI4u7C7sgZ0/St5Tyh4ygtIvAOl1NmWv69MJo28rq9F5rOSm
fZLyZ5u5kjxlG/zrc0A1z6zewPrh7VjGVqL1w0Tn62D8bkptRSfHX6fWPny1jDGgdFAQ0Xa1xpSi
5voGOadMdd4PBEX+4VRypSSzrYhUrKRTzRrGRPqyFAEZ5T2xQSevky1r78z4D/4JNp0tCYgKxR4L
vlZFv76sfs8gD1jxf28o9uP5MEiac0s/aUr9DwcYpOpARnHKM70KoNYBrp7U3a2xmQ3hx0IWAITS
KVd6SgpF+QwsN0Bdxevs2k54FhIlJ2ccXUr/xlhb7h7fpV8CiBqoeKMsZlN00mSgHJfdLNSmXMsN
8rxO7vjGdvLFa52FiF7R+O2T8Vn0PVg/DhXAit/2oH+VjG44gcOZDmkS0n7s4tjVULsSC9Kom6XX
3xoJ1dKm3sQDnu0nAcT6fuT+9KaFZF/owF0WFN86U4A43BI/GW9/KzxIlwrsWe/Qm/my02lC3dVx
oAZj0JH5cznPiEUxM6Pa1zClzehASvtjHJaxnhkC7BKbGGpQNTQdLINDJdWsXbJcbt8ErLjpkq9Q
foBjKut787DKNMGh70cR1asaqtvRj8AVTIND0XQbJfFoQyVl54ZHrfF3WYnX3NfAj7ekZoStemKU
kmgDaAicXtldxEwtPg+dVcV5oUqg1VTnOvCkLXBG/j3gYdca9O72LocMNWzpG4XsN/8eOHS4FIPK
6sEj9zUryQ/CdLUjyRGf5pTuHsVfQZxktqjZKxWRpSZfwWy+QeuaCkKQjSHMdnEUhQDW6nopfa/M
urCAGbJmlzcGnVXH/7dz4XS895NiOHTGr0bh7aqGQ25ru9nWti9cbuYeiiMJ8T6BDoyORfcyH4rG
Nx/CwNkouGGNG9k0HM6/cV27+10EiRm1QISzsIk0xGYhjLp3tOEpBe1Yi0bRcisTre3U81gSHH6Y
5j/mZPv4ANE9rmEs+t6fMCpwJp+XI7ncdG7/ecXsx9Z+YqDMrFPCkzuyE1dAbYfGK+yLKO0ixFMO
n/qGsTxbbsOYrYmU0TeuC7AbTXKsXKHetgBkNuHbMEGfUsKFsYiR81dGA2+NKKGxbCdsBe2iYY7P
QxnktQkiGpYP/defdmuCeYAGg7ZEj4vFqtPfpbDqqhPCErT6vovGAEAUUIGkV7uSlScWIdHzf1/Q
2Vd8Kw2feLDbXiSfIs6F3j2+Qzw1uk+6VDsCZqk9G7aStt1Z30efIyFaUvDzkvtmTszp1Ug6qtSP
KLbfKpTHmC4WDHtZWN0DYXip+vR3NMpUCdcsBf0yPTqk5Kx/ynApSCYDgwlK8T0f12VjFL35Po03
tkPfHkLMNjNFVmil7GYq0bSnOwTBL1NDPGHQSFHRdUmBdrp+QX2tSbrzA8dnUeT+kyijabTHFoS9
pZ1P2lYm1dJtpfs65u1agHTgWpcIRj8FTcjLnK50QafjL58ZaLrQExQRsxQqgt4Yl3+WEAQ7aYxK
bcJF/beEjGXnVrpXIITwaV2ZvUrTvuhzSQ42aG5Sb3oJu+vk+uRbksb6HbObsQv5dRxsljC5/Gzc
9X7uJsWl/djfptBdvUTkoy8EYrblXpbmkJU8GAdykI7blCL62meNg5o5NW4ASPDlt6Yvl3IxJwC9
U9T4R6p7wpMCUiXcWnRu0KTw8dYgOc5eEgfWFVxTzNGy+FVEw10qWPu6z9WKW6BYK0LMp5TNDRb2
ZL9RE5zefCRPPUsPguuVjlQUSIsNa9upXRfD0aan8MewcQIJK6vtpYEhmC4zbGoaB3ushTZV5Nz/
VPzLf553g5n4i9ZFFFi9OrbCNmYBqmwTfir5wL6sXn/E9H4QHx82IraOHsG3j0FP07URbWHBhJwa
e/EkAKPl1f5MGfFmiTD8B2PoURDDmfexU3/VXSvsDtDrA1HHVohoDExoGRgmSgMXLSEDaT89/gLK
oysao7Nd478SfaTVDzjIaJUqKw1OJe1RHl/22rJU9x21+jvEt9TGiPAsG0fXeUMVY9b6FvYdfhDs
27M9gPjx5sWjzAZzSzdfVFql6T0YyzJZIoVHKOopi4x8UoxRGO00cFTEoq7GG+Qdz+IXCrRBkaNm
iqPwXev3u3+BHuJLLDouvwWc86lzsMSpnMCiTIUnax2Nwd06kf6ymFvm1uQoN81Zx8F9mUBRptCH
ISkN/ZxjxSovbS24j1eJcxTJ47JHBwQFmwZo7wohv39sH9gU9wTDiV13Q54KVh3iPSP+9rEac/aD
pOzGpgToijl/dJQGsSQuFCql9/HTnOW0wC6AZoCHeBV/IOH9dGrKdLME9EjbOUExQkcDAssQAwxB
d3Pm/c4t5tLcFf7mmFmcDfO7abGyVy4ye206ADP5Gp/hjpDkuDGepYmH8oOy5agJB8Yzfkc8ZK7F
drbtOCF6WfAh9PCcE366NUTsvdase+S7aRMXq89yDMKNhrdGfZCBopYiJe2zmp9HlxD1J8Cvcyez
Osv0Ibuvvh8FdJd6l3D22ikMLUTiedShjdZ4wMIKYPvk4TeWJ2Zrvc1e0/5cB4gcKOMGEBWlFTOm
Rxr0mVo0DU4EkwmGullHCnXFgt4SHZyRGX9PcB0qS6xUnoTdcGJM3FhxUsZ4cQOSUhUZkFBU+r5/
r3ZNofrGPjwK1DM+aeqjjZzDKujkbqCFpUuyfmnamL/EukabBhrx0rY1K+pgkw/C64nBlCnZWAY0
BNq5BtOSkb7i5kLCS2F67Mw4QX9F2knC/481h84jGDM8lhK8UMMTg1WNKTQbxLXjyxuv24VuGwSe
/SkTH68idSo3cKfES2SJLH9cdVnCU2/2kfRCfpNtkUwc4CgKd5oxSZq0V5zvjA94FVyM2nkIxTIv
FxxZdmIY1Xf3s2K/iM4z6flZaOpnNI2aFZRz41I9osRXfwfAND8bECLAWwS4ayNOyHyxX9Z72mfz
Y+D+q9B4is5ppZsRV9shOsD5o9ZUxzLocYFUu60oX8TTsxZZ0U5wNFKuAtU4nGM5eQGhLPLx5Uws
JgZliGFQLP8nPH/+Rad5AXoSTj+pHIJp1HyVdxAKthUyn/7AzSwZpP+f7S0HqLTkdcDazFX6U3vF
3V8l4z2MQdA9D6Kh6O367PT74X6Ta6HiIZOsh6t+s+KlNp4SDUdxZ3j23kby2JlUZnRfDFlz/44y
f4mJKaWTxZJDQQ+jZCDMWkVKJcATzpj/8ggZdJHGZFHAiHKAjRuXvJLFOm5Eje71zsfgv2O6Cw4f
1Tp18A0+j5mPGT1PgTPojQOByPnfXO3qqySkOSRGvMPMgyLUbM6pYmQ/gHesoSvmcxbHf9DrOx7B
tZ9voz5scD8tUmzzLiuhFo2E86NrOcktjb7x6rST/T6CxyeK10IJOeJVo921BY3tu9OphwZ94JTQ
wCA+oXbxYrRYiLUT0P4cm63E9pBcCYRNvH2xCRVmVGmnoCzGlWy6ygH2X8pM83l/q/Hm1XI9OL61
BS43cHhqiKf9Xcyt/ybFZJXTfTOgCHk+sPNJZs23Os/iQbphRvMYcmu/OEltNzovU0KGFYjPe9eo
XkRDSbH5xow1VUcy169aZQXLtcXGrUVv7cEAqNL94h9qr0nOFu+5kaFtYhMe9v5MaD+f02dMIQpG
xn0Nno7xxLT+6e1LrjsLHGZEHMwnq2sEOLvGi1J9xN2MeauG6EaVU/KViaFAmHLMUBotwrQUvFLu
9oYYuVYwsT5dw9hFdMs9QZu8Mn2F+U+hiAw/IKwJaP+FKrD1nXZ/3JmkS7EPcisDPz7ptrpg09fU
YCjz/MlKYG6LEO37yIgsMgwWzwe5TcIjcGWC4ZJCvcxxoFnoZ2q+3ZSuhtinbgHEm8/OO5o2syA0
9/8Us5cqchg8Ma5v0IV6tJp8xl2UzzIkZ7Load5OVWIZREuondQdJvQE29TtT3ZhzXbygt1rL3bG
ArOmdHSGyF6GMfWKFKQtB4us526E65P/sz1YKhNIkDtAwWOOqxu78twh27U9h+bBChVmVqKhK2g2
SVQigebmN1IZUu+mNn4SdKhcgJwEQijQnJI+FBCoGJjCxWG5Q40EkEdbqDVbSBKlvJK3FQnRw0lO
IVClv38M52nDfBF6/MRv5MGadXdTJfIjKkvAXitWBjPaRnU/Mq2WZ1eDE/4KzSK8VrjDn5jy9Bc8
SnBeETzpJdJZ1pta0v2Nr8KIn6A5hufRVwDEMajreMXmYe/OR6u2q4Q6vVol82OkDWd5yio2mK6Z
VJe3keL4blKUL0JIdSqyBaRuP1hpH+1gJAhwC7zOsj3fVBVRSTA7UFvAx/mqKOAX2cZKZ90Dq9Dy
T96lwyHgdqIBkXujSQaAEPTpWXYnwLoMzyQ04QiGe4HzLKGcD7ctA4a3tO+ReFEynw5wXP/oE+sv
jV/eG0fXij17+obUIaTvE3oUpqCkdoZxp3AhpdajhR1QnElDj9ZIe256UCJ2eTLwCLM3+uAuoaE2
HyJFBhb+TXJ2mq71VX4Y0zmW7Cb+3BVtLsANtCvg8YcJrfwGsKXb67ulTl2hAZMMxNB79U7TCCs9
itTpwL3poiWAy/Ddtl4MxRQ9X7Wc8ZR7WORCEurhfWPLnabiLhz++4z0qGqEqpF42UxMUZfPClSG
aJ9PX4gKyuBcgw4jwpuqf17uTv3DHw4v7HIhoC2GnOkjmGl0tbZ2rzkT91yqvGq3X+zpvC8dzK1k
r+70mxbrq1olb+mQFKWb2EKNvlIqg8BE5XAcUp9rmyXfgd1rbLGrDO4bSUmAnz8ITbtAchyGNnjT
syG/Sz7AbOSi2AnerE+W4TCyFvBPxjYSwOQyoQcrheQheZynedptqvvhnUpAaNHix9obobFE/2Hz
jxSI46aEsh6TaTy22ufqnRioKUKWCES1FkL6Z/krotTUXWenNFwUHI69TWG3iFPGUfjejSlU/Gs1
91cfeIaD8reAEK/ssoMlR+Z/YwheJArI/j/scpXvIMraEWXG2NogSa1xEvi7rNbxswwgkUeFcByy
5rSHs+wSyDHjshq/NLRftYOfZmFPMdicEQ6tquq7GV48JG12wIgdZobW3nzspSpclnEkoiE8IhFw
UH9/BZt3pjaUNAJCK6L361IcK9HtqpdzrdxXuGHwiuQ61sfaJe/ON7szetMLlH1LX1WEgjYkprht
uOaN+w+slj5vmfCmXNpM0CVZB0JAkRywg5BGv7JCYFUkxv/914HJnnADR09JUrQlbD5le7E98jEb
gnec6kzrN8l9BMdhbls7nmpcBNWwDBpdiE6T/4Xnw3tbzSCI54OP70UjSfcpCsI0HQ80an6rHjqt
MjDvp5Vyy2jUxtFCFDhV4pdLVO7QZWv38tBCzum0LqHG9ufCsnvDwvhE9zIsqmpCqmDQkPfQ29Q5
Wq6wyAXVSFStPQTSuILAPvcYGiHkb/AH74BEoxFsyrSi897gTEGGF5zRbfdOzUrPBjyvVKQusdir
3H2Gk8P6WaCDrYTZdMI8Cgkn7uBtkadVDBdvocWCTIb8P7NTtS1JlgAlWVTT2aIJCPpFbyVmUywV
RMzYDqC/f+oND9yRqx9Rn6/wfEj8osm+MqbDB6OzOqPg1D/aypl3JRKGp2GvwCHk2OoksP2U45Ay
VQ8lyhmo1fiYzWz9j37VxMIRJVlaF1k8qtbbSFb2WA7S0Nf+aopod1X39q4mXl+WgDvZAlvOG/G7
6RCJDZtJX/1Z9FjYlJCpL98syAFvPNZE3IXeX51NFtpn+Xctwxa6CQdfv9CJy9QOEUQZldpdDtbw
otxcIli9wIi1jI40Hz+BAIDo370XbECBK7aJ+je3ayZTAG/X64EIwg/k61OeYY8wH2WJk8/KzM19
ucfVqkKYmoY6rEGa0u4ETETR0iMMkpNERIRBOzqeF/Zf52YeEa1fE5mZwwjlln2uFq9RAOEmfl5w
OZ3lhcCXz4VThvpcnN3BR/TT/p6EN3L0BD67drin2Opn2BqTR56kL5W9dW2PqCX8gKrdijRH5hyQ
/BY1jmeN5s15DNvAGwchtlP6dTFxcFT0ERZm2GA3GPsN97WLufjF6cLo3yVMqIjjqqqTM7o50ss1
VP9sEIaRElEtpPj2y8Tas6PEcWvawWtCnUgdd4bvMd45g4SCW6OL+TbboKAYt6Z5Z/aig01v8EeQ
dpARMQ8f+KZtoObAlvye1IdFhIXN94wcxcHm24gcdUB/bZzLVMePlPbfxCfu0qNFyfgoPb3eiAXp
5tx4LTlhy+1g8D3iz0mRKzxHlQQg47X/Qm/YM4/EywJHm6RrYw2+UZngnQFcVsarZznpPXmk7s6/
FYkFhRFcACG5HrL7wkeKM0zi8+msGu24ThaIKzZZIfkRLLk7VmWcoKhCwwtUJ+kieR/L3VKdJnAN
4TOakv9NKtQlbEXaptEZChmbs50yhUmX3QyKz9RMPTw58cZX4iDjx34HF60dci+eRJsiU+ilI5Zs
JdTWSWz/NCWQU5Ua6LC8cgp6ovQhstVxIJDfoiu3sK1lir7WJRNiDBYgSsL+S1DC9C0qIGQK6ilq
lDYuSjRAzDRhfJl4zxvb0QB0Y8MNZ4/ZxRCnEkNRCCL/ptKAC9XjOx3iN5YlfR1aCDxHrAfNEumx
MC8JKCOqiUYYQgAsyYjstGarzJmsyrYHaXo28NP7wfKMzxmQlsRNQxFqt9InKL/hm7MAidPeuiCU
UFVSesXtN7VJ+OaLmURnvErwCk7tiiY552WBOUVAGMrg2kHcgC4zy6Uk+h8Y4nKSFz8iAOPa6/6m
2Stj0fyPkCFvVmvg2U/i8MVXbb2jQIu3JIiigezRPbsFn5uxulh0IsWPBizrlIWE00jDRHcmEcXG
WutTb/l8u/x6sMzyiis6QVelElkSsbk0/rjD94fbqFg+9a5EuSXZRHC0R3v71qKz/COU9jaNnyCa
A67RPkSXSxj3rLPdJPLwvpzpokSv6JZ3BfihVTFDuMYn29ftb2sNxPiE29xCeaZkJDsOfv1u+3eE
vLWUHQPMtab9u+8DV+hwzA5b6sxt+DOtkH9nrduvCzTe5TjdsC7xlfC8xSz/ql7QSI6QHpe8v2n+
5GuwI5PKSSZ9eGXW1oJP2U2FKyi7gXrkQUuo/sbxxm5xyrraGMYcvCgIixWK2sljJxc1O1OFQiaQ
ejaFUzguqJbsym/mxAXaFru7z2V7IJHPrYMpgtozLVULbtoDO5EuPFFC//QFje8Wwh/YGzMVdL32
K1l7iihJNQuK15KdGdrsl91lSgA3BC0uwi/MQ5ZulK7RrPZnDfcF7cBtZcdIJf8xlJe1fdhVyozd
0iDJNNiWXqrtfyAMqmnhBgryVlKypU1NzHg49uebOORXnYezXE2I4SuY6pD3vcVcKoAhdFMYodNZ
6NnF13KAEhZZ3rPC5JiUmD33jRu5yl+sAQNAmeES2dapU2A7u+R3z5xy3JD8yxAfwDPyyGzbtRfy
+1uDazQ0D3+IhY9eQA5wui2M/hEEyYU1Qf4gdW6IxejAQQ2MfSJWFPJRk9JQpKzPDNqp92ZpnQ1m
Mf3c3ewaEEHGi6ILY/jSpAKZgRzPPpAUfOqqW0hsNb5XGjMcqoOvre7eceDLDMAzG2BaCQJ406pe
MIneJaecR3ViYeLQ2nNUQ31L0NzkVOykNRCiVlMC8Yx4/55jSRbb2nIdm+T1RRTG9fRbFVOi/CmZ
3FDPsZ+daVg7fPaoq3Sn+vOc02A0aUuGzx+bIG+jfGKtUS96udqZdwpW+tleWMnV05eZbk7mHoNn
k/+Rcl3543WXAJq1bH2rMmjRrGWRw6M3Eg6eJ9OQ56rtamqaemcorsJ9DNh4hqm+lKNspYf76YLn
rhCMMN135yTypn5O0fhJycENlIxnleKSEH2viI1mTQ3QePUxTKqXtqxuAxTzgP1rI4uwlW31TWgl
ZDjch0B0CsGvqnn2RlwOnKiG6E8Yk5Bk+y0p0Fwbp9+oGpOaO91B2Q/CuPDZD37P0aDKqhw9M7rm
Dk7qxjZvycXblWRdcBsVVXYviLtJQx8mr7XVo1h7DvW2xhqI1FhR3i2b0rU+RiH1spvjzuAvHIiC
B6iLk55tHxNNZNzu9jvqW126i3mD8AO1lvOrn9c0eOMMxGjmVqR5BjnUISOoEGm8jFOw5HwHgdoD
PkLq1XM0ncHK2TaU0y2uXAl8lTKJzaJjUxoqT54Phpvx1ekHziZJ2QMxNHRJXHczfVaVHRaXNQwp
qy+MrQPe+YpUyGfw+nhh/+YbJccaHPERlEX2XKSzxLLcg+Ll0S5ahD3vqsGNLh3VfiNV7VMeVX0+
/EhxbLRTAGShuDWLHrLi0yRBp7qYm3iBqW6tpgNXUvNJvldK5iOZg5uIG3KiF75YDyjXWWdvWBPX
PBP4IZYnKcxezdrsEtysT4o9+VVKpk2G3jQruyn1KRYZyOz80UJx0GHADcu5+6fKaSnxWvd5sVj7
1c6YMqA4ZpaODIqR4C7uE5tGD1pUdyPI2f6jKfPnqjXxnDjdXmexZmyOPam4FDQ9kl7u1AxCUM0D
0BVFVPDZFwY6ioIsPt1m7afLsphpWjorrL6qddMXc8IynHW+ObKrYB1now8zbfsSVhCCJfLJ74rX
gxYaaQj/i4NfNe/00cicezFcVEymKDTQVR2g/FY5LD/MEOM5P51HRAlLNpd1vBY7kNQxsbI7ZqCt
49TwzaqXM6IFnR7yt85x26UUOIW3t4s6/otvaNUV4J1aWqKUwhgWBnc8p4452nNb5H1gMaSWN1fu
yNzBATq7xjc55vgO0psIPp10FaQbqyh+ubO2FbAaAdWidTixormP5rd90eVfA8ESfvdeKXsmy0/K
hNi/UkjckgAE/81GQ8eWmRjM15m6hnkTgBDmrppoGnXd7WRIe+rDx9LOJNNlOEy1yf8olhzaXENs
q41pfo+yVDDvaaSv4TwzJ2XnB9IOghqBI5TwRdckCzuyO6XR1h0TjeoAO+wgaLDSx8rvgZ56inmG
9wM54rN1ShfZh3itTQROokG3fvRF9ZDX32DX+s8400rRhw0T7k1fCfIrIzNUJtoBRrYau/X3a6A/
/NhEWacFTEAtV58gByTjmjmMY5rzjJWkODCyH0zVwqFOFC0XM4zxeDEAY0zDAna4RGSFGT5Us2PI
1rQ0rttGK9fre+QHMxFfleAX1v9AFA7sm263Ite6nIGwZI44In6QaH6r0EgNedeV1ihhLkxifzAB
kLwiTLo4/Th9a4ytbKNMCUrC8NldI0Y6+PukXbZTOWWZqfGsRpokRIRsZj8PDf2mcPX8GkN6b7sW
i2FBcvbI45smXTCUz+mT/PpOjrT81QW5610oXkkFGnp4p1d9foYWGVUFaMvAlyTijp0EfhkoO/v0
klw5OFICMzCuu66iG1fJsYVPvmBWbD1ch1Jjj7mB+00/Vn1r2VAgecEy5XCshIusCGMgT7VAcCie
bNKpQj3JemTFAA1RkAE6wRk+vOolN2P2wDjvqbX8JAZINt249wws5ovyl8rG3JFk2z8dhuTORfjJ
+jhHPfmvjAJaHQKzN7KU/BcCDVPikASnnCoD0BRUBY+IqawhEwGnhSPmQ85AsOtJHN4DxZm8D5pf
p3QfO0faBajlepNwzPU0UsjehLQ/thNWuc1dQqH+tkBYfbjIecdFYQFyvl5iBDWMZz3Z3fxheDyb
ySIrwxbVoN4EpkwkM9ZtdZCksUlOcvPY0V5QYtUq7TMlgbaLNbmp4+ifP10Hmch4auCjLrcxtpjW
tW5OrmqIebjNNQDVJdopURzK4WVwzvfDzO7n29MITPdfLm3uy6f+3h7rwzzoFk8kWn7WDTS9Qwtp
L1LgU02QrgQv8YeeKfHAarF4KU6xGyolY6rFu5Re8t+pNN+Vh44T1XGSMeoZF+Bwm1g9hsb2QS6y
zGomp83zPsTiq6JkLvZKKOBlZseI9t8DrbKCi+pgv6BZ2X3F1CPTxf0IfJUGAyLGUqI6a/40T91h
lFqJS47fmotG2ydQhcmIFg+kiz8qcTKXIc5LOSOef9pSjY9RAGtQ8vmVSPz6VDBkzBDQ4UwjrJYK
C5umG3qLRuKOzakq7YM42ycYP2NADzsmgptbg6NHCpXtML7kUDs+8N8hSqK/jyRl0guP2A23zFwF
kq+a3swCSW1z0jbFPuoYi/SvTWujlgpugxFBTKRIKYEIBWdpCV5mhMEnwRojft/Srydf0Yv1DVBM
1sgnNviSzcpPF4QUkrDtwYpdP9UL9Kv/wvt4MINQ7i6z+jhURY3iUm2YAq0v4Rvgr3a4f7jaLGxI
nNOr9Frd3tk9eeCnm3X7+b2QzFYlX4NM1w6MfmaKLBVVidfN6BrzNUTfCPik1+6tdl4DfuwzZzFK
xJg80xxV/VkivkRkaM8VJ8BxAUxO2tqKOvkAoMLK9aQp9gJqCBr1AFfAEnaXNN23ge9lMrqOWHep
XD+LkOYMWxpOATTqWVUhCRsH96H7seLuAc0LHEdh+/jOn/ltRRtBtLpUNWOaYjrNMLaSIOm/AvOR
U/m4X6tx5HM3XPXx86WXz8SM+Qq4NR897QsZXsyn3LURtl9ss2aC8iRpnoXOwDj6FlyChdUhWyYr
imdUwAdSSPclDond1iHnK/dKvCEHPsURxOnOhEuoiS3eewE7a0gbhp6zhmPkLcRKskllQ5e/eMz5
tL23HXGbTbrkZjZtoXJIDANqte0r8wmXjBkj6sDZ4oOcSoC8hDdU+d4kcIQRvO+fBBrq/en+AurY
uiLjkg/FGgAKdS8hXRHiUcxo62QvEOdm+lZRx8Sf1JeCZZOjOs0hu4dNMW2H0eKONNfsTYENy3lY
BCM4YH90oWU2BK41+6aNtxyZenEeZv2JHRfmYGwCiktdw88d6uL5hMSWDBRuyWUOMZQ/mgJSgC4H
biaWef4skZbsy/GHQcp7dClsgDYYL68aaANoatUK9HolvHHz3CicarDbPA+fHcYNh0gaauGVIliU
8Kp7vC8+V8JHsvSLvyLZow6xSxINuRBOelSG8Lj1D1WCX7dpV2ThrzGd/HqHSRYsQCzdWNBSkGuo
eqny3x5M0aQInND64aGEDH5nhbcLArfTeoWatpmL+tdgrGCW6Qdi196mW9mFqYPjXi4wM8vrOME1
Y5x9YXVhfPvSvnmuPRyaW2rvA7OuAQtIvQ5FIKRKbEuusTV8jAbLT3ib400O078DFUZdQ0kOwi2M
D3DuzE5M3XNIbSFOdX5/hbBPKB+3wmpT20lxw5wxa3HbS2cRs0ofM4cGo+HTJXMbYGJ1wItOdkHY
LOPCFgsSqZHlx8oXJNDjVmMSl21hhjp2srL8CYtP0XwgGtk7DWTYF8oqTW2+JlI3GyrxACAUsNFb
58ucOWlT+nj1pFNkyp/gyO+XtUqoRdHq9zz7+XPhreu8mpUZMgovqhcwhE0HU9TrwpAhIuG0tsf7
L4ipoY6pmobmm3v8tYQZ3QaO96t+c9eq8xxA7a9IMz4ZXZ7AcBksRcP83+uV3VRJfxZ7O6EoXrZu
PlnLIq2AnhVfv9jdIQg6F857EDVbuFxh6S0P3EtuGuawrkABbOnoEK5O7jNUMT5tt3Iw9y9U9ZMu
Q9LplP00mF+k9WwjUsLLZ/yl40UZrM+MD1bRjf0o9+aKcc812onaHWWmvjNipLRVLAsa77HHqIxA
ZfR+higoSRf+rMy50K4iUugpfGdkXMVtNOQh8xBOSKxNaB8kLfbyxA2IZblb4relXlOF9QYQcH5B
IM002hZqF+tyW2QQOPtBhcwZmf5bRRMQku3POGPl3bC1Y5SVYN12BcM7ddBldPVEyO5zwzmMuePJ
1VZiwgFfp0QyAn8AWBR9886WvYkovj7ADxaIjMmEREAiAaSysfJ5hCJoY6emmTLx86BEwayIrh6L
anPaIHQGmuh12fTtFU5U6nq0YrcgSTuZYcwRG0wxdTC+eyYfwMsOmnuZ8dleQIvNCF8gphtpSsoR
R1fiTvZdeI2WIQ+wgb14xQKh4jIF98AQzDBtmsEsoy6PTO7kcTLaV7X67OoeLI9z7ii+mX3yD6yY
GWzRWguxLb/amvUzW3UZ/dpaJgYmRRx+shM6CUEqYL3QSrwaen7uYBtp41YmY5JRfqnbDwbSfkPT
aAEf7yepAlsES3cgVc5aSSw1LK4HkLFp+yUfYuDjvLM68fvsKbnChIuXY8kZkN46E94AbnV25UzF
Y4xING3/9eY8OZPJF+pVzSOWeLnoGab6133c5g8CBxObMTesQUrHIzibRRrvv9bI6nJh7B5zad3p
qWhqNhwGS3DBL33C1PuAVcEENreY8OTmCoKh9POnPAxtwwn577dMZV6kmkcG4DAL7xve0hn4T1Iu
o5WwihrvBSyurdyVV+JbK89KZXXL9Nm/mGZ+cqnOFuSlTQx5Px9gBFyiQNR/YwVEyr5FuTn5ok1U
zExU8Z4NPpAp0I6IqGclUkxxWENUDNCtG1HOQoEVPvxzj6RnNB+U0dhJnVunkbVl/IJBAT6wN5LQ
en1/yCYW7e2+/5NYjfN9E7/JrWFJloRZzDMpTO9B0n1as29MidecTQY6LLMt3RWGtLh8DtR9Lk7c
Q1wfpvnsMzCXqXZZOpQ/O/hZ/DJR4WV3MEgAUoaNxPubn9uddnVLmTT5OHpzRzJwc0ZF52IenEhn
LcnHuhFCKYq53sKm8aKqOi+gsoVYse/ByTc395r8UldJXlUICeVrk7vUkkGBVd07SJbZMNHwYNPQ
ZXNSowTctwQVyL3ocRnufPK+oqOoa1iIVMv5B5GXXnStqED4M0QpAMIC6ZPHAi71yHqZ0Nbyx4Nf
scwDBADnzgqr21enSYIXFUGCCr6tL7DEIO1zEApJ/Aztyesrn9uNRp2jj1IchLDvVn9JmaT5gVKB
xx1CNNHJQonxybaigHjWnKe2xXbfOVeLwauJfY4HywuQXdwVgoKz2SYpHoJf7qpKUJveQwo6WuOB
mGaAmr9y0Nn+9A+ih1EeBCc37sP9vRdVTfwQ+DPzPEBI6KPr9FmXLbEbUwCcyb0mwovHF90rVIQE
fYRg94/3GUwQP+0y9vOWHi7jkIVtJk0Pzxa7OrJvkfxLLt9czZVLjCLBjPXSB3oHIlHmnGZupPcy
18SQu1A78C0W1SOvo8I+QNEiBYmnmMo4EZJC9QsARH5JMoQqNgQ4Gs4Ox4k2aJCLmOixQzyfichJ
q6D0y+wl4GG0DYhSjNbRn92qoOct56C/aYUj6zH8VGtf+gIxc8dy3iKOsOKeM9MMuphs94v5wj8z
IVlAKqixGjjLNJPrpyyapMkne2JqbUZ/761GXhe0XvserPIhkZszDPZzLWGi8X1k7K8hJuCDm8qI
HiBjFfD+wH1ZmQ6uL4/DyHTII/Qp7wliJNJ1JWH30+UV0XNqSLa7YMLp5cQ0dspLiLAWb/2o2gOu
JEBvFrxgKpH07K4LEqraqg4Yl1Rai4JssCw3gQGNEiOwS0IXuHfxyLUdP6xhOcOCO26RNqDu92FI
9OEK5QGnjuW13SUGeX/E50n1KMJLJ4IRChjHc+DnkLQWKVL0OQxMI8f9wStAtUAeoooinjO+a+pD
9+naYTGl1HUA28S3ubWOGUzhwQjJvSJE/mFkUBx/+otIwa+JaFun0DFT7+AkA5FnQBLZNyaXJMqS
WVyXOaD2d4jid0TuhdUAKETnzesR+9owh48b1uC/aHKfpMz8jlm1gAf+TeR776lGQS9vnIHO6zgp
s0tzAw2mwoYEVrjSKbMUs+mpDJcLdZ6nsTwQTf8L/5l0tU9ZJlh2QFu0uM2/d9pCmpiegORpkdfc
89rHWxI0bRx5V4updOOITyHfyOIzTRdQgDELRO57mL6EhwCCq5xMchNQ8o76SmItH9LsqU5t35+i
WllJnjYqg61JxCxMh+r+ATwigIjWA3PQ4p7d3CmuyjSiWpRrB5pIW9sE5ZEMHzM+/8rDaNb7LqnI
ITgC7zOwdL742dLbJl+Yp6MOP8h+PNS9+xcDC/K6wlhI8QiWHbrw2jW0XEJshLGREtt/GLMgTatM
IXihb0DdYVwbLsjIot56WNU1enmh/6ogFRUlAkAT9GcKB8pB/NysIcsTIvXdwQvNYNyLSpqL6TZy
r6v4E0O8GP5jUu8wAtGtciSuAe+ZBXRE+C+25HvpfTipgGfHZ+JQ4wrBHY4D9NadW7nzKjnuoWjv
rnDaKp/pd16SJgkl2W9bmn9AVk4CpPmMXq2rX29yHisPR+Uqya3uoHQd4vt+c+uIbxE1nIBu0FxO
jy84gQkxnuzjOdWKHdON6dSYrgldjN6U89oUOnIztDhR5FR+FjoEbIPKJpMKE97UI8N3VIlfKzED
5TB9XMoTo2ID7oFjVwQY84UfxAf7UrFAtJzu9pDy4E31KEdYZTyWsR01eWsMTDg9eTmgL3y6AbOa
QN0p+fxCYAsn582TDydUainE/DjkmaHeBM2kXYXIEndHVSpr215Dzdy+F9hcdcH1jO1xlHukQMN7
C8yq+VkrYBJbDSmLWrH+rVsOkz5ki4U7Oadl1zT5yBOZV+M3wDq/cXzh0oO18QL6FFRh+hvaod21
ui+mXckEIU9YrdWeov8cfVizG2s1iImYSQAY3EsxEtr5kvW82bQsN6dxb6ijOnx3ZZPC9XBhKSJ8
PECrc3V6F6u4N4gglYS8qn4dG+/7ePcjMURp1tSLhyJ71LXaxmwhLOjA3AYlgv9TrBD08zzS6LPP
wYtEvzx7ytFHhuXExBkBPyUYqJLVvTjVU0EPhfpIwELjkwIcdDx7FfQXCGOUzDErkypN67LDgkVC
HJUrrigqMLgqAHvdUTC/cbm3cZ0X2ITL1gslSAbC65AyEdZVZYjhVsBZ7o1+IsjyQ/Ahhlmn0IWr
nWFyMs8HvZzm1YWj2elk03LB76O9s96r7iMKE0ihXVM+7HCnHy9MXd0KbHQyr8JMBpWPi8FJbaSn
FgpT1tqFKXVE20SEDULK6nBObTky3dObd3myrPLCH2dTgyJ2L/L4q6ROhrWlP/jF/ku9ryiZ5Iy2
twsvhBiCsZjx05Ja9J6UPRY8kjScormUUrKhlmUyOBofSrGWijaMuuiGX19qp83PPKMaL4eydxkv
+OF6xP5fDjeC6HdRIRqcezEHyFM+mESRmRKkKFFv5DLBzrO9ArnWyFZyBZjIZtsSZ8/EILKXB5FJ
4A8LpTjAcccUl5VEjD/xfXgTEBf6k2uXIRldFabAUMwgo571OwYjM9OVfR7Ma+SXeynhsC9jI5fM
5gKRv+wcrqo1dwWGqHMRDapI7p8TCErxN5nQL6dvuS8KEsuKCpuOM4umUXpA5nMlNdTZ/2dwYtDQ
6/01EUDljwaVmhYP3HGtC83lfUzOCOd1Mr6b0JgvzvWmBoCdYI17+4QGbI+i5ImOPWj6tLW2Lkuf
lSpjWuzQWxGhPMyr/DOf8CdCbmeaIuGqZp8xvI0LDjTMBrfc6HbzMxIOBsG/BtZRi9nWwNVyEYrv
nr0JSAS3ZtSSS4FbeTdb4UyqRyQPVGtiPX8RdrtTiqkgl/adKYM5SII4IG4akz+bCbqOurf6sLFf
SvnUfSZTV4DlqUkffTgtIv224ehZSAqDxAPvRnLbKJ6ay5qavSK1JZPhGmTBPt0e8Ybl+Ja1Ddst
/1aUmZLjDIL7WZgQs1TOh9JPZjTsbZQx8zNffX1WZqWYmNFvtTZpcKGZoMX0CVyBILOuVIVpiy2X
DgtScmvPuL31S4XbdA//cuz1C6GuITXKJ7Yn9ufZpk4+KQ+VoJZES0EZ0riw/Ibz1SeTijpA0tFO
rmatWLVKAo6u4DtEaFUhBmbkuj74GetEtxrxX/ZFCS1vhu6XEXBlcdVG1IPahFJv1ixrOR0BfNjH
Mn8mNUA3HRk0Jp/aV5AtoPb7NxLLUyut8pvzv/Iyxx6Hagnfg7q6fYP6b22uHWC2fMBb0w1OJ7k2
myMo2dX7kbe04ZTotxYLNjczx62eHllDmpc/xv/KTDpvRxPmdIZzIXeHPSlewbniuDRJjWuXgeLY
up+A+OVKYBeck0RyCw5kXCDpRQKxUQe01Lt0zSxMNt81XKdNR7R3PIv9ZeVL4fVIbIR439KEJD27
Orm+nFFNqMWsbNhcwGI7/w7hn0rN+20T++/6miTTfAtoWXOWstDnrgzo+2Mg5R12v360pL3nvGfB
mBjcmRhfR5b1VodWHfeEjERdLdHvOkbe6QehW+b5cY5GNDxHHwUkGU42NVjpNcyUmZsNmKYstoR4
2GP+aThUJN36GocTDkhukFzW5aqkiF5jb0zYe3oLTGmsCdpk8GIO99Det2/TxUTOoIUzy1dU16aY
A7M+vS1GohJnJny7nrzrQT3X8hQW246HoXPefgpDyjfDSm+VTJ+MWHUZaR2NiE3V1a1RxmhRWhei
zH0WSN6oECveaT//Q7Gqssju53hzypE7gzVkJrXBRbbomeL++2bw/oPrdpzIdKhUGuPnAcoRqr5R
wdwpPvdQo/LrbjGUvMhj/5nQto7Z6fiMQyb2qqjqFuH/cV0XzJ5Sn+bS8mFp41fWBnzP+pi6xWqA
CAbTdzVtGPe4km5PsURn8Uz6FMvXdTTLdvpGDsRVFszsur+41ir7vv8fzi9xoTiLxN0oycArdK7u
6X8RNg3bBruajApeTCIeLD81bOU6UkxJxyVU9GELBMauOk7Gdp1QdbEmZoqus6pe0dlIMT7VCRo7
juvT/bT3bU5zolMwnpJ8CXwX2FfbJwOa+wkyDGJRlHPkQ5S9nFz4/w5wXQPKllD85UiRUyYunNU4
WNWdTKpIjDPElkFZs0ujGx9zgx6I2vk9W4Rt5Poggtzf9dZjSNKugJl+RXb9lAutmTHO4X82vcMV
JBO7u6J9Re7kpRRWhGY81PBwZEEvgJiHl+pnFeOjjprHlMKWPZ2b/G8LSJWIzFCnLO1BbFZeE0Jn
+qdhuDc3Q6g54LsPIySeV83Q0i6je/sSUUtFJn2iW0lkBrCP9kNI9UZ9LM82j0lSzyP/Ui/f9Qo1
GO9FjyAYIXE2wV4/n8MXEu6ZoOvyGR2f7OvNIs3HO+JHHaB0OKXyYTLlDqe26ogAA00kdbR8th+b
/GguvSotECcskYCuAepAtrWeNW47bnIamxvRAafkOnKbF2ht2+2+WWLba1MtMUzQ1DDiq0bkRX4N
xkkp5hb4ftoCPBxRSs/Nl9LuzL2CPlitREOVNgEZLacjI2SwoNY15SAmneRwy2aXeFD3niLLdSCj
Eoz9Q+Z0/3x4fVsDebCUqUnkFPTKR/s9y7nFyvGY6rcFRPjFkaHvLGQjl9L/m2XBjXk2LVAO/qYb
HIOFk4XV5NtruqKbmR9NbvbKFWIFMKfaYm95BnSmam4RbKJeOrvd4LRYU4SY7YlLGGrKHNFtPhrX
xHih84SEEwWLstxMWokLHW5aV7xoOApX36eWwG9Js9lnnFAcNEiIHhf7BGdTePv9TPb5J91XQVBi
+aaosm+ZGV/9D8PVDW3KYNb+A7gQtMvPHvHbJ/bIEEDTdJIaNC2Wg9l2RSr6DqhoDoU0aRZyPagk
voS+AjxPsv1az09BgjdG7Y0oTofyO36MeirQUe/SCC0lvEcY3glIloB770Zg9xlnutvUxm8/5HO6
B0oJ0qMsluIB1aJNt9lsuG4pj4CUr+7RAGLZBY5nwyr8/0FOQVQsMNdjd6JQ51/Rm0m3dl2pABlo
4s6uRW7MYQegwKclgNanNwzydT6hJ4cDG62B+EQ2r7L+J1MODIliDWt8EATRW7vM1Eil6jOBjy+g
GJseKP/sDISL/4LKM9Whnx5703a0XAv6J9u744CW80ioGSXUm0DgVqkDwliw8QpFxghoE4/I+SD2
yMKdUO99t7YWKdZAXx2vqWGLU48yKcnEsYNXvFdIS+T23Fo7GJ36v185I3vOF++zVVwT7kDh2Mqi
Kn2844jQkgARBGXalSrc6DwiLPA5TtutiraagC640/8rzLq/TLNabVAhHbk2+ItV38cVdV+ahJxc
868mH9JP0z94v/JhtyTCpbSh4Z0rTnK2vN0VGI/z9xa4ReOsYtrE2yOu1RrI6KKSB9vldjDl67TJ
t6Z/ClT62Wmo+eysY9lehzoA8Rvr1Z7D/4rnPVvhbQZyPssnYpvgmxLE/zT5/oJyYBugrZLz20Qr
2rf39XgkiG9J0znXArYCCR3Buuo2APSPnKzDR/M0QrTrcxqG2n8k0OcZ8sSbK4Nq9xnk+ZlSwDKV
D7ZfcsTOvZhzSmlXGFJJxZMSM3+w/D7kozy90PxgQ6ai3BI8busLRgUij1dcXd6SC864WUDjhINS
ozLRgMN5iGFe+wivREleuCjFi3imynD/ElS6N445xquvBnJ66rr516HOp2HnoM8CLljaPIL+/QRo
jcy6gidy1pQgskbmS4YqdoRBr+IUKDSTcV/889Ugg1+P864UtEuU5pampglgqBlKG+Z4YRW2YZED
QQWWyJl8nIFUmuZ07+pR3OUYKRFxezUNfQkbrsxTxF2jEazSmdVB2m1q7Ol4IgJTpdHKF4feqnix
F53AC3eeGmC0RL4k2olYSPWiWCvAkjaksesq1ohzlMej8Bnm3MgQ7yrlxfLQ9qQ3vgq3sKuTx68/
8Bn391N0WDtnzEtwte5fTLBDK0Hshz68NEIoL9Sv/6Sk5qdUgwaQvIq1W7cRCeEbS8FeSJoOZbUJ
FAZhQa3hi1xWVlXDzhP2In1lZK7qOEOEVJGtbTE4ScZCC3Ljeuzg2DdScpmZL8vnTPvww2rwlIh3
qj+dN1iO59jyF9wcOgFxXJ7cVLQuETWy7IfGPQ8GNIDFuF5Pdm2s2RgXlM+VPHskw+NJPtnwJnM/
2j6B4fWilFtAt4pj58x1tButdGpqcToMBhYm68Bfgb2CB5V5W/DTtWAQ8AfduFA+vWCKdq/ClXZz
2UAyMQojSZHzcBUjoKXOLdwj2RwpHhfFkwhYsuTvX89JdABAPHrTb0sLKE5nA0NHHbdGONRdT/ol
hTMAxd9D7AK8l+T8Ahgomd1pEdYvcX0besQeD7DXdbOLfBlnCneSMuC6PgGo7+a9b+ZrH44s4W42
FUF537YVYY/yEZOEjb47ai6pCOEsK2FAZPnmhtoajxHPJp0W8Nwa8DTwGthOOjmhTfCHyVGjxU5U
Iqk1DJDTJJBRmSi9jo/CWtZi9f3RiqItf6QiNoBgW/y/+IIUycBXyaVLGV0JPy+EYoBWTrNkauoo
gQW1W/lQBb6Dw1vTpIE8KFf1nzFJDrt6idQ/84wqb+ukvlItCGYCdoPqvYTAHEqWtSjv4gpbym67
2+1vdgfN0Ir2WdTeGlK8RxDf7g78p/d7zA+XK0vI63XYlhGgfRP1b/Swv8m+7sm2pYbyU4PbT4hI
6bmvfQVzFZbpKFLaZ9aWvSbKBo211E/DLtVqf+dZW+3G7gtvLR6tZMatysAI2/ACJqbeDwyI1RwC
BMPbkXkh1TJAnppFoegrwjBfRPpl58ydtDiacga2slB1u8RXaAof8J8PO4bzCEY87+8iJaV29jwO
GwKt2gTc6M4ikkDq1cn/n+id4hhpaIvlpCdfRT+USSrtAwuVIGlSIJzMTPDlKoehMgw14VEMau9N
/OCYpkv9x6GYdpwfrVgslPPw/rKkP4fUm7nxyqA2oHGvnQcxF8F9607g1+uRt9fDF4KU9OzqMeBZ
4B1NY8z991b2Q/7bbqO3loqzSndO2byFXsthia461AmXFhU4H640FVDsFY8gRzzUXi08R6uOuq6g
IL/7G3pmHri/eRPjKE4YI2yNV9augbRU9oAL1VQ4+ysTqizhiu4EydRNN8OE+lulgTMlwx1g2E9a
eM80WPX59y81GJpxDKh5wobQkIjuQ1i3yQQIBZO/Q45zId5rjQzrbGr0prI9DesDDjSV4RHBhBll
fT38aYEzEgyf0EOs+SY+4Me4Qi8HZBDlesE3CENPkWg4HQA3YcS2Epx48yQAMt8NeXUDBio+o9K5
2ktPSOzKN4erBKbKaHf15E3Qz6KcSY70jX/EwiMjDfqFQ3c3fcf7ynlaCQzN6yDuv8KrNo8cNHZx
YC1GaKojadL2lUHgSdCudgt0GIlIV5PZ7K2bbFh6RR5Y1WVKqQPD1MLtZhoGo2sGBRvLWD99mQa3
nwAbm9R8cRBJh+Q6XbhWxOZcOIpyqmiwDFlDm+r5HTBI1WFr70EHMkZ+8jf6qyoCWrGIZfH6udSP
ZqbZiBVsHQgPiygw+9ywsD7HHIQfp2YFOGT8TRywltfqmeMLye1FOnrL7GSGa7QjEvnTJ7TtBzij
6h4qWQKBehjeLqGNxTndqJdJSyfvs/usSZt6mtyGdEcljrKklGT6hARzY15LgH+N2ASQ6yUR0TTi
ODgPWE89MpVDowGUFhspk2kpMWfL6YP9Ubsm7kSLRuZGj4xr2T6FKiyy/71TutB/TtqfQPVCLq+A
pOF15aOYdroATDwAyypmggA+x97866RBUc+8viJca+pI3NPdZmgIX7sbUk9RcO0jWZqDTG8Nzchs
TVthxx/17PkR9E37zLIKYJg5oUZydpTvM8zddvYEfnLW+f/MhRXqdpcLKRMS6727U+6KCcapKAEZ
NIwlJcBDRxepSByq5LUT5LZw21QggSES5Szxye4A30i1ARNbOiK8DJITWK9ZUrFsjIXzHDx9xACS
uRVfmMGrcGXWowmyIkLPQCwtS/qo+14eFvOC43KKFzP9x+SnAMyRPTH5+VVJ0ilvF0G2Hr0EOirQ
PmAJJbL97VI7JW2r3+4RB8PbguDc4c+xPdNYBvaEDeolzHWluFps4NehBNz/PBl5uUm+ehydukxO
4+1IpTRywQTyBW5oBRpSH4w9BQfiISgD7aM0Vl3PdAgtkzSNjZ/525SPnyHdolVgAn6ebom2b7uf
rJhs7zYsGUnwK2apMWl87firdIyjHOC1tw7QxQYKUpz1MlCj3wJvY7mU8ABsWHgYtHMX/OPEBUaJ
Zsv1nseJWOclIfZtg64KCvqSwsXeWOzsCvc9BrFJrEZerEJob6BNMl25oMbMV3HYG/jpAFqBmLDu
AOitaeMf5cxWPK000AFovr99CoyWep4ARw8+fE+h6pO4CqWEsw8243Ach+IHgEBfGdn3TCltI1vl
fPBvYFcgZsMnW6Qmr5Rg6rrnP2fKBHm3BaAIlWXoHDb7p42ZoPfnXxWCB6ntTBXO9TtVJ7jFeTbq
7s6mwTcTQxpC4NP/WL2sWzVPwm4VyvRfrDPk40L/cTJedkYCraEp4Qs73EuENPzLTxdR/q1/sa7Z
dKfDPkbDiyOQOZErkgxQn1Ko7xsZBY9RE/2E3iAXsIKqNhqVbnr0tbLxHeLN0PrzO1orx+GO4nyc
oFDO1bQIBGO3VgST3PQrW2M5SDOcmC90U8sVY8cy4PDisVgZh+3BqIMr4378NT3qC+AA6lmE3PLj
jQOZTeosz+morlDEMzWsXyxkfAInyTC7oLFXkVEkPWJEW11NEuVuOkddw1p6N6mZHViYxmjmEg48
rgRJJSqSoese0917Fle9YaXkVMn+OujL4OlAP+J/luoMhuqVwCLpH04Yu7pKg5VnbjIiuCyipZIf
Kb0GPoSnf3wwnem7+cdCWF3FRDvif8/mHkF4vUNYCBXgjAIcU5IvLoDHv7/wG43X6zw+jVElIST2
g0M3V75byo8LT9DbXdLOytNeZFQMo8I05XO1JomDzivvRfbYjH3bDwBrwfyMOxwCSRvXRBXisykW
1REMuztYpkgAaGjYxvmEryTZogH86l74y97e9pHh0diP7fBkkrmhS/JCicEiR3Bgz1KzrpFDEDkY
CoVCKO46F0BMungcM8ksBKa8HEK/fIKMBpL9Rp6ekTuOQuP6t8XxhizM7YhJjYXg099cgITyxeWv
1U/8djgHK8tBGZDBGXxnMFwjpSSN3oGZ/lctjuTNKTKn6GjyNw6Yy9lGXHf2EpL6MYhJwRWDIQMx
qfjNUDi6dguxrzch/6g7+85qXZ0QtLbAZH7PNJIlGuTCLfHIFl18Frjy8zenUl2T17tf/Y9Sgem1
yJq4CPuY0CgBnd7D+aPVc0CJIB/Co32B0VNTE+ecA8ZxuaETyKJIw0c7jrAI8I679KlDjQnCvkcM
SqUj8L5Y+Wol2o+ICqPrA8zxc8Di1D5+0wl63tXkDoHkArtmGdkgERXpkKfZxX2x3KcprJIIlNP+
OGS1qIcwtU6pO4AmDZ0UKeaNBgWybB0UJGbI168uO62Yh5CsRc/H68wftHca4QrbNuZ7jBhWmGVp
sMzEUw86tMP7ewWionXhz6QSlSyKZy3oZKVV1PHaNgvT7/ymijZXuWdJZClMpDIk98odPjZkJwat
BTDQrWSUUb4TKjGq2G5ehUK2pvXftsAISQ/wJOlwXKaOoSo9+7se27ssqQPcLp3qx2RvlKZpokMr
5a+Wdnzjxy+359cLJeNvvxiJmftMQWCzGd/Wde6SU+D94yOow3loEfUrDCrZXw5AoYVMv5A34HT5
tjw21to2DvSvloa5AjvrbEpjWrp0e983fkl+qGepoHYySjv7azZh95HbNDxJZkIIdKn1IjdZMyJU
afORiXazupNQLpekkNbaIZtJVKgL1jZdWxET0FDNMjXOQDyzeFrS4049zpVYVYmYzwg5vm+egmMr
pqu2d7riRJO0Yixe+q5TmQjAkxdQ8YnqYnOTq64Um8rkcryHEDon7JvMstDDy3mcDmo2et0GGLQm
OBzkcn3XqoYLLZF1s/jq/RgJEorYKZ6Amu25Fw+cuaVV4vU+HgjoqO7emQU6ktmXBsrWQ71tMM/i
YB/Cd1fK3A9nP5dh2LTQPzwx1E3SjzENGgIovfWrb4Yzl8gTp37FUSDxknVe8O8zbaCEldkqwZ21
sfPVPI8Aj3yscvs1kSCmrVJKa0TLCeDezvth2hDBEhLETbbCiZVJ1bIy72nfvBGfMim+jOAJoKRh
+5Yv3EL/9B5+TrHpfSznEWcY3CZBJm7imT58Hk03Q1BRzzV4fkEbr9dospqrrJowfGaS8W2xmcT2
OUPNgG/dilCcqclYnvBx0ar0Xeq5DFFMViMzw/dy5DuD8xQmZ2J1RNTKrrGj9wlb+Bf5bWpSgM6s
+pPl0XKfgwB5/be0xTBHnJvaImlXHRJvAg3DMEG8T6XZLiUxGM5rSHriByPcL1tqOIRQrBM+rIfg
4DGnTkUap3JDrjsRANHpVHioaTiDfIT9QllKFmmYokI/17CXqLtrsH9CR/s6e7bEApBa2r/1YAY9
U0JmAiqw9wOrQOFCeZzJa53mEf2wCIe1fy/hPPi+jpFrdS/4TrY+l6oALfvmqkYa9otEUibIt+q4
FIgyqxCEbffQmGGd1HbdjnGr3Ylcpy2D+DsEaiP6/2SwkL9A+dDMY5F4InJZRUmnrM0GmTlQt3ns
TKb0yQx65khY76Fqurqzo81DsockdYS2ZBQOjlKHlcN9nAjy3wzjoaB8L/YFyhdQRsOnWNB1IL4r
0T3HOIJIlnIzBOXDM09FXPRwParVp+1GIxOU8aohtcf9acb3CywNPGvZ/M/E7hoX/ejZEijYHW+9
UF6QoIoglNM0H2897yHyak9g+F6ETMKGxYVVp+qYC9sT0yk4y+0ZRBbvbMp2PO+/fu+Mrm7bDs71
4Whz7tRZC3t7iHNc3vAWFd3WZK9oRM7IYiriayIw2mcKQ1mwbbG0Cj6nH97hxOvER/m6+MoNn6d+
BR0VX+uFAQuG5uFkU8bbqNYaS1wrwsRmFuDPiTqlvXkXyua1sqemMAuzpyLNOAPcva7k3ON+bj1+
lN4TpNzPQaU6FEXh3e52DrLkJ4odMO5tosDocUp5ZEK1JMZvLCGiWAHraQq17RWW3WxkO1BSXJO4
BZ/cDtW0MxW/h3XDj+XyEQhxIvE5I6ETVXEzvYqLVpewDCBj6HGqHuoG56RzLG7xCbxKTJtUqCMU
tpqObMoYyL7psUrdXP9/ozwLAM5FoHcYcryW3x5glkPsltDqUm3f3nE9nFRwKleN5nHOl4lvF4Uf
srJGqIJd//TdUtXcjqiOTjXzxInnukWX8ZMsuf++lrv25in/jeTTyfuwdWgP+jChK6lpgp02mVkY
cJdrtVkGjiFe/zmu+69nIBXduTq89SEGGRGaZ4PzAKI3QpqOvsAg4RQvcE8RJJsxXIlWu0nGkdk+
beUC+4L9luDREO+iem2YnRGhlZmGruz+R+ynbLrO8SqT6TSR8iT8ORUGGDnOIenjcyrK4UHlawyy
nhoXBGDETUxPNi0BMHOzKxNXL9cKj/nBVS53WXR5j0UBp0qQysNsLaSNqpTiVbO/wKVBNYpHv323
EQtG3j64rk/ukOeFOerRVWowvhmgveKcLwBBjOlTJYijRlPoI91wI5dQybGbmFK1PmW6bnJ/T8Er
nb3a2e9eAc36fiyZoKYTahaVV3dkVvHlunBvWGWsIbjsZyE83yEda9XKG8xpbYJ6coEOoho6Bxi3
850qP2t8RmZdjitd6cL2qVnp3Mplr/OR8Hu4Ko/Zo6aGO/pOgZ2TbiBFKBfwgFAOsa+l9nDH9cIS
HibNEfE/9LffuZcXyWTbYbjSqGEiDrB+nMZwcnDu5T4iCIfY8biJpBYJIKJhBMjJqcw9BTSCYRB9
CI8yzMMwT1QXCEPbz1WMHeAtLx3T1+Vd++NpWOnBxgM/uGfQJnLelVRgQAsnqG3xJCKImY2CgpRJ
ME6GcN7W4mKrVk0IRjIKSUjUCIHn2LvjbXX2z0ML6eCokudPPVS08FR05WvYqP3SYQHAtK5/loJU
dgpbZjnEFw58okgz8Sp+GXpWggm0u/RW4t6VgRTig0bUdhEBRbwkSAau58f5QMW1+7h7MypaiYk9
2KNjtwGJZVgtz2FV1QqnCx7O4k22qBF6yzn6HGWHblWlbQ0wSp6Rfzcy69gA9PgnxOoMLR5xqd+8
L8OCf+WkH2Z/sNN9m8NRUzVynZCzasvcjR2h6N2LH06jMbZvIkRraJrtqfQUFsqHRdwfCCpUr+ia
8f9y/IkwbMkRJu20/SbdGi0KJmyCMsHoBvXvhKpqmSWMJxM8h8xv6VVv8h3sCCIZ9v2BU/JYQids
o6OmJOf54Tz6R1fxCT1PxVkU0dfPO4c22Lhv9F82aZ2l8VJsSnXX86p6Jj8VrV/SU68c1Vh5CTpx
LUEL1vu0QN/ewt0vPLKqTNlA7qSDDOtqkSd2fCI1tDi+BjJbSKNAD8HhmIjARcs1FUwTAu2GmoV7
bp+8fak6Y1zK+9TDn5MH9Zvtr3G+nxuks9pz4ChC/TByUC6e82ayd6OPZVtcalT/QDY5rv+6PZra
SvvbKZyCo1DJpkHZqKb6soPhFDJt51JQpV7kOWHJnkYd0AX2+IMM83lN+IvtqZ9uMN7AU6Z6mahZ
jgQobfdhaFWqZBuY6uJnfcGExdKINSE1PcoKFT7E/0DbChH+/XOGT+BF54PXd6+ySKGbXIkIktwH
a405gjK0b5Ik4shTc+Xf1yf5EeKDw9EEB/otbOXoWIedpIFHMTfGwuuCA/5GVDxmLkOVvKV3AgJ5
2qnP823BrOpyH1u3rLsA4LY2RbF+KGzgy9c2KcBRFH5f0hOXKOw2Jc5J7pGf4XOC7LU97bokGo3P
JvSsE/BJnpy+ik4soURp0xy7BQIWSnslKelfOTF9xh5Qy1QwtjoByRJ8I35iUjtxbeXO5Qrkb36/
JtJmnyUD5E53hkBhEdQaywZfbSRFF5iozXPJzrzlDP90UaopyUtgcZIpsFG/Bo3nqxpPLFEawoVx
BDpwr800cvkcPYsovgDPQ2j3xJbhpNjFMzyPllIGFqtt9GBLyS7J0HYPUwfdz3VHUke+EzcbxUxQ
oMdvlLg6S0sfCIg4PdJtdkXuPCNXcT+f1LY8ZnCm/YMv0yJ1GFao7i2WmE1duDT+3r9WdvNuwcGd
JptjrNgxLAE0B4Ibroa+q1cQdf2/KDd9ujObOnNtUUg7Nbak5cNdjhRjMxeSAexzvYku4BjR2cGT
g6j08XuWIKC0vch1PPXT00z5nZ8QZqh7RQ46T99nWdb9V6EpYa8ivF1xB/3j9AcCghfzlhAoWh0x
wt0LYdH1LzUnvoENiAglkcSw+D07EGkvCR0U0YRo5uQEDp568ChAJwBFJxzGib4hmnMAXYILMwQa
sKvqfnct1Sv6twbharjEZDokU9ntfEV6eUyEbZslDs//ObniasoOCrjT1naoaDhTUMSyJxGMCnAw
kT1jPk4ZQJq+XpvedKrpBcrD35/XHq9FeprgfclT5ioBe6Eer8SHlPMluNxxvz2JPyXQh0fN2E5S
FgLNyB9kHQ2G2rjcGnpkyypLol6o3xekzO8kF8IyYvUfVpOnCO3sVFoG86vo4uYhODzbaMdSNwMH
EWOTQ1u0RUhU4/huKdDEEzT+e49Z8/VV2PsQQuQGVybY4jngqx9MNTiaZfk1gjxKquzIGEY1pJ1T
AUkrjKrvli/CerSzv/sA6487SkSBBTZkumUYn3AZ+Odwvkp6UB2h4luXbb/OwXgB/2PivpPZaKgF
4xTrlUWQLcwnKzcdiwNxYvR4Ql5LNTzmsd4ZO9MGynhUsvvnkcOImcai4dRWBt4Cf0tTfPcyii1b
wEUb1xnbTsu0gxjZUsV4HPkkAFVWgv3tU1KSfxC9lMiyQC0BBOmVY73GcS9vRTd1tGm6NBt5x/h+
BrNoLH1KGyCjL/b2J3Gow9qlTbFe6Ikeqw9w9UxRlXHatEb1abdxE1iYjHQXDC9Gwd2TdJmzW2w1
CzXyUKhTBjS2MU0b+aExusrZZDUYheNHaenBi5x6HvbV6ve14aMgByU2OyRLHpLgSKgi9n+RIKIt
KpIc2/+0+60VNw1ex7QB3o0voXRTYRLtlO6N/YulA3CST/qXKNNpFYqXQCDzraxQ7eDaUPGGxjAh
LwPu5PIfvtCSls1L1FadHdn52/rQHQQAifkLYRhq71ySca8dilvwqIz/D9tk8INYNWJAcBRHRvlu
rV24DYUhv9ll70a3Dm8buYGOlB51b1DnsASnhnhNQ8FlHOxDmOO9mH5JzD2YQxDCVw6JYjMeMB9X
hUr6YjS6/GsbizSaYbU/SMXi0KwRb4GRV7ADGvigDc2xwMZC4QuBVwm1W1TIYlPhzINv9nrxKKld
BZRQpuBVXidIMBYU8DuJSpGdyXm0+Kq1LH999yC3c+ALKWOIG4K9F7AO/ZZQHjLC+743+PKnLNyR
9QB/he4M7L6xtJzwc8GTzU/ipUFgChdAq602JvqBmKuEFu1ZCfl2h0zafmxndOAG0EG1zFyPZW+H
8/DPD+/tg52BpHEEYFcSH15eDFiIuK7IyAK6sTgN5YlMynREJWNWcE4i969NoQ92erTSmD3Mg4z7
pIQCFudjm69BP1b/X1gMyglsIA5m0gFnG4/G6Tnmxq/+kE0GdJsRxPNUOkbcGbO0DoPzDCOR1Nyp
jbJUhl1nSe5oy5FCVaRsxvW7SWOczQmvdNdMspmBgRpaXUYkDOIVlxYX+lJ/7RAhr2rrVV2lQ3kd
lQQXk9gJFrAV0vEIC/bJb9SzDeviCvxt3ROzMNKotFRISNN35Yam3rRbZvwhiYKN7Wgw63dpZ8v4
SxbeFwkUXFdhW8tSZ4c/P2krX0hO5j3MNuotDhCZLDk9GYt/Yo8iK/U+NBJqD6wOIm2X+7Z4NIFP
pXzpQedNNk1ERbnfAXPF1Y/2Oop/PlpLPLfnNXboumI7O38JnAs18E/+ts9s5hKFiiXW9Ofec8AO
coPsZ3grhwA4O/99k5sLougboFMV7k6A1lovRywEl8DWPpXnVE50bkzG2oGM9vzFdWHiHq8z7wPk
bqWs9SfGlqlcXiyniVIxgGVbVNU082hYiqOYibXi+jH/jdwx/RrZ4tZoIJrWtvlnMS6BQj+AMRKj
JSGz6kDYd2EgsOwm0wPnvjjrC9yLBoCbF7cynqIleVL/a6DDfScF6rtD1fPpMfFGCIw3AaS0GQPH
xzdKQA/y7xf7x9p6OILOkH7PNKFKOWnUiFU0JYMf73XK4g1+rFLXRA1630hPn285rQLLzcCTdyrG
3QOTQ6DOm5n16vzwGamYXQXpwxBu2be8kyuLJKwK2KQicP6EcX0Ty+520GM0MWbdG/PWWOR5vaHf
wYZOnwuU1KzijN8eVUN00Q573zmvvGZ1A736NkU7WC0ujfvUjFyQ+pUC2KJQdzcCkjpfM8v7xF1N
3GLFlbaF+cbX3F2FvksfodoQNJ5w7iyOM4sbtUtxcYZkANoawVdM8aG3OGdGct8PYGd8fiVEf5Vs
ix/i1dWR/TkTEl3ZUtqDYrTfZCFdYSqpfR95kSTwj4p7EVKV3Tl3ecC3fv9O/ojaDcGKj+kTWzii
rU6RD6Sa8R9ymZGLTUaGCyg5lyqkkNzbTBfBL8D4J3HpKutPs669oodBI2S1y88KGP2O8/jLL1dA
YE9GRkxuT3m7lb/lCbP/XdHyrhEVL7FtG1FoNF/bxAlTbuLOAn0wEbKf10TgxhpGmrIVxuDvhRtS
70RBstNJ2GKA8UYRSA7iehT2BAyVdj4kYBo3H/WBh2qlJN2bVeVKT2nNvFbdwCFygDtDTz2V3Kqi
IyL/ThDkV5Mg8f+iDlklNK6jpf3LLxbTUlFA9EkBlmVDuD6DbxBX9VSdw8rp+i5JnmBTBwS7dpR1
ZsF6H6Mto/5fvGasJjhRdLy6Kvmw0vOpAp+zz4CvFtzwhvEGmSFypjZr2go9pRkrUxhqwWcB2Ll/
Ef+oLYXhlM901jGCxkHRjX44Zs5uQqpevun3e18pMZ3Nte8YAwUCk+tzvALj1vwC8UBRO0W8q/XW
EJH8mqaqvBj0N0E0oIyqiL7P0a7wCKWtx09j1sBNrKssxNtTK5dC/Yd+UWsOhpLr1bWsst5Prvqs
xNH3f89XxjhrX4rC2PB0uZICNQvXtou8gZE7nhJld1oqWRo84ZVnWOaLtPMLhoXXOeUTQY83+AQd
Zb7qKYi4b760a3fClsrOfz2+3Hknh92XT7CwjjHmaBIXHClw89LlAt1ii5Hn049lCLnphao5f//H
CEAIaljktBtUmNcNSUB17hIkwfxCJg4va5+/AZjIDCeRQPjG2ksdjaLJftCNHwDom4+9+SCwFH8c
UJXnhCUS2XJmL3n5wNqfokqvxy4RptpZTWV1+xpRO/MxMa+oNRcXRRSLhFVMttUZsIggZ1vps1xw
Jlb3wIIF6B7rSHegL0i3QjbVySx/eg3Md5lB9TiA3bOoQkok3Dnvszj/hwe01jEKpZeyyj1DIrC4
P1xe0fItvF9fWGehR/UbKQQW3TkAQoR9qxTqte5t54aFBoVQymR+6aOCC/PBjiMhtiXNzKGF90vE
YrVURbDG/502VtYft01AZpFpHTVi+ZyCVM91KVE+2VAT1vKLafb1b1xB1yt4jYZexUJuv4xGi89t
1qzwxM80G1FqZKay2pKdlvYiTQlJgPZY3jo5LgZqMo1ixQ4Ay0itEnDnW9LZ9XzzEqiNvzBA3i9O
9d2FORfmBizcuMszZywreFcNSnToeIoZKzQbpULtMVj14plugZTtjKNbdbJsJyp8N3eEoIGV21qs
Mhm1+fS1k6HvH6hVv3hdgcewd9U8SeI1jk3gFtU0kjuILS8eRSoCHY58RhrsR6EeXl0x9XDDLzZ8
hgwhBtYiGdAFgmk1nQLRVQ0+dTO37nYhKuqgfa9PlxEaT9dyIJnklGda/gt4FASKs3b/QtvcNdj8
y6m2JKJ6FlpXZJRsgjK4/I9EToW7ugaR6X7hPdgGBo2S+zh3t8TcFJWGa6hSzqmNKHfJ9FuJ55gk
JVUja5EVnM1ChPc6J8z4NCN6/88tm/I2l6dTs5DE1iEJyM7tzVWwfZd+tnEVhecRxxQHsDl2t196
aCOpFPiCPOS/tNxYllyIchamizGLjyoSHF6yljrPXgPKgInDWUajTtnANbm4ug/BUCQ+flKLHP4Y
8mIAvjDGVhtJPX3kOujGHzqB9WSLtHBc/4GA0nqO0cBT2y//wU76v8cI/xAuYSP+eIjxfYlMNyni
bvGHrfeMS1Gw6gqD20fT81LvPQNlrypM55l5fPsJ+VIObgCAx7/bzTPES82f94nD8I7MK273dGlZ
KFu9Xp7yu82vHA+uPDA6hMu/XkyOiFtRMyXQPIrYeJzos9QoiP6doynPKjKfKHQHcq+OMDDPrzKP
OH9j0lYPcDk76LRjt4Rud4K40fDul01Q2hgjO3VuHR5BxF9sXxFFG2Y6tNsRZxRMhaY8ap01rJ5P
cQJDwoSiKtZFIrUe2DLurtLsp9kpDT6Wc/4xg92/8bF6dbYGo8V1bCQhec3mGXY22jF84GIktbY+
orkXGo/H3B71oQh5tWQ61u4ngkfGpyQ2DtNxFxZEM2TjeSvbivFW1BuUpPy5IZ3JyeS0CtKxXL3s
0UD39YRzFMpK/1tovzVuzTcNWeOWWyM2IQst8QotKvqo/W2FBk2To79BLg4PiduDzn4zqRQlvlQf
WC+RiqC06tX3hpuGmR8C0jdzmqKCEpX6MnmK/sFFxsGNqg+/n6omuhCtrZKNPP0XSVhwFQEcpecH
RndjSzFZKSC9eoW+7zvemrvv4OuYXbUDh4EUtZL9OTXYSDBdSdkc/+1dHuOitDMoHCPhcssnmNFj
kqbOaHEgcRPUDaoSaCE+WZgooekOyAjquffzLV3lurIUd4RVa5brsG/0SJP+U14+cwJQsO/gVKYu
5wiVKbz4LNCGfmPGfoAf7oknK1wwR4p3fOCxO2YuJGYFjgIhJyyX0i5Qq+KLSP/6ogst+ArqS/1c
QTKq8Ln9/uD/IveEjhsSwccjUCzEN38XS9zJCtE2QGXbr/1Hwa2NoXa45Umt8xSlNKaQtO5UlozZ
D5c0AMzXsfToRqHA3+8pwmgezYtQiYDDMd6Ikq9XrPimx0QY4rBTsJBGEIooPJAhAmowCyIASh0u
adB6AH9mvx7U5fusKLy/5KbcnLgKguRAHicX50i9rbK39HbGmpLbrShtLW7TruWutdKs5KQAT6NK
ikHBbjcuEkYZzuUNcysNK0Bi2JYr9rKg62unxO3Amp7QNc3cWco729jQE4pYED7FKhTM7XUs2Kk5
3GzAeyRRehVYYjWVpoQHEQliQK+2L36HZDpLvRthkpHsvmncp5H/bph7Uyvts4rROT20vcJZNYLD
5E9T1quiWNmWHYCrK2rE97o7H8zwG/T+5oQ7LQ3TZp0titgWynHkQD17b377JSU+y5D7Z3cenjfh
AXo2f/gXkWlweUyOAMYWgeoPIiyTwmUfniGv1awLFaJIWPz3bm4cnDL3krvgSACEEQfVUbg/r3Fw
xOSuJqIrvmHWod8DRVukgK8a3ChEpivAMKssIu+t5WxYsIdkjNK1sGYg2JxX9ImFqEJyGQbYyZB5
qkK/nw95/wGQFnd8tAWh7znFOBSPe6PyKzpNh9go52lJRnBby55upwZ18HtF6p7OM8QQV9ZocmbO
dKZ+FOchV3z32UgcDlYntVg22pTXA0YNW9TMtfLZQGzw3Y84c/rY6LqBdengugjG8PiivXXTUS6r
FnSPIA59XP0rBT3RFSseJg+mO0JnjSolww1zYyC+HOuxJkdScasS8eEpV70nb5nsFNZLLd7mCnN2
AACVAJ8J10rN1B730u7tYYmevCupV0X6EuNaGkQ5+oMGgnoFSIA7cUYpjYQ/PdPuCMj7ycKL9JIV
CvQfmn/eoNUaQbZX2sjhFpjoDM4tBKmKLC3Bew4YfhmE68nTJPoCtpvX5GuqFNwYGddGFrXQ8BmA
1P0Q9B0YMQyn8DRIUbHxnkOEBwM6fPDQN3M/nrolGwVNvep5fLQCCcOVa+3e7/eTAkD6/+BLtgwN
jDLuIUiOAEJ/3ogY8apWXa+RVT05WF0V/h67rt5tz/oUc/azBYGxtpWYg4MgvyyH9AZKvuCSviMB
iUMv++4+QCLIGGuZlh51IHXA5zV9u7FzxFcHfrW2otSkewWW0XWkc72yhYS6sjKRWkX1d0b48CMS
1aJy7ZXKfum8uwKDSuWCI7FBLB738d/YN052JAWXqh850SLL1SVLlqBpfWmzXluTx7x60VZXHtmc
uYvC9/tYFnrv5YI9Zk3ziGmfC7ja3aMl9JNqXkM/EOvzsG7cQA2idEzfOF5mYQAe6azXLmobHoeF
k7RliOir2xxUlhEw4FGJdvsmf/L10wHIc+8QUCMoqfEXfYNKcwd7DRQdblEQIcD2ZAhc431Se1mh
k2IMlM/LFBeDc5EYnyc6nT25aLz6crtupLoe6Ezks0DtRkrrG6ARwjwq3PyCrTJVHqtxP+kiT92l
As/nH23rKXXtowAKhafDHdcQTm/eMG6ufL3yhCai4nrxgxm3DTwAzSGn72d7dXYUtqpGUCn8MBoU
X8O3pq9IbRQ+mcwc0ZlqzNOSdBtXM1Q2nJ7yREWQmLdq/juez7wFjIaswBt8OdKzWe01Nau8Dg+f
o8TJKoaNC0AcroSz4bss9yOjCBrN1NwoZi5R/NEiqeRAiUwp5WO1jmr8hds/vlzGAkL86J2t5i5Q
Bw71JVcoX01IveOk7azFC0CBjff7tt7gaTin7oiMqVbU74JKj3L7gtCy5CHS+9WEmj9P1FKIZomo
oEYhEPd3UGGIaGVfXhp6inES/IA//UNIihqbaoghAw2oDVQMZTI4BHcOPdMTdj1I5PQREeqodjyA
xQNVmAn//m0P2NiDEaBFIw9wCFIUL3b7U5+VJWGz/nvsq1OE9d8T41/CrZjMWrQoHbTB4qHnJG2e
EctD65Ym09IuIQBhvlZ+H8Yyw3VQcHgxcTSM8mZ8fAMotzLuNE4twvur4PtLruQh5kw+x5fNCn58
chiM0dbiWSs8PUB/HGNzVWZI3gEG297rVyFzJA+3m4juZXUCQYQrjaABXf7aV++3Uf4Yylatuk4N
gugdCf7w4c99JXdR6gyfGyjuDrQOWdr4WGqhuSgNiTBhFIat+zCpgFKARrktM1RRDYCC+z0+/uId
eZeGC1GTr1yVsFR9G2YZPtirBOrR3+a96FtbUKXd8G14lFKF3mvVTD9XHhU8TMyEb3/t63vRXDUF
OVB69eJp8mZqQE4zUCiZaMhn6Zzugl9yvhw7L1g4vbrbhHRLomMgrB542UqjwtU/QNFcpGBRiuBc
TjE0HTKmx6CfnC9l5BUu53dxKV47b1aevceIntkp9cxyEIYb5CqAXOtmPOsf1o3Pc8tlMcxbA5+0
n4tNEXC4GSdPDbMSVrKULAfHFONjAUB18Bxak1pLbF9aKFazFs00M6khpTP2/1Ve5zK6AO5E3z5L
XCaWtr2H1gJHgXB47VmcmPMgO8EsVaxI5b1lNxUl3dUiyni1IqZZX1ue0Oqn8EWN/CgGoVxPlyH0
G1ayJCegHNu7OiCU8ZHlLqrK3/DLjeYbx01CnYDlXtNUnqd/eHuRx/K/pXkZDgj1+lqb/fBb/otp
VUZvMnoNPgpwR5qmvnHS10LJmzeathyfYg70kdhNV1rBlriFgNXiIuUdMmbBSwzW7NpnU538K7kD
HMMzmFqSvo1CexcfLI0+fKvDg90pciHP/iK8dCiedWL+U1s6MTG97PHeMi31gQWcr3O2B1h4qjlW
aOzwuzf3JWLEgBhKqAe8L3giGYzU5uRdWdS83SBEjmkoKajffaKO3dbWhPfQpE3Uh8RLvGq3T+F/
GlyHN2zrn1AqHxl3wkZgEyjJQZmCEB0vGgZjZZD8NxOGao36umrhRxyjqDh8HvszMk3pecdsbsSK
xtD/8i5fH659p9qnx0IiERL77yRMIEzl9mTo+Uempq0SO3kjDwDqs817lV3cePHsBMo5TlEb2BwS
Ntrp+olfa7ml65fS2CJpavtTAYj1lvqR8HGxRypKBorSRidy8/gr8639+6nXrxVdghTN9SvvUMQW
g2SiKAxtWvk3eDmhG3ktbDG9f7Ne4V9JqlAiX+cRBedCArDSxBYn00PlMA1q+pJ5EQgagAjnlY1/
nF+UIhQ0WfxzPqrysKfae9juP3TqvZsJl+ckhyPTbgWsArbo7E6q83JGE1HYDsc+glbCk5Oi3FIS
CpHgEnYorIHiouR77u4sIGbQx5j3OSeB0AqgCOZI0y4wGTLbLHOGPAsQjW9tWx43V0vwa56ZcKmz
NSMOyIXbRCDYhKnW4slV6w/PcZFYD2lYqOjOQ2BPmOlj8Kc9KHUnxgekp//V9Ox//SSQX5MnDaSh
pC9qgFkmt7+QK15FqSZggJ6cUa1bz/DVGmdlnQDMMwRRHzWgvPhBvtrt3Bz+oZ5NKswkbg8TaYkA
5y0umyAyt8RiQyYu82oRzL1UbtkhiErhgQZJ2h9Am8+bUkf0+Fx5mj1tsZX1hXz4FamsU5+2IDYG
SvCFbAnAfIOIqjKqAkuQ8IpdQlm2+LQgREY2oYABducBb3H64p7MT5gusGTGQAVbuqpRwQGD6zJ0
R0byQV5quxWsVnTx7ogUcbhOXi9lvCA5RiDsXv0y6baaypIh4piEOxEa+KlWz3H1f9u4s6QpTKs6
jrEj6a0KcICiS1oOcywPmiSPq5c1ytoLDCPk3PBnYPq6PA8f/EaetdfvXMQhmRL8/LooPb93lZuX
/NaTgNsUBfX0LjXRSu3WSJN4T4Equah9a0ZJYCxdw4QO/oK/zwWIZQ/DVdmP8xXuYXmdgYF4zA7/
6chk9Tb5MEazOjjQq5L5lvF/0zZy9CqbRPb0sO75XyE5JSsZW4P4mERToHdrHCFYZq60D3K5EdZb
fe396x6neYJHH5ACmR2xORS+aW2ju7OVRt4RGTBGGE69lC1BY+dusHZmZOs+TXISvHBpqXs8AwFc
tJz5TMnEIzP9KwMU48elS5srPbeApnLJYuhS+qZtyYR3xDOfLMoBRK41Qi5X5XSv1YeYO4JEWXId
UixMR5TsxQ1fxEuipGqD3MRr25leAfQlZKcvZkgsTcKcDDdX8NZ1BCSS6/QKM2f5pC5QWCRKuqY6
B+5PlOLg1qPygqzFd0SIYgIfYk0AtqaZknNXqCscky/AAeUY19MN+itxl85cpD6ZgegPFVxrF1az
1MJ5WH4EfRV14g2U9QC/fIlLZZXVigDwabA5ZH3clWg2j8Zr2QvNfw6s6bCwbeS9Gay06XhnB45E
ZHt7V9O4VGbD0203nIuFixrYfTsbGLe+waJDBSQDZVrSZzCqMDzaXt6B92eHbVUAs1CCZpTYh2IC
8+XACE7EhVzNF4ZlzSNRG3vTsfe9fqoW1/EJPQ5pfDqcf5owLqu23dUsWY53KveqtVVCaQd3zoQf
3fd9vf3SHVP80GlmIyyn79Lc+rNNxz1sPwSWIQBbYnAqkEf4HqgaljyP40wgSt7OFcp93csSxLw0
ojSDpOr3mpLECnt2XGml7tnQx7DU79NQFbyIMcE4ve0FVkvln2JgzkJTJKNQ7VxkJtqhg2tMrrz/
MT+ACb7c3fopmo2w5Q7i1W03pjRPHgiGnZ1wfywRKjqouuVpawG6or7NLOAZ/aPnVcxVVCvQC+w6
iZ+Adu/6QZIWOoxjTAGwGKGcIPkt6CmJE0kh2h1u1hKDYIyavE5gWj0n5p4R5LzS8Xe/hg+6Zg5v
1qpqdy51OfGdEz/nvYA6zQDdwuYOGiEu8/KIBwHrGweNgn6sFA8OghGyJaxqtzX72f2M/j52PziF
USF2G/ZIWOsoWoO8psSqqeybj+vht7oFTVOXBGcNTxXyT9QAvI9f2Ouy59ZBdpbCAlcCZrstCOSq
I/i77MzAQwh8GfVRjxiNbf2onZiy19nOLdOGzmTxETxKdEm5ZGtPJb8jXUnD4lUFJAL718q3z0e+
Ul5oSo3mmWhkh5Kn3tLiNWn3BiPvXvWwxKWfjef16M7A7WKFKIc8eE5AiRPNdZafg5qk68C9qS9+
rPxraKBl9pCJxTlTt8w9/Xkz/9kJKyFiUAxya8TQk+SRNVpUAFA77piXf41N7I4yx1RdcwwEM3vj
VqzuD4Muj7O5yH7HnVQpnGDuAPbR4dVPi7tTKmrrzL6qsb5AerKdANFfFD48skAY8X/TRji6yFSk
9gU5mFL1cA9M1zgaHzWvKtYKB2xduJ6x7bphDcPHnmZw+4nGW7bXiG6ZXOH3RNBwtIkqmkXbU0Wb
iO+qUxOI8vm3iqsSCUynMDOXp368nYDGOhNLFEh1ATQQnyrsN3bu3LLCPUTpabHZc9YqiquMfuB3
uxr3vvY5pjz3F4cYNLhYEfCLSnYrUaO2+NV5FCF9aS8IKWEY8lecHGRvZ7A/Lbt0r+L5WVnVAhqg
q0cxOCZ+JJGXKmFvViAMP0V/LbmszWYdPsEDXisxOZQFSZFsB61Hc9VWR/Vcx2Uhqcxku2qjkBHl
ifyIH5b7+W5yAh5iOm5u0kbF32/pZT65xkpXurCxpSWhIzCA5Zj2SRx7Y10gReJIYzR6W2QFC195
VsbgIZqvrSOAeNuB/imfvYuIxYMiOdTQrALXjjZYQa5nFSUkzUDwwC0CzApjv57S1nNyNE+jCqhr
0Q3mZ6+zqfQYKhGoFkQD+MdkX3ZLV+OzOwdPPZdia9mArONWQQ73DvCCsTBmiGuDaNztqE6QD6Qe
bL2zP9hBPpuJ5GgnKSGN1QruxFFLB/GRNtcDlweurBk/0hLRWnQnuXympo5qynfQXtGv0DEMwaKK
u+ba331+n3peM37e/nvKCzC3cRBU74ItAfrcoeTekEo3C2YrLu15rTDUCLF3n/e0SryTgRfUHR+c
AgAxFoS+Ed+kq+zHq/lFk2zSPdJUGWbNxgjDzXnX1/YvuDn4pxKzpQAIL1yrIGAlp0Vcj4gk4DBA
JF2YrarvX0qVy8pQI1PqOk1HS1hywGfu2s9QUs/k5SMcrme6mK+jLc7b+nJEfge5huwZAyJFnmHR
87SptdVWq1dTIblYSrUiyQMAVfYe+uw9mpCXhpVOHQagFMjklXCCt8JnmQVqNyfyRgCgE9v6PgOs
DnfOiQM5o9pExY5oOE0bR5jtDlm2IqFokL4eZ12jbhNkqRLhN98EElc34thfHh45FGAMMCbUKHhe
lPLiahl7gejGeLP4qJMdFmh1sPF+3vBACMg958vTUCKQp8ruzOuW5y8xOC5rP2LrCihULNsD3lDH
NytOlThS50S/rZXj7XGQZa7WWq2qi1k0RtNqNa4IS4MZURq2BA5DUK92IoJAaDUy21Sz4QQAagKZ
I1kupfM0BdfHVIAOlkx6oYDA6ZmguzYtXTTIThihZvlGe0lxdHwCVvUNTbXcTmwAupi+SA3iqxeW
Q55B85PZ+pEIc6XAP4H27MaOtWQySe7eQWcrkmzLWaZcPiCLpy3ZB3AETkk7khIIcMqZvqF2sIWC
vRe9gY7iGon5vufyBtOKNRHPA3X0hkKQKrCUUpPkmlkYHfrzgyK+PKBJnMeofXiNZ5Oga9io3qx0
yY8IJQ3gvLxJmhVxWHyLvgOTBUZ8AEOI+cvxZT+5TI8nCwDEFOK/o8483X8TWuViupz6rvNFh36s
C3mTT1Ej9P/ARxOAFmGsZW1jjJaGh5OXK8Y6tyN/t0OTSN86E7IKI+w+GkIETjhvb4+pXspyCjBc
42SN4sAmNYrvhZiCm/qIk0EEqBrE6BJev8gN634ssSF14amss3/2ek+dze7J1UXJ1jBv49qcJJBG
Zp+zvCQDTcWvnmjdLIxijNzLKDwXi4Bgn3dswXoSdZOhm2BJW7aKhyR4rk24VfP7aPh5Uxb9nZyT
u9hPzh7R4XUzJU/HCPlDMNrdFSZfU59ajSo5ECfTwpmLEnbTyE89rI20x3dHCe6IBuGeq+qs3er+
pYQ/QnmtElzljm7FNF2Qe84gcz2MYlB0jZBfDMKfxbXUgtgcKxZFbqb9/x5y5twsh9DXLjhVNjf3
XUDMuqQh+xL9iPf6qgAz5Ply3xUM16dFJr8x3KBSucN+KiYXGvpRMD5UyMtX45RfHj4yPSJr+c/f
y10giUuK6SYD1lMtpaLjB3K3G6UKvgp2XnNfmhwA7dKVMcKQrTGsYhB/93W1VBkhMB1R1s3oZDJL
+88eNIpSbznM2TSE5R+w0mFrtlvFhCcZWippSIyTIpV3+hRYlDUD6B7erhe/BWcRRaQJTyxV0ud1
wD65BfEvhrgZuxaUmGdZSEtwTr5vCULrFkg0DOmYoNIUcyJzjo6pj+ig4JxQvloSYD442tKwWUQW
zKWdEDjy0QCcRNbunitYFglM61nDsrF7P/kkwfs26LvYbKS+okoSwiy4/jV98J21TE3WwQJWewX/
pBUX9KBeFy+Udml0agqaCv1pT7GeSYi/LJM6b7oPIBXhVI6DXpgbDcMluJJqtdUxxBgqCktDYTXb
w0t8pb1mqSfgHG/2mzt9N4IUHsUXX5LoblfkLM2uPdxx3yer1nAdGVt0FGOMrypvvktz/jp4c1ur
C8cKX4w47NImRYIBr7jJoR0tMJJj51jrDlxTHOYSB6SwpTwoQF4fSr29R2RfUlUSPTFe2DVlSARk
vptfHDm5+ARFpAoDlif7KMSKRIJF7OX4MUPbztfnkFVSbnrohLQVw4ha7M3u67+ZgPi1Wt7FjBGn
LG4EvX68fBJrQhACwldM4ku40pRarE2Me+IYXkzleQxbSA4izIiMyNr2gdFCyb9bdCI5vV1L0/uI
BOPXCYP1vhhtdQgbulx+dS4bhkMV8da5rbFc6L/0wYBBnarhBz0uTi8n0XYpnxGGrpGeiGNhM4PJ
6nVEBWY9elTnfyTMWBYz/RBYA+F+5YITpKf3/KDyBBkC6VE8q5Me8Bx4K1gf30kihfg8Kz1i3VVI
tirH1/pfnWsGWaYtfqwniOhLVAYENZD2tzQUZ1EOOGNC+OTCqJLp6bMxDczvW3MXoVtcJz9+EIh4
+LPEL425TfU6uVq38UmmEFCmoeUQesibsNlvtGj37N8vDqizodJAxYIT0m4dSQr6Qyz+Prg/8GQw
NXwYo42Ht0tQakK4+DoSkhMtSREWcXKoXBLYAg3Y3DLZjIlRlsqJn5BTEAQhflCsVADKASyFSLO/
a2rPUTe56Ea2W61JubHvz8JeetWzDHys4mGJxh4L090oZCH9ifpwcJfSxkGJEvmFw+ti7oL2sMPf
3gGywtsbKDFeZSfrEs7GYOHDtyJrznY12AJ2NlN7gfeRvK38lUivggrEb8QBj9RbxCl0UakxoyFF
zeVSNxMq9FK9cn2Y+N4VUW5gN9QrYTBZmhv7TTx76RaODWL6B2Y2KwYUgs77o/5FLOv6yhouf9cK
wA9lj0TqGLiymtcjJN2ei/GjxrocPNrSdkezvncdKYzJBmfaQgUSNPgbwsmUoT3heZzcwzqTYj5s
hbqPkpmVVwsaXXGqoQMozJMuoZWGs2QXGmNl+KXWWy9gv8VLUhZYK20e/ubYeCboYB+hhfr66Tmw
KpOWs0JpH0vuyiKgY7pYubaVoWtJeLE9ypRbGsFkC+eDqEHj9u8GJSpK1SmUczjd55/iXYkFoiwz
sk8LGdMitAdOI+GjDrX5xdA2nxJfr6/HHQM4emzUpVXgOB4J/m6cWx80MJSt7iVlX9myFHzHut8S
kW6LuIdkBvLlKHz8AptVxGtQvP1wpXWrS3RiHNoIRj34B4+qIPvgk3wWvFcsI44HZLbvoifoLQH/
w/2EaDInI13/rLoyQ97+v1PgbLgpdcQjoDjzBxnn6vtolus+ecAp/xZb7imYSOIr9gp+9oYMJ6wj
eSyh4EP7/soKUfdpi3rlIse/s1eZYZNgxwA2Lpc0TivMGNATsgab8xF79v8MMg+M+nDOH0uRlaMY
qiD+j29Pj5Dmnz7G27g4IxVxX65PjDrC1fAnA+KDOSR2dgH+ZTCuLBgwjurZeZI/1zThV5hG2YrP
6dAdKog5kF75RG/ODYwXEWuNf7EeanAeLPA4x0brZ8PctEslCsJU1BRLLOTDAwtJKeMOUkmCfUIk
A63aeZolWWTQIVj2YpvQ6fjX4AT90+R+UzE9Cycd7odrA0pag35OHGz/bxwjp3PwXguu22Yc2wMa
dlx206kiWhBsGxWRYXO1C136W5HlU6Ri1i/RP9UKH1Ori5j37rb/38KKyfj/y4oKVUpQwqyjXsUa
wUBaUnffcdxufuZqjRhzfsh7eCrwGQLH+B2Tch+u8J/scrK+EIzbIedI5+7uhYLXqf9yVvf1KXu4
9A+6RdhJ7556bOLprwS9jxzXhma8cNvLN6ZmT6U8tWu2ZVWiNwOv3+DQ5l+0pPwlcCWiNRv3DwSW
R8uRVe56OH1QlMKw5IYPtHB6gLYpCd3DxXwD4WnYyv9MeIurR6v+82M/UcF0KIyRPMJSTl9yZWC4
SLOI8n3mrnRRG9rcCxb3MSdjV0deL9qtSGs5+LApcQAh/47ZAEHQ+kdHWOpFxE1ff8Qz7SrA5ohp
AdZRIXuFycSgRlTzx/aeB8j92Fku0gFv2xq1dNMJAy3v0fnzS4zxq1KVptMNlulac3eNhoScvfnv
NjbUpmiVWkfdASzERbaOHU5WrZ7HwsDBpEK9FgUjmalnVnMmXLeWsJjNugNUBEuQxsyTIDYvdmxh
W9JnUjGGQmG/3tVHkDD4fn+uf2mwelKZ5fEP0bUtZA74TxAHvYVCNhMc1ZCyP3d9AaeMF2fcmgef
SldquwOldgUzzJGBEyOaIc4lIPBFMnJ6CGxrs9piuTpi5TrhHumPfot3i0uf/Rh397e70w3vRpTn
GU0cEMECt4u2DOL7kGkdOBkN1GNqvjI+mQJglGmSIwDTXfgUFIwuqR6zHaEOsSKSxsPAAeJZnPvK
vqzd0jTvTJdi18CbmwFGGjPQAcXWB4RODWECMe0ybD59tYW6qqaTUMhfJJmqNROWUXmSOeJ0AALX
K5ov8oDvAH8mme4IacyahlRyzkNFveDtuqkx2N+HtfMFQsU7Ef6Qq5Q1pB6PYdZycfr7OpJuO7ck
C2L/F7Y8t9bMpQknGNvE7KKSmAC33DMA8TgCssglO8SXXIYvle7RprlTarCh2aAoRbSYfH3RumQY
Q/7eRecUrmcpatE5vMHs8MIEDhgOltPZBZ+dK/EW5NSGaGJtrUuQwYlaOmIX5pNWlwNP0kQYDqMU
HYhY+33F9z2uGV3kTU9NJgJUBTlT5YiM+qjOUSWjgO6kOLlUoTzZnBB2f2CDHSv+cuRJR7yIITFW
ydGuBB7XtjIKgscbPBaomCQhNXE6LWuxyMf+P2h43pYYai7xOiPMzbXD6npUfBFMQIs1bCTySY0S
yOM/6o51IEujr5AmTv+m0wORu7sEyR1yhCBeIRjH5zi2Nk2n2F7tegQz9BYV9jWlPQpPTELSdbrK
QWAabXlw2YQOGqjxmX9yUBzIt9k/aVukhKm2guFrM2NzFxBf+63yLKWgYIZ9x0IeFr8uAaA6uO/l
5UJLI+ZNCURnFJQ34wBlODyQjySCtBfmta43j6hV1/LM68lcqhOhb1yUPZknaDktPNT1Nvmv53Lm
faYNTWiMGGuTV70lft92eg3V52Klm6/giv53p7AlNa7o68mVP2ZhpfAWairh4FUV3+iS8duftuD/
m1IRm4GlIZj3fNles5IPFRtvWGj6OSdVTQO9iIqxmDKkKoZY1/zQGQn1DpfH+fOLDMWgcRb+k81B
hMMOdy/bBdfRR4wrfndv0IG/OoefCRwyg20NsEh2882jJtlyrf+Fm14hCaZ4My/pSvT5yXTgUNt+
K7v8nnGuK2WaTdd2XUFkwy3/vwmGEe+nUosUVRvSS8jhH7T3GKEidiN8LbDYrEZN+sOWmCbr6Z5H
POflk5dA/KY808J66DsVLzsIbT08FwCW3P6qGFa9aRblHQK5CC8BJGImjAkg/uX8uCYDuudoEwV1
0ODgqTTtmmqs6vy3P6WIeQoZvhu7lVoPDWFIpdd5i3s+nzn3kTyE9dNBBTPcZmCQH352+89WcCSA
bmOR5BgQeL6wrY9KAOdo0H4QOprUWmuddmv3UV+z47hU1R/+EGXMyvmD2eW+yc66g47okfnpSLVN
yiRYp9cD/9FtZ9o2GMX1L6uQ9CN+vEzvR70//inXDMJ6qK6QL88abQD8bjFioPnNinKwn4gs/HZJ
P0DzhJfFQJnfKtd14PdlXc1Wbe0U4bAohQCj0AwR1rHQVOC4wKjgA5QkEGWRNb4Rwl0rIom7kVVS
MHgmLdFP7JMQffr8uIGqJC8QBdtf5VruQVFbLltO0PbAFLVOCitee51/WyK6HRt7IELySDPYzZH1
rXlTVvWWYMo+093iJ5kMQ+yuxHL2gS6RucSarLmYUPNsXF+6x60N/N/Cp+eprgL2TTKi/lRGCMaC
TggN/JgISuhMv7kuKUOQUNc1edbEA4BRATirJXGwW1mjSRe67AIacugAfWE/aKWR21ztg0qcbaLR
9NGObus62qm+P1HCdJ7/S4CNrRfjycq0TsfE4w3IHqRZj1vgD5Q3D1ywQ74jylRNfy16ZaNSpBQY
/vksgldGwQo22mEQuh7uQRd5MMG0cWQjAkq4MuCsgSmC9Xii4UzHOrNLZIZ28MCvQamxzUYvijsV
fVYZRklonsDGN2I0qhFAJJEFyhNP0MzvVo3dGkvaoQam5WTXFX4/aCIlfZ3tu2HWE0g/ujoMBtal
i+FOKWWU+pwtulVhceHorjTkYdHOKbxaCuaaUrUk4nUK5OHCsCYZTuUdotX380GhVe67GbH89wxf
bo2cQkzy44IkParyYQFDPXNBLDe5lAYtRE5bxvt+33WTlUR+iXMGBCGL0pHr7RKhnw8C90yCt92l
fM7vrrDNfQdgYmf+9maPGFAMOobcMWbH6ks+VvSUlh8ooegzXLT3ac3sooXmy9ZPMDTJvQ1y9tIH
wVweUfO+sF8Xz0IyAZCyZKdkaiuYogrSDMjGX/nW43pGimLqFPA6EzI1b7L8DbdLxOhnviYhEEcV
Pb4SqjK77L7MTu4t2RLeEXNy2lXPbg0IaVTf2ezeSgNFpMOcULDVK1mZfoA0/oZnyeOLQB3aAh1b
qoaW+xSB4Dr24BmWTyr6ng69Gu0omYPmxhCruUyB2Y/rcg9KRc7vZc+6kk3JerQtCh8ByxbegyV0
K4swjzonqiR5gH719ZWDZchuXsSoxosSCQ6a7vmnG1i7ANg17to0yroyeIMnBAdulDHEgbbkPBch
+r7JE/aWB3I1sCcVndJoIo6yzdcJBnSGjB+/9K/r/kecb/xmDa31QCMYfAqBPLXsHzEExRJO4NA7
IoNEs+3UZPDB9QmHYy/Q79Seg6mgSNN5d3cUvW7UOIpqkLjT5mWXGX5YYghI9IYvDwE+f1UQGki1
v3tcImD8zOEhw+2j+JUnJAxZBRqjGSbQXsB7B6eZUpvYEoHslQJHrc1RhWZsRPwninsQp/SrZmt7
OcYoT+EJ4nM+MRDLu9RgBCa9HBGHNIg1RlFWHU4AjzjoKNsTghXBlikpD9ENndHOd0KqYFtfEtXH
4E1Ue30xrO025wBgAfliL8PlYjkYYZPf/fepcGDltWSVma2+wl8SfCv9Xobzv5uPfqE6bTLsbBg2
vOekJaA634g4QtWJeP9VArcg5n5WETJS3r++is19+Z7iGd4gK4HaR0rOQdzJCpAcxHCwcTet62gC
L/sNoC8A4wAVdyeWS1kzzRtsmez+jGZwXqREkB+MV6yuJHq2zPV9TxRw9biEapb8VCVpg8DtHphZ
+nQZI4QyXb1ExDelghmlnzT+Tmx8adTjEQmXF8DuYrFv1zadrFclerFNEsLUYCGKgQxzlf6y9zIX
SyctSPanFykle5cYI0yniJDLdpFvmqCLTPFHdDL6a8ftfnT+RhEwRcRdUKAQ1XB1fEZRRf+QAl7H
R8mpj9JyqA+W9WDxQsMQf7VwG9MuoWD0KyrViFqsdU15BynW97OfXJJlrjNqTPLEdIPAWYa7rPEj
dfF34spU1S3ieeLK8OPC11oOa2LnF83ZKtBWE0A9PkdUuhCG6RieG+yuDleDNN3fNOC/OQw83GBS
XmXi0SzY2Nq+bctM7MS/4m6Si/2CdaJmRm17rPUie+8bTCttygiwegBO5Sz77W24tC91KZn4aBiZ
KeHEM73EhUD3Gzuu4mERn0/UxpEO2sJJFMPyo7WTna1Y4EoU0j6K3v42gIETY/f4BA9OZVkUFN50
EoM1/PQ2fyJUIGLsZLITGPPXlr7uR5qUuIc0GWN6ei94CuHl0tLuhYLhgOrxZu+6GrKPj303L8kq
Q8js+hV5oUtVdfZP22deZPkRvr4W+31V5Is5OwU+dFvKIAMPVpoSVTvzyn2mCX+MyseadaMjcWx2
WwN8Ff8vJKG1Oak1sZAZArSNaGYa36+SI8JF52LjbI3D17qOwJSorQgdtzoKTkd/V72g3Uf9cJwU
HYhh5KxSh6Y9wPYiIRTXh+LfOMbj0mE7jSw5DGVnWQCLtlXZC9kFaGKN2/5NbXmvKsWnSMmq3CaY
yQ0j8scYviYBkjKiprZFs3X6VHdgl+ddMxbxyyNZnShuSkPzlB9Z767ZBYMnXv06LZNkuAu8glgo
Z4h0qbXMNKtg3a5cmnrsclSEQGhwUQQahwBHgpvYNMUN6eRPpfpENS26+Iw+KJbOBc56v8vDSLfu
+2Y29qDQOukM+LQSOLcbpD2KSJudqgO6zKARUoWmmo1r6ABTHZKTfiRSgCzzVEXKrT5iZDRIH7Xz
KrIfSvyicfKYk9FsOWeXH2NBc2Bxhv4duvMLDTX1L5+3o4aU6bMlVTap8diTRYcAp7VqHu7kglsl
/Ue+q4IRdvOSMfDY14VnKNCFKK5Av6uY8apbHo6lnJYqAbLfvhEYRv9G4NjnGK72H3a6DudXQw/W
pxEv5AsqDTh/ITPnlszAW+0jlFiXS1IM0xoYHDGWKv1ljcLD4jp5/ewXLtMMiefk9lW0fwtg157f
plKabV/LQ5MAGtOZCh8nOVB8I/c8UlVXChRIG8bUdKYTd1IYLcloWoLRRUuaq6HFNLY/RhjxKn0g
UcE0Q3S35m0w/50c/WJcgK1d29BmZD0rzUlEQc2xlLizlEBb+NtUNpXtr7ajZ8k9E04hCg9LwB21
WCAtHRXB70vaHe0IWtbJrfQo3NxuRtrWJQ6GgKwKZOkKgEkR/GLkVSh6GsLTvM2nhZFw5fCNrTdW
tLZGqMWfpBNaNuw1IOwYXYU+ZSAMORbwcjL1u8QZ6GYOQGcnmYdWU5rLS65qavbRSCkXOuVPtyGo
wSaFmCUvWaFggDzGicGhfcpsBPX2T/RRCkq2+YQT2aTwW9xhcZwbRaw+nBHBz5Bi/fEl/jd112AH
y/fd1KXKo4XXpgs76cHjgKywUe0l+N0vouLbWsROuRmk2uKvpBNYz/ackJohZ45DOVguX7gq2WID
Wn0VpHWEzdFvfhvE71+ApZ8cSS5v6SKWdIVKAMEQYxh+C9Owpjk4Um3vX1Vbz3bzdovIXR5XEgRr
EJLgbfI1JHTJoEWyTC7c/xloY9N9KL7SUdkbcxyiYekqduazfbBJPY3BdR7PrgujCxrL3VqxmlCu
+6dtnTR0gv0TAAfHzvf5elUrtSiXS51zMKlMIGgJEnkUfq3FJQ0+mFP7xU6yT3Ws0Mbi4UXxGlXd
VMQ0HXw9wzIQ3yoSiRXjHhaGZONgNd5z/F4hDCct9SZTwKg5XYwwmohTG5znQPK8LVf2A6lFa9u4
u2EzXKwCvFAUtc18Ejnl/iWW3bFRAeOJJGoQUJBynrvUYscX+95R17mwub8auxKP6EzrjGab0LWZ
2JLpZPAsHhNpYiY/yiWdCxr2KXO/5I53XDXTWyWB/x9gEygDStVkE9qUlGLsy1ohGD4I0obA+wng
ii9+rAmYe0SViT2AiSO1euQVcyt/+TA7OSML1kDqYmvuiWe4pFGRrHA+hipbR30WrqrCyLfFMQvD
KVPh+i93AF/3sRVoYxRepLlp+TMvkLhZk8Lw6kNRM+cbwLrFxGfsSPlAETrnVZMzd8qnoBkFuEau
8hD3fKLNpCdCgDjbk20r7xq/uxbfjFbn7aOsw8oHRiBfz6VqnBXNXI5Oexc91WFy8hYMFmkWpAp7
xxC2Q9QyY6DcM0nasuyh1CurqlHZAqJQZeFtJV/KrKgJoml7nUpNmn0ZedAUTwivoaq66SK7ncl1
lFS6CefoLBTnccyM6jsKNQfHt/uI9Vk/XwQG/FSjPozsmjp/7Cs7/TF6nDLtfVlN8vp3YHm2Wfgg
QvfM3Z/7njEVduwMc1D7wBh1d6jgWClwk47/z7H2Ut1GKnsqetfhCAhyIf/76WrHNteAxoznoZAP
LA1j01pujMUlpqn6+SWWHGPHUEsNvHUpo3xbJMLgBN41DSnXHbLXqwuK5H20wFazlnbJpjyQA5D1
SaVgWxXTIqpDU9UmKtCxJgHLgGb1b0/LsByIUXfNPTBAJ7JstCwU6wbqWoImKNX9FH/kWso7q3sg
k4yl6KAVC/XTPHtMsHB49DYjDE/eoH7JlILefkNuEJr4YUuUHTyzkJYNkQ64COztvgRoYAyyvxUK
QkW+zRledVgbu3QK5583StLOCU1USdq/yE43QmnC1te40LtLez37fAIIgBwNQvhb9TPL8d4JMZkL
yILzxKkHjKiH92XCXyTajOhf+U/wnt7J/tPbW4niZHH8Wfq7QQcWUBRHjoBCF6jyYmMQSyYZWW3C
Q1t+iUzDaFQlnr4lfe7NrltaoT0cyXs0kmZrPYIaVon/NhnuRFMedwi1kWSRFOxRILT79WmFe46c
X8qsaUKz9u2YHjAo9d0JvFbNef/pMJ+XnwsUdopUT3OAkBuEODugY6KEjop704gGb1xTebmenVsn
4aizQN24tA5LwVDboGlL56WvRtwSbOLd6SKwONGzWlZAUC0Zl73tWnkALPMi8IpsEhKQByH9oFOk
4Dn9GTB0obPN5ix64DMXxuiv02JxBql+fY/SKYwpVBZ4sBhEe1lJKEh1L9HjgWnt7rISTvtxID4Q
rAUpefTKPN58zEekfsZDryGhDwQK7ex0DuUqRV7XE2miXJHAJL3+uY6+QSW/MSte3UcEE/Dsr50k
oDjOCMrUIVfdjUC7KOGi8nfBCBQ2E3EwzPhyVe+R5ZDN4Hfsx8lRQpe1JXcAyRD8oWNKlIbESHS4
z9bRLQ2pJ36MiJNAGhk3S/YuDHfKeG+Y/HGyBZbXW/smq+1OBwTRF9PcEmv78b3+NFtf1kmYQoJ4
syrRuk8icu7QBk/Ji9XbIqIr9teMU2mkqUuG6p3ltXGkvzgBsMH+q/Jsj2OEbN43FvWd7WWZVoH3
H2uLftWp3vJGmtSSHpj6j1678SStNAc4Tc8oakbB6muEFG9WIQIkocLZU7J1WrRvqGFDDB3qzaTU
edqP3wBUMTLexKCUJfFuhZE0QoYGYhtEeCUz23yMjPcjMzaq0z/Xt1hyHUCnPWxc2Wt2WxlsQTuF
JsbsL5Ybsk9p210Q5TMovjtr1O89BVAQdv9eMYshNYbhwAO4kbWNpb10g08lbRHa31brci7s5I3E
pPaVWW95H58mWdYCLY7B4UNtW5gYADdhefIwQCxwI5xSS+EG2lFPNzNzG/25fNUC58RBrGWqHyfn
FNG29XOvF9uTUUgh5gvuKUGAFWhl9mP/EpzV10tpxRp3+PQvf3mZDF78Pjvtf9RULki2rxkQlHkA
Pvgzvt/VSuQ9HIz3alvRAQtN9YbZfGEEFvD7C2nwyFQHauAXSJ54D1EYjEn5kYjoRfvrZixq2o2n
6sRsa6ryDgptHmLjT98N7KSZ6fB3im8iUbCpm5L0LGnObglGCqJ6kHPMqjQtiYPtw8CVBJUzmoxE
+X0TkNTNDY1+5P5fuW7qMxtX26ZFz5FnQTmXeOtDybOe8Oiyoi+vGL+7VVWA3K20A33aX0AzhzuV
wGkjO96/Zft/Ew/DZXsA02qAwPMhn33ojA4yRW3wdWEC4QUTqBzZ9bANdky18OW3B/aXKtUeEPMh
TTfhz7LO1eIQMoXPr5QEg40QkGsSt9ps8C7GJSp8wNDqyfXDM2lk7p8g/bz9MgRojn/LW6mSLKPO
ETTZi0FBdSw32VUI37KRnZG2Mu2N76/ablNp4Zmpe0QuFSrHkd/xbEKKks16s33OpbSz2oSuHbff
+kDyNpZ7UF6JQ0/18l5adVYf6SEwmr/l+/v6SfPzS0elAtwdfAl/bFHnyUsgcONApxC9+H2VUnqh
SEd5uCjL1z5TGyD9430BvDyyQxLzDJPGU0zZxksrApsj9hHNbMK0Yqy8eZvqJDWyr3hp8Dxc5f59
p6s6VYcnQsedJteMXNQVtDEgAaTODuvGV7j5aLh4ManGBzzyXVsvqlTxuc+K5BE9GfogjVEPz7hC
dXKCCzP59rAmRvkHC5n1FxmZoVjDEIyIQMWV1tydJpg5c0kQ5VlR6+FgMQxl+J+24iGxbxH4/yuU
m5peTOzZtLBBceR1SI1v7+6Pl+WeBnJsGAZze3nGJcC+Efq5g0d50eHp5FdpXw2Z2Gqcb+nlIH+A
q+BBPQc4MZ5KYJt0sp50kc0JWHvlf7mEd5g47IdrdX8QF9GQvgE3N2djS99oxBMr8PfeFT+5RQBz
dGoHdt2KXWtsn+yriJHfB52xB2f+h/ZV97J+bqLJpn40GyDvNJiihUhFcodWG2AqxiC04jYKIEYW
Wc8JAurTmno4nPX21x8TNv9LwirTYfulk5xrsFd5OLrv71/EFLMbw/hCetM1R5h7CizZJuRyDRK9
G1+M59xWpbh0VbnYx+B/V/oVffCSHV0Mf/5hIBGLMP+1VVcklVgG77g1IiOqvXlqEjPfDSm6h6pL
OFFbr3AB7EAMeAal6tzzz8E/K9YRQok4X1yxBpjN/YpbjLkUAd3bvFpT/flBpzpaISw5ibIf1Q1n
ZxsWNIkcwXNE9LX2MC+xJ31VAQKCZKvCvBkmALG/46A0VwRwwp88ADY/ViSAHWJHXQKLJvspmZZy
OSK01dRWYv6+r0bEr+JLLojXWH8fvo8SJ5psiQ6AIOBh9MQUTR+jfk9dnDWyG4NRmDf02gZoYgxR
pcBL94iWOoa66yWMpwh5ijXa7v2zwsipEN4fyeZdNvjTEyJL0Wiu1N4sSL+y7TmDlI1BC3jsV3yh
c1ZIb7uAqMYLVWmkB5IQ1REnvGnGFXix9gY3E13rrS6Z7btDC9Yc33ci8wHqG75FgugULq7axq8d
O2CSHVwp6IZhgGn35JodYbEHA4uaOzg8jXyackCdPm5d85nKZApPIW7syu1XPbLz3wptKDSzol+Q
MvsCHYe4CA7svtg7vz/g7f72VQkS55mfL9Bihtssk7Xw0kZq43kf6qGAI7hsFxtQk9FI1ysV2Ecz
oGC12gXMaI74GubjNJSS/4NiqItN41jVhulqwqd4Bks+/s5eIN5xCmof2pVpSt++4ZvZF4WfH5em
D6XqoNz3eIbgwY0CXHK7iRaTAbNNVUPHyEvyjQRbHT8UX8ih85j1qIAYepa2Uys3RFl26lbC1jRV
FU+l1X8sO2ABhoqc2dwjbse2kBPVtveC+GI0SUQpG9fHhiHg8sln/3WtW58Foze6Xobnvq4KDklQ
klHDb21VQQfS7GI/r38LGdg2jHngXyEHqbpX8WzJW8csV8/FrkapAFcunXI6rnu8UmsuvR7lEPYb
vsV1sx14Ug25pPev8Sez55e7VRu2zSlW7lWCCvXpBlLGxmtYNV+RBtYYamqG4BsyWJInSHcyBYuH
nraPwfHnw30M87mPdECmggcz5417+hlr/rzBOG2mzgXgzCHa4vp6ubqsoztyZTg9MpjYigSfqEv+
VExYw5h01NLYxRm9nuFpCBUO9n0kMvi7emNGYp2ZBzaabeh/aH3KMlIASJYibSa5AybvFxq80dAq
fyVX66WtLECBxqIPbG/Q1xUVhc06dXYDoKOIBaWtsEW9KYBHuuCKJXYq2KAzTy6sTl4DNz1PvzI8
IjqxoPc6QBE8AAsT2BPltq6KjrszCTnuTZxFzYt8aDCckdLfOL//asFdgVJ6rEfs0vmdjc0E6pgg
8mEAb/pZqWIeKoEwBIEuSPCmOMjVM39kkrfp4AZBHpolE9v16qN/NF8tqIuZQ+NtY9EMNHO2dDYN
f++prCbQ0XfAHe/QWZGpTd4phOH858kaAgewkbNjbIcrBLs5x6zhW1AfoVuzZX5bOsNhusQbwLId
kuredSDfhpzgk/DuCY6fnvlx/T762vJlDpHaX8u/EKe9PPXzfNJqGDx4+YNeVJQjvRcAzLEq49yC
WxabeGGuthLGfH+a/QbYmBnPumut9DB5yymHqm+3KPfQIPJHb2wY7RGzpqZUR2jzy1vJ9HMFuPEA
MxfJDHR96W9SyioFphoJ8DNudvNcXDEKi/MyFvJcb2m+kT3ATbpIzf5j+NtyCdZorOKPA/y23awU
CE60TNqspGnETGDcAcQIK1kKNp8MrV2RCViH8qXj1dDIphL5qUmr8TxMUs3+nyCIyommZ59Yp7Ex
ZSnhH1tcSt0LWnQYspmGSKuiYYfFkJjjO8kQw5kPw4q80KSnwOKGI96qwFiWg/GDI+23ygGG4AlB
RRpfPuzGCdjGRAxAPiDyAazCEUxxLsN4a0qtMhVjtBXFHtJoI64KvRg7faqSb0omNXKRUWF2DBTX
rkSLUnLST5E63qmLj/Nwi03lT5CtAbbJjc+Vh5Vyxat4JqERla6CY7nsZoB3oUpcYPcMWGIUcb2Q
PmAJp+Uumsm983EKH4JMSSoBeeQjhwNdDhrMAic9zDZDaZ9dJ5wKx4wKpAeKuRy1dYYmtYXz5Exl
twgnlO2QGxE9rvSKOa1y1n+GMWG9+NyBh63AQepVENBZYol7j8Rd7Z4SwIN8UMC+z1BexFnZ22hk
It6F7yR0ZaHStXJGESZ1nRpiQNN7AoXeyXT5/YT6qaU42MQdNi9jueN5WrU3MduXLxJweI5BhHXD
C5iAwUUDuhjFuZOMmrI2eCuXo6WFj7xDUrlwjFHB6quKyZZxlXwG6qQ8K6IL1rG5Ia0al6eB2sm9
AOpa/9qyuOJ3HKikoNgrRD58el2UTZJw8This40rNiuDraPhxBwgDl69fTL7TFA1LVkns2MfhScJ
EhnAjAq3c7n/Y/ArLCqLl7rod6Xea34dyiYwcgD18AVoI3d7AFlV+QFYcJzHsrde0ZYms89yDQfB
4+47Uj2QlBPoSzT1CIIYAtE+y9U6Wt16c15xPEAaB5xlCtBpPf6Tz5/Qf37SLQmy5FyaNzXzCvGK
5yHkkDwc35RM4eKJh5cVDFa8NU+BvCawyHYUCyNCRjdFjB2I+cIB6DbEbYuePI+xlNolrcnet3qz
RwRDj079myHBzxj4ycKFzXjBMgwucd0BBy7n+AMey/J8G3G7krmTBKgsfTt2kT8sriydi0OYJikm
rpX8j4d4RVUkwOPUYf62aQpAPHr7GkRV0ruhehZnBvDEfnYTThjcRzuGHBEZ0jwUiX5Qf6pbvjM+
IynQXDGgMoc7Najk4s31xUOm8JrbqHeyqlJK0f2wv8glYhyIVRZWIfhPUkgbKwJmvUrB6EKtlKSH
dhvD5n/O12nZP5V1TWRfImLJNBocxsMDjqtPeBVqKn7Yk53H9SjIgFN1Ji+VY5UHWJXodd25IZbS
4PnS9gr25OZBmMzPvFV+sbvUP3zJz3eVKqLgXvKzdoVFOrVWhvYLJtHonSiAKPWUUDM0bjlSylb9
HH5eJ/f28819h+gF1KoyqV8hiqDiJHHeJ7tcszi4WaS7xiapRafeQKzG0WCgCgUSCaPXZhc3h8l1
QvR4ipQALCLgOKN+wp5MoxlVWtQHQNP6sPzNOwL0pHfR1iXQV9fQRrH0HZltiKzC+waTkJ5Vdt3w
j6d3+HpNqN77apE/0M7fjXYiD6O1AkBEyfvPrRpgI4mXcy3qlFmVxPJtg8oVWwK4Nlfz2oFpO3l/
QfXL45ru1WqOgSjavGEqrYswMaVfzfnN/J/9a93eowHLQjkM2qW1rXAGeeas0taZnaw7z7bSJg/X
L3ytdfETITnzUsFrk9iM8jo5zsDUb5h5gIGU/nyYydw6nOfHYexzUnyNYdICMsQ3bxIp76CNCwrn
LAJIyWyO613+DZKoR6o+QETCemAyvuTLkwxIipW06+3BytyW9WL8uLgKD8dua2waC/2CmbjH6P3D
pD+VZ0gNxXjjGn1ub77tjoM9LcfgDw1Hvjme71YEndCQUpjU0X4ma0emHI/sFnAYVOq82Uvk5DAB
G6zxXr0d1tCEdF7D/9zgpG035GHMbKD8B15Oh1/Cf0Ig96CVyWYdJBkcOeUaM4QKw2jhRq+SPSts
P5EwKsYbUeX7gWJYlfVDxOgEJ+DWRGFIMxMOAZ1+MOOvsqgg1ZLBsd7B+RMapzJHVG+FESvBWywG
1Shx7jNkv9fu1eY2HzFUyvT7zsXfaeHCR8l90sTfoOZE7I0aVX+qvuoqsy9Tk8Sd/CwcZFR8cE1Y
H7IAOq3SbWB8RcYJ+yU964Mw753lJLqej3EKiiJ8kh9Gd8uYWN//ESnBnDuyP1OK2Z2VzCqXvqmW
Z9oGETmJXxyKeyBDL0ohywxvOIMZmyEA9657ht9HwiwXd8+WwbtBkoD6PBVO/6MBwdNmPml8TtKQ
UyGKeA+nQgc58MTjMU33ZKrdj7bzJGUP9q4kSvYYw5qQsT9uRmMqjfVwg8xmtOFULBDEMFvUBhpQ
MhMcJUPad8MprTws2qhDODYb2bjGOH90yqpNKYDHQWNKXH++joWz1fbonFgCKTiHEQQWjslAVnkJ
tj+yfrhpco+zBv/mHL3H+JRnJ0BTGDlfesnufDY9RZ9k31Z43cqfh1PiVkOuTOSfvw8u5934iRBo
2bkZlqRBs5GyqVOlXgEtuJtHwwE9v3bnr0xnb05v+srYOmLS8qcdyWAkKuEIaGFdZ+gcQROxdNar
+aqr7vo96fGnFkZDla50wXF/qJJZ8STjcam5nvDekNVk503IwXkmz3xyntFQfKjzyWJU+Zd560C3
ZfE0zpqBYpZ4E/u0Ww5Me/nty94K9S2Hm1JuGkM7eEc9QaRKik7EcISA2j5i0d8t2oX9vlFe8DBZ
0bc5HvFcJOybdFqFwL7sjJl5NFqUiFcxqktBz2otZ6BeOhDcZNA9kYSF0P1DrTSXg/u8JeNaSooT
wL1Ja8PhS7WFyFkPkr+Umci4hBbEJ+UhZ0s642qIse/5ksaJlTUYnn0c+A0Dl3aaUIZFqYWESlau
QAKwuUCZl9EsGkgQOTlThO/Un7eywT7z7+NBw9Kub4VQ4I8PTNV04r0GMCaTnnfloyOYlDiAOwy3
xINdCKHvj/sZV5V1Ys8OcdIN6cXcjrTASQvjJn82ldxRSiTrmN6h7msTR9BZkQ9+wlg4+QzvGoLg
YlUFWbNCRwnl5hu1S1b+eGijQk6LYvziyEmqagMHCG6u43n0HQms7qhdNATOhxRlz6mTcRGg8gNo
GEyZS3x2rvbpCvkneoiMPRYWz+8+EeGNGAKFRQRkyBy/hmTxU7fGepcPc6pIigLzbqMCtoJbXY2O
xl/8EC9LC7URTJtOM99CZmKWOmVZjQWcK1v1cGpZfV7uGAq2KD3zBqKmE/sPylJ4wO7MBJ72FWF9
hYc32cs71AhXcfaaxIHTyBNn8z5wf3JsFxBc/EYVuSbISirR00xUXQcp/d4KGTOqz3NJrW2y3oAn
Y8UGLCey9CDD/CBKHdf5oJxZ5z2vQ3kxP1CFMVnplsenAa+euWg70u2mVBfPeaAc8dy666PanbFj
c1ohASs8xaqCAA8wyDS35llsp/CQDcQNbDLy/ZspNrbWF+/BoLpEj5cWHdd+L5UHRDob7iGhtmL+
+DJ/VlT8I4NHYFcFkd7S4zcMmg5ktur1ry7jv3jhO1sQ4ioySZLhRz/ksBddoRXSOY6flol+x7DA
c7CSGCOMxh5M6a0+rprOf/ZtbV50BUZrmFN873Ev2DgnjalPFXnIqwOodQbQS1Z3DZ4wUHvrvo7r
LBi7eYjgDsywseSlxdgIwfn/iF/q+4FrWrU6S61MvXxXrrDadBj+jakdkg7X4DU+Lp3oo5cFICb4
ALkWEXFqxwA7XZXyu6STIOANrsNTnCm8CSE++XdptWxER17RLcLhJy75DkFdSCgPLn1IgbsidxwK
UqOTofeIQQ6FQ5FyLC4Pry3NHPabm5ByCynDE97RWq0QjFXYp9o1xa7+GSv7Ui8uxRhojj2t1Dq0
hFRiKA2DHzKCALd6EYZM0DHFn2mpd9HdkI5Su2kDBfbRKWaRlz+jFe5lkU1SIPEYwfFqvTXnO2Gn
ga3gt5bFJiY7OnKE8hoFSuUPZj2UrBc6GF2i5ajIGM+NFhoS6GXUqtjZ80j/YANffD2Ue2yFK/nu
8HDKFkWOCXM/TI/zqyCF02RiQy2PA+MMaetrk/N/rs7K+3zf2mXrwcqaxX4aWkpfhhnhMs4lC9K/
ktkhGLrtxuIiqiYguR3KyVkWwcB55q1R3EeHf9bW33X4f3dSw1GKIddY7+ULHKawFUxG3zuNoA9M
2YA2vzN4hjfPzWwUvhlOJIu1F6bco+c4Lgih3CTXTmVvOcggtaWw1anXfNxAZOZqn/DOztnl8hbA
uNlmASwCo7Ix6xJjfxNyAdolCYQV3kflSGwrFxvKptb36WQRfUehbvh6wcf5VO3Fgr3JATyvYJ7j
INnSm9ExCo+HYjj0jX8EJw7CSQ8gvZUGa4vUCczHjJoQSC95acomQOVnTAhT3uNUdKNZqnBzlqa7
OzOG6+K0boohlci30ADdzDNJ5BfcCNqfI3P+ViVv9KWd3IZA7JSz2WoS4VBPCnCJ684W+q5r/Bxh
QUq5ofx5+21aG35B+Yw6xmNldL7dD28x9zZ2D+ux7GcI1um8XMqCLypEM8bZpmJNwdiiZZ5UC7Ld
w5+xycHp7j3UQny6mZOTmk9N7X3waWJIRuucyGAKhOOacHcKjBmneO+2M/tFPDA6F/JpJRBWVsD1
g/mbwWOJA0sGnIxcUpXgwzWakSziAHMz7GmZo0upln4DXCcQZd1sJfv6EdKf+p3rKvO/YUva2Cq7
NFWVV/b1HBNSA/IBdD3pQTOMTsIQxzI+nihEusoiu+XlVecA8EX6igalFHuVKPQvJnXCIoFyAOqj
4tmRt6YRyXBFtZqqWrznm43T92uAZJqgdpMqmYn5qmdffAA7E78dhtUmKWM8IZLJcPf29SyNddqW
PmdqDD6BQqnrVSOgmgfznjfgDnhMe2gmjwAO8C3W+Hh4cj8eanNoomkIZtLEF4PcAfMpPEYO/epT
/Z8d/wSqwQn92cWxiK8MLqBEtDDreu8Vuk8uvYUIfjwtmYXbnLYIYFIL95LHLIP3TV/7MHzvlwkP
/RQclWveZNCW7g6hiyzRLYxEkQwx6WemPC5VtHqxk1k2gFzBAKMSVI/sjF3NNcHAUVIQv7x7a+kg
GGfLP8u54OTuom8qQlECAjXm0tx57ZAFfmSfUjLZ1iWzyMOVU/i3hb1qlebqxdw9o9ZLduFRMSdV
IAIErAd3UVK7L4MO6zbaICrpNiLvHADKNFgaURfngmrSznPh41n+ho2+l68Sn03VzHlOB0yTH0gs
5n9ek2Lm9Cl7GIiST3H3wmLKaDncIC+1dXCfhtuGPHEtn67pIBQktQMOFVorIMz403l8SORqR/VZ
fWQsWf/VgYSv8PzUKgIZFkjHIYPLKhRNdYiWXLIdO3/HBpVMapoQYNMP8t0GVy9OAUbJBYbEkOj7
givB/Dos4aRE/tPE+b/CFWvkvKs7A3RwcCSgXLIhFgH0JziUlkz+k3FDaN27wBNGOkuftekJ1bwj
5i4vXjVlz71k9jfIN594w1M3lMhreyYGWLKAmib2rk7MsjXX7uJk4YmQnt2MMnBR+a0vkTohvb5q
iSrGLM/LDCEzYp/sB9oJ9o27BRyYFEQGbJi4L2aqmggKwGBkoo4vWRAe5bTMfMBuwC4A/io7KhAq
PqlNzg8VWMqSL4UbBtZePtpYz3CRzNiO0/lPiw+Npc0cSCL5S+0aF2y3NTi79xhtR07vltczTAgG
yHxj0fZcEomWGbfIgr79GdOzdtf74sC0sDNjw7vlusqD/OD7p8sPmp+t4IaTOye+oxGiIWtvsqNX
xI1sF3dQwJodpZ1egpqSJr7kJmpapruWL6Eb+WoQN+y9g6rtw2J61toT2viOSNSSNo/C1EXZgEds
/bZfqelEfic//FhoOCj4WIlYrnFA0C3i0wAf22l8m+l18H8uiIIWp3wE/GecKm2mLhjgFivOShnw
6yq3RSxid/PsUP6v8ZgRH4SQsFnDQLjibmlZ4Yvkfmm7xa0obMOoPrEvRYBog9Zk54PeBQ8bLtFQ
T5fJZpx7YrBFt9xorWyDAgWRBzdvFxDgiw2e1Bwt+EDm9fGIyXqZw8DMTPNYMvaZMM1BcFQkB7xQ
n94l4+2l8SO6qQUjY69+RsXCr/wl5dKMVUx/G6Tc9kSLEoTkaqGT5zkxrFp2qQmnnXv8g21J8U0l
HiPg+ZsK3URBntBGFCf67HYCxoiK9CukNDd3cUEtDzfYLHy7kwKudxK2G9lxwZNHEJGNhG023wmN
t6hZcoNNSGnbF/0VIqsu4B7Z1oZB25nGae9z60Wz6ARGoYUAuJdnslOfX7YObMzfCP4ErOB7+aEx
LaQBYe078ia77z8gvPsI7fygjjop+2F/BP1Pn6RuMDnR8L5XB7HkYqhukm/7020XGalga5mahbnN
RlJryDhcymwvAo4KubL80kgxjRK3xNdc+J4tItfHorL2dpPLzz91mhTqpCB86K9EEo9XJciOZ3Q1
4GTsxmJQpvfeTRhptsWZEkOPJfh/9WWMf7FzRYVc7wFKAFl8YZsSHV8knmuxJnO2BscMY7bTqyi4
Cq/jBOwggrprRthBfTqO5Aa7j5frppBBr+0lCEA8B9nGFh6qG6zzb9P0+8XyanOjRRSX4t0LSF78
UdfQew/hhYqI4RH7EfFs8mlSeqVwQ3SbPkc+PbWvIkLhkfol0lJvfIrgq+FlvQz1myISJBi/Hztt
W94ZxXUCkFh8DOojZgO+tLiZcxZq3UWxvcZVLpu6u2UTbElKUZBRf66hRKQOp5/o+gf+Z5WtN0iQ
mHzgDGJzDC4Bi5Ynrcer7o/hRf1NFpONafQzG8kXgSHRbFlXfUecZ3Ej4h/H0oJPQwrgoNbJwx9L
O//zYnci83UkV+Sjsdq+bkTvZ9hHHBrDRagUuPk6FeoUVZGG26UOw8v3biOgw8MW3JxE7GbXM8nf
rD8IZwC474Dd0UPqexqWG9kkg02gED+h8HgykOBfu0FbnJ4RFLzOsevk/kAY3yJj2Sn9bDvM46BN
Gz+e9zn+3cd3j5mnhMox++Qr8hpBplZWoevccCnspY+C1rv/LqcDC8IuU7pD2kDYV3+aAeFoskKI
ECPcgTPWhBUEhrL154kE4Yu2NBC8PDVLAo0HLcorJw9xa7kt1K4amJD6i7FENidVaySzEPihWO3a
me/GfQdVp9MWP8jxMTg8luVqPIX/Ga+/oTPTUWiq/NzaW1kgC2Phi6ZgjVyWmKdY71GPUjovXH+X
Ls1QnzCyjwQw7EsWLSTQQDntEcPVB+asCzU+/q4tN4FqvTCYwjF3zl9Q79ULl3C5N/vjUW4eAXD+
7uwsDyrZT5h2Z2KerNTYJeOcj2d2TCK2HgaUJ0jvuTCieT6VZBQ1zXbvy5WyeHhkIWt/9lqmllXm
/UzudtJHj0D2sDBAh1vkm5aZ36eJYAJeBCWSGhaz4h5+ReQbP4ak8D4L+Gf8KwC8LzSyqjawx0zF
bawIiOVdZZm4pAgmSOyNCULsjVmb5unOZu4ES4+lLV5bo+5/sJTrC+Ss31izv3L8dddPKjHaWN9D
8O6Ohg7nUvf/dXiAk2FW38Ik8Kwbkrw+L4SJh1gMn8lXwoX38NNamJX9OodO1jCnGcXWQO10YJjg
lH6i/1NJf1qvM/D6tAxI08jno1RQSd3u7LQ5KVGOfMUFKfoKSzhG8JC8HvHqtcuuaZ+/xVRTeGLX
UFSSD1iNvD6d4fy9T/o+vmD1L/Vy2+yIYK7ZETW9CGJkCGnhfaQnZX85G3mnxhhW7l5NQy5AyGbE
zYvCM3xVXHJCzmHDa7CiSwZbezai2vg7T0cY1aKFjYN2Nd3GVWsMlSfeLKLnP4VkthT+4MpWgSZn
pFTJB9T8OiGuLB8aEMekfeQSB/Nq+KJIfTt+7VXaOb1fs8jXCRslxH3E4EjhoMuFsvOv+QRtImWi
lzf7V6ttQKeFrFlxkrLYSUgbe1MS7FM4XOklCGgItOTt1bznqkJdd9W3Vm8TDek5XHN0ysIV7Xrr
fb8Il29GZD1LTks8ryBgr3o4zdPBADQe/IrHbtK2HLnLi6l+7XUNWUW1dPf8doLLSx6KMU/2id87
RyHP88CqVTOXD7cPKohMZUZqLAmEQb7c7xsPruf6BkvXysc+A1rc0tsL0d6Ps4sBzBeZEfjxmRDi
ct5goqTodihUtFei5GBPxw6fcwnd3nEHQKXB2kayMyCnSG5rWE6/FOFQG19fB1uVe6Z4VncqVsvl
XKzGsfRhK4vwS2dDKqy9BrAC+ZEWEpa3qB1iNvvMeYunDd+OTUOMBT77X5VfoTGNh0XD6DL1H4o6
+EsMSpQyGe0BrObkRsvGTJnxOEi9QOdp1w9crEzaZrafyNJjaU6ojFVT2nfng7Md71zYRAluF5l0
22mv+ooiBKOnrMar1UrQDi8ZZleLLB0MpsmeD1IRJ8jp8A32p8Xnv+gK+yIKDygEC/xJFpTZnfb6
6/v3quYTho55D6w0kHGd4g2AP/rh5MMzKj+goWtja6igom7KdxHnvQWrZsuAtG2jwtdmn1YZZ16b
JRmY/9434gQoHzhufpkrS0ysHROUgURWgPE1ipODzA/xnwdRVje5Ye2kAW1kH+L2BCpMYebM4iu1
5uK6171IIc94roF9Coeo2NKjEWdCQp7ofbHuemLGs1wj8S0UDjY+WCGSdKaAa3gI3x1D+ov3pU0U
DrgOQaEsMjQIXxA0c4cihE8zz9oz/OtAUV5ok2Np7VbWex91wdhJPrfiyz9r07K8o7WsmjIVMzPi
vE5wPauu1b8M5iiEWV7mtxJjMCqYx11pBAW+64x2gyTfpRje+j7Muiyv+V9M0yHf6cz0y1zXS9e4
jJ57K71Ytwk0T6GZFPvjQXPEx0jXeL/XFykLdhtgrTqtgqibQcTuzx/oCSNsfJgBjnQ04DPlA4rA
nxQH8cevImPNFhwCBptmZPr9jhxq/Ya1+42lDnE0EzqrvKUtRl8ILSXNy2J/u4cJ5Hv7UMkeJwck
qU3VkfggGJH4fAHaaK9wjU4QB8mBCGlc/cb+VxaK7fvlYCtKLQXFPDgnSrvKVPTT6ocbV8d4AsXP
4XuIAThfqW/A9kBzqlekt+rijypyfGIAoOHiY+X33nudIlyukJx2UvjPkcpSNcgEGGT4LUUP+t1s
Klqaoceg76vXQPZhbHhuyhcVktKltTOyZGT6vrM/uZq2AilY05jcukiTx8EMnjbERBsqzCbvM/8m
WRVHlVSmg3kfOLHXm+dvmXNZttFkqMSMpV6mMbENXtHabksV1BSS4/Om9h9wHb8NO+zjYhclIfYg
774B2eZ09QSeURZ3pyZeRR7kSpbsWLLJFG6ug5sfLLcHgSzuHTXWJaYZav1fFLGubXqieSTwmFJO
tExwb8smqZ06P+y6CHLf3aPLbfIxwPjLsltE8ZcyNPwuyoHhKBBrz9VuFmarA3cvnl8Hnhi11Wgt
Lznq72djUURjOJ0wa8aMwu13xaDfg4F4FTkgCfIeBRKy1alkbuEeJxyK44HsHCEtE7NWJO/I25/C
Nih5ZHl7hXqxN6E7HOT0wkmkctQ+bZwqhN/ST1z6K8g8PtZ0+RcJREJtGZZQh9jSrzc7/5sBzKgM
OG6HQMKNEfcb4IRr2T7FLT4jfhovRCUU2gMpl4hgL03gjT1aZSYldYVCbyEh1ekwEEi3CpCbaIiM
c06UbcGOwL5RuH2iEny7LqMWsFepn9642Y3Xjti0PprrlS4EyKCmUKpsYi4kv8r2nYtlDp5I8w5k
jrU8sD0Wz16zvrILutnY2tfaxzWhjWqx7PE/7ZEVcQapr9xCX5W4k6UuZMgtZF5P2MfHbhNupRB8
zu8txjZs1PVBnqgjcVLcR3YSg0dFpB8Cv5yCwh44W1JI2nM73s+3peDqoKjnul3k0eCWB1KBk2PQ
EK65/79wJUnWwfuMBKBJgAYzXt3Ar8+9Z+lQQRBGevxmguAwoj2cmIt3Sol6lUic0FTsJ9V25wVh
EDqkshm68HsTw+a+y3UJpimzwf35Evurf9RBTCwy1M9r5jgGy0d66hWm1Qg9MYyaWfGaWIZhzFQn
AKTMX4my+WtMwU+DlfLkEGd8AxCKMrfeF111qY+fjb68PQ2Q6CP2Axrf+LXdqwxtClFO9yUGoB8j
VhAoPpEwhizOe/r8vMcaDzdc+GZR5cSTDyPTqUn++OlDnhUwSOPJZ60fsnma5mTyVzlEllpBUsml
z4LXhESOPUee74Ghd9Pkr0PNmHCpPg63guOQcMWa9PCzUwfzIYwr7aLtN/G74vUya4+leXbPlM91
wseIf3c8FYh//9X0+c0agcVjmHDP6lunymNrUaIyhOH0Nylyft0fSP3ajnFpQ+nQLJvb+lmvHJK8
C5upFVL8pbNKaAISTH2sSQ94hNQgbvssXhUpcoQUuDa3BcerW4xG2pZhWYoKzyK2L/3tH1rHISbC
PTGkLDqYVV4Fr9nzL6bHvviJju/k0sm+GI42lloY87o0NRTJH1M3vf3FlCA59s/kd91Lx9aAKsD3
fMRFQ1UHkdheS89Py7Jf87nfrjrBNgIW0RtV33gmCMWl1qb4lkGRbVKrPItNePlwuCAhifA+T198
pS25NUVrgZddlZeXJcCnw44h79FIESf5thfnW+1bczxJhrNOAKBbvIf1UGb/DNYcwIVIVonfNuku
/AIVd45gbF/m6CE+sGfbM25pkwDi7roDo07kjviMuvkgYGABMP6r0Ozqs0mO+nZSPq2Oo79215av
QRFD3RqdvYrbC3m7iBjkeARgnnTTPCowjn6afOMcMGvhB0fmU55ho48vEib5ibX7jRcBrIUm+NhW
ewPbl2OVYEce+EG8rdHsO8fX/qCCd91XQvSxUbQjVMS+nF9fA0t2pXU04wmhXlaDyxc33QxuayMi
bqCseTsSsjhnYbjJBnsg/87yqeUFGiBhDdOvIPWMuBuUcBAY7PXlw6Ya6lpfomIx0xCwgkGfilqF
Ve8hYC72nKQsDBnfWHy9GO7kM+tDpi9huguIiJpJz2HosNtV/P+hlcev/wLrvg05stbAat6MEFoI
vJb4OM6kMZhyttqKbuYxGGUd/vwvARMNxDtwUYWOPx20loDU2x9jQj4i9jLE6l88RWKi5BzJnxGZ
QKD89I004ToO3bDwnAAyelewpEMwvWI7Wqx71SeoYx2A0XYhPx/onf+h8Psn2br7g9kiiwtBDUWk
GeVodyiu2YW+yssr9IAMSHpg8tGYK88chYVDFJhIBlXTnzNpR0eSsIudiO34tOhBCJ2dGsflzlP8
P/tngEBLfYJgzrllqPcVBChLsjE/a/Z5bg45O1pvu7ukLwWFSXhKez3gGd1yAJPK4yiNojZkpneq
rSg77/68LC7VeanxqqVCD/nDeY44EW6gQYRHsikBRkCLEAW+wtblHu08fcmULj1rKbbE3wcjqO9n
6TMAALKS12KbijnIF7kkeLF4YC9l78ZZ04+4vODF7Y2flYOz3xt8ujGcuf4MpESObXN8LIe8Ntfu
SmpG3L3+l01PeZWe98Z/rn+rfrEeLHIArTZd0RkRYFJt8lMUrIN0zAeKr9DRLlZST0oBifbbB/Hg
hBRSSjNGSiCjbnwbnU071ThDZ5BlGqXfJqEc+giC+EiXu5Or/CVrxFHtKiYByqBZMkgvGemMI5ir
BcJ+YtgX4HfOKaB6Xfq9ErMQAyEG5E/bK0WomqJhVllxiPDoOKz2V9xersKxKgnSg/XxSbDgbmi4
oYakcV38dSB8p2eHzKAOGwoQ5XltVF3uG5z81uMbPlvuAxVOFLPn2p1lqWKDLetWZi6TT8vdFtnz
IpSIHO5NVpIPvUGle2QR4gtBngEhQcGZ9ioS9IfesgBlZyh9pyVCxI9YjA3AKzXHel+OgkOZje7/
0BmH4DEkPavbTSehjdKSA8gM7YQSLwsLDfBs9MIt/s5BhqF+H3SFdQ7Mil3PwYhs1w2G1maNof6r
cbvprKOwCPTPLZaT2jdJKFbN3kIVlyiBkAP20XvHG9zdiu1GffWBXGQfxEUUbneMLFgAR3KGo/X9
xtMfSRsvKZHB7MYTpBwdgRzxKgrb6fU0g9Vw+gEiMtIZw8L7/QdDMpVoNgjbSZmyaXm6Omb7PP8B
ZO9UbgN1Z7Zoxs03Tlnes4u/L5xVgd8yrtn4Im6+v4YkwBtae3+CSlHXlXu+xqP+2wJayHvv4frs
Cyj57cQKrY2E/Isjwpw8jeAqY6Wm+6hU/N2PksB8V9lXl+vMChUYZbxUXaAfs4zeBEgC5zEDglE6
QRE3tW6EqqtxVsj1pq+Q44q8PujMd0AmyBK9Kq4N5AMfGOlOVGGKxfbEioydGjVay92VIomIwjIn
488ant1u99HBznJvzh3IEUbqvpE6EoFPCI8d6EkXSYhqwRBkXNBH/6i+rU8oGZJQczjnK6Eoe2T3
Od+F8Br/1o4PIKZxESamyacc2lP357tCEGPfhbFiCgejCfSsxnJsXCKibzhw1dBsfa97D/hiIE6y
r3+tgZ2o0YE0/SHsGDJLOtgnLzdvtObkiB9SfBq8Z7iVLJ9BUVvILqv//nx23al9t+KoFKKkY/uY
mxpfkqJ/dHKdaC1sazEpCawNjiNg8hAfn/tz78/QU+Sta/mBiXc34HvbCeSNr3EuhHSfHANcgD1f
DTYrlL32J3oGKkzQUOMpyZTx1yAWt+gyE3cswlADO3IuAcHxrCxzCKZjVDmy3+SjSj3GWqcWk6aG
HYjwEiuvP48sTIXmplDGIBpNhxuOBA6c63gj12BQAW2+tqNT213n30eMFSxM4WJvL5AZ6Z633vEc
lU0aYxva5bK0SaChZCFdQ9gjerZfw5xybCPV7Od+3vCrIXa+iPAqMP3iSXHY+xF54qTGM4yR+5LU
igzHH7L1Tfg89qRvn+2ZuZosvcQjD3hMaB/razdsGadg1Ir8EP02i5Cfapvm8fJELFcBeSsl+13f
zBWXN0meTnzGODdUQEWndiFTQau/gU2QNtsOvLh8ipKQkjPHwC1xdJzj2+N0Jm2MmnNmgTuTJaGY
z9jnpifjfYX9+qh0mwpYJXaPKr6J9QSALLHjYhBFo3WuzU8+kQ7iLVL/KvktRBMOUnKO+27hwbJn
DhGChvCjmy4zdKXCYL2PrYu8XHS+LNEcnqF0/KKJGKf/FjA64bkqb9Bpnwf31ywDUUeMjXpYm/RC
sH5QOVZbFju52fh8Y+3+/oZnb21RPHUt0GpAtDWhbrytg3SC+71k74lXjsgwMXddJXrd/nkLW0g7
7uXDcJ6dUEUzLxxAgj94pQ/lWch/uebxQ17nsrKIMr8CO71WyZgzjwc2EjJw7XZ2FhGC/+BiWWs5
h07lTTQltSIgz+oSwBbETRILPxsbWkKAy7UDvdM/zDxJviSBR5i6gV6jnEfrjfzqGDQ35JMJ0T+B
JWTTYhvgeanhS/xEwcN6YtciLuPB0s7levhp9qAq9yIVRZp+VTww8sL1zvpv5GwwGzAQYnfIfekM
+lsxL6w1sKEadytE3YkYjHFfO76XtJOnY7/1aJM4I37jgokCfqahW6D4uL6rnOiZ6B7vqWkPAMEp
aNrMaXAOWh0EenlSH1pvsaZN6KNH3xHVdcpy2nsAgiZ2H+s52ekobo96eIqXMiGKWWdLoQ0N8qLt
/dapJ55NffvIgQTHlxZrkfZUIeLVX/EGrTBnn+/ioF2Hq0F+iHj4qqzhTa3yzRsgCvKjIWizK/sE
e9mVFYMsLkdE8MvWqHKzgEH0gis6KFcPK/5zTSh6NdHhyQkVKa56iScfuPHU5z6NEkczemQU5XNj
PvUeZ9cS1CMfNndZYy3o9xdGpa21ysVNcFOkGg3AT3Uh6+QpbHZZCzy5Lb59SJr3hl7WBYjig8SW
/i1nTq03vugwmrrBdI0NMUJ+KpYOEYVBMc3WI6M5JWUvSbepaG6EiVQHNB42rs0ZHcbZux5+ovxM
zzVpcncZkZJee49Em9BvUr5fVh7k3e0F9Lv6ztgkxIfNS+ZYUh63nQVF0+/Vjb++FS9DJDmTx1gY
QTeHI6dJb87JyBaSxjUHyyJAP1A9XKDrWE4t7vks6HLTUaN20VtjcvQXP9EMAXKW5xOBh6RFW3oV
LIpw1zl+rtzLJtZv26PDf47RKT66X1Oz1QdqWdxysr49xMDHda0lhqrkIkVMPTgb/0vjd8JOIo9R
ToFBY2Jpk6npSiQSCmK7j6vwhH8MluTG8BlbxI2CYcisNjgP10cWKyasgzCVMAwatSzNXZSjxR1e
NRvqgX6PqAO8OupJPJUkmGGDzLuYVuM2fp0GwNY94e0QMpO5gb0245wodxeEeSCP0cexm4OriYyh
kNS4D/aGDpU4F7lLVfV0WOZcm1YFZ7AdPRh+Hq57LiDR1J7+2zGGy+fqOfzh+bcXW2SRAnoGqIDL
6pkbTAX6ZUKu/AkVUESzhGHaFgBT/u6jBhK8ZqQzUl4STkZC8GT/nPDvGHh/56WPJ/+q8FwI3/Tw
N4orIF3Z2YHDwyTbvZLvv5ouJWReZtzJWSQsMFGesPCkFcw9rDF00ybclbjHn7KAtAg3oAMQ8wRO
7qIZbWglEVw7/pz2C8B1x7woT/Vtn6oGnhyfuDKleYZ83g7v9//BoHTLwEomU65auujYo+/EbT+M
pel5IU8yqqESpC3N8zXyys/tIQ6O4S0Ail47/kiELUhuijfjUWPdeEicTB6wlacZGF3lZ+KhMFse
9BsDzbkHyJanb8/wLCjhgPu40cVZomKQCjmuILmYxrRLpC5izzA/MI8IL3oY7Pnrt5NrUNPUWiOO
DpQDaa/IfeT3SDKhOfntiCzYAoSb6kGH+AsmenSWznD8FTLWN5Ff3Cn4NMNyo7CmNsDR0jOd+xFJ
CMJxg3Zc9gD2PbiF2zmdiQQNC8iLrl7V3K3K9VC3fxHlJAkf2YxBUfhNoB+8J/aglmcwxQ5uDVJp
zc3hisez2L7cI8A7IOMUTAON2c+PVsLG+oEjFsiH3Q4XUvQhhTBvsz7QVL+MDZYWDZ5E8yfOJUJv
A72KzZRKshxBnRkCmyYv2A9ZACrYOmXRq/Hup0Ivk8KJvfjJbustZdaYeXr5QscVIwzb1QqiZhHr
onYi7wycoF8GBKYskB3jteid7o4CHrgx7GSSx8qXB8MS+AG8FbGg2jb6j1IaNt/4z9kYeqEIGA9u
V/77bGZz0jHR3z1tSu0JdwXzXiws0yyH216wbURgQ3RQweFbdHGM8O/wGgkSPbqIc961PzsRiZZB
ro0wUWEiWdeuEYxJhSZ/A+CQ6HCVpc4X6R84Y2mfGyVU1rFXfOvyv2vsDo4at4PUhkH31+7KjE/G
OyqlgmbYhsKpQx6Fn4f3OAe/TESSeVInm+CqXGmvlPNIUgT/n+GJ0svGJdGe2jHNvtddnpG4NF+b
6sxPKwourEHkhAaKTbu60BAvzZG3J6kvYu/G3svlCjm8qhTkUe45jldwe45K6h3bfD858eDlOhuy
bNr6pYCssVMVPKQ/3uO9M03O/sLLdxdGxaNzJ1BZz2LZUQbP61tTqpxuHG/JV8P9IwHgTTnEDYri
XzZn+dMWSBCLZcu4LtJNFRXupd4u/PkbSTHSGx2xdsA3Pro+ekn5JR2UtOothVvrasqPfivr0QfQ
+1PQdGyVJedaIVZabtDl6L8PfL/S1kQGxYYPX0Hws58mgKjsPn1iloC3FFJp78inI4wvUSemBeAf
URriNYE4Ig1vItrc5bCHuWKNRKZPT6CM9pa0BrGE8nR2Bzn2IpbXVUZ6qiN4MplJNSsUo1KNKidK
4NV3fJHXuryJ7DYWLJ6g35qefrrnyYYEXVVCS044fWGOtkN+GIE/H4joqNyhzUqC16Vz4f2BnHef
MRhnX3x+6es0lrxJftG5UFut+DqXlduZ3fq1q9CqxkI5wVQuvUYa2cvUxd9+oFqEshijeveGl2OJ
HXrvfTjGihfiHBpMOSRwbCpZtG1jIpB7GVyoROnfa2BWOMA2j0xhVOV01oOWFH+YorXLeXnX35XW
0VL7n8AYgXdpHklu1ljmOZksoF3pFU8+WXcB4M/tl9cFm0jKbnGI9qwWV5U7VKqvCEaToNtHN8CA
KFYECaW4e4eYTKOMQ2AF9HVwBnZRbss8UbjY5A7muLn/xYtuvbWTNEpt0o0NUc700ttPvu5QImFx
B0dV2HI8DWgIqHb7Q60IbBMA+ItsbLFkn4JYdetOnyNyJtqiSLXMQebzxDZke/vZ1obhnU7oHPav
y76rYmq1ExHJr/tACMJIKhOAscL2l0r4y2s0w9OQvbj/u8U1Tdb+eS8e6tOsOdnWDIZT+q9klJ83
Grqvt+Y9qDoS40D6/gs2Y4Sns5Kk1zDE0RrpF/nnAil4vxiLNrstBA4Ol+jpQ0A9KJrfoumn8iGm
DfqI4wpNAmoKUlr3h9uYZFM79Zc4Kano/u06xnS8Rt2+7Vy7skzHNkCyyE4czfDfHAzuoEA9aSrx
hOfUpcGRc3BozH/w8hBSeUgDf4/lPV9KspQHz05r9XXNLoZ/4bx8k4+2+rv+kNcq5tJc5gW2+P5S
TcCzdOQTOeMU8+JGUwm8mZcnidIeQ5kWy5kz+MENPBMPRisQHJPICX3qHlguzWJotsvx5hzub32s
6ROm3y0+gCWRSDDUqGz5vJc8OWFoq7NQH6GF2TgzIBktHWHk0OjpS/WJ4OXwjvNuDyzJZZ2+q38M
cXxTFuLhiTtTFH1Om0rTmu0opKziFztxXt39qqYXjxq4TMOVuCnYjUPL+jZyIcy1fjgqe4BbOEPp
0nTrM/wlq/irkTe4Z5//r+tpSZAjECDDJUcUP61APiq9CY9cZlGlxOvr9GRSAzFVbyPNxNr9UNS4
Cv0yjS2BvKjiLl5RUwIpUg1fmx/elypmbEJ6ovv9+buhqV+l7W9nZbgUmuBPbm4lXfQewoeaZY6B
x2kq2C5fpcyIr4cc4uSEasA+YFlnkRmRqi62gRf0oXGW8SnYIVL56yDQo+fZ7w2KEK4w0vH6mkX8
78CuDXTcMpRi7ymXacxXj1KPuZHvEtpVbNI4mojHXaKqYwhOr5juk64UM46mk0GlPVx+xSaczapK
euxnDyg+p2KDurW9dZ/r1jwG5N13gNT+uMSL46mZZtzJaAotuJLmPnqmmkY/bHEaK2QUtCas3I0m
reTafJCpI1HAh8eG3vYOyD5AAHl3Qaf+rihxV5/HIfvLGTCBuleuECbcIYieJO0Qu/pwTFg2CWjr
rr66rF47jbewKDKAfDZSEmShJq4476RbnGnpIWz57X4leERAgiHmgM//jU9FuULl5IF4OaLPKXVc
ZleQ5eEvdBqUqyMDb3fEBQn13Pvh5xk6WsuijVWprlolMYMCqaIPmYLAyDqn6nzYEsl/+O05EL3i
vHsZfZKu4RsWC9Mgo9UkQShK1ef1j2B+MzrfGml1tmIt9ywNIaH4ioRLsV95tCjEwDK7ZMG9bhSk
AB+yNM6TO9iufz6KlTbJiKYrsf3Y6OHEoZxgzyyMTWwi5uho2teMaHgel3YUZTW/+ZuWq2bCYx1X
h9qAD31B5abia/FOrleW+Cv4Xm02xz6W6j2ibnDTVTiNJSixc7Q0k93IFVDl5gS0HfMpaHlWp+rZ
1v7gBwtn4GH4jF1yy4t1ivvwVoDO2H315TWeD9LjojQbEn9a4QpqJBqQWX07cwQeUVkh33USD61f
6UnZuU0mLR6jOfBIxl1bB3PYLrp9cUIx1G1XAoqvyl9wrVEMfoKqSO4KaC6tJWbOCaODeUckQQbb
BI6NtBcSqTRZM9o4hFUtQ91dG257trsHtlw5GpOpFr5vr42vM1varuSK3bozsiimziERgowq3Cpz
X5kSyjt+3P8LEQC5ileWrqhOfAO25o9EcDOXTZ5NfQwbBMABJxZmjhnk7s5EQjzoHutNRV1x39OY
+14+Ny9NHP7360HEWL/VlO8AWt4N0iu0ymXCeaXGsy75aUC3HEGRCbEutOqVnPkX+bhbG9Iye94/
EPotf3m3km8E+0QJFOSp+194TuR46b0kj7bKN6oYtlNnQS1DgZhKwGNuGdgx/0Vq9Rynjrnhdc/O
Io7YMQImJ++rb1txBTOEfSJWAkzORuKrgIOmdoPtfkgoksMDiwkWg+RYdGXUKoNzL88lN4mLaHjQ
4uCCsxy+gX/p6THg6fToI0LeI0RLxozxZFOXOi1dhMO0qEOZEuUmg1EIIlXgKO7UeUTkD1BDBC5Y
iVt3GsP2mUsvfkmXZ3h/oQl/l6W204yGKfnClPrISYfGTkJAy/SumTZaiDU1dw2nFg/5sn5JZM6/
u4qvy/Sb8YdUbzPPpjJ2kYsh5b0ZWTjdl62QHmuABc5XhLqeb/REpXip9sFNPqpOH6CXqXXAimAF
/f3wo9Jb3VB7wB/FDc4OT30EVWTVy8eVmAW/S6cw553q3CeeKD0JWVHdttAhJfwEK3P8wmkESawJ
/aMz43R3AZOWk5Ublx06Bv4R6O6cOm9r7oZwnMKvfTNjwq5eubcIgS6JE+FgUElpnzQOaoHmu+y2
V9mgGlM1Uw7vJmAETMjKjxcTz6RDU3sD4vCKPcl8E60mvlXsDTkMxs5BK6acilSPiRIeJIPFeway
9pC0q0MpWa5Fz6eSaA0ISmDXmACEIG1Kb7ikJD3i8zOc+/0sKVYQteOy4WDj5hF87Yi58GLDsGxM
0bSG0QGrXs7s5pZA+TJT6+h+oOWBv59P8gki7pg99xMG6ibqMYuiHcnIYv3w2JlBKkHVEV9MYwQK
ERIRMgdGtv3IdZOdUir7eZTH3Sz65HF5HuegTQITvZqi4Ij9pCwmdEq9IWhJPyZYHlvT4YVD91e0
K0jZG/ri7YJriKZ60jwaTOBpt0ZJE1FQKQto/jRTbin4jLZKtA28MArofT49RGzf4tZcQ77zPDgj
+I3NuWc8ATJw/b7joz8CDId9oBdTSaUCYZSuine6jPz7kN9Vkgwv0YBRs5NrkhrekJyG/3d8SgpX
lDeJjwF10TnM4I+70PbdcO2QwpazmBNQZCZGOvsvrPCHda751j1f7jFvleGbxMrq7gYqgNOCE0ul
dpidax6u4UXbWfu140hpyEs5BtQ/2XoB17ekju8bY27gxAUEyQnmAriamCKI5HKFSSfKNxSVrhdm
FLPL3zSl4Gm8ncuN0Mgc62xqF5SVd6f2PSuyEsTNE42CyEHxgYh5b9L9KQmMMl1Du2s5DHGI0bNI
f/dcKc7NedOO7lX+U6l3MjYFKZGrGRXkSheAHTSPgK53XJRnmHV6UCy9mwO5J5LVmvrMMqtZpodN
93neFUh0RFuPcZu2JfSek/Au65QpKIxWa5Ssy1Pu3U+qI3LITLto89dE5TK8qaOxL7LWZ+sf3TB3
0mti6Abyx/Vv1iAN2x577NH84S+sL4Fi9jh2visHazGHCIVAugdhEEaHge4ARF/yixAWMrRUnOKZ
NUQmLoE1I+NZB2QlHZWClvSC7DCOBdWR6faKZs4Ip0jBqcxc3YnaOVEdpCRiZi1hkXY1ZrORasV5
i6wsb8qAu+enR22iKhh9u7wor7NzFcxuepb7bhsd6JmSQQYHUle0ZUZC1+ypuMxpq39v90ViHlGS
qFrXmQei+VpBCozpEDsTUkp5Ox1WnNUe8Vj2c2TI3Bm5W01Qa3xqPJcOIGKO6vHSm/8oSsDiyfTu
7kKz8JMfT+k0t7rBzgw5/I9JFBnn5gZCL89QCLqzVqKk7MubPBJmhwcys41uAuCfXX1j2v2TpLcV
pEQ9v3DOu9GVC3eER3opAdKaPaGf+pYMIIQN4XZl7zPckcuVZzXA/gguyLBLLr9CibXCe7v94r0u
zd2mzU03h76z18Z7djdDEJxDK5mzG0WR7SlmmyJf7J7vRo1/i87ZbM9e7A2SVNPsYVK1ypm98/bY
d8QvWQ0HHABxIUCy5YSMLxW8nhmNgHjov1PvtcD8o24kOad5a0PVhui0yLEMhn8yw3anifiipR73
SVVhdRbVHFKdElZRD0PJit6AdvRQh60DXBLGkaTlOKi3PE/dODHz9K0GGW2cM+7nYkIYb9XFCH5n
hxxlOb9j7l8qV0YGTqokDL1u0N5l2bJxjD0/Gh+tayMRP1s2EFOZiNFw5cWIBikVFS472d7axkZ0
khglxxsuypYCg5LNjw3fiuy/mWu/FaDpllrv94GGxAFNrE7CpKqZXgj7svdKaQShJaPTs1jzlcPX
xlFWiPGx3+S+VEVk6at3stCxsivwTvq3v5DL0/BRfNaOO2CIjzY2yLfEKmTkfpLREf7D0gH10+9A
6nCaV44qQo9IM/ioUGNDu3kS8mAdpxf9LF+GGwXoj4zf+GbmWT5jDBWR7irbrt3RFZTagnzTZyMB
X2Y9razmX/G4F/ohC8wKm+A58/wCq6DxqUWtVjXQJAEDaVXfECvJQaMTXxtF6dyoSu6QUu2VSPom
G60uc/+u5sDMl/Am9N0AlnC9wMoytwdul6cicktA7og3opaew9edorw8ixVsh562anXfh4RrSJr5
VA/TXmNZx7gzKhVDT56FHRVq4gEYs3GbN0VSruUn51EvRF21YFlkTzDEHjs+yy0m5IJwWZOioQ/E
jK86FRdlipJ8MEjX+PBLzBC+FmA7b2KHdyZlbX4qVizSn+udEKRAJ7RsyLZ5yJBFpC1/b5bAdas/
cm3uSsdOXLeG0PBMJFTUyFbt/vF+TNt/q/Q2Xx+HPcj2/mbfBpCL1sioWq2fVmLde42Yc2ATddUb
KczZRlTuGJ1Jgz0v3eENWZ4Cdu1Jn5/qdz6310a2DDNlfa3lDT+SIy5WXDnA6IK6nNyKWEv58Ttm
1lQhOQEcJTGPLLFzyHzOCQJubR71lrImdq2HAAt3atUT16n8NBc7NBScPKrJlhPcxNWZ0ZJV5/Vn
hrfxXJLqdHsLzNZfuYSuEWNGW9K450uQ7ddGbnBsnebQYXVtUZSzWTHxn9TaogSxDA0PqgsbD6j5
kxAN2blM3GNkTHBwTO6VBoGBc14ShymcHOFCRZ/HhIkCKm7S0T15p+tPH/LpE4aFNZDRBckSundQ
DnjK8Oat8+nloHIBOcs8sgKsXIEXPes1FryUIu6l+5gOmkPvuM2qa7PvrIUGicwh5/CDy8Jsk0pH
bc6zwwgnmQ/zz/U1cYj5fQp6xS+cM+KlueyXlToWA2CW6wdzIul6kH1rMmHmMonry1bNfqxYMXKW
Xt9dJ7fvr3xWd8zdn88Di6NdPgZt9GbYpxDvIsQjyxHhaxeSzPnNoksnSBQ5mW12wvaEXaL5EHCB
TyOvOo6stjwiAB/AyBtEg2q1Pn7p2ss8FWH8FdUpGreYEzYgkk2uE4wvVpbfsMqCXRxFF2Hb3YIE
L6YHeit8EvaQMhdvwzwBz/m1br05iLvUD3usViPQPL7c8BEk53Xyv10fr3NW2GU3ugrbYd+LQg22
ZwMslSGg1lSx5hm9wzojAoKErbNAWMH2C3Krv8UmsPAWqMejwomNddv0C353v7OOdifFwFOL/hB7
2EmsXFNaEWqwQQ/gDCfLWNBl3014OUkbt6GOOe2eXQ44uhrSKPkbigbPgPKHzdBnoyaDmMZDgR1E
NfAGbQ9bTZ4W2B3nMDIQnZ2s7tUlrOu7DUlryKANOj3tVvJawQ0JiCDNubA2iArHQiIrL0cV8MEH
/PWZBjDoqifWgIAxywXKNU+AxWxIP+X5vlo8npttbI0fi/5j38Di6HZ9KECmSmZpjU7UD/1jYLfl
pv6eeeCcZqOvNZLLwUpvlrNzcNrRrtoOjeaipKFgX7aJOVi+3zwZcUQdFCnG09zxLHMqwxDMkZok
neAVbXXPNnuGDRB1I2MJArf40A0hwZvJHtXcAUE3exju02LRVO/XQr7NmQN+6eojdtUPJ+n8b5D2
Jijr8YkenKFOi4w6jQ59G9OUl7B6M2p18sKwSFh1eHAvNHqxgjo8JnYkKlYjsNK3iJTjlruU89qp
1/CAsOz5DCJpK2ixzAO82MlEw0tsdRXuhlyfz4WZztNR5qrB9LPhJTn2HlTF+k2P00PiokfAd5JI
Mrx5FSamhE8poxgOx1+3VTEKYTjxDda9vGa92GBTi+uuofs8RtNR8oOEx72yET0bGBftMfpoqnl6
8okACLYMCMy97y5Ntc+GdiE6kHXrQGYG95z2CJ8PMZVeo0JGjzq68CNA04IRKyf13/puYIhm2zTb
0R5pbFGeJS1NPtjz0qTPdMV3AgyFjd265UGE5Km0bOSbgKDfW9j9pP++0Aaz7sU7mTU1jy1N7Uk7
jFFRewod5F6jg0S4MmmujymkXowykdQEGkrYz1Gw8iepGwA0Z0adT4lzUnBwBf/6XMgzWRgVt5kP
4pWOeTDhDlwq7Gfdu7YjWk3vyUy5DElCUrcJ6zeuAw1+ZlIRF6f6IPOYZY8K0SfSg7Hl9M1hdoXZ
DFfjFsjxjOL3PuIhrLONta2MEMt2EmQs6Aw6bg0dwcQE0X3ogOePZfdw/JXCkY3YmjO/y2KAa7YF
/mawe4qpHgPFW+/z51p1taTJL5r9j8sqDd0gEslntPCfogeMvrKVLheldg4nKpvu+cmboN4B0zzx
1VNi7a8fYS1HG6ehNmoWaaj5M1uNOSXXBxTM+JC+rpzvEMda+cW4or7pcOpMrlvWSYGIdfa24bRX
9t/g761h5Oywez5hvv1DATAQwxFZXIP5xIIbk+VZCg1NZd0dEhlxGljNx8dMHaCvEOFYPsF1hN0H
4kdZ1iz54eWFu5jlk7lR8sOxdtmVgdnTQKzMKs1mCy9kOM/vtLwNreAJdpVZsxoFkZjxAQIHBR8C
NRW4tIQ93tayrD46m47iftXQHNb4bm+1KS2kibTnIAx4Q2FR4rY4QSUtNDHZGV1ImhVsTnvb2wdd
1zYOx+bTMW3FR/dya8hteP3bqp55lAAvrE+DrSxAy6kzxvEbT7desKOS+uGUq7C2/suylioj2kbh
0pwBXLRlY4VUAMh614RhWB78opAAbLkKiwepQxNsJGv4Qfm2aCVShWO8/Vp5ENZZw/tFtqyw9u5i
ykxs2UcrhTC7tigMat9EPW1D0EkIq8USl+5e9WtDZly3ZYMJnm1w0Q2mEj7Lvfczjpnw6qUYa4aD
q34ot0TAgdD0Aabq9H2WR+1fGceICUy/jk0cXnmPtPFELB60184Q4agIn8InvtxfqO2mfY2XC57e
6HYsxixUWvXP9aH7ylavweNAus35Hv6hAxGBgFw9QOPnhEOqgqTnB8Y0jPd2Xq9GXmNdVUNnwTON
b0fW8s00dawYrXPg7I6hl2t33YPgj0YTWoEdMiWkt8CU45rdsQ/KGN2Hkb8t55L8iNJPgyZ9ofeq
JPRNmcOmNm0exlKu92fFv7Z7KmUSjOmx4y7rTDhIKbvCDLcS17ydYuewzQ+N3Ya7hrUwUX61TS0j
s01hao1/obwmAfdKLS51xSAbxYZQvQ6/pfJKcTHB46f3b7epipYJJGbcI4U7ScTk2/UClWZB8VNp
/0gokp5BcwrxEISWzmTRoIGy/PoDEoEIfppMNft1oYwA+xHeMn/h7xF+WgSJ8w9Nueoz4YEi6igT
FecKVCfIRhaYSdQWJYmCdEVsxllHkJ9ywC/ubR6FiCthho6iaj1kmtD7DpH8sTO0/P9cv5x49/eL
gvVbiwGnMXOSbKO/gK7wxB7ryGPSZZgtI4Jgh6QgmrR7tuBHioMSD13vhO4XRDH1fbaVNV93HDE+
wtmqaFpmWG6OjptuIPfdJXAhw1AsTYp8rxvZhJ3txRpqrchSV3gUqcZ1bGgxAm1Tl3BvlsQnZrRg
cPB3zvAoYnwifqxSCLyueZ6LYJsu1BIUsYD0PlNleh9v17lv3ymrSFlo2n+hVBXsrHTfaZi/i6e4
vBkmtbhSRoXW+bseJK3LcJXrtc2QP+Qv10h/cCOlXd6V48rxsFZnYlXya/nikt4REWJNRPGat9hL
/E3flyC1KXruHN5W5bpdD63E+TWDl1jglkh4v9IQ3OVVRl21V1N7vl60kR9DreMSLJrq10p6KZRN
9Lgm3eOJc4obXGrVy1V4N8WI2MhmxWHdN6hi6OWvQIQMo7okDlELekfMFpkdf8LsnQuarkGqOnLO
cUddZEendcWcJCGXlXbPNAVpIlrU5YUK7r+ht234+Ft68PmWCpZcKXB8Upze72vm6yGmPZsmcwTv
JWrEQ1AixNjHchemPS0TxEKBzw3AS8K9jREp+RMju+oH7d7rcfkaN1/npBqqa0cMNPrLek0YtFgq
Z0mWEAyWS/jSYdurFE0RqZGpweNLg5pEjpL18na8wD96hCW4zum88B8AZLl1SBlsFM6AlVj+5Pa5
xinUWK4ZhBJzMFK8s3egCEZesn0fzoCqbWHEb/HdjsuDquCDr9cWahJkq5HTK+sTdT+nx1C49vqm
gJmknmAGXH7+3jbGzCJj++X2U4hF7LNEprQLEzEtkNfw0MMXImimtmR3wNH+yJtVZAQKEPDMZmz0
ZAJnQJzq+gflcreV22C0f0Z40xvsLtCE+Cv/YTz+0zw5zoFVvDqavxtKZYmNZqTK4iwkznLfTVit
SeXXktxV6SSQlBKdZfXWoMV3ehhc/Xyr2hBSk3KfXU/SqZdrMI9mkbXKjm2b3gz4baBkzW8mg5ZT
qeSRajx7maWUGAVV6f+ZpATW0hzjtDUnqJam28/e3rqzgvsAxg5Lw5Ugg3febqkkaCinRrVeRLvS
deBKNNncW0HOVW0EH90nVk4mNqc8z7bll2fsvsd0DZURykw8plHA3cDIe2deDKvKcNCsrs+VliNl
jp3xZQyB449SkONc7BsVUeqx+C3Y0GdyXMHWPcci+MRcl/x5b2ECTx85Ha61MmX2WKdB5roKipGO
bUtvAZoeRct9e6hpFylSMcnWaozBe+2QiPTxjVpWIVyEM0V3dbTqJ8GtdtEtzv7k3bnewuaisoxg
Efhg+MpcH5X6qVatRL6HZzi4a3SjYX2E1/rj4UUr3vZWQt4GPUt/DbCFEqe1I04tBiQIyyB47p7H
nVw9iYD44s5sp33OhTQIzCDItgjkMJS1W4mX2ayRh5ia8+/2XjctGX96c1HLbQxMP7sj394GfCIa
+m0gXhU5x2Bqx368r+BZoEFj8//8iXFVe0GVDesIEUud3RZ7++D5oOGWk6uuC5nWX87MB9JRNBIF
9WMEZmaiBI4NWkOBvi9xtt6SHbN0knIJqjM6jInwHUiAYbgaF7iG3cQ+YrQTE3NraRP+G4VeKBdq
/RGBe/BRbxgsA3wvZmR7eKdApJ3+bLzBzF8HlKmJuWdiqf7jG0A04lYDzeN2u2pEmRe0NzQfw3+/
rH5tCsvQ5KvPPJWkz23kEV+0ZZUuiwt90bTa1i3hVfxebOlcAR6za5oMtea3ktU7JDHF88r5xe/v
xQ+bcYQYWRS1qNiNlsbVN3iPAjpdLX5326DWLK5S5HE918G7nk1JHU85Q2x8exmxF/muzi+hPT8g
QGDENKur75T4S4qqpwmYDsSO8JLVu9h9KC6fRrP2hvGukjb9md1LpwxHkVW2FQ7XwGPJhvuE7P8t
PvWD7Ieu0JZZaJNYxin2SiCjpjre5t1yTnWWVlPSDwD7aUlW5x23HPQcIlHHxBlapDfmKeIHwbeV
Sw1m+B9d9xv44Oe+F895Fvw1t0Qs29hng+rLLX4CZscnPbFcqNEzILNNLc0Bk/FFB7htuZf2qO2j
TPrrw2iDhy+moocS6CvRXRD+zenYxlRl0bOiDP5GgqxySYfd1e6rrFQfCT4Syhu0DRSS0eTZRSr+
hUFxR1ZXu46amIT/IbE0PWjquZ6NtwmxlrigsMc1waercrmx46bd9QINeDb6rFYwiEBfgdZ727MO
+Gw0xWcozVKKuSWeSr9vtLfwl2J8pjdhXhzVMwQonJolelmB1Uide/dEgEiyzUibmm2N096B5c4k
Ao3vaNAzrwhkV2o34/620l8mUcs0vi4Bm87UkSPoGHD2jEpaszYIcfjF46BvxnMP/vkhek6AYuni
tO51Bv2dmxiMf0cEytvHQ0YxzGIdJwVMS1ka/X/z+tD5qqJJyI4zw5jcbuWd7nUPXpdZDqtA6BfP
ottU0+kh581YLr/HduFVKYnIOI2JLtSonrAXGnM27Zzs1Jj64Mlg2TqR0nPtqQ54t+Q4EYcj+3oX
F/CU4qwD9ngQiDKA7bckEsA67MPW2NQDLY6rcYHVI0uRppCLgkPP7ZJKP/jXrZ71aHr0j17ovqzV
0XuYgE5H8SM/MuK212STs1ow61s1d65LmbPJlxRSBS+qKQFn8IZ5MpaXviq/Megb4VG2eq9llBNl
YbJtzD9d8iTA1w555hSgpzxUEnxIN/aq428VEohaDS/GGW2ZgeJv1HaeIIQLJmeNINh0a7DzsC1A
Vc8KjGSVoZ7vLxTCG5MN3nyTrIwMKkKw+HaWFjAivoYo+SEgH/KDMrAqQuSh5Y7IGWYG9O8IS9hY
IB9F3MWJWY49WdD7VsnJPEsv15+0++LWBSvkgHM8fk4JT4Uu36Or23bfm2y5H07jRcraLc9h7u1z
ZMZVtGQLaKjM8W7jHQCP3XNFA+qX7RnqswVY/eW0qtzDmEsAfdN8AFIguLW/qiP1RXyfPQ0E7ssQ
kTdp+d05BIdGukmY591OKQCRTbSpOnqvfdbZNWM4dqRVNLElOKjopKeXEsHWXJRSFN1MZE2w8XCq
O43NKxj/T7E04IYbiHnf64r8/LLIKX12jryN30BqDZ9nZGnQyc/IpG2wk4B0LrzkbEWCdTxf3yrx
0IHS/VaWhs7mYDyt33fmXcAUYWUxwzZfbkw9XVGV6wtG4unAizzbAcuytu6EGvUVK8I3GPfgk055
kSJfKR0bnA+8k+9IYr/aYLiQY3wHTFc50v5OVpfdS/H0PW2rtCCC+0u03M8QLKjVhCuVpAdqKcbP
YLydhwKIFyn5i9KxBxt90VddIKNoQkNQ746IqmMSfC/UrXSGQ6DpcjgsZI/E1qHdv+On35DArI+7
oDPMF0uhbpf0qozs2hYM74qrROSilX80tA7D1v7QV2+qIhvPAJtkBU4kpiLsDcIKs2cRFam+SZY9
mMPQ9A3RoWxZ+vA6vsn4gL38MN8TW4zVuaB2fathK5u9hRk0+CBTPf/Ni3cZisydZgqLhFimgVzk
AkdnKiijABxL9TGpyoHl9++lPuGLuxDqElvCmqRAefH8vhfu6P1xOYiELNrJAno+hTsEUlKZAAXz
8fQlZPenTlgHnBERyTJfnynWYZePByeGotAeloXm544YR54LheRQoA5KUlnt106GCcO75kuFIlbx
0KngO71hMHgYizt0QLtqL0BAXd6rorIbboR35YRjSVLiWKSE1yRMTpjA33UKOHNdM9vFFwiurod7
97HWWl2sTvvpZtXs5KCX2lnLGzfi8V4Zg8yQZAi9cAUxwppPYtVWp0Gxq7NzpNPYqC/FzZuZ/uxH
MYlasE2aNZZPPKMlCZEwU49oyxUhUWnZnVdngq5K3wqX66xyMr8g4P0XxD8JjfOLAhUHQ8xwlY3V
4Yhp7B5q4/irJvsqjbMpWGL8cKBgJwF56j+Nyq6AE4S9AyYG6n2a5+AiVeK8wOazBJwpEuGU50Ab
e8JH2DHcp2HfrnQVdm6G2zZpn8VA5O5zs7Kqwc9v0O4L4hmQwZOF/S7O2e54cB6CPw5bv8PChgcp
SejkI4bBaFjJYx777InwoyXkf4kULGjaOZ+U2uj7QQjHVHX2zn7m0T/1++m9tpZce6cze1Jr137C
rsoFsruPyoRgtU2lzOr3lIILyCdZmaO8yQ6pjiuYJDMTMjaEzBSThJ6XKRIdHdZgYYgTTAc2WLAY
yUrWdTBb4bEtl5Ja4v82fO2xpuVasxPTX5C4zuS+qejH5ahkCbVHsEYIlpZbdG6UWAjcaZH3ckfi
EIN71rdbot7E1lO5m4YCtTm+2dNG5SnZR23Dn/sdXCdwQE8iI+8FAdge9Sl2M7SkevnUS3tTdrID
na9jdvsXZs4D0WBbxvt1MvH9dK2gCxbUpDwhWXDtUKtLT4hlm/1hf5vmVJ49SbTCVovLUm769CxI
QZIUulorHBotBl9+galCLZjYloXo6ODxq6Vh7YXBYrXFi/cd/UYviJ6rNXTOkyjDUOROe43GmZH2
SA8XFmKo6oN969snO6DlYpj5TSI+qjoNL6X+2Q6BSnqpKb7d1wlNHNpS4adg47VK8ZU4I3MkfkuE
NO8vNBG0ujo0kyyCSNnmg3vB/VSENDpW4UtlGzsgy4XLkg6noqxLg8kfoVt79tGVAM73+Dkzunno
8PmCKYQweaaRREEW2Orgk0RPiMxDhR4ada/0Ytlfu07yejDfgdPUHGdbh0pr1zTCbbZtCoFiojlL
2rbnutPdTXuNr/g5pTDuAL5aXKB+33yd/iagSyWndC0pkd1h0x9/4UTS+1FoLdzdxDjpZO9uO/IM
NQsMFLDsLnewSVtPKx1jhkmsLXuSBTsQUuHwYf6t87tEpmmsdLrvgaGU2IynC6Y90ryNvONz+6NS
D3hN6TzSpHQ2GRunuNMYQBzfK2zk70rXHFaI14YzEGip5UPRrt0kHYkQGKC+hw7hQvnnCvOgz1yt
8SZ6trkfSfrcMAhX+YWkB/0BWDY8uRETFiaSHgMJ9GLWfByaoq7pFh14aavWIoWxaORl2CmeKxJp
oGynxmaQeXqZiL2GIx0HtYIIzMAJagLKwHeTEOXMKV7EXEADIXTb2PG2xZ3IFHLnUIApF4iTeq7X
UCcGEMNL8pPoTx3c0stB5fF0Jhl4vUdTevThBp/Jut99W//bm+pvyewal12aQKPZ50YjfQ/fI+G0
M6eU0MWwd2C4m21JGdv+y+Lp9E+YdKLI+shvVGL8XsF0jDfGmh9+2m/AXHU0cJ55bqSR+u069LWk
f+qDEwdZ628/3eVNFE1BL8OPZiQCqQYS3YKpHWiV9yAoBubZKlFsmHHWOfOpO+DwL/cbCbQoq8jH
U9+KF1hIergcZFwYPJW957G1WwvknPc9TKie5Sd58rF1TY4KumC8jArOPY4xQRNKKmk8Dh6gsgDe
HjncjpT1w986tMWfTZawJ4VV0mf3yakEG/WH9j8yvO6V59vGPo9PgtqGQc9YczLY1Uja8kTdnlUK
ROG7YGqFlq+NHQL5GIJABOwOpPGPMMOdybTBxyO+FmZqKVep8O/1n2WCcen3NB7zyUW6dEa1HkWZ
Dbm9sXEzchYUGgzqSOMmm8/P5GQ34W1Kz5OEYkNNul2sLV7VO65bN56YIbMKUWH/sgDpFtgEyOvH
hs8pQUWJZtpx1RLxYHXrqf5gF74ec2O2uTkdOIKwrjD1GW4fDSx4trAwKR3w+g3s6io8Ia48Mfn6
6I8PrGg05U7leu/S5Gq/3irid3BGmE4v3ftFx4qpSUfALSpvzDwFeHYtg95fm5C8KdBRwVGHRHWF
lF1FYuHED9QVRuqONbOzew5bGYQFXB2+ZldyWJsbrNXMX4doqs+esLSakVBDGKyOvhJCuKAI10+j
1it53uxB9JTaB+vH5YtPBOzIL/Aqz6aFFQcuA/hwesyqJB3ipnGly5RahM7YX63TV7px52CYmHJI
6ZXhX7DR8ZvF9Ufyu/PqaaDBqQK1LrUBCztsasjLtt7qjWCqnuQsz2rK+51LBKiDkH7u8dl9ykrc
pChB5U/LgZ35zbWtI97sq18+CECPZxPqpkeWDlfDUsrTKxdcPm/DYPikw9LATN9Pm3lX6jnDn5Qa
vD9YNcxZcLtTDR5qEflfvX9RJCLjSS17Uda+h5GT9TZIeExkDWsAH1Nw3IOfgi1sU8ZIrhMwnUnt
XzZyTrDw9r9pZU3mmAN2Q8P4M0nv2u0ZWkX8kuQyAa0BMCB2PNzTscu76ChtcS6IpN2r/nVe8B1t
5vWThNGZI+6t6LnXuirg+szMmCfcv6RNRRSka8abJsv5mrSZd1AD6vEdlpVH37K9k0HjhlcT5HYh
mqGOvjkqvuTzqeJbP93UZcnDOjDxUL8s7fr59LFpCSh7FxpM68mjIO/z0q+Y7qU8IiYnaAVYGHUT
jlllGEMJjrL/Ke9sQfWElMhxMscRVP+IzkY6CoLCSCsXrnjvoZhz6cEzqLWsyOKYMMOCgtL4aYXL
D5WVyHLuislXb5/ZhnnAIkzQePHQL7oiYxWSQkhkkKfnLeR5h25IoCEJsHVzf4RtMCRy7k4UOV8I
mbc6OToqU6AVfbqyeD8ohBpq2L8X+hhkWHtzQP6lLa7puTPMAKmpe6tPVUhCfPLveO8mrWM3eGRs
yMeHeQKWqFQk0XV+bXFOfeE424ewLSEB+/APBEDaOHCZH76pHqYa6nYhB7qviq9yoTrG3arYPwb5
6TvMDtvH6yejkrrCd3315DHsYqj4QW5FO6EEE6wKUVau9osPQIbiCFOXeN/+zO4G3l9SoWjNd6Bt
rwkuJAx5rKzr5XxaVmcz8pSSI9VM1n3MoHPzSMrbskNZo1GuRG3B+mPaYAVWmilCd3o69oNpLJ7u
2hKm+ub+d5wfGLj39kHEm7qEi6RCJpjCKhTua146m/eWCIrPkfTBEf5ltRHy11rwRRRsptaElB6h
3rovbMYf82Rl2oglm/9IHJFLr7juA56+Hupl0qd+YJhPX6+B+5xPmvb4fbtT1NaMDjYZZuXIf6Bq
sOd50LpgkUVSH+xsbm2YqJGbmZtsJxCLht8Vqlmhw5tkwnTOnWXFT2n9Kbjgu/K4PXvADtTarfzh
fmK/fILIwGj59Y8ufqIH3xy1cT5qesmKD24ihZxHULSTT9n7gUIXiCW5aewXgo/8qgYfCgYqp2YA
Dz7G5EEAPruzSFg+7mJJkMPRfc0nplnyxWRMc7Z1nbXQVgUoMWqyygyF45LAe/xHSzL/GKjT4QKh
5Ku0pCwRhcea8piKdJJ7diuCj+fzmPG3qsmsUfO/mdskmHnwd71H1ERWeySRPl11RN8C4Gn3hB9M
+e95M8fJ943FDLvCSTtKXTsNxKMMDEGG0GVoHAYw7vBTGahx82JsZQBfY2Nulu/ywpZhhdJLsrvl
s27OXb15RU1GcwyB+8QOLpK/P4LS1x59hjKPu92vsFg/HwHDd2c61kwkgHenmmBp4INhDvshkl0m
BSV5vZboI6d3piDpikcyJQgSrqbzianvQrzT9ME/6QFMmkRLsKPyVtOn5HwYH77EUl0ovqY95chr
MfNP7qZUnhLuPkoju4hjIhsU7KK/9zjRbXJNhsqSvWP6hbuvY8RmXVCO7hsnNRl5C6LtsEhftaI3
zIY35DPPcPFwrf0bD2/84X7a9dXS3fpWYVqR5/xT4gzPTOpO8c7GECT876eVxm9sbTLhn8WDsEKo
twoI8QBHYIdVEbB1hlagcXCvkIu/F9U9LT2yzrLvmgamAorG7o52VxVapZm09CtpaKpeXmsXd60O
VTDYYEMrP0+mTL7RHlGJ+YRp7fNh7NIibpgo3EusPo/RsgrHwprGKi/h6+rSS3FtW0r4j7W4MHgP
3i6g/mA6dpquXVk1RF2glNoJ1L02bgALkrn+BFx+vCkDQ4h9anDllyOsbRRsbgW+Ht24ZlVjkok/
lIViZKtlulFAIhmYGNRs5n9iCKUjMjDAoeMHs8GxUYfL8TOKkckf16CJ0sd4DnOwaMJE391oBvho
p0eIdxH2FwjI608NwKLyxNFrtAf+3U1nlde060V+boJJx8rYi9k1NZFjjML6yzOyMJZIfa2cGzYg
SWJsXYapC7Vrcw1livvZlTUnW5Oyno9neFIDcM6YwRqyWr8yJXzsD89EqPMXvaK3qipyJDjxIxyr
6rxQWAUR2Tnc/AuceZ8HUnN61A3PkjkJoxFM1JsjWPTQrPyjrOxZCnLhxM97B2j7tVBLXcQWMHYg
8X86pCzdEw2bJANin9DkcCcdx0LSfrwQ4zgudnwGz23d/0kYPZe2ZDTXKRr/vMgbxzKjLjjbn8nW
rIE3W90aCQBq8P7DX7KDCGlsd2Ie4lrBzUxbm/j4LG9Y8yLcBn+d/ww9lBih77MJO8XtCAjt6Umq
gNkofZLKAIu8ue+Ui5Bu4tHlQ2q1EOZ+jnJB/cBRsNS+YbQKNr2SdCz1AAH/o3gm59OOPtOkgiI5
UwCicrOtOhyeny7qN/YP9AK2TgFIohzuyQd74s0jNcxDLxMKxKUupOiiJMR0n9+L2ylHk+FhW0J8
jXy3s6+pRV978kc2ERkZHJNYMXIBkoz0iYoz7cAbSWSKUGhnJ/TyP+eNCmvT1hS7448N38iKQKfY
ATVWKcWsvMSnDh0J3XAqzbrny3PwMSUP/PrgGM6UergAibQVJWYRC+w+2jSsbAAHx75/fRUPKAIJ
2OADpL+wiZtfCeZre7mKDm0EQGP4BQfoNYafht203dciDc0XyDF4tqhK0FizpDYXgLOUeBsBz3iw
CurBpELFzJeWTBFKGbur3vYtu7xr0r/q0u9Q8dsdNkQgesV1xKVrmocRrXzFmbKLvkGTrCHCHg0B
dYW2n9wdLIffBjPK77oFb/N7sD7hzDTPUKYTW0havWLjeKYJWadfzBYRiZklNh0+IKf9y9ko0iKd
IsawlvEXQjNJBDQ2niqHw6Ova3XveVwCnYitG/O/YkBn9obRyvCKtH1JhJHmmQI9gp7x0RrUk20m
RRlDEvtRPIB9EKzRa8KyL+xmDx/aWLoSXngjOQ50m+y8dWoFFcxh2uuT1DM/9fJxtAxcpfrgDF5A
LqEyxpqikQnqcFzyGRaaFNGklbjYTmHkpHD3eVSqopfiagRiwOaX3UZIhiBf7U4Ja2xLY1adQyyu
kobeUAENq1ZDeuYOZN5bQQMpXBbYxvDTm/tb/Xn1si+AQLd//whAVoNyvA5CgAixYSEzxOB9wG2h
ZxKD9fLJUodne/7HTiEHvrdmB8B/tDY2GQ7B5oEieWAHeicMMuHQ76sfcFirJVVfoqhwma6uv3GO
kNC8zZj1Q/PPfp4hwby/Ce//EB6i5sHYhiD8a5AkTcUQe9t6tsUppTdOvcoML0cHF6YFLzasbTnP
tQO6bhYiQ0y3EdLLdTTR7jnSSRWxnaA0bGeM1nOBW1EQ2Wc/esC6FzY0mEhN2xeSb1FkrLGHrS2R
SiErLb0TBaZbRGlFZhE/8TG9exch1cUQL+p1LTpX2I/Z3w3xDobRx3datJ/AugI5C0IoAeepHI6n
S0+Bkd/ne310mQlZgntap8A2A/cVWcljqqALNlzUznV7h9cR0F2YUcHfvO8gYXoJWxCAjZuLePUm
I0jt4koIHp/nSIrAqOZTdiKCjYHfMXDf1NXOpSsJJSRS3IIf+1DCLvBT70Rdbc0c5TVPEWQPxDWv
8WOggnkg7VoExLraSslB+mtDct0dpEtOBZ8HLcT+LepBx+LxQcGTh5jMwKwFC8cXPj236Ok7G/bP
GHW1D79mRXylGswvz6UQWZYqIVmYnZ1eAgprfJ5cGFM4yYAx8bNhhLinf+oJ7QYDwLMSGK3aZAg7
RTrh/54D++ctm+Cz5RZzCK4n/Xzh7Gb6qYlLeIF9TjPqE/zt9n6vEd74ZURV/8WcWvE2Z8qyPxPU
zm5pXwx8P4EePgBrhEpt+LXSqTCY4sVT0RoVoQAj9WGkZPwjP4GEHBGqqAyZIwH+re8L7I9wFSuH
/SKy78gjg2XtRIub1xl4NMgFcobbuwlNomhGI/0OiPiXzKH2WqSaGYPNxbdBAACKaOZ0H/ebK6ve
Z7gVXIQTaEolX1wV1DNce5r6hM+96nwqgUqOK20fiYGTtSshQdINQn4WqWJ30E+fCZdFRf8u2wf5
7fwLHS0SURtk5X4dAEDZAEgcIOvCr1twXybpCk949kJdkUuR7yG0gaxZZbTDUi2bRdWZNDaz4Cze
yyMcD42pbtXX3pSo8vpaYbmqvNYNRC9JXJhpaH5UiZoJ+KU0/1HxGhpv8ttY9P2rMJ+vfCF5gI+f
kRqI5Bkay9b0NA365PZb51pp6z8/s3upyfI5WdpsJ6+RH59C/cOm/BK1CEAW/uCfmcjcGkUlJUFH
yg7f5wklKDkzfR9Tm/B2Fa4egosRd8AY5ft7BwZDhlrcSV4CMHR1BPBQPRrnY7RLVnrpWUtY9A0r
sjYgEEE3Ko7jLK12l5Me4tO6Mpg2Ndh1r7ZoOj7Qb76dBk1C+FNObs2oTOZTI1JDRtoTvvPfABqL
qHIfXf7OSqsqlxzpStwCZf/HIzURGTnwSFeHUKGEj4LKBKho4O3o3v3ck60KYA9eA0boBiX2zL+7
GJNsDNfGXg/BENR38JANLhreEF8bvS+xqQQevq1/8NAe+EGvUvZzkuVtZmuT0Tjphimg+uBkypml
pUG5DlasmcBFfC3Z/ZS60NU+oeb2lOy9AopfHiKsSNuqS6JPYrmEOZbT44SUU/GZaJUyaG0b9TMf
mvEvScv9oZCRK9uIJuGPLIFw3cRf55EpEdrGKtX74EAhPmdYVK7NfD2da0mdqYHkgJ8b6L1aqw1+
XRwPbxtYA61nfeo5wbW+ZR3IzbwBYMfUxtGdJ/u0HktPbCFQg/3Geq0xWctCg+UCAjygn9nPzJ3j
Y3viftOVjIFbsBp0G02oCFfvmV63xoE3sfWivTnSEu/FkrPVc8Y2sZyPl9XHgg3CgF0pjZdl9Ii+
8B0jvclNnxljbbfNnUdEtaVxwe3wb6uezFvzpok1DgLE/nq6DbMbKl29M/AzFkqn9lud83NkD1fJ
0mcFrm+c/L6wkcBTLRuWivSbrKYgnaRln6X1o0KK1dMKfwqIjTglZ8zsqJY75PongjRUHcRkqY3H
7jr7yZ56LFmIGLXJfx64DVsxrZ6bjD3RZVKUBPK7qPUs4sG+Kfwt2Ou4YBg+T9vVCNbyHO5aS6Mu
iDdyM9LAU6R24YK8ODyXBKX3+KGOkoIyf1i2pn4IlhKdWm1pHOxqe76GA7VN0blUcwltVSLuDgP2
TgExEqirnFIZJaydFbntJkeu+SjJX1FZkCQ2+qDac65fSddmL9Gumaf4D0o/acDIKej+Z5eggWBl
xBMHBJ/YBeacTyrXBmC1s9FLeM5mgfv8YqFC02sGJA6ZBTi5iwSP2xjZrCnMCjg0eo1uEl2B59XH
Qpjn/lLDrL9BzOd2W5p9fXy225o/f24dg+flnruPK7AYVc7NhXp4bviBdHc99k0+hFQZQEpI5Jvk
rnBb150Zs96Jak3zwc0LvSn05eEZGPL7wRFnWMXotvYI2FGyXrD6osNMRGi7U/0HxHERpa9XOLla
RFwmDRcu8HsmA/ZYtm6nmxN623kRbw8xQ7vOG7U/YV+tQLW1X8PC2HHEOxTsofs2bc/3SUm8wZKY
YwoVDiY+QhTJKWZnro2eCjEfwQWUqmv1BidDsOKNed7WJZECr4JxK3XwdOiGDloLwL5vdRxyW9fr
VobryHdSln9vdqFWdlPzTcCK3IRbfigtBKqGh46SeUxi6mnIN86ZYLkNvHTbE370kJl5fhDZB3fe
QHRRgC6ZwprxQhcYNeeIdKSdWnZWLnwOw/ykLne1cfQZKXNd+Ek9PebmW2mlJzfSNq/ia6HwfV31
T0siYzerIH9KKktMUEweF30ZDPv+FHg5E43M4L3i70tu1ei3RePOCQek3zDn7U87VhNltKddYPBv
yUZMk1Isk4Z91zMbtEDRxTctdqmREnjKmRRLLcg8Cew+A+RNPbh5CJJfZuFW8zlXS4AnEKs28I3X
0T6vnSw02C237qiyzBXPSUVfFYuz669TTuRR3eTasY09jP3r/XGsXr8PxbVnaahIVa1I/XFnzdXu
NyzrL9jnpzQ/JwM0HeCLeEX2MWTvDRvHYXkZC4DpW1s0lDb6hhrkMyGurTuC8E2w8ZCehDPbCInh
LxotwRFgP8+oDrQNHBUhWwZPITD+BqTuEjkqySHCI7Ly9QwamRqgn/LTrkqUgKxIIU2UKWDIefEi
bsPZKlUow5P2FIMBnjiLr8siSQJoO/OnKIPrR2e2iqV60++ySjAqXyCEoHFhIeEEQ/ArRWr6vTET
PEWm6JW/WO5hLOntl6kJahrZ75H7UfQOO8ZdFxngCVg9ggjYJqciG9FSA9WAvm5spPd8AFbsIpET
w81ryrWElPBW654p59/PfotKg3CBjGlGiBl5D8YrOgN9eCoqdvc5mSZT15Hgx8wFo3dWpQeKenFO
KrSHlyHq3J55G7gRk4wKwlK4uiUaNFlYkpsAe+JToEz5cI9rfedLmm8Fkubsc+sq7BHOnVQMncHC
ss2P0THNIWJqtl+2AouSQqfBMvNSrIrkzXfFOr/xK4X24KQ1SfIbi3octrJyOzhj0/VONYDw73RR
Mkci4fQrQopj5JGBEk5FkS/YOGflnZNkOv/sFuGP/7/2mHb/F9Jmfs9a4NmAW/EAh2x9iFvjNfoo
P1AcNEFw64ZDOaKIupHPxXeIXoTMZ7pcJ7XzLydpnOVWBvy0IAUTJ+pP0jsgQk8HxlvZ90csQvjk
aJ52Hc+S45e9cWOAgRnZZH210cFVI3vPm+wpAZ93H2H4TuNY/NcUAxu2fs0onzGY7ddkJsFdpNjS
YatDT0BeFiMtLSs4uvAOMpMcjXe+maeFaHe617/u5FX0PLwqQmwIsa5vV4q3VskfyLD5JdyL+L7w
fSOmNd5reAfrrMB9GGs5VrvDUKM7twGFQuf+UcV3kberzasOiGs/JQSh0iuI7fhha+SERO9U0isV
rDXUi9qdwqmI+H9EEh81jOmWWjyEFwHySlPco8AkftpxH8TduV3ugpxTkrTe5xMaM5XAfP28PHx9
e0e7dKDAmlsutnF+ayND7Vw8IaQtNGXbgefRscw1ZoygQV75uXyeCNXOam3WJ20nlNIrcFLtFl3T
JvvMfsrZGu+KM/3WSZW35socPBYcbPl7fcvszvrdZNHZqUPrIb6aTNVjpaA2sQd3mvdM824p3Y2O
t2arGu7dPWp35/N1azJmcT8hRMxPutPzym1tRfJcsOtKdZVqj5sEdC8+fSvtw2Zcfz30bJc2tmtP
3gjM40MoRN/LBh+EwAmoC2Bu6oOyY4TWRh+11QrHI5k0YupzDkqG0Fhnoc1gvLpD3GYKKs7BwzSf
nvC20A1zAFmg9qqMrLoGbySPKJYQI2YeDfGGp3FSMlS3XB8UOGfqFG5yndwvDzYCQf34MKKSvc6j
/ixIv/d7RwBb8zyaOzwAYr3JkEX5WQmqiaz1xN2Ruab87VRrX3IHtcSGyry1zhAEeXbyx5AEHk+s
GlZtrprgQke430e8bYVggvKMf401P/acnBesnzgSVFbkftgyXQ7sKuNCyGaQlQdfEz12AkYp+TWR
5m+wOV6Veuav9k3CTI5ei5Q2o0qVMC4CCgJuZjqSCnQlCGWkeOsrJm+OafDH0tp9v+IYUrctqrLi
Ur3h/khikdoI+L/Vi+BkRNz2exIHDStRd4IaEQ5xjGtsfIUYSsYGiWjwNb6Gc1CowbLHmdEdOYJB
U9XngVyIQfl+GdjZBHsklQ8xXgEPIKNa+Tvk0zSwxDf/l5Pii09uiwmHCDnxNTSJoGQoFThRqtEX
ROpHt4vbANZ5Q0mhkRmgHrGwX1fdcFD2ouYJaiITRi57duEzO/Ri6CZpjnV/rlCATZs3QwpTBCfx
qv+Zwqg0A8wlpLiRzqLYJ1B+OL/yqOOtzmEHKmqxUK53+FpBEvl+q83WIfIiEP9uV/z+2rf6xQ/e
tcoeAAMFtmShSEhK2wezhnT5cTF8jfXQpHm0P8I7m/iCQOUGxYiq2KAEZeAm4BUewCTZ9lJnmXPm
qvg0D1ZHVMzGInCpdBmV0Q+msQRK6oqLRJ/90Rdh3dOCvD3yVSTK090HQUnqnDdELGyhZGbewvWX
+uayLM6f/LUimcg4shqOIKVvI220UPs/Cgf2zvNQZJAPCpKVSiAupKCyzT5Km7pvUgYAbzNuYXT8
UaTUGGs6eIgefhzNK41G93OK+AM6x2CFaPiInkRpWAx0SP9XRuMEV5gR2Q7dc0WxTFJG22oH2KAr
kvq9fZbDlpYpa4mWHgWH5Z3TPP2UG6/SEL8ajaDZRhsPXeY+p/eaeIDcU2Hk6Niv/1bynBb0jzRt
Oij+wuvlskclwdy3uCKgaJqqryHJrvoSMVkYtPOTX90ZkJqR/tQXz6LP/JCZ2b3wBUf7l+/RbOBA
kTk72zM3PTx7bckMuLsRAukXVeNaGo33uBlTT0/amdqsj0lKg6XT5YNzYH6FsngOQyAtN7R1HMsn
wFApbcRAP42wm8wJEZAwh0foOMLaVC18gP7L2xN3j/HtAMDQhcyiFawvH70fhU84k2y9vYLMZeXI
HJyS936xYKUgaro0ieYt87TrBN8703d99Tm1IFKzjHpngXlINXJDQxm4OIGs4pdSOWMHddiGjBXu
G9HdfBUhLYOBPjHiPDuSiMoxou+X+XJ8LNFhJUzsGNpUErMevNm94KuOWu2NLGtD3J8hUEHTJOhe
qBTmBcLRidugt16/tmZn8O6FBBUhPLbovDFYmYQfP/s3a1mbcEfDC1KOyBTRT5laTvtVF6kLswVz
kqI5C+DeVtf2ORf3RC0Tc+dJvTQ4lOMRaI0Ik3721F0PSSxsHVDkCbkACoKfnwOZht/w8hFgwGNE
is4nIeXvHXpwTawsF6RIIEH0cxal0jTPsLMNK9akHb1ZipiBNowKsvqzYg1xR0iqsRQ85kd7ViFe
f8B20Yxl7Y6dvK+lBIKVD24/KJGn05qrIhRmyqW1GOX8Z1ad9OAMkXTscqUU5EgOj/VN/2zOBNiK
9Da2A32IUOZPEo4t9gzzIvrJp6cFQCTBswA5Jd4AgE9YNKeSocT2bpYaUtoXEVMRAO8hT1KXWcXh
vlLP6/RsEp2DG4V528tWkjPSWwat84vIKiEmpDR6pOZqBC9SEr9KlWmdvXN38L/lSEVbOiDET+bV
BxazaC0xasILq6fx/QPOknGxmWR2TSxdQWtp76qrlouZFnnkzroinpJ2sWO2X0T5LkqEjZ3VWO0V
eFOKlvg6uSK1Xmmsmm651Cu8lYiypuHXKJ4+oOXoem6mRxJAADyCieuFNhCfr1HzYy0VhV2STCOE
4v2Q/flFAVpNnSzmGXmRHKsTTAfSOkY3ML90rAW6K3AaEdvy5n4FG/cyxd9qzAplBi+3u02NPIgq
xUHkw7FgLxajBi4Bf3xf2DoT3/fDJLp+JBDEQF89onfsJCGlwHZuPSO85iv3AUPWYJadp0vYtxtO
D7KBlVbrdii/8POZ47yYzAzkSbNuyOrXFVSEH3K44gXyBYs3W05XSMJ8ewBj+Sdq9WeCMVkk5BSl
OBOVfCLdVyTug7bx7As7cCwX0ie06lBW+mIK2EwYGGWYVLJp6QMu9vBIWXs3JfY4eOwh4DxBo8RU
AKa4sxR+44RTgQ5QGeVQCmnQ1JWoHwVfoKkcHRg+Xe/Tz2IcE9BBziQBXj2cZM1Ib6dqjFkUJh+D
zRULzhfupsNeqxq+Q9UO7+mUsnvZUYTWdhVwuboxYXso45dRU94eReneV2aRwPkkc2t8Kh2jYZKq
0kNMxxzExj3CynHVGv1QiGJyV1A7yWxNe/BhrS7MkJYJ0rlt1XRwAx/8qInX3nZa1FIyQZJdWjZZ
K6iyueedRENMY+HI6F0RCU4cmFJ1JpH0cW0DEFz8Geknpk2PvrtYr6XYSje//9B1zD7PUY+AKfbi
NFE+HsWdDBblg0vV9NVv77gcw4Euu84IjUm0AwzuILdlktlAaXaXS9upM1E9uoAgR7K3OxCYtYfT
vIkIybrESriNtb8h3vBHDcHzp/qBuxZhd0OZ2sqi7gfGcxxjdN2oRJGpi14/NBGbusWSgosxg4uW
SMiiOPauUtZpBjByHVU2EGj+pnRmL7ng/5/iTOtQm9xrllPsZz7xuJl29amWHyPohYLf4uWz1u9T
VJxJ/Aya8R6plt1EqQKiyANkwd1VoTm+HX5DLFlg69qT66jCY2B5xUbDkPwX/k9cnsz/h1CEZ+4f
MH4Ofj6KP/PXfC5gpAM3nvsXCc1Au5IclNqgugTw8MSxyUMO6pk5wGJJfBIfHI02TUQ1b9+Sj2iD
DWVghCdmMZoBqFQaanpg7DgpKuRqUDUyPCjBThvZ2rel+UJ6Pm88PW33Wj+Gj/A52TijAeaK8tUt
8kqOMcGGEoAUQ8XOHoqy7rXmL3YBLvRdVlaHkPlglXjL0ZA2vGKT4oU5ig9GzdtfeqeNZ5zFH6kL
O9vCp7EZP17bSVuXVZs4NWDWBVS6YgsUncVm76tz77uIs0vZm5aoa1Wb6z4cDvicKmHag/qXF5kN
oQy26T6g4+/UT9iD2UbeXzoH+VrFFyPCsWAxeomaAapzxK7nvmc1qDKrOpPlb1iodnMiGxnFfvfB
lNuKCCmjmiimbFr4inqx2vg6LkK74sAfMTZBryD+K3AFWz+FNB5gvaWbwAcDMWB7jsHbiTgw2B2+
PJ0+EyvKxnVmY8r7FK2b6avMddB3t9TMpM/nWVGMvZAqZlbswEQEI+gYIdntXaTlTpRhtEJgI0oj
woLpFtIh+xV8M6BU1OurfUO8rit9q+tae1A9v1NiYGXLOQHULQGTd8TpYPPCYRYV5zXtbWYxMAfn
KwEjkI86FGkYznS58jnnauvQAAJhhO6dwwFmGPw/fVsGgw2bUPd44dvs4YPcBFmBAxqM2ZuemnST
GrGyLvCBRP2RiUpWM0SyvtIqL20MUJhBKcc1Jr/vspQ0xRJtNTEBk3m8rhrcPocJnlfZ8qcCGl22
yuLyxhTK/tTcoeHJeu2NPHPS3OyQOhBNd/ktAv5vLjSe69EQLsd3bFyPCzdF74iOBN5ChIVEARKl
IalLHUw7j2zvmV1dgwjTlKr/hW1lsL60hylI+Ao6qHp5SyZYN3h1rI3TYB2NguFA7ceHCgAQmuA6
Ar1f69BRjm3G63cM0OSN7yG4rz5n4ZnFk8HIA+8TU6sGvwsUsHR+y8TAHyPOestS2fJC0Y4dPzBY
uNTURZVgEHlPQ8ORRnIKvaBnhzYiFQ8HFD+hRPGCz0mGaOPU/FHgxhNPaT9DR4AMihycmK6NTpok
rIQfaXhDV1Nlv8i2sjrr8kXoNAJO8SXpOBYgiztlskjdbM3vzXBDz6FSpn1ior7rwM3Qd49kXqsO
BN8OsvjmQg40NRMfU6N+BQfVJJyMWuqfQSboeeUO2gxOkKWyvaOvxnWs/QbFmgHe22m0PKsgF8qj
Ilj+0IMMpkC3O98BMjGYtp/Xpcf7vTP6rURDd4Ey9lkX3GZECZBspXSWSCT8/eBd0e3vjyr3vuVD
Bz0PUzZq7xwR4wSRre8dh0Ydci81NJ+V39azQwKMoicpAD4PITR5Vug/sLj4bmVCSJ4HNYpPpOV+
PKNGaBLnQBoEFlqVLbMRE5M5o21/UFZer9+MBqItlvp92xtpeROYb07rOX6meXyEDizCxy660Oit
FEByrlhypOw7rxMStHJD1cgWGNE4PQ5Kdi1eeBtGOz7udTq2EEI45Eu9otMCYfWfhgVVGCb7f1nH
kgPx5S8gQ4Zbt4szkZE52G6bkK1/rt/IftbEdVeo7IzY3CMyngJVFXUYyympQpYnIxYOJ2K/90+z
muHDP7lxxfvmy/oS7psu2sDTSBLs/H2YA/tceV1W81FNzzX4zc9JbIqfO9ip1fJKrXFhJOUS6Tn1
7dcHUUlu9VOon8iT2VC67Au9c0JeTNX4scw7fpJsu8OStDj1wWI7LRdbW5aeCO+5UbWjceot4GR4
iJKW9N/ZCAYmi7IUY2/I9kYTp9dZfmMKO/VPJBFzd1a+Gwq29c91UMVQ7CFqptofwUeh0G7VHkMY
ZWvHQZcWpquxvisswFQdU/ySX1wZ1TeinREXY4nqnYpJ4XzKfFPgUKm2pZp/fARzXyuJf1f1D0We
oBu6yI2n7ruCTKFeNjiGLMe8lO3I5ftvZzCFITkIn2iF59cL/nYiJs3/IKi+LJrmJW3DyEbI+/uW
ZjuEBJqZ/jOypyAJqyN23dJtlg3PNNDrcLlcE5iyyI+hqdIt5ek0iIf4j6/RD942YOdjT3KLfLir
wgB9An4TUOCQIKzgXNhyQUDnIXKdpW6ijMNXWYMpxGR/P48zlQEZ6aSb/O61bgwxm8gMWDmVyfLD
l4YFxc32wNLAQwejaZJpqhHXtete+HXE0Md1AF3ISYpihFSrB6lLdCgCTKXds8BCX4IwKg90FO9b
kSiX62UCOi2YKNY8me7JhGXj/yURb5o2v0Ak2HXBMiNNQCOYv3+C1+KnCjEhvc22HGQfpB7EUKG8
gcwVq9E00Ud5uR0yY5p3u4TTWMc5nS9mDK3cvZeu+auOXdM+FGCfpJeUUIrZSWpKiIoiSfZLLdag
cYKjtM9OvRymXo2hD4uOd70s0P7IUykfLnD4KMt3CTvjiDuJz4ca9HybPX063zPh7NdP7LSOzoSb
n7denBL5hZSA+PQYEih+9fsNl71JXYcazddirXlVBvE3byJ+EN98IfG2cigpJ6QPLuobJeh/26J1
vSivHrK8xvuzwb9Hy0QpB4Y26CXdgsYt8ekPq6/snkUz/NchSjXY53pywyJnhd+yaC/n43BX+8aq
Mxovl70kyt1t+dz+rzzj7/YI/9P9/+iEv6GLg5FhaOXJf/cDaimeLm8WiHIkgZ//0V36V2U1cyqf
YgamZl76wXK70RPkM7vZm9p31xTCYZKhqzHpTkbv+G/dwxlzTaWxI6n0VGCg1Hqp/twhq59pL/6t
1QKnj5R58jdf2zArMDATVLz/PrFtoUxOdze2+48usD8BaXkeRGK+LF3I3lhoZY7VDskdwPwO7TNl
4OB4yMbbFVQRcUV/1vNUD4OoM6sF+wJLFg03L2397ygPRhiERJ+oKXCvlkJcjjyvpzC2CiqYPFW8
aTT0ZuprVQ6N4uhuooWHiLEpWGY9FxvZHzX5OMA07AfTMs6UMS54s6ici2fRsS789oopoyJmn2OP
AmrQG4zt6xRag2AT02/fUYR4HY8wz7doM43wkfvHaG+rBqyCZGoGDGETL9vriAnoz8Cnjl66CqvC
u83tq598tfUjkdnYPuBPxflhA2tzZXJvWy823ujaSUYBi4mfYTavIBIK/GEulp2f8yW1q37k1zZt
HLcy4M2CkjNnK4S/cbkxBdN1OkIT0KEfQdEvGy4VNs2Oohv2oBbXiqa4F4CHGVyFTaiepk3dDnRt
etLb6zik4ISmvF2odDGklskOZMJLqxCo80sgDrpwe0dXwj8zV2pnxUJpYFyFceOrjZOF3UjASH4F
CLG3wMY0zv9RzyWkqP4OUL6AxRphSasPz7QnymenZPfHhT94ttqV4pGDKFJt1ZgArzA9upEcf0+X
P6zEGARne0heqtoyhYBfIIVBQlmlji3OdwoartGqKbjjSe/Akng4TpGCGVfxq1dfs2wEesniN/kF
OJ7b24PYOcDBzO8lks+O02TxTVXfbehQpkH5GboMdRevCJOkJzCt2rs//bAaTrVQJfJNSzmT1HC7
qtjxe1CeQ9oJLtvop0waWKEz1dc3JaguZ/Zi+0o5kIK3rXmQGfNZo1dHcRF/bBlSDo3tls0rzV/s
YnJNVwse7vwClcNl/zqrWS/O3bZKnI9+XEII3h9zcg5D7tkxPMTnZzlHbuqoBppApLe7Zzo5NkNr
nAi68FNzq24rgmbbcN3LG49wRAcDzV8D+9y6NwLRSuE6G+Zx9Dy965w1fD2QhUpwZAbsYiPK9qan
9WurYVp1doZqOTMQXIf4RRkbdUoZTd5+tkuhjNmF2+DB6lEVCqQsVM6LfHvGgUGL9rKUkGR7WO4v
dkDtrpgs+LamA7Ov96YRq78qAmUx9KvNNEOXYalsrhsRIXGVkwCDoI2J5yHa/nnMI5SkuPY22w2b
u7JdXWbKsCgE9EUiqkOu9eSihufLszgMzq0/J70dRGLKYxhNOrLnPB2plP8HwtR17kmtWV5xl781
fH6auY5HI6UinQpAy0afaMNvSSy3Qugtmqph1pfG6jAukB5oluanSQ/FsLVuXZ3k8uebH3sm+9S6
yGFSF1BAT3A54Gn5p2dt6M47m7wtops0sg8LwJqUTj932RFJ7t7xRpxCKPvF8trB4L7LHGa86HJD
hjib3z0/dHcyo5YldYCk5E3Ljh8jEx1zt4itiSQNSTh14hqC1kPBlfTrCBTrXz/rg2ar/t9dzkuE
7c7/NLN5Og+cdldXDaywtLKZvYbO4IzBYq7smp39FonK8/YJHFUC6o8oAZSbFz6zDOelo0BD1nIC
YGoRTUrSOLrLBMOVIW7+lPKI3MbVSDQjsy45N9OaO/NYpArlDOuAPxK8uWS41cr3jmJdNirE1PtM
t+ds26PLvDyaEJL2FjK/K5JkEby3GX8Sg560jhCbRDNKrVOxgLPzBhdEYqwnj/mNGpgfsk1YHYDY
u32xLRdVA3K763SoSPHrBZHEFfNrMp1eiAhcqcbBjNCYwlRsvV2fnO3ZAh6r/iu4GgjiT0F1eUj/
IqAMaM94ahtrlNR1GsOCh6WCpvbEphLsCxTz8RrsJj068tobrPFnjdYfFQTOTELDJT6aCS5YkM3u
nhbwR1daGy6a4r/jnIeaNmvmiLxlz/8gNTfYJjcDLygzKvhghlM4yncy9cNw5U4K/gcZom5Xk/AQ
GQYheyNn/GimVqnTxConD4ubNuNk9Nzzsu25PCb67+TjBwgRZulITHEVZ8BiQFitMvxykBRiFdGX
gmciVZRVk5A4h8EOx+ZWlqdE/aBTjk3LfU3x4J4KJ7Qlm4viJJHt92FLVHBmHvYUrVRXywu95b/1
q4ZLT1OJiNax+DdS0gWmwFIbSm1sNUjQwmJxt9eBC6zMVLwK4pGiMSjZNG1UXTvLmAybOUb9yozJ
cu2cqbvAxUfhxF7O8R2vVticqMDFmPLBii4g4vY0zs0iO8PlZtCPg5NsMjMJ6jXo9K5gFnY0AL+Y
KKQZ08biLZskSfdwD922WlESAiYHG5LtFJxWexX7OwbcAq2P7A9KmvuH5GbLPS3jfxwjS7iHRq7S
0/n+en2Os94ltpSzujlSHrIqBEN8699eOFVgSsmhyCo+q9flyMVZOUPPVXzkjXfRBPwopR7oju2l
9AYSjuv7zJ7HXXT0UzwCFG8FbmNPn+tT3sdwAC2OfA3cLOl0WNCtecBmyPy/HZYXSc/mqaQeNjpA
WYO7cXcq9krI7Fj9DbYD98b173W2KrdflItmvyVuB6hGLNgqHYvkOPWw3ctANSmxIIFnsRFfZ9xw
Mx/goeA+uBnobmLsItGDgaAxHosSxRM057jTOZ/PzjCqs1qzhLN0t6QmVTOwCkF5G3M0yTRXXAbi
G5u7Ujb5hEMZ/Ak9/8a/RnVZvQ8r1/vqCa/LfEMgGTM8B/+OgAb+kJ3f6R5unQvDP4MXfuC5adWi
N9/BeoDXKKkf72iccxREzkeM7FLziubhUWLJKE9cIOm2ALHILd7rsYvKKP9jB0m5uSJH/JyZ2VSo
bLnYV9/rV0KovtzXgQnghBMuY21bR9Tq+DgHM493SojYX3Zr+ES9ZCWae8Tv87d8oG7k3KgxsqA5
EofDbSggoUbgaBblg9NNt7nipojd5KSAh7o1B0rBm6kmuhqjKUC4DZfqKQQl5/SpMS2Kd9lJnOOQ
Uw42QcvGUrrYHBX0MlLLG0XfDLyE1CxrMo8IcwVf2roQ8hV3rfbx3B0Ky3nsXYPz44vWQqlaA791
REh2lRiKQyOsIGirBQGvczuZf2vC7SmaDW/s991aq2mt9kT+sc/kIDR+DPOL5pG2bAdFhDnHX9Zl
DX5EP1nEJn3wNSKPlTLsBVvaXqjiwZZ6yrfnq5E84Dy0KfgebHg4wdPt+JSXSXLyvZSXk4gvJAND
xhPs+R/b4vdDUc5BKKegRP6LWXu8Kn1L2Hk4T9EHtnR8ijeajA+h2zj35lR/cUJvwdFkrnVrOgLP
qF6nclVhlmJvwEhbSw682XXjwW6io/FYjZaUlX/WKmBF4nbX/bcm21gR7q45jxBQXCzhAZ4VqC0S
1823qUL4eQtcG6pepuut4fjsPvjLZ2HbDbHh7oNrhHo/JKPMJLkJ5uUhuKd/AMYf3j8R5Ch9FuWj
JqHVVXXTCLCx/x6w7xu8UpeNsOW6EbzfMZhz5UPqc1fd4d9XgqgWTxcuzTCKw21egavdkKLGeSEv
IHqz8r/AGvbLQeKFfIVm6Wqu6NxMxnNcJytPQdgyKYsZiQNWas+ys1vopgMmgkuCgt60EYgcLwuy
aI/MVHfFUbM7yY+oull4ycQM7lqK3k3kDOF3K3UQ9rwRU06SIg/qz3hfcVgG5hyyDXlBvde6H7YQ
JFPf1GH2DimTH0P60B0Dgg/xUZmD1AgauUTkPT8lDTpdQT5SLS+TW09OVdFDJP3IbiWT/uaXsbq2
bSPZDfgOHsXilPOvNAvJbplfARsK2PUB+V7UFd73UP0uJZ9RcOwRyD/EtoCt6JvvKYVUpaZ0x+9B
TzI9aI3Admk+7TZ4bV8kxIZ/UWkDw4/J5/Pp4yudaNiRLwG4PdNKxQ7mePoOhHMNRb8tlvxtzkuY
8arhPdIRDwYVSrSIFfBWVEnt4yKtDScxJA711MZu3zjFM1ykV8+zCQunUnJ+BMcNcvjHiCWaDybo
Lip8DBVVpNlCA4IFwpm/VGvc3QavEB9Nt14B5M8OiJFjmnW6yMnqw+rWL8mZRwzSLa7lGQY6gVxZ
aKgl0XV1gItRQXSttI1jvwxHvhKQ5QMpfmsxR/+Ww9m5Sivk3qiLsIjKRRp2YuoAd04NWrOYxG4f
3/WZFliNsvLC1xY2BO+mwIuL+m9JIXZkXDVRd+tB2uQd+VxPc4vn5WcruyBUGZA7dgz7W4SbGehG
yuN3IbDdsbMACFME283+zzNunBQ8pBQe9YrfIAEAEKS5DSSKJCjEtwlvCH33U1bAwF7vnYfG284S
KgL2EwxhOKpPRWHf0RygzpwekCGcHGa9YcaawpkxPTGaGhLKBGh0ET+uIBAkW5hRaNyXIVk6SrDb
kSaT5RPP/YQRy63XzjNSvATkQlR+GB5iYjqL0eG6K+8/MKcvvrO9sEFLgUjXmlfmMvu2/rMa+PNZ
hc3zQKMVlgpZj8nknGyocOfSYG8Trxnqucdm6Jl8lrsGpJY4dPJcMbJszSrjpBygmnUEsMUISv1T
znfGmdC0wfkVBOkiFmOu6eG4FUh7HP49ocb3QUflOivL2JqqiD/buADM9lsxpiUlDFo9K3BTKZTX
AsSjBgVngUpWQGwsWVARRF4gyLg0bPLcRXAsxkdh/nPn7EdlPuLKf3IXrJ6WVGK7hj/YCUzVC2Wh
sWV4/TCBsGDqadR0OoUqY8koXLy+xFNnLLZnejmjDiju/TGBbQhhGaP/QSxHYjIegTYRNffAD7DR
BvRSBOOr5Ayue9sdLeRDSS57DRMxwB7uTUKVRl0+W93Cii1W0rbekseQtpRbjjZcDO677UnpDnGw
jRzawQwRcYZydsi2tfHx+t4alaOWW3Cpm3wRFAZtasfibrDOQ9L0ILZzbB0pFdj5zwo4yt9zImjO
XJB6YHXNiMHstCVRhLHBaitVt3b3agSy8jXf+vRkPkFUQ7x+y1qaPxeNsYWxQ8sd16jF1kJcN8+T
Nztuk/nRix1loaXM4jMFPz33A0NNRRIXG4cCThbKOG/YMErHaG7MYjG4Ra/h+FNNAqS+Zneo8UYp
+JjBD+4iFNm3ODN14cnU3ojOCnZe6n9+ZQ7C67anbU9Gxi6hd3eKst+Sd1jYXQ8pRPwVFKl2ryUa
g0PdWnG3wBuhd1en/G6jn8k1+QtrZnbYDAqWjnuZdkaKUq6PY5ZQxTouS1DnZfwJ/7XFmBRI0NuB
oyIQYdKkmoAvwmLhtR22xBDmQjJJSjLjXtTcxns3Kgsj01T2M8ttI3io8+OOwi/WoejNXkWgfWRK
hS3RCj0OtQ+b5CmgKMAxOfG3j7/v8MDAO/DKMG2R+KuraXC1MyQuGGciDk7/H6j94cU8UgIsGEV0
+YfOpRIi3zO/4d43gvphQ+Q/9Lj1iljAasQ7ZeSloFdyr2OL7hCqVAGloweVJXZ39Q67S1ZbtVxU
HXW1Ln7yF6ht9FX2hzGwZ9lOpEFYIC3ri0T09s4C+/O6vhjNtW2/4iTw9D4IyLIGHGK0z5az/sg5
476rCj3vWiA7A/Pq/WeU0szYLxAcB5YNLpUYjjubFigCOBMfmUiW6zkVprT3BrfqJJtj0vcqk9VW
noyy+PWUujVaCRfG2ZBfWmEUhg/YQNGktejRVTXMVxnu7wUGaB+pBosBDNUsgRqmVW5iSIrX+Nom
7bP73/6KnpVDZ5hSVgwgCjmvtGBWzebTu0GYSFiiPG7O6sSRYu1v7fSEPIGi/2RLc77MvAx+THxM
V/w/owP+5Kjg2rsx5LAMu76zwVvxY+2dpxtvb0XiQeMr971GE0wDryJLgGgDBqv2VezaicGeAa39
DFt6rK8gqcVdG/1Wepr4xWB9v+hJek1ZqpnU39/lLWtSvy/yxSwITB6EkFnAq/lz7OTxjmJkqQM4
HGgyPsZ7mDqoBylQeqSlwxfAgcktezxtJ8EFBbq8SNSGp2Sp40aq1dFqoBTAPGkyn91+G7j+fWKC
GNIEtFIZ5cieyZ5z4CrOSWf480UmnfRJ1oY2kHcJ8IWHKKf5vAhvAOZJvszvU9PaSf6RHxIAJ8uS
ZSo6GkX52vdWN4g67ZAWs5J1Pt28DMi2lbYaDQK6HVnFJdM8X4G2SkrwYJd4Yz1PNdYkZu9Gunad
BY9+kjR1+Z/SgWDGcIvBYg5lZyY4Hif7aKtigVtd723VKdAgzItsSAl1ccLveULS0uDjavd1WUNE
BbH+dMjeoiPj1SD+UcvE/jIRVEiVxqgON6VudO3XYWjg4HIbw+vFVZJvQABv7cpAa+qaU06ijzP0
iRApaGvPUE0+UH4rjB8Um6k/mVeEJK12ZT5abaYGdJW3BSdZTUqJ9lzlgBNFD6T1UkMHUlc3cMbu
yxu19GCzfwIxlzap8o5FVjHRoAERdpCXKLXifw7YmZqiVVjSfIi9F3kN3jDte3xw+4VHgDUdTmrM
Iuv6TZShsf+3RcFMOMcGuIhRaHHP6ifWql6lMLvdKC678/ofky3KmB8mppoe5mlT+lXJLpGkmM6y
yxfUq3gAriPs/Dy9iUBu0AgHt0cyozmyt81+8P2COH1Rj8bmiRQCJrcSI/4cyTv/qVXJgUJuanI8
Q5AFZEze2CfSG9rUh3y3K+ny6MSCF2RZU5QYzfcrSzJwfkR5xMq078PZKYY3F5yMj/hJzv2Jfikp
NC7+Bbz+iJ+2Qxyt06wFe/iNCJ/Ov2Ep52gvZHBWJXlbdN5DLYtzJJI4nLaqopqGkaK8RQnRvJAY
Kg8YvGDFn0wGPrSiCQhjC0CrcbpizhOALDMn2f8+6Ww3R89SNw7CKbWa9oXAIYtUPabU2N2hOQ61
nBQ4JaSVkV7I1Mcl1I0ZSFGsY2wbmcfwsasHSsIrC6tmCEeMcliw8AZnMX7jMDyQLbleFs3pF9Cz
Z2BDmLPcmyq2ZLix2GURghHclTshoysXDsVJIExqDIiGwTMtQoJ/KPC+s6pMf2PqW64BP67LiGF9
BTdcpS5Og3qViNfhUxY9yZFcOsHnj+8FSzoMkFlIR5+eHSE3i1D5Tlr4pQq0oiV8mltvSfPGUkKY
ymY6ZVYjZ6SW92XYppdbHD2NmSB5CE3hJt/KFyNSkrblsQWcfR5Q2AGNO3t4GJw4EarBkts9hY1N
bYOQe+j2KtIHEngJ2Ji3IleLAw6FqnWZQX+zNG+U03/Pbr5AvITdz/ubKp5tU4mwHCZwTcIcLedo
EyNXcxIg5/6r87ERyTIh3qpxFgTVH7LgiYiHGAyDRjtitEBVeldRTWGlK2LuGC5Nc+dN734tM7EE
54pAUXNvY6/qFOJOyGX9tPVQBSNkiehVrBTR9VC1UAp383i5CIqMONzukX+gDLKj84urtO7DluPY
n/rUB4GUpPci+Q7fTsNGTvv4VCvvbZJdWaCpCkS7aaxJdAFWU0HdAyMbxcwnRvMX7VNrmj+oyF3D
mAOCj4YW9R4w1APLr9XztrSrYaXF2lQyMPlJon9nKqLAGW+REUI1T3tExcLQiHt1ws8SPKoGvsdB
D6XmQd1ChL+5dl9AIQaFen6Qb/mCxanz9RPcdVeRadsG6RLHT4yy6x7M31ZTms4m6DXykYhw6Vv5
Wyv9ZtXSWfD7FC37urHRut6mCIEbB0mgkD/ikvTwZ6GATwvV3zkeyqG8PjzUX9iWKmG3bVHCb0+q
P8ICZBCgW+RVahkLQPeolP8+71lxUg4Cqisa00+BDaqyI5IyiUMNpwOgHKXsO4B69gi3UX89bFD1
wOlu3fpvQXFAkY8dx35FFgbIOK4YZGrEy7UZFD3LxDx1MQ+Cn/yeTD73OPuAZNvtWy+3mZqB+I3b
E4UBNy2mNdtrkXwXXMWTj3DdyiJIsMRy1mzRZi8s8gBJHhlKJVpvd5N4xAelj2LKeABW77dqa9pU
QyhzOC0SQxudg3R7ZolEurUik9xiCxQOgGmVfN0luiYACus+RqNmgc+DKo74CUoK5sD30ySknfhN
dnLeKL2TB4yOUytFxMOdm6xcAImIGUKPtJNeKhsX42romBcZckMC/TS1I9LUP5m+eKMRwsV3/Csc
3uhPZTcKwDDWNTXYOoJ5TWn8CUW7BxapqDN6BTYTgmF9UT57HRjtdYQLQZes4Z7mC9kQHducqLic
NFTwLyaHcfWi2ZwdqA6GXmPaa0dJGGM3X5Yb2XMN2leR7eq50Q0fyKpnfHTENVM/pgTdYe8+KaR4
zObx8f+0yTs37OihtsQ5XM7AgADdrqk8WhRyRyNdj72+CduDvkTnsSjF0Qvej65UARoaaMVoH58D
CP3FQCYaO1VL1AckqvM6gNEuChCP/gRotlHC1vOp2ffFeiRG4pXdqFgYcNOqi7mxqXTX1DneRagi
nliqXJnplQssfG2guqwig3Vhm6CRSTkiMuYUHwmc/5Pi02El4ljsuCndQJ8JGQZwfwDBDVtUfsN7
GQh4ICvgxyvTCYYyjwvCOon3t3hysc50g2pRgDqRDHbjiyURVbNL1KE3d4qR0J20GrMsrddzlNF7
Dnp3iL2hzr1X4ljPWFe5IlKs12nCeiMfqdv1re5tviZkaGn7cIIgYXFHFtPLWoOmSRzT0k4fC/Iv
02NbG1p/el1IdMzq+YsA+VzMcLjdLina3ulDWEF5sOSjo0XNEQYRQHfsFGGlsB0dVrrJyYjaU0h+
LpXJst77QAr77KPXpGtF2aW1je7r24LjSbXWoLbYZ7xZxr2IvHCdw+j4PNPLTpAR5Kj4L+DV56em
V9zrssuybhURLmDySLtmZ6mGZ0tsdDIxJ5Odsp378Xt4ZTCA1mw4eSsxbqPXtFP8/2UTtDStwtFu
27XLUK0O9srqWWq9mwhsTaCA9htPFJIncP0Xo6aWGm62ZC3QtljjUFNcyO83G5aTbkPZhqZK6Hpb
0/oubZL3NQfkVDIg6XAhN/6EBUqHIcipI9VGt5FcppJmYbovCbNz/Yl7wW/WA4Yvu0moEA3r6JKT
TTZpue5CsvKQagXO+f9THJTNbTulzj7jKNVbg4qJgF8NGDpdcgldPUd9mvXq0jwEJUQncTIeoxkD
o5HWY1S2fMSCa8bBuSRaXJQ4n2K5YCCBqX6tZEAB8mXayuO3QusEnL2eswGKM2JVi1XwP7gnjqBh
rJNM2dnyc+EOVISpEpa/8oRwIduHs0OdQPyu30p5c6sptn5HXDDrySDN3oNkqRjCXhfYLM2Fp0Pe
MAY2m7LEqOCDM/BZkkGjfrx3CTrjXsnM5mT7N+TYFHtPUMXGKwQF8qiIa0srohdQqtN+jH7OGXnb
dwOSJJowSJexg92/0Ph5JEaYsD5kRFQa3jqaW6Zt9KbrW+4IGUxjjiIvFUdmP3BcukxLm743oFK3
Zk8HJN9jzQe9cYdcg+kHQt7RMbrs/Hqcb2gKSAgzM4Q0vwp4KdIt645JNHCinUtcw6qBJso9vEDJ
VpYa6yhduxDhRGJvJmZ29P7OuSOjPcz9HfDLKV0WNX1/YO4i9hpLszKoVbsVSM9sReGYUZ34OcWR
03ihXdwhLCsgonCAKrBLb0v8zh17eVPmOOb6ZTvl2+YiiEHdonxdtspzmtNOZD9lwHl13FxOsWtF
SDRGcEk2xNvqFe4IFkXzt4S8051+zJF+KCDn974GtoAL6T0HlNiSRUnXM87U4uLWETG6E171P1Dm
73s+YJZeCGCYdxy3ilsqxqgfhxk+pbNks0cV8k/2G8g73cFEvxwMmz/8ThGSPveWf93SgPYW5egm
LkexV8EOV92dwQB7vX9dkL1T9nMyp9HuemeNuSgsVpLs0t9qgHloSeiAc2aVa01DMyWFlKFdF+tm
Fw8R4Bbfrv9lqfFsWj4b+SXcn7F0pCwiRqXvup5EmhJIh+1xX9cJaputP3MJ0LELDxSgcbgO3Eo8
vYBRreG4kPoZ/ffDRABbN5hhYEMyqu9yYjstYJY9Myd31TzEZoXS3dtT249v/pZBiUQdN783kX4u
tgcjLj+CC+NZcXNr5XhmN5WdISIH/+RNLq1IJQBXLbSlfbzaV8u1aTDo6FdewMhEI2h+b/C9Hlrx
FMq4kWV+hms5YTlSGePghK9R7KH/s4fTTHMNy1YDWVIQmSBiygbceJLyw1Xe8tJz7nEudojtvEWq
PXJZ2BHxQPBsvtkBGhi18ZBSMjCmS0qKVWAR7dMR27w38DaFFM3kEbuJCHfGln9Ljk9nTzLRRj/2
kllV/6iFD9gDXa5C8bF6BKCqNb9S8f/SzXrkFBeWHjyvYJLzb5BBy6a4ZeGBOcTImikeR7xDSFgP
Lw8HDQGzJSAJuz205maEzyvVH5gfzj8osHFFvp9UG2BH9mMb9BfkzzvjFbMQbHMSAUaf2p9ccXaM
i22khBrCnnnHXw4P8maPFnn7eK8iVcEF4320jXvKewCHYUTNx38V4/Q35IFzTqKoV8L7icdG+emX
G0izbut0breVX1dB02o2CyT8o2QjCZa6DQy2W+/XeiKFntoNP8RvY0AsG2rP/OLOTMiMZFKfSVGz
m+R0ikLuFl9k90XLkiiC5exnfGHF/UrqAI3ALgMBWIorTfIPLYfiBRvCTq+LIiXtgOSXMjrx5dFr
0wJNRjjHqAthOEv+Py6+Pev/C5S1/IjxKw8VO5UHzRs6k1wwYdWtjgLYmnGZv9woxCkMtxaJZkJB
ZMfdFX9mELB7g0F3rEqs9ykWMPhJGJ1rU8tBH9ESHcYR+TjTYfGwOQhUv4Og/4hHe7GoPMAjftIy
Bwgz5SU54149lMqmHOHw+MHdt0g/5IE+OOBmg/KZ57uapxjeEpqHVaUsitXvf4fxqJRKyu+R0d1P
a2VVEmyAgkC1GaOBapYZZjlhQ1o27hrCeaiC7W0jHKM1oCxiVHeiLTBMwvXToWU3qbeyPjDqHIiO
bniq+vf9lz1SY0BfVZXqiJ0lWZPd8dyQiI9dFoH665Se+0ZebNyGK6+e9TgCn7B8KMPM84E+F0AF
DxUIxf0xd4b6TbSLyEqsBWm7xnnAq3W65RvBEOOE5vjsRIzwYrM6SYJgijFqaHUAtRe/sM3yIWvB
kd2kdAeCNgnsZCHxxmEDzV/rZJe3uBCQO4Kur9ngBOqo5u+ZnUj+DMDblDIi9vnpMlnr/6qB2RAl
KHZGu2+wPHJnWwJNAJG2SRzJ8b2aOf7nakty9SgXKPHXB27WPSQ5MU4HuUIuH9g67epqxSIAhN6z
/MmbtstWkSpXKucLTw4dZJsoqwllVBcdt9OTNgeH5xcGPZ+WRlzgmWodzF1ZicmNJq7vlmkKKvLm
w9gsVMgx5MLoLStoG6CMsFxpxlOAeynQ+ZHvU7N40lWVgsRWdlw91SiYp9EYDd1eqGFBQ9NXCLYK
6fEK/1QZxRcFctNxin9/fwO0h4Xk3WNYpDT5FSXjq++fLwvghMWrnDchZZhNKiRYYpYWCeDQlt5F
25BmMd2cjP+jjCpPDCLKUCx7IGAgYEHKTC1mekyke/7qSLgoM6DpmlCtivvDXCcMQVQw9OFphrXk
R+YRI/8RBzxr4EJHdzVESQKjBOF2KECxzaSi5BMOEleAveBYIjMMKFR88D7MDDoThb1WNmr+GAdc
r+a8ElKZw86WbYhP4sFMicQBq5rkGYzwvhrrram7mPvhr7DDRgxHVwATGFdS+EjYFZcxLqRLup8U
QSith+vbcn42qRuF0c/3PpeTQVxzCemqNIdiAmJGVHcTsv4JMFW0rrVC+nhEC7f9s84HrcPWtLbU
U8B5ihE6IkSglOiPTfc8JcYRY73Gc4k2KiDnWChakTiyXwVD2c/Rgn8NmeOl0vMD/IZITLCsVJyr
CNBZ+jlYCY7XryrHUO0wBOvfOcf/g8H+HXnvu8JRBt4+1wYmyZ6DAuM8s40na3xF8Yymc9ZC6T3H
rQ8GkQoHs1fmJ/RO34cXU1zvxxOSdguqDG9/BlGcKvvKXX4QjqWIBX2RAKOdX28SI1P6E3IrfdP0
Snu/3EP1uUtOoDl0sy4/X1bv2O/gXnJl3xkH4vXXsmynNZYxRuB4yeFV40n28L0fD/1wXIp8DCGX
KoKvT8hHQZV+WKhNtphexCVkSiUtAji+eZDsfCWpfQLof9LG/IAXFfz4Dp4TetIrwEiGZC4YiG+x
Z3bqQrUV497/YhsZqtmHc3cx/X1UwuHr2JvRw+rlfEn9nFWN0RvE9/rxZy3V0RDx+KAJFms6OMf1
StQKRILF6z0DSxThnV3CpyQk7dEo3uFJ4pNESEj0AypAo84s1vLMtoniBGDIF5B9ylKtbL//OnVt
4MNFM+8Hf1jV2rUn2euEJv4vFa/TTgkRVd0eSCEhUgAEkehfbLh8+wRkZdypH+p27Ngt2PUGYxjM
cP9V4FrOQ3l0PytPIzaZUAtYA74JcW2zV4JbrdkzC5mFVJXosutP5LMpFl+WrkmO5j0cmTVpH4F+
i0OBzRxcBGpmbHGiYKrEFyNo7C7xhmcxvuUzYLeGjmU9XmVJtNaOiK7C/rcXraJ/cOnCFB/wWykG
Vi6gLPRtLq3oxDERhsL7/P89xOMmai+m4cJXSTlmyxePN5EZrEzgg0mOsbAlvaDj5H5AwsglqFcU
hCZTHoyZF1gWAcVmOp5Z6br0iQDCsVhwsXqmyuzlqU9sRP5bTajVHGvUzJu1CCcSh8ci929ewbVv
wYgUYTHrULlj+08xi5S1/EVhjyxegt8gJfgzdM7mQRrv1uWwIvzDCMpPE2F/1eo4H43t1Zt6mTzy
NnCdtVr0n7E7oPasLdAcslYAfqjMT/ezAa2StRWP2ZIn9y4Bx9AkxTBFclkeI+WcHJIUa5NFuGpD
1vBNBDatikWF1jeeiSxfdVA/mK5N54tEg3ejbu24L7fc62786Utobd5b56C9WLpIDw2u/OvxvkgY
UlcVE/VgGVHsqxmM1kt7H2Tg9Fqg547UaktJEasN12/yNjJAboWA7NDjdgeQGOoDD1r1DBf3B/lw
DvdVws2XNlmSuyB4kVDKdMzbX4ap4KFMsYW8XTd0c16hA5B6y7hzAqoz/PFrG7Jl+4aF0pW0XUqh
kRJGlkcsEa9OH8vw4KYHtl6YXl2bqLS8VkUMPG4ln69S3+Z53uurff4byowdTcudMO4hXP3lgIh6
XZ4UEoEykX0z/gZNjPs+fqKvlxkD7yUfUudC4uI1BN2Ybt5tqTaRN59MI23bX8awGCRmWL6Z/Nyi
U64bW+4duEcp2c3rEAUL/jgwiJCk+DRwUBzWTrvA65jxxGwboGcCZhJCj0Gxtwjao4IyYiYgRuZS
0Xa2A3Yv0JcubrVNRaNqG0SW0WC0Kbcv/vpIQcb9DB8xYJ7N70hI948eb9ZzwAD24dnknoo/uH/2
R33O6DaS3dPW8NXWdR9QcZwb50ZCHVnVj+0R3wuHrtH6wg3gH8y31KZn0nclzh9ecohxlG4Ikxzd
5//tUtsLeTOjSMJ4YyEs5mRQkcNL0tBzk7e+FGwS09WqLbwDpw37J+7k1GjJLkpDveSlwouavrh+
2LSnRcxSWJHNiLMIqnIbaMOyL+pLgGSNA/BfwuKo8jPLEeAtln7LF0t+ogJ0aNfSNR6h5Pnl2Rg3
Lw2mqg5CeHfB2wOtixVkqBe00OL5atqodM4ethXwibvguYYXs+WoscugRuqsMl9hTXatDJmhrbCO
Bc5iZtWQR33CDQT2XBUb3EXXxxKu/EuQRdfLw9oQvO36VvU6xhfXrT/5h5doihiww6ZvTGZivcxq
AVcyUa2tgl2kTM9kawQVQt0ZBn8m3u8I0XM8Fnl3MpbATf1QChEgzqss4pJUpaM1Djd8AVT2tCp6
xq445XKZUfAVMoGwnNZ0z00JQKU1OoDJ9919jil0o2d5wE9jTb/o/o0deVqMcZnk0RY/nGgzczZn
C0ls/gWsHDXFOyMYKnoc36ovcEiDSN/Akrs4WuLsyLdM7mA1lefKNnIc3H/KF6MWccrz86iA49gh
Oqk9Eex5u9tO1KtHqilIbBN2cIweZ4DE2zUMNzPczfhS5hB9eFG5ngqs0f+6+oQcdo+jEdPT+mND
r8Bis21wrb0bGRPzKcthhO2Hrxo3z19iSgvNMl2+ZG3uibV2Fe7gBzbuePQbE+CYV36YTBx9lSfE
0uTdGiCcqUdqudehOhJKxH/7UXyZFd1hKERMyRg1w5VF6hyCg2vey7jm0gy3YWP6quq+744hxtpA
2vxhV7oqXwjIf/9zuNXq0tioljAXebww1A0J0RpdIBYMi4ZPLFCO/HMMcpQdmswVPPbcNlpTXsG5
iJ+/hktE8KcnOqGc4N8YipzBMX9CFrwPR4rgqonrNKb/PHjC7eZaOF4THU+otQTUhYrt2bco0TGX
YoyPhAxst2pMNlU/3bBHC4Wao2KylcqFFrCwI5YBNGKMafEwI7DNmsqbgBtakmh/MHnH2ZYyLBmu
sFqPqeLEU+Dm2vRam+MSnitIuzsrsS3I232eaoPkGVAc/aw+Huwic9rC9ftXdtZ5W1XlhFOxsWcs
E6g4TK/0VWWwuFWL20M8DadM8E1G9SznVJUifAW5/wDTfR74ATnxrAOsatki36OsVQNlQHmxutec
L9Uh/jLFMVTOgZ2D5+1zuvI4L2TlbvlVo78eljlW9wDQQtvqJMdC/zKNiEX+u8zeFM2PsQxfJE7f
9/iJn6DuKiBjFpVs+9RJxnro9yA3Ni7SGuahE/jDvhUXo39sJnz5klg9ly30psxc2lzRTV7xaBjk
IRb7HsIEJs3yV55i2SNFtsJHJi2ZGevuBol8bQL2B/OrJM45tf8EVjxsTT1onzOqzVFCysEEsXWl
jDEXodSpvm35uIHHvfGr6LuxQSCsOZJd0uP/NtojsB6eeyH2i7HhuQaEEDUPgPXIDBbK8/gS43N8
Qxajxy5i6+vVJ3zBKFcDmxNhnSkD99QbPHAQRQPT33Dcxjhg1q4HseKBfT3yvTDoSVOuG7A8P3Lh
9YvXnDmrnByvzGXS9aoMORKg6BdlMAdTqL4am/GBbdHUomaT2az+Eg+nuUJadeZx23NjtBSHxD9c
icuZ7otfkd4wiBjQ+YYbd8Vfi4DBveUCVnG/Iyjm73uXsiFL+BdbbFb+gqKIiQnit1kOOF0Kfm12
j19+suA0BdY9parqSisJtTyzQ8DbRbS/6GDSP9ypCSUwlbvX9Mtx2D8skBLUBnoQy00HGo197eTW
h6Az98Dx1qdVl6Oj5cEu78uHTk7VBk6wWlu+OIzz4Goqc7wSRiAQnwZs7/bmvqLfuiQljp/s/Rbo
g8nXW7wG/Zi2qJPnmkuXRzRqBX1llewg/S1qycPZ2wJwi4L7kOEpfzHCnLey65Uu+ywx4xwTyeZq
oWHi0G6Zp0ON+Ve7mK2dKMnu6heNjOnwz3Hs9yXKdwT0Iuopw1cJCe8Hp31Ykpsi9rcWRFw6SQFM
Cp2LQQKY3TmVuv60Xnj1P8JF1oP/gizc2mnBYnNeinfu7+MSEet5JYFCjTvOAx4sHUNcBvDxEYpH
rD257xEYPObpXkBM3iqk5XzsPCTdhLL6BaNzUM3uNUEk8q3bpbitMCzdkKyJDyn95d+fEmzInAxQ
XX9tUoF/CeL4kGVIGnEE9U7jLZqolpiSihqWwBjtc7mxqEXnBjxjTHszcrbC+zKgmUKOCeFCFRth
PInNtWWontN0S9qsI+ZFvbtkZow2Dvu/QF9wTYQHl4xNhOBf6sk8RZRO+j5E0w0s7hs3fL++o3cy
zHJT7g6bdhBV4hUdlDPiWP1kRufUJCFXvTSLFcYjrHRBGDRCHDKVUo4REk7T7tyeGcLUeOAmiGEs
GOhA6KxLtw3mg3+I0U8+cSrSSBb11Ov+IBBN2udxWdPC/CftCy6n8h6hX02Br/tMd2vn1bYtFu8I
IoqsxToiPNaMvOibZ3zWWZOp4M9K0ATqaUO3A5sMIUz/SCxOTAkRrYspZcVq/pxaxLuLAmgB9gaD
aLnbw7zFz1KzkL2s/4/hm1Ei88j75oRro3n8s880Maj87TlRAgC0zAkfWXfKLlh4nmttBO0f7pp9
exVthg+dSZpiZ75qyCvb/iUGVzp6dy0EHx+eDwIs37ObUmXb6xiDg7tRtoYSpERf8PKiqYbmzaNy
N1UBQbyZpRM0mdvGBNN78WKZnK/Z4Tst2oOAPA+mT4A08JawmenS54VpcKtCX3uMmQz5Fu2J8MP7
IlxaQoh78xebk5mUroBneTFvbsTnPUggwtZCYPNzwEaMnM9MAHtMVsE2ZffypFjZDQJto5Cdi07t
gGwVMSYWS0QNjQ6EvMm5206Qu3D+/sf8kno9sSfa2drgJcAigB8+gSbvru+jFkyHPh0vcCTaAyub
nEy6PcTeX+AzGxbcRC9rfvFtPVv6ToiCzqdsQ+avGi0Z0UWZe+YFlucr+ndheeNwmCNY6uI7QKRP
+QDHjkUK20KMgzqtwzRxxo5EJeq8pMOyxkRpSK8dg6Xo60HOBuorkDv0avoZt0P+mYICpR/bra8/
N8/f1gI9uOWmw1k6SGK50c/c0VMjY8PrQm1d67g5E+h/Rq/yt8/ZFyJzKcJADK5JKKcCy787vpKz
mZC4QYDbSaL5E+cq5WnWJpVtxiBw/dp4XBL5t/yysKJMm5P6PaR+/xBtzVHvL+0JSp5tmAUqE7wz
xi70n2seo/U9jHljuFY61x+hd5AM8Ri1KrmBLLBat8dhaQCuRB70G9kUzmLoMDRPlA8OAFi5jpTO
i9eOetv88M62zd7Z5vrCwSd0dupnFOkrkD3FQ+35d5vE8RFVZeaqjwxjfe06y7tTXNtEfyNaaOvN
nm7cwIrIBBs2yiSvm8VZlBYbFexnS93BxN5kg64ihj4v+Oc2rfjUpAauKo80xpXYSiInQeBxnspZ
OW/v+SqM0EqW3MQh1DtnyfYNBc3+h2WXSYLTJqORDyzIT+MxkV+OVlrafNTEU30k+pAlFpiXs3uS
NXutnlUuz5RIMO+8SdYn+CP+aSXiV71k0AyTnYUvNKoISqt0Mb5sq3ZXauma5uriqxj6B1cuBDc6
BOPoykFDccZ994S6WYwJSrYiXTxux4SfQka9A8H97i4UMEAtnMPmGGk5yoaLimxjJcRIIrpce/p4
CutMSoZVdaDjLOzjXGX1x9VD0wI/1tPZ6b5x3L7Q2UB4nv9R24c8XSiTUhfp+kr2ZbVmiYE8cRoD
6YWvvvuh6Joo2F6fZ3HFVXnOy8aica1tYo6bOj3YG3bZkRoBLBm99dHgh7IC4EPfYgvNbd8xAeDJ
QrVO6FpM+rr72eD5I2kv2/1bviUzMBETIbn0VZkvkpu2wMlQWiN721UcAIbTzqlcbqdYZJAou7Dv
4mA055WB6pUxkOAvaj8ubQUV+jceHdNUKQE8EqRu/QYKUA9ZfKxL5IimnE9dQwKIlZ/TkLo6PqI5
qGXXMqHTvFIg9YGpG2zxjzkzJWNp1LkksWt90fZNKVf/dZlqk9fFfNZrsBpxmYgOzlHNJnNF78hJ
3Z34t4f9zEcha4U2Ere7iUoopkcrLR7skzU8XyNX+S39mi5i4T7GliTEQEmYHDEOqc5r9mIB3ZdC
t+nXYWNEvs9SBYRVuwrNxWi/BNRs/mH8/j7XG0stFw9mIpL1QdyST8tIlSB8+YVt/8ikXVsb56l4
hf72ssnL+WtUYmfyD+3xDJVQyzVYFoCZe0nAUyjEsQDAz5L7Zs1HTDq88FLGw8Wwob9qGHJBvg12
+lp/gXG0ZW0HOGht19ae7fhXtSHIipvljZ335gGZD+IndUU6OY6XmIwPOUETvCK1LlMQlER6hWyh
CsL16ZUiOl4ETWt90OXG1YIdLWL4ql/EB1+vDYpV5ksLNrP/UZIXl8WHMFBN3As/PnmZCjmyEVaf
TmiQG/ufEcErFAKV2NceqoyQv3gZ+wO+tVk6/jglT63Il+2H+BhHrArSniEV5eK2+KxbKJ/aut6Z
2YQC89fcYaVJ4TCibQz8KgX0/1JJxwDiFEI8dTEgUJA6ykBXbBW+zu0G3mJOgzm8eWCh9DNSD93H
1E3CkgTMctao30ReVBMxcIO+O+wRY71FGIvIqIT9lXmd0aKqSdw5ZrtHevWmAjuebae9AI1ZPfqS
KH2ehWB9lwLjtze2eBQ941s9nRg0OlNvQiuGwXPxewOVLZDyLJ5FARs2CsplShjWYabwYahrWYfA
yqfUkdnJoW8kE/0KbShREBkQohcD30PN3nzKSrVQCd5nt2H5+q5tMu2dVofELJy7k5N5OvaRt52q
KgbKRrnyclcWBawCGQfPA33+gmwmvchIq/UOz864zswN7Kz8UqOPDl2k9uldmfaVKPjPyElHmKRE
zHknQ/l1yxFJYaYLSyg61f4p/I2CwuXfdFSF/H1hnqqeked4FzaMf6/jk5hIAnZW0fvMBQKVEVhn
+o8TF3Rypuu2dljOFEDBauuPkg6AF3lrd6f9ODwdFxa+7/qgoD1rceRCTw3OtDlZAWaijpZ5kPpY
A1o0aJmIohWX+JZknm8+uLyH4akmXUO6egvpEM/ffQnCR72c1zyAnOYDncPA+nNDrbcoqVaFdNdU
8TJwI4EfImlWVoqLJUgl7epgXbZ9OZOZsGAja0qbcYnVoC/yFDqzEeEBnVjoVEAYKlyv72UvsjVr
rqTyP6aVmCP9lPCeh4fzJqtf8mZD6Dw23mGZj8fQppO9re7KiPie+DccTEJPQnowIr0oTXLM7ub4
nB8y8vDnjr7DdGzZ4iAcnVodzZZLlqOh8zWleyfq/YgRSlzSex0wzGY6gIlPjo9LAL6l5PKQ0jR0
FXcjtTP76pJy7+R+IRPZyfFHPIPPP+dAJF3UpLWy5Ls7Wtdh9Lo+ByomuAFr9RRiuqbFJznkUlgy
U8WjKqrH9QoaGfVNIUI1uTA6Vf/IngZ7G8u66UcER8fPKNZRgjn+NdeUwbVLXXWg5kJJT8cLjB6u
NrZi7UzmFAHVwSqGG3RfYahVFAInFwrdWPghg62ALCRXSZ2AXjF1JiRSFEXQkC55JACotxza+YYb
2iunnrYBIn/a0/pE4vDh6SPDixcUsDF0izfJcME2/brwUJrSBeci1QrPbyU3DWTwCM2pJz+kKEh1
VbrCMZBThpDjJ1kD/4romkSeoWwWvJnbMjcuM5gzI59BS6oZoQA/vYEsRf4E86i2rSI8jipNA270
Gxu/oBP45f40cPOKm9IFV22I7Cm+EswSKI6LMFYYLn5Y0osNyVH9Nhy3dwRf7NwxYGMDqqL1KlvI
M46GcUsoBLmEmuPssXHcB+pm77G4uVNWqd3O5LbcZVIFPari4cpv+yo3J/Kdmgi1Vj0Qt2AbnDQ7
ab4tLIyxtXPXH+pchIybY+q27lrEnwBXRfoxtmx8NlFc30uvamPaZFGxY1COwgleZW4fwHGjBlkt
NIRPQo0Xpe5wO0Lut1BhxbbXxYcE6j9Fz4xuT/Nw1TIx2Z7qYxQlx2FV6zz+HU5XHI9OWSlspoGo
439x7+1OGurcCG1KprQHWJJ0Upyaqfyxv/pEwQMQ+49Ktc2/5W8gxozdxe39GL5rzVqAcvA8nZay
Bg1UBMbLM2anih6xjvZEff2Si0C9pTJ37jOxJ4BDgfnw9FUWwKIrKl8j4ijhnbdfEg7VIvwQqHdO
B2rfKvdjap5GBfl0Qt50fn8A90mzgFyKTy/iuEu5ELYo3MQAMnDyeguoid049RdRVGMJGW7JhvFY
JHto+O4GPlWNXlQ949+r76SSDC16VuqO/snNGVCLLf55RdPvrX7DsBrF5WGCZN30gZpo3RF0CLDy
mruLCGumGPB2k0SbRJN29iHpK/XlxJr5cP45r6bTH3E3l6QIaRiznpyc+CSb6CuywMfH+p5wu249
Qu+5fB3IJXcDmDHwKc0ShGticcRMRoW3KnK6KFiDMjIyYOVFyS/3UV2bJYHmkB9n+S+g1U5dAXNU
Jol5nKdC+o5TkgFK2vZAlxjWr4hnlRj9wpEpMrWc7xiszjpjQK2KsORHH0FTmm4HSeXTXC6gOi7P
tsdIy1guepkaoMz+NrZ25ZDgsFgpGQY7k9AUo0yHZTVXVIAIGAKfL36QWsk0t+MjaYZw0siySUOw
5I3T095H7jIDwFMlVA/E1UMOOM3nZgxfsokSUN1aCxqYtOvWr4HkILgrFWksvyOW8KsZEN8FSNHR
nzJKzViydjPQQ5vkywi+akEHX6tXmcfnaNQSNJe8E+HDMOb7s2MJPT7lxI9pfKaCmbL4sFCQK6Ct
Afi3iF3F1l8kkHef0KtZm7cZHAcOJGU0bDSdJiRD3dZ+wyc/sH5Th1OYzRwdLi+Pn+HBDvZgA42V
1WOdvaK5e7zrUNi1h8TLnaV4Uy5ycFk9BBETgAfNImXFYzaX3ZsCpxVOilyKpYdybQyMssYWUWMK
dJdSvk3FlgM9a8eQd7UsROUJW0adR/zbre9R2RVaoTT2EykfOO9jZRyFCYvPQ25i4Zjew+dpJ/2A
fgz0KYVqow5RfZgeoJtvxT/YWt/sXoL4VJTyrWWMOogdcSD3+RF1io2sRNZMbWPGgR//Vki6upvZ
DYv4MB8MKMtDElKgH2I257P66SCmwD3pTUovggInW2FarvwHkB5zMgLmJkEC8ue9g6tTD4yLnSMc
BGl4any6P49SqFmfNqWIhGXf+o1uLctnvA3sgrrXAZfW5IL+j5IFIMPItGJAMAw1MXsKRcu2RYa8
4YhnM7GbtHSvVNWYls4e9x6BZIETYKBvAM3n3+hquPTMihDJLPTvKwZ8/2fXp1yjS9jeORnbFfs+
w/BB0MfRLPKVe/dXUX3fu7xfhvtJmMkQHj0owXjE/qUUnRCRkeGTBigHeahDBHdw1EXq0LfcCE5X
L3ZJxx4IuxWaLq3hfopUd4sbaxVhCbjoRNiR/YdMgLviti69R7oCibfgO7LCRfV/2RuggW7wYQL2
5BqhwAxYtSXE0JMJ4KU1/lyXH3dFVZberUNr4gqVsYnEkVuT0RB1mJEDqk9BpnHpadksG7/p7M4i
tjo+TA20L5G5a3aTcEarp/ksuiiv1kSyeBp/Qo0ATkHGkYdTXEmvqG51c/RirM+Cb5UzwnRPwzOK
SIV32XtunXTCCubPqDCM4FceeHb6ch4SDZcrqltjNEonFewK+Rmuy6EAlLoM4atb9cqF8BPYgfDv
kxrnsh+x2dYE+4OVhR2c8Bjk/Ldg5hAfsnHV6/NYbZc8iosIqEN2pTvuRcL1/nbC8ULJnzXHEc3O
0OdvRQgV7SRVfDcXYK3CpjyMnMgqm/xnUT0zt3DG5J0ZWgJ+XvOnlyck7Wz9OoDWsTBqFEs5cnfb
S2n/HdY2l8Da4ibJuWG80WLd27LlylGxiDXZosI6Zxzvf1p3a5NhkMBZGxyBOc5z0wvJOE+5rg4v
gVCDMTaTvXg3FE33ApvFtsrcR1+GOem1MYRNalmrs4BINY79Vg3d6tFicstmivAlXGf01M6UDWWJ
4bsLp78Cvt8m2fc9/GB8C76m/MXMilrMN0qtCO+ou6Owh25pSdJ4fboh779GmU9DjJewWt1w6qQl
1qwH0lDVmPJaPYvbjOQh7wL3Ykb9ErnEMJYB7dSgIYQePxnG3aU6Xikq8hMtQ9hEJIZqAXXjYYsh
+TPzeZK4GqYfCdi8W8M2+7x+5r6x7WXe2BxIfEpdd2ZKcMQXC/Sl47Bo7UcEk4/eKR4IOgUNR0Ym
M33mZkGR6duKNm5wvpG4eBws64sEWTJN76+WJkAy+k+HP6XLoTbjr/lYyPSl2VsjxiMgoM01CMSJ
kYBcyLNrusr5FPhFyVnCHJ9mzOI8moqU3sYxSO7TmY3ArJ4fqsIhti7DDpk2LwgZ1tEo4D/PElcg
jG6c/leEeJPmkXQUhlO9HnPuq2XAIogOnXffAWXZeRDmNdAUjoesp2Oy0LCePQb+aneM4kr2+vuT
PWY10MYR8tVWfN8RWHD+aGuvlM8vR10/Tf8zZRm2Lf2T+uyy8ABL8CkBBT+hQUb8LIHCKmd0Ly+P
8+0jbGFOc2LNaeS9le83nJ65qiwkKmw2iz4xuc9Jo0t5qEBnCCRqpl3ZIUVrpzxrqCruothlB5n0
dKUkraLKb5g36Tur8DHJoOiY2SdksepeT2B9lSsGtHZXrhewUaNZfizezO0pyexbb9TbnAzx8qm1
M8UQIpS/Xpo40AKbjM3S2ApQO8X7R/wQUsPyo1HkmNB5c45bXtvdnLOVDKW3icdqEtMngTr1dreC
M37XINy2JWB1L+lLBIfrQv5cYhVtokOoNprPTDdKqKMg7MfLmA7h5B/n88X5PGyjoF/FOzpuhKhq
C8tdqvTb7K0BdHCDRVLm1h+BJeY3B41GusU3MWvaBOLy84nV9kAPWrhvqen580tNOuc6Im1QuSlx
rCZVFsbmZxlJ5PxL3FD13DlCFZYoWKb5akkGi6Q2GsZ+PzyIVpJyklLCwMmmPAi0qspv9Tbg2KB6
8+2qNaNymWBQb223yBOAVNcWfw9O2rdtKfq/Wx+swYC4nfx1e2hv+YzxkByxYrzs6gmePzXsGQ4G
4C8kKmFe3qk5ywWta/qrWgKBvnM3ZOQIwW+aKo/n/8CDk6LDttIQM/Kx6DiM4kIn9PbWBcw73xlH
LGlwkGT31GJ1HVD+Nf1+jVz60/a2UOfnmcCDKU9LpBtbyFjCtbFhEjlMT+wcxkyXwZ87gI22p+bn
mbTSY4wic+Mh0IBmd3zNw7IROtGa8mtR0q3TWK6hh2V3SVPbdRcUBBSsUQ1vh+gZFMKNYgDOCIKZ
KMR69hinZBICR3Yvl5jdrbSwwCjzbqA3NWsO+cGEYTdYDm/RzqmILtAGO/ndbLaTIW9n0duhreAt
Nr/EDrbwhbmnFLDjz18JJdkw9alrvJnXYk1TBBxwNCLnKiJax6KkD6Gt8GmCSWpQASUsQhyJqWLl
C98ac/AHw7aXypH9c20mJudRr770bGHe547MkQURovE+RdXOds/z/v4mNCzok78Z7CGBPfPJ6EMo
Xft36FAIJH/fhu3VEu1AWO60XCBf0mAuT3wxIC13ZpTsriU8wy1RBDHajmLBugHFcRBLHpOHi/Yr
YziBrB6qUG72Ol2v6qNBoTMprk1GRcPQbFsp/TE8MRmYLsvmCPKWkK7333l7rHAYgS0R+KdZYQsQ
4S2C9BQpM432iNvKXcUDy924TW+/yG3LFbzjwztsih9e1rQBqTsgdNAZZAtdoTk14foQ3M1uXjTW
t23Z/bviQuBMsLchnllr5PINKR7am+UkiFUtw9asAv9raXwuFW08yqFiGEvtdac7LEx8dxiUCYjo
CIrtXB/fjNvqA8av9Rh8sf1KLcA+yVR5zCFIPA3/9wCpD9nTwO/wEzGDbaU/CVIoz2diJrXfOYvB
d80U9YC21HD5WqO0Qi+1SEZ0oZ5uKsZ2kuSTdlD6WZL8pEvxKzmNQEnXh/KoyKsp/7chA9KaAAeR
U0Q6Gz2hCcP7LDIZwBroWN2Adl2G2HmXrll563ImqC71h57b7pYm0po4KSOtSI+8+IAYt5+115yK
9AzUKVeQaR5h0RvpxRqX0z5+w8D0KX7SK9KPHDw5fyAv85zCF3fDZQiD0ol1bfPjWAEg+Y5erSdI
SsTNVQy7R7jC/pfBlZSmMfSAvdu7yGxrcHSAK/iCPLoEncOCXTvT6AM5k/kM4Dt15x9qz8imiIc+
Bf8bziKRTlOC/7/4w1F+2AFMMR8EfU2jO4dQ2W7yyj1rFdCHnvnGOQ5uVScUWN+T8Hpwx5SrLuYs
C1i172vLoePiRfqWA/K5QQkiwFglxw78a2OeEja+EFQfxFXKp6fI3CB/Tc/ESrAX6gZcOo4Wyh8t
46/L2YnQz/6phxfa256iXU53a6wVPVlqSCuPTU8K1Cx4zXbafVO5/8djdBcvVDd6SRPHnsV0R10H
vAV6bHXN8faDDYp+86eS43p1Fqfn5aym2ml+3HKb1r3Lkc0+39tO0KYF9lwFiy4rxPddqWpyR/rc
DlVs8aipUGFb8EOgM/oNPrav9sMRWaz5Se9WT8hm9YRy+UwzYv7BRni48yy4zxi7Oj6opIu5arAg
F7TrEl5oKv5SlX3aJhCm/uakI3gM57/lPdjNFCM/KYDC8PYU7AicnQ/3UIw5PLL6gB/8M1Bq0l4u
XIYJseARCyBO26XMcgaxDQ3GS56asqC509kj0nOjMIse5JZ4g+f5bDZk4NkTeTfBi6OoNurcTm2R
cHGR4tDV0AeW7JccuboC0bWk8P0YxZv3JhEMBzOVUz1sBQHQZ2Kg5tz3rGQ13G37LwTDMd/J978P
Tnt5bpsc3VqtZixx6Wft4/u9n6xM66AWx4bTzb+Td1n9Y47ajUiM+zVblsV/u9lhAoW4XvSPH2zL
Jpk2WikXdM7BZzwhrzXsHAbZSgvaZzmbKC54+2nOAqjocW/fIk6/rkWAyeIvksO8ZyqCNLGUMmId
/h5VE12FpsSdlIfmpoLd+Jgi+2p70dH5ERYkSmxW9YrZjTqz2eXP8VGxFuCgQaJD8x8VGV9qdnii
uIL81FggTDEadgXhf03yQmMFO1YNKJx4CS7NN/UuqPYZUPtCmLKm83A3B4sYGSPrkgFqEzW9OAhk
xQAs/A8OKLAd4414MtEQiTjYiQ85dxYSl1e/l7wXZXCetWHC4cUTYbMU7xiNHYa0LjFtTK4UDW8S
g3HBRlRYLaWliC7Ma7s0z7FMCP35pvKUr+AAmI6ip6tZz0YzGxx+eY9CC16sSS1bqSwkn6WKCJ8u
UM3O2a9PwFWbZUVys11VHTgE9Tg5hHvVvl23JCSldTI1p/XkHYgyNclm7RoTt1F2/NbprIHdapO6
wAjrl99EeHdXoHKnPY69Yv5bBSUOKyyKklCmxF8gqKAaP0a9GAyV6q79mx/bPU5Uy8BLJc/XbGmQ
5VaZqxv7u8APPmpeWSJmsJtlDN0Asxs33qRZtYCEIrg0ih8AQfCI8Kr9uR8Ft5YwzRExGw/3U7H4
hL/jDz8SApb7zLZzI/+02k50bcfCPA0laWhA1sAx9VWMoHbxDWxUN0lp9gJMWzVSQZORztfDXYKk
Wa7JnM+XiunGAnFX+bSoNCWTLIXTUz6zVfDZGNCUQEFidFaEhu+L1gos6A94W67/7HjbYV0DC5a2
N0lGcsHnGSMsGH7EDd1vkYQ2g2Bs60xI1PJ39EgIzJzm+0juUmec0+l2G6hXKaUh0d2QZ4s1wwH6
2Mm4EvdnmGOtXNmYsh0q8sNfAGvwAJEzxDU+NxeZYy5h41J6Xc3cRg8pFPJjj/g+Rk9aSqeYNouP
cjadS4wWKDdwpxJ3Le+kELdu66cin9BTpkZnGBJ8M9thEKA3QJUEk/AjNfo1lHyc4V2v8tEPGbuW
2myG7eRG1fETlnj/4TBJVCb57n6m4ydxAPbr2s6dPtqGjAs1Tcj1VvMe8iOnvM4tYZNJ3ePWX/S1
+AEtNwNvZrDQzacfJrYTn6titB3Og+1Eld9YF1oZIgQNiR0s/Z4zz63oASdZK374hXHfLTM1YboB
kuUsjaHeHdMFCNcJtJIgnOLlH82z+aPHDLF91DJgkVFvY7kD6j/fS8TcjDRX6W0PZ6EEIj0ZIM3o
qVds9sECaNs4ln3BQcrvu5q1Sae06Qu/umohblXAXFyaRI7HDmcblud9l3ea3RHR8/nkOMB44qyX
VrtcLPHGvyyRkogZBZUy9XBM/GuoWX3GkY4GIG7ntYf5btiJIsrmATiBxvwRXaE3Yj30BM9gDxik
7UnUlXULUnER4bTjKUczJJY8v1ETk+RzZ2ZbpS7//hSVg9vUEt2//4K5X/WilCccLGovIzqrRRKJ
PZH+owmwss2qz2JTY2N46vUWKH6Yw1MGNTrWLcidLZY+e00tLo+rYLZlLuFtnlDcP7kKGW2tUeDA
d03TEq13E3yNmLraoUAJKzsYWsxjhwSRtpwG4wuDZ/L5Gkv8/E1P3ONKxviY6ytjgMwUlZxod2BH
9P0fP7Ah6CN2C+HV3dSwUHgRoBBb5VDLIWysiNxqs5VxSMvIHsEgrjH77Wy5/duXLAhrYC+rDF1L
aqwgPuokO4m9/68Db1bSGgnfqpTdyICFiTsDUUy1FoSksFrjwHxrFXnmlwH5z50t4eQLbxgZEGWO
hrzsXM1q94Q4eY/8mbpBE9atKufibp67ThlW3PDr/z5RQ/dKZQamDSiHyBkQ0AnO3IbnfB82Itim
u9gvZrOWsVXEsTztrleJJeixxUdRKcVtlu6punEG3u5i0vsNwS3RaCHf3Y3iSYBLdKnOSmp9S8eQ
u71nOcEVohlRzWG887JeaoRRkwQ+6Xt/1m95shQrOs8Ku9utSStXZJq9ZsqX7csqB7fODDOkU//L
6JH7u2Vlc0ORozv58xP6H2O78MOVVKn1l4nN7SAWMYpp1sX11/xD/QIfgw7c5gFKiwC/QuRFDQOk
2YCSOHGXTgDT8WYK3lbQUxVdKebylakvLuENE3BgY9ZUihEEcnpi+Oe2EXeAtxXZNHkcBkapf9z2
ekal+0miZByJD+MbUDGfUTC6f/klLv1/DpKpYH+psMZhYJ6Z276bCuR98ElvfHlS/G7kJLrEK1wp
FaPVgeuKFceZVNOvs5dk/jyENmHZEIcFkzG2vHTbhfqEldwmX48xHmzzy+P+XNatGqeO/yU+tpiA
QsCSO5tr0SWZXgjIor3bN69AXCexIXagGR9D1WGfuKkxM3EzhjVS9K5cJ1DIKaRBbqdhSJKq/dRS
qxP139VZE0lox6KPHw0AIMqx6rtybRW5OwDTJgmcJ8i8zKma1lETmErfcVkgrDsKOyD81ezkLRCn
BlSiByBhm4zD/2Y8EX2s41b3X97qtGVnHA59QY7tkMnsWAqEpZxkDdi1VuykCHig3Qz6KbHguMLW
m6iYQy6JqeREgLJ30FytHWMfyBNvEErudHWuHsOnKq6DOrCZ4vljq1486nprPVwfSP5vuECMHC80
nx2Slloefq+SJSuLbPpZH9p3f8ZMB9gpaQjM+ezE6l9gUXHhSoxieH2Z85vBnbIXabxfHS9mlUPi
9sGyGGAG7krlTdYdZLQvtLjrC1kbkbJGheLA4o1h3I6RnVD+3mQkx1GgLvxOKpF2Zjxs8YA/FIZ3
Uyqnhyeg9b5f+aHV/pj0DbTvcPG+B/V5UNnGAaXozzgBM8bAJvrFmxgM8BPmHrvxr0LtWhgE1Q+I
sEds8eIuUFGG01IyzoqYlVt08pZErD77gcleyiUl9X9HiXyRdRVBnQtdKRGFLCiK+dXW9O01VWdm
79r/wmnlbEpFCcFYC+Wx1DkM3sRpYwkLJJg3bISNzw/WhnOztkhywZ/sNoeufXNnu1udSk804lpN
Wmwq6cTm3l1s4fFfOkCluOSzm4j1MIQ15rwL9JV32jQsqfh4DuE+7dU2pNPRLEpYMSOWzmxbCx8l
SZEKzmpd8+sEIY3PBYp1Ye+YUXNIiGZwOpSta14jJ35CkvaAAVnhNMrXXsAHgzpRpDBd8ndw5xyW
DDGboPV9cWRccEaRUJY6x1B/4iOycz2ph9Y0Ndqv+JcVONo/AkK3QHwIXshuk24x1cqozMHLcd8Q
qNU88sYZza80a71F122fgzIgd+TiY7a+z+0SoE4NGl1rOPR4w1rEDoO4QHH6y5iRinuTLif1k3Jd
oaTmHMKV9b0Kru5QuukN5O/7DeSc+uljDO0zh8ufUL6XELx7vHmT2dQ01w0ua0Xf9JcDEFY+VUJG
m3HCwwkX8GaAtlNO7x2ZueTnxPYhhjbnURfsRY+ezV+ICw8hGgOXBMlUjc2OAF0HfK6q8FXSw8Vn
w+126fuDDYXgvYg6jtbyBeopFQRe9KaNv1KbBaWSeEvkq1ZctbNa/v5NG5Ms8nT7EWbRuB87ruF3
u/nfTfj/x4ibdAbrqz0QXNO0FmMJCk0uxMJxSQebZ6TML8husM/dBZ1ktuHPyiIlZCe/RWKKpGxE
bwtaENHK+Ys+7ASmvRPLTvdyWJzXHppWlCzxTt7P+NEgvW3wtc+opREiPxoGbVTkV3TycX8CE8R2
iyh+Glj9+41kg/0o6wcoaYxlQY5QMy61NanevmpOPb3OJA96Mi9iA09loQLZMby6V2m6T9LoL5lb
FvF7rClUwKfnnMSBCKYHxXs0oH5MUyiEdqdLqr8ji4PSjzhxrbXi2pAWi8Z2uExmcWADiPDFtG6j
IeFoamPJhBpUA03AKp1fygV2DXdhsVpbewDquGFDYzqRH2RYrW/24Y8oC5N6qSgbdy6zw5Nd8iFL
myd/R/Jm2k47uI2sPC2tlsODewVu2hCjMhahads+qfB14i9ndU8Tyj/j7wK5KhjrVwjexIGQteQl
bEILgub7No4m/j+Vpd7dGvbfLnkrnHy3NHLvbhHxa4z0mykgypqutAvchzmaUUsLDISET9cehTtp
09aXdX66TSIAD+qpU1qmUZTJU37PBfc+yVhD7YbvbKtUhWqEDpd0WkhvKDACYaVQ7Z1JkqW3HwEV
IvueBib22e64WTTocFS2YRH6mPJu3byXBv9xF9YbfdA9G+MPxmIk7w19zqgBzzl/jiEmrDmKdOHP
2WRL4f/kFX6InyyCWuEWI9/6AD1x7w8JF4H3HUc9Q7U1ULAyCaQqpimFmvSZPOHNv9meXCKpruJU
YRYairZHRYgwwDir+k7Hi8Qspn6Gy1/6gkKJjX6k/Yh7g7Bs7qj5aJW0tv2ydB+cSk0pn1X9DMaq
CP3e04x4gDDlOgGvBLYtdORfwVPdl9RMY0qk9H90r5CKKvUWufhHdaAsTIHwucR+BqK/Xy42TNgu
XUSXy9r+NnQcw78e41mi1Z9FcKQhdOuPP84y2F3agT1I215FdTFn84+RtYQS7l5ngEmRC7sxpwpY
P34ZtD4ifxD6glA5Vxom0UwQdkXsJfCIvyhOm74DVliodktpknWQdXFsJGRnv2hKyRHk/f8BWzRp
IcAWQolCpn9KhQ385PVHKZfpBfq0zmvn6jVXSe0Az5eYwZ9K3T566QQKZ102nDh4OABE1Q3RN7EM
nsL3+tvmgQSAom/4nx1jFOV+syijusMLhubIfjErVpvJ9+gvHTveR95wLaruaq+S7iOx0JG8EiTA
4Sm6s5nds50A8vMizQOzYQt8tKIKqsf8vYjazlWrgaZf817vQ0WSBzphbyRhBVa281MTbpSJYoZ5
aJ1g2dmj8swFP8oQDRPHXay//XAplQvDArx59TKLTRvxREwenyInbXxzhIW+izUWkroRSROjZw9g
HqWFGrAw31k0irnFjF1oX0r5JwxAcvRpBxrCXfGzFZqC+P3AMggZbxg/8wmtH3AHP94C/BYQ+XQY
cevy8g7RLq7scZof673GxYwf8509FigqqRsQSAsnssl9gLjY5qtNecvCd2QS37i6xOpmLiMRYeNv
5pfuoCLL1xI30EY9uciE9Sd7Ti/+CDaxZs0EwlB+0ETlOL50AelI4peU2VrvNtw8w6Yvy2dzEUMU
NkLddC3MWIp/PKeMlEBio48VaZrjFfQRM6AfVE4RRDmqw9yBLQEVrub+FrJmhK/655h1wfpL9INi
sTyGdngMMuYB+vcPWpzXYOoDeP0oM8UjmeCmF2KwLrg/bpxVouY2+cPZwQ6eUej8DqWOaVkBSB48
un3FNu0Z56XQ2EOH+V8/FQtiDNVFOpqgrQZeu6Ow5r8Lw4UTx9/L3DfPFw+4VxOPnWqzVDx5eCyt
vDsHf6jJGWTxU/BOV96CUJ0uyWWBUf13dHDjliMX9t/rYaOKpyCoxTSEmTAaAH1N1AKLSfq7aVYi
X0dpq0piLA7sMQZDARzj6jK0c62aHy4NIb53LT+mhLK0Hf58KC8l+3CygB3HJlm8fSTqH5fXgHKo
d/qeiz2JfEw6d5TfQntMvkObxwr0KNZzj7sPYTzhuqaYlOUoWifZlSYaeKrfbp1/CxZVHt2B3ajx
48Vw+31y8ZUJQP7NntJ1yoHHclg36T64gJRA+6VzQdoqY1ebnkhm9a09XTZyA4H9M/MnVSC+ypdU
s2dGmG65boXn/lcVyl/RlfVdHkfpaSFg3a/v4vOuRN9jQuCxi3MHhtZArE5BfGcV3igbb5F16oNq
+ST98CZgrjWllhx9qdrziQTaYejVlyCpSmueAkXq+34YRJBYWLrsA13w2uP7FXUPmE/8+hS15k/7
AsCOKlAS6otX8ofuJ7TPEgpJGzy9QZuR8O/zIPzWS9N0o2bCjM59a+i6Z6361ssIIxqYtKKA68FZ
D/h42c6lNYw75VS9ktQxSJMWJgDgxYP/8Cem+XLE+MAZxpfzmiaSt6kyGehuGmdd7HUsHsxH+5Ge
XEFBbLbIjYmMvdd8Jank8pQsOIe9uxgfZvTJyGZKZ8zX8zPFOF+d5I4gRnEnyJoi6f6IEBusHH4A
L9eCCVPFh+6kQEGOnYGC07HLXdHcB6wU8AVE7iZB4m2nfQUfv1PyIbPGS94NjxDovnfSoDsnrxgz
XOmh5ZWF/101RuTz7mt7QPlCoJVyRwBQ7ktKHS9jJmFOmI/EhUZPTQo9tqm1hjt1Pwfq/34Qv7wZ
evGa4RdtQJgAw9UANZMNrLXLeeTb0p95DAhoXU+x2ZUbwQYc5Zwd2VCxV6meAtr6Utapr9g961zd
wHY6bZR/fJ4h71P3Z4e/3k96lLkaMSDqBRVfEcGGeJCydOTtTNK3FY6sxBuOUFx4WGrjjCgZoaqG
PdxgJuplmOHurgV1HDUGDSO74E7cBCBWBOT2k7BcisxbrSlX68HQPrmNmTgZHsnPkBBG6/+fTMD5
8Hu27Shjd075re99BWD9O4VXPajjnh4sOyGJNW/JlaHIQ4j7/ibve7qw+HULYFoOR66BK0OR7FUR
faSuQrDJ9so3U58dTX6BpVqGRms6zrQg+ZcXq2nUdYAxxVYkmIal9sKWqXPG/abJFuiXGGlkyzXE
k2p7J0dA/W3jYoaxnRXm8yhC+Q9f3SIYdjP6wris+UjMXMpXzVA3X3nRH4vS2UdvBHvsgo3hWXh5
RyT92HxVVb2AFVxrcWaonCExPBVa5+x82ei6fQTG5nlQxFfBdE/xmCYzxS2VbI/GHWLi3N9u9fsW
0WokNx/3UMEMXoW0e2vB4pYOvt1W9dH5zAhWOIrhKyU+NdWhuAsbCaLQsLSxpTfKeVkeBeYkZzs5
zlDDWabLYfaUH7YR1v3uOu3mvFAwuPv9orxepOK3twmZnI5I0o9JFjkjuftH6b6n/3GOYQ+8KI/a
oioPjQFLbVHiGiWNmSx6iSiS84cVWDGAxAuslbQ8JwbrO4vEOkUhNTyAQu4ljsSvy066YXCUCMag
XATSvVI2Fb6MAs8aoQXe6wu20zLd+LzcQ8Te3tGjhZMMCkCDo5nbKipEyMn9GiIO0BFWkumv6Sko
8LQaZARKadyCEPC4a6B6PEg9kwHbRg977gC6jKpP3usc8CFXj/MwIMA5ecXnRps5ZrO9nIotiBpO
rQGEUWmn/LQKp4MmAY9SkAeFNP3jyrK3VB1ZB8HRyS3ZTj3ggic2DsE17j5xBEDwHV7JmcdDdZaz
IAp0RQEYCSX8tEygMB66tAfkbxd8c+uvzk5Xh5Z6eK+Lr36e8xKGxhinjSBVvo5NpDDHp7Fx5XR9
AurKh/A7TSA4pAcCorHA55cA/GrDBsEqYhdClxRkHoKDAfR9PKFrzpWC6zWfIBPSBRG+KY0YVynv
yKo4a37hYnlU/XBOyJld33zp46/KSLzWWt7jL+l28dmF6Fm0slxpPlNH5PBhhNWQBT+dQcJPTan1
v4fJg9HSkeqgrJIwmyAYnd+FIp86jx4vDNGRvnBMr/ZTnnMNH08vOBfuhDk5BKK0r54R4/9oGnJM
J5GpMV/LP8WATw2QxzKIx1aP+8ktqD6BSj6uRy+QqrCEeP3xzag2UL7FBvc8c7iNWmmR3oX6mgnu
ZEVWj0Nqd366PJUEb1ViGyFW3wZk/r3PfwjfYdXYiXPtXuuzW9yyQ0MWnEpUylQ0KFhvyQ2buwqV
FQQ7vN7q75a1KhKXZYltoag1bjhhaF6hiS63SzHnL2oFNFeGbj8wTHlfggg7QBx+LrXQxLtI8zkf
DYPmjylMmQrWxnii2By0KHSBGhVCHCJaX7X4C+RvAk3TYH6Kkt/6e8+qyfSlSny8AzKzokebbZ8m
iMjNNgJ4TuQUzv0fOriWQnSoYY6d/jYvtsM/KS8BYqwsdnwCAUlUsgZyUVorpRHSmG3iwbR+/DZB
FX7VBNccQgRxYUldgi2BPfdFjRlI7AZ3CbVaB8cnlwebiAY2w/Td410qV1RUeogY5inFJik1fCUW
cCTLGY3U9dAcU+Q/g2M4oiMHneXlkdRykXthw/qKbYEtz8sj0xjVCsREn0q+Jau+3BRIK1FIxUhO
9D5jfgP4GOeIU6c9ePFNhi9+RhAGEz9BS0LLWrGMBuWFfd9Ri75nYAWLC/18cXwYYYLgIkL8youd
B9RdiEJ3DuSP3I6x7v6dhvzr+S2HSji8r4ChiSDoxcl2ktHcGh9/FRylPpIP7ADdGpbZOrG79/a1
MW/Gu40ASWkTxFQbON8NxCK50WNdtd9qUkv86xicrAOcmLBKdzu0grqst8xTiyrl0fCICDKcnkI+
Rfbh/VzwEX95ER+j2ACNh1WPTfbvvFE/J9zJH51/YyZhUY6PpCH8a3qEn2aKfjtzQdBWG3AaJB+m
87yoMJzXO/3WYQHrIZumie1E8CQ8Nc87uKtB6ynFhLyqEH0f3jOAxng5HPJGKSIpKzRolUw3Yh7F
H0TxTZOxlU1O2a1JSoUS4dTeGWdkSThNf1ivM3vjOmZVf1JWacdqRLfHIZX6KWIL+XlnGus9mqBY
NnROLHULfnmpZ8Q4x0RUQdIsnhKdML/ilG4sc9mc+y1EqKP0oImYSDWAQe+Q9wPkKrUJvaGTjy4h
DwBHfpGXWdVSKQMrlZ7SRs7OZ2HVbEE0X8wU1XOISLELN/fqIBuegaBBq/kcsozAHa5N5WpAwQbm
llfOgXxs3x/6gBbsb0nC7Br08PoTeOI/bjAGEyVTZC/ketdbC6S42iGc14+i3+0OyFBetFLy3KKv
Em4hxcTE38SBIakkPxdNEnKHYR4PpNbMpop3ncvXtJWbt4OFPGEwqc9MYYstFEV8J09WAKA6ceBw
BmolCF910ipvhoWV7LiwEOFuaqYaSMCp/NsWOIFd/LJTx1mIF+1wADSDKkwg8y4UO+fVBzbRHbBu
zALPwzqeo1a4zoMpBWY3SCaorTcRauDsICtSdsc8GuZkUGkLKVHfjggJ8+POme8PDIDrlKPVSU4n
sESdFlNIklbvREBLA+wDBpnencOHp8L/JRGWkmWvfMnUpjqr+1dSUxpY6a5TkCgGKyOVgNiUG2Tj
Vq3e5orPrAa9oTEofaFMiDy4qZK5mJjxJCmFADLulVJnvDoGhCON/jtwpSN6eWofS14jkYeUL9fs
VBPshUNIpuiFVOTAXRhCYTo4rxim4I/Ya5KDmmaXnQhJkcxIfPmtNu1qd7C0sb1Aq868rh4/BbXA
CJyoSv8ovK8MDk/u45271KxeA+s9zYxLHsnJiZfNi+06ojVXp2evriiCnF2sRAChNklDAT9gDjHw
AvatvkjdoRPUCcD+W0pStuAC6oV6WG1hFIiPZ2Wu4ZHVFfF+DprUE4AcPPDRSLGVr/umKv20weZM
pXrUpnHbkW2oMMVJWiRGj8A61Z7EEixnvcYM8Xnh6gsEDRA5pV0TACsirYl8UMJSfPxbPpADYcDO
bAh4VmJ1IN8t6Z2iAAWsQ6fjn3t77W3kXsH/lvnATmpsmWqeK6HM48y2TcyAGrs7Jfsfsv1trLOZ
XgoNXRloS3Y97PecBX38Yrl/ql0X5/JiSMKI+bPOe1c+Zy+TpGk3uzlnu7zzvG6R2RfWBzlpz1YL
GQh/OQQstubgLGS3sx+W/bqYlWWUXbhnWE6K4fwRrMGWqoHvLPfreTgp+CjY/MS0+e7Yvt85hcd7
X+M6QsmeB/xJB7hhQAub8hF4UtiR37/j6Cx3b0cBOK0jV/EijzHp1qrD6gBQjXZjOBy7GvzrCWRD
Cdg+4np8molcNS0rGTXcWjJ6Qd0D2HYtVl3rv9U+pSZmrHZF+TwDusJirMU2x5z42ZnI5C9R7/O0
8xLNExPshscuQ2CTUZ1sJTPGd/EcyCby5AgdQlu4m+bQkeNggEWvkT4cVz5tgbr8CGMiqAaxeX/l
HqJ9SA/y7VemvocNXm3aic3zbjEs7va07OJzHHl/8gVeVIJylh6dvc4ztpSTBs2WpNi+7GMs+3nq
5RTbtU6xyLyYBRcRdw7SQWAVtCvYqonkJsjkEU1Lrfa6YPAs/uQ9TUZpwE/bPBrXU8MWm12oVet0
w4AOgpv7o/34GxyoSkQydTZ+9sVi3tWYPsSo0u7GPtSx2yWYaCLdvrM00UN0t1qPxDGMUHFsBVqQ
LxQQ0q/jzkhzc2e7KBVqe2B2MwSiMuYLRYlikyxqoX+Lh44D33/RTA9zAhINlYbVVa5Ico8OCk5Q
1BglMZiIYsrSbU6zsj8RNQmgiLwtPwyG2ade+HBmCZHuCN9ODCXvSLTooq3hEElQLy+5by94xGK9
KKppu2C5PHQ356RlILqvK+NzwJtDvXysMFw6iFCBWDQ9lm52z3GNQpcaRFP8ykMof+nH/G7jmefa
pHy+WdfPQirXVBBs3qYq6m8nE+XNSmY0izyHgMoRw+SU6YTPsH7ZzDZMtda3bwntaeK4sVw0glgV
QjkKO5xquDtSxeJBvNw++bo5PFFA8yhVkD88yeh3Dnlt3rx75RRaSt3hMYv0QSqSqnf+cvzu8ryy
eHQ4+Cjn6W2yUKorFNTGj9akwBhxduxAxvg1z/UHV5MC/5/cAyEkkk247cazXAgPAcFQcY3gFDrw
5UcFXPw9wh7LjJ6og7nTttTFOhEJpI0wQpLsy2OG2MIP8GPS8SowvOSI57bLR7s8bl+jCGE/WHrl
T19ufCbGA3SUSVHTa/qI4eIXhfcU5qEIXR3YGlHLTgD+n6c9sBjEl5GizQacVO6mIzlt8VWaPDqv
+UahGjgIIGv/CNl5ATQOBibZ9n9CghTdEUlgh13RzTpNuYqo1lLf6IuQKsHrRiMeewYAeCqNZiQi
MeibL05f9uzB8FoGNRZzccSwQ4KlS4UCwdR6TyEIdvrFFy8Cu/5ZVjaw3E4wRfWW8aoGgzx8ELfP
iHs4OYSyt6hpguxNFc3UHBnEytp9oQBVA37hE7qtQrRvJzr8HyDV8wypAz9VxWi+5AKy83RvLK46
1YVNlgrFexuVSjjl0/Lrm3hsXRtqmcaSv5V97A0K081GQWGWYJUfiUN04sqbn2lb8G6EZtwUtnxd
dwOgNMdF8Ef108EEuEfw7OaUe44yXR/elpbZ6bkziAt9TvPU6g0yF6hRILoPgl7uPh4St8c+E4Wr
8o8UgO3zxR7BaR+UVDOObKZEKFOp2MAeDkwvsXZmzCS4JccaC6tdU0qiL2Om5RG9Q9PFcgpYtM8P
/a9ZmJ2+nIwXuq+CDt/+gBmCjycZQPdXemuxRyOvbs+xE/sd8sLeP0I9xM+xShVZUWO4wFPhj2VI
iYfLq1yufgM+hNbSWT0L4PqcZEt2yroEuCwUzL61NZ11Mz6Bv6DZEaYyC7oXPqknTbZesCxVROdW
tHJSY0cm086XxGFvFgpHccyrciCuykspJ4oCNk198C/x5w8L2i1xqxBRCpcle+rEBdL5+d4KhT6V
g/F2GZS+JZv3awL803r65uOZHnBVFHOZ/em/0A8Njy0Ix8SoN8FQ6BDH5cVR6+4U8xL6ZAoBMOKI
JsWeskKd7mCdphHGgs8Rj8fOvT/8vbME79bUHPHwC1Tqbrd2MjfKy/Vg9/wU1qvTXf1t1H+lWSRd
Gw9xe8ypSTkDfQe6tR8nscVLLN/o5eP/+TakgjSu/Lhx2bXuU4Ei5USimb0YwCRD/ZTMjgrA1rN7
AEfp9Dcd+bXpSth8m8cHCaCakQJVGBylmmoNu2Ch3kWwalUKe9kOdT2xRjc+GVbOyVaWSYCKHPPh
HR5/KPOMNJNkXUs64Wopd7MQyfeOBxeIVvurNFHTNb2vf7lo439bALwk2e85snz56eYKg+Y8ds++
/gi0ePThEMwmCnHMQY7TMFkeypJ5Fn/wiT3m9rD2ufqtwYbPUVXMBNPKZVqxC0Vumx8LYkP/WF+Q
S+iU41y1/t4mXb5Rqm7s/mdXz9y5ZsXRNr2cSnBah346rDYWc7CjdHG+uu5ifLNuThO/QJAJiVcd
4WTypHn7cqgqv78eWz5yWxes3Qv/chYMkALHDjZ07wqy4LiYq4iJ+Q5PLGKquRAXxl9FimiEQt4C
ERmlCmp4h9601Jqcn/w/pHHDscgISrkXJujYqEMFNJwluWUmb/bKdPeWv+5Eg+2V44IneEgxw44/
Q/AThrmrdCwgX78UPXttShLO+zzJmbpcUXMpviV3rR20NrAsnKLhkVFgN2y8Hmd9ZG2E/cLehhI8
hdUbXCF4yMLYy5+hABuZNzcr2JTKe+JXmlnKt0+dWWyvJafOnhX4Pn9uw8RqfeD6QuwXPL+x13Pl
voDEnF/jSgWzzeqeeiOSMscJ3rqBEbib5KO0epaZS9IgLIwJ/nbphOR8nsGDR8NnUEtC3Z3riDnK
CMoViE7ET84pbdKEJtCV4HaRM4N133ext0VvZg4teHvT74DOPiit7L8zVS2ncC3PlonmzqR9/SxU
U69z03irJ85em+4PMaR2D00DHKTboHahav/Nc4670o7sjqAmylhsWNXdr17wV01jwmECv8qm30bM
b7GTVrpqWCcZp7COMC5TgtZAofYF6MnZUEIFaa1gvBK+DhNMuYbUfrSwyPB56sqq7gnXQVyySO8g
nT0nrHwYom1lm722CEPiVt/zcR4Qv1rco9xgokNuYM/WSAqoW2WandPTGSRhUa1aKd3TDVMTimwP
/fXyds85/UfJ8jlPYFXeNGyR3d4AFAUNXZOKJf3Xcw5OYuRF3PCxSBcygDCl8LusqxAfKBJ1vD8c
vyvuS5v0OdRg3C8VDs9CldQQMTtJMuxzUNQ3vBQpMBIBW3ubBFX+zULXDziaLaU9kFlPCFvwotNo
+J92ZyhxMKySfbLrKQTOJ1hkzQqxH4VVZD1j/CbuW0yzeaUq6J1tWr1yo9OrsSkMreuJi1YWIi9+
MUclGLxblmwnBVvDdK6Qa/vd+8YNJVY9ZwFDgjlmCKKqiJrOXrf3IUdw+ACKCqz6ic9nrdfoGZkt
KcaHRkAsSzfBuTf/jQPlW+WroEFq6SZJKBqAJ++x3XlckZzDpJhzhGbVwlPScK0wOYbqiEJylPhI
LpCq1gEruvIoiF6vbvI8Sk0XR3PU04tQsrZqESQB+iI7NMyXn+TwlAf3w2duhuK7osv3/JO0XDVK
J8MsWphBRQkYGz2mhFrX0CYJdm/o9yN5/I6Y8ASHTbWSiNI/RmSw6RkEOJTNEPWMFKYmjvGGnx8G
gYB1iBqKE7YgooFsSDa6G9L8R9upzx/KG98dpUleAVWE9xli8MS/lM5LPGKg/WKnsC0Yc1ddnoTG
9aC5OCxXhob9pZKkWfIw7StKQGYbQf8IyAr8hj73/TeyevsIkJI/dTsvajDCMHk7DdrJRidrVYuZ
z73Xj/AzxDtpxhMUqsj0h9Q+80+5UVH0BrKtN1dMH77vQcmlr16Og7WVvbLFr3IerECtFoFLXb2B
Gq1ZffoGGa5qB1+VZKiiOsNXliq2wRd0iWaJngWf7xFi6JNxYmc9pwbtyTVMnIAuNBYI+LNJQ+Yv
6+U6+03IlaOV2NYC7TmP2Z+jEP/e8bPf1aHx4zEfILtskSkOh3cPIE3QsxOmkYr7Dng1ZIPs7hHF
JZJJdqpgYGIQMIfDB17r92tI8CvHi2Wtq8D1sfJzxGvqH+CCcVWmNSnSGkBVj483jKKuuFx0717d
asZnnhRh56Uf5N3uitOIZ/T9KvO56SlDQ7/f0YGXHYHMJSwxkDmp0cqFh38T7bwS7KIJlDt+BTLS
3vXbGC6A1YDOsJiiQ7ATIIg01u3XI991/RR25mxHgtOFDZNvTB0W9Aih8DiPmAXYPC+m8UxQNFp7
J+qUVupMSPG58jggUEa/9oiO3sPpe/kCnN72+Q8zc0Wwk0eUrW4uPk8I2WhNGQ4kb8MHOiVgZoF2
yGFQepUrtUm2Yj/dwsNKyWfawcVuFZATT2Lk1kNj0GQBqHiggvc6N5UcxyUE//fDii1rFtCsjaFS
pOBHV1SuJoR8CZpexp9Dsakx6iaCjY3Ztcs7RqVmL34oUfnfGh/+pc+kSzXdgetufnQ+WhceFShm
uC23YDGs3zd6h89SHPVkpqP/8L/wb66ZpC5dYZdJOhREtiE0G2UJUnoOKPOpL/RXRrN1SFE7g5Qf
WVrUl7ophjD0M1bclAlOgv1miIozaolQYVqpRKLK0HF9ipsEmZJHmUqEoWySjY4LEPXil2C6a5kY
YrOdAt4U3VwtHUXHs9NLciNfXyit2KG2qO3kr2vja27L/KgOYY5IKqkvngbkSY+0BlrTx6fCba0V
76xZaf0ly8BiFFk4S1Ag4ZirBuV6FGe+giz47DmG4sBXdWYsVScrCaxZ7P7Go/GQ39wqAHINlpnU
oZcTlPrNAMgcEal+3p0wWLecxzyut6v7OjsCa74aGZZRnivXrEIO86AtMnNymbNAZiLYaWiwfNu0
QG43SHnaVUWNjP1dPseJRmInpBOuizzAzzWiPR3s8K4JqoAma5V/KVE4RWmXkJ0xly1YsOCJNfFg
Yq0FzmAEs2dibdyO0iz483i1hTjNLNMi8BCUzXBmIqqXX16EuXp8TjfLtZJCQU5einx7uk9oHo3Z
d2qyGauAI8HzvuG2RPh9MBJZn0lub/z/Sm2ARxdX7NU8OGmtc07zUuzVUjTZc90Q7IxkRkftzrmf
In5uxqNpHf9afy3FIfEH40OrcDz0aB9geeGPUUhMq/2nKm+wK+mrFaqAZ44/ZbzL6A0uAK9kBVUi
JrIq0GHgKKfRzl9YxmXODyO69S1wy5iuMk4QR7BbMUlZwilQ4RHo69pAhgu4T+C0NUI0/pYv51NQ
zJftqi7np3bq9REdYMtyvBCZYRN5vdwgqH5mloLYRi58ikHc+j9TTdUaXBo4u6iUY5DHG7QJUf2R
Ksw1Js3gzYSliqiL4Br+/QIk/IIKtY3IP5bPODOP4SvtXVZ8bv12Bglir5DfaU+ZWptw61rml59E
6auQ8dBcmSZ5dXlm4qLbWqmAEGm/g2JbIVLrKHg9CJckSBC5vsV3to35rVdf0KySqxBbbjra5+3l
Uck5snNEkTercappRF1eccJKAeAAVVpG1rQzYt6hvPvDU9Sc9fU8mxEjA1LRCEp9g8cIK0j0MSgO
cIsNXg8b9HZ4/q79+fitnab08wMXnRC87x+McBn/Mp0uhMHqo0SZJrBQXoQPodaYrcuKqqhUeprB
K8kA3DhUZoDKvWesojTmrR6xfOM5jAVTmWv2K6cHT4L2c+eXMbjwZ5LELDTPnrh60aM4J5M1y/S3
5VXT3yq+d9RaEbmFGAGqXGEuAqHCV4SqZSsPr+BEHpm0MMjDe9JWE+MlbKjskngM/V19f4BtaAOT
OKA0dJ7BxTrVlY3PRxS+SVy99UdTKO+uBY051cDPw5T/IMuNpDiQzCJIAxzkieATRxa90hlh3ioo
TTwyRil7T7H2thFPxFWOZOCoAcDmDMDcZ7fytzzhnzvsnrYDS8jWPiPrW+yoEw8qWEoenhPpsS86
8wv54L259yxWXVtrNgPOGm+pORx9CCl0QV/unDHgpboocT49/IruMgruSNqxVzP8xoPtoNB0BEPT
ekMmktt3RYEOqHF8qF1TIfSB4wUrQPULndUUocE2y8As1E1282soLboSExrVd7U3uaz6SJvbW6M1
QIg0ZmMzhbIyJ5RSoK2Rcvp3C5iXKxMMHlyptW29OgANxmy/xfazAFFFd8awCV9RbO94rubN2kSH
u9R9gLvSTLWaVFOK9dKDX1lLfCpHGQCxDjejd99weLrSFsmhw7/UxfeaoxV5mn0zs4tvB4Bg8sRS
IPsPNw+vR5RoUZIztjk/x0unJloX3O/zDS1qcoX4FEAmF9AO5c1kENaWHKBxwjTcaZuxZIpPGEx9
0zPAF6L97AG9I+agnFVXSyNKFJOxx4axjWnMB24x0sODNjTnOVRb20WEK1XJ9iu5Hh02V3wVIyqf
QBIcpliuaUXK5qioM+Do5ckdKD1zK6DRFraZ+Jl4jA3QtS7WjHqzE+W5GACeTpP26skuUxy4RwHA
GtK0C1Fhl6R8vC0dGgvhj9GVfAGih+ZgeOa8iXPNBtElak9wm0Ov88/CRlpvejSzeds/lWuQGdbp
ukL0dGyOGxjDW+XsE8kOkp7d6KpH66Pg3mTYNcF9wkGP9Ejl8r9n4r6RsgWJtUj7pw3alMNKuMuj
DAK8OgeNmvRaByGJcLMjw30VmNfNDXAYku/Dp24fuEsZ6opdoc9o5Mw6iql0bdodqj+KELSn94GG
HPTxVgyTS+OVzYDLblXE90Yi/UPgDSXDgMwoERQlwgi+liNNFeP+PHI19isWRNgZtt5u8R2Wk6CP
3wEZYMqxj1agTXZzIInDbMYxR+Rvn0m2cFCzxgEBUJm7vnhoR/aCuiKK/D5PFLs2ieJFUcdRBsXF
EE/ZQGFrKWsgithIfkARdX4cKZfamStQnkocMeAUzdw8cyZVuxF34doQ5JO2jLd0rWDSKMxkjMLS
Xu0x7Mn9FqkohuSaArZoly3gvBHkh32n/qkk1/6CwSd1mg0zv+Lw4JZbMXC0hgvhLqSX7CMhkzpU
TuYAgbxwafcerjmwRQ4m2mFK8XQVGMrD6fExe9IN+v5KhEPXqQx4d5bWckEEVZd8TGOBfRvANpuu
sRN9yuODyY98nl1vUBhgISiF5BdJfoUX3l0fna8BbSQDUAVlrzjN5kFMCD3ikpvWkzqj8Fy3TC9T
qewIFVCM54JgRO8tbFTNP5MKYhA8l0t2pR+e6ObS16uKsUqtVmu8/gvRdm87F0YKHXdAVai2VwIi
OOo1R1memxOflDvslua+cFLk93wEpHnGR/g7V+DPUd+LSAnsJlV+B/r1iLUrGXmmaqfoZ8Cicqkr
DZ7yYfSng1j959udd4AFUzLxBFDMwPgbI7duwmB3NOBjTOknbQgYIg9UjbTC/jLOLg6pAjdO3z4e
FPNNAQv2YuTmG3gRwuwaYibPCQJN0Kar6al3+MBmV+zIXfJxanJkWJhFq1dn6I80sdMikIZa7LWw
KxEBt4hA4e024Xn8k2KpZci97hbutCE4xt6pzcLzVLm+0Fr3zdEsZuF0MgZslknP8dvzHMQdJDi5
8GU/mC0aR0ZUjpYgxRSYNrxg+Ky3ztlkFhWO35siNYGu5yf4r6bawH9wLPJToveMfBwcraFymNEQ
y+Mdm4Pr+XSARVgPuBcECF4dbxzn4RhlpGBuBAwf3LakLiYFAL1Ds7nR1vmbWkKRjjJetWexP+S3
WAjc+DNeMLWSFpqUkOIc43luNqWrGf/oZblZgpT3cF2fZB0p7SIswTtgbj9/NIlztVXpuNiewu92
ymSjlm+t/EUKiq05xkGGN3IlhKkFxrcFpF9FIt5pmgVM2pyHuMvup0qxF+MZ6iCZwcF6PN8ZOOl8
7DFoYyiAAfHkm+vGSFPmQE/aW6mRPtznaiWQB4z+5koJOHIUvncj1ZYryh75UQe73FQB+XcHd5SR
HgXYF6Z4z5CKZM32PZi9njE+jRsVxj3jfYas6Q76sgjGaxUhDf38QP4QMnPpF9UvFiXMcmvgzE0l
xZ43BiKYNNC5PCFPKpEkWbo0f4brfjb6GXrQULbMBleyViFHHcUsD50CT5o8DN0xDY1y7/MeZByg
IbKSCBvEpNRiz68OrPEysyQaNaTuFyeiDINuyvSOgyQsspV8MFRwSUQo98iE1Ex/ONqt9J1QJCda
vz9czlyyPblS6yS9428j0SIrBgq2sMGi0SrlxlWqwznLE6wDagw0zHn5lindh2/u/hoKOHY4BeSU
OuK9JfCdgGGzUipNoo2me3VeZqySB3flzeqGEQGgyK7ev5HKnueJQcgDeEHQeQh17QZn3km9hIva
g808ItIE1RhQsRTXxoLgTBmVrYzHHbJhpingqxElLnW7QZCJICIN2d0pN979qYYHOcVPSME4Ptzr
Hcr0nHdARTy9nsYXM7Pd1YjMVuI4MuQMnKMt2FpuMK3R+0/6EcFX7Lc9IZ+Nm8qSQH0TLJCMeXy/
+wuQB5fCGJ48xGsGwlOO6EU5YsiMjea+EFa1lQVAIBRjPHS0Hc7q6pfQvUexyCrCdgUR61pBACj4
dpNX8r0N3cVM1ZJDjR2Z+e7XQ1KR8aF+r0DMeQ9ZmgSyXmz6IjRDypWJPSYKDnihJoQNiVgdXL2P
hykORlj/YnY0QCE6xpLi7cBgJClkIOOnK4gjhLKaXP19kN08JB3BC9g7jJmw5s/Fh0otIuMIaRWN
Ys7gJFV9xV2XneFYT8yngRrTFfphYVr97HINFGSU3/Cyq/Yb/1ZyQG5Zd6/Ykt4Ti1WFEhRj+rH4
J1C4w7qkacB+iS8LEUCtghVZ3wDLxvBKADTQJA1CrW+YyZWbE8F8Bc8DAJTx2JxN8ETewFhV0zvQ
xWaH5ttJC8tuZX82rCpBcNyEqRYUaSgvpIgL4WPrazWXkicyGtgfRtR9xgqnLFH8fPhB+IaMeUSN
dq8FhqQ9DLGUab8OrOG/o28LxVBbHRtt44aYBh1gQetwRfsTPs70XhBzdvbADVy8LDTQTIlzKuQ1
ofZob2P0re8TZUG6f3pUB6c5Eay6LR5fYm17Fl18N96Q0AIr5V+lfK0kPc2nVWiMSt9SNgcw8CxM
ffa60mZE6KN5VdWWLDk9QbnZYaPc3wq9yveeY3hojBB9VezDiqHefXa9s4i1wxjbdsYCjMh9P9VS
0hT/P5SShlRYww2OXDKsf+wqfnuvDfrkZmQxuJ6/wcwYJyEK1LWulK4pAqDRB35wF15d5lNvItZi
geseNRgQoUSiK09mOykIW2D/gQo5EfpapI29HfRH1MMGafs4izaGHiKSelbBZYV5AbnKvui7DFVM
2B3zPEPKVDteXj2305QoH9JgxT63244RbU1BM7nsAp5wtOfBOZo3FNlZQF6Q5qXgxSdlaQOsA4qe
GLtlQBfN1DKX0m3wxx168hLBbfC69ZjHAYWPrW+hl4sAyBKCt+BymyxYvnzejOk0uajVKa+hZW49
BYOz4KhZzQ5QWPNwhF9X7zVnKIzzeWjuuihK8/rRnDXS6zniBn9rQc0HTwOoJt69X7V0yvoe7xPY
vuH89ZfkzYkp/lLRsIf15qxQU6ziwAQM91UzSOaSBPWs+G9xd8H4LhLoV6IdLQcaRPuV1wFc9f+p
QPUnaM3UYwKlODM+yq07qu+q5SWHL6jObPuKavPDvtcJ/EUNQ+UzOeNNKcrF0ww/LZFWFHEV4Abq
Ug3rd+9kDJbpktQvVChTG3zgvF2+SolBLnUxHCfLkaVlpPMTbCPiUYx4ijVx5QPq8ah6x/4fivsM
PnUdZCo2c/WuOhrj8yX+cIihfy0gpomOHdXYPu1Qejut3IssV0H2QZxDzs4AaTEi9OtnGV7KGCqY
TZmgzhXEbU0DwxrlJSJdNCnc5KdYDJkC2mJKdjIqW/RoMiRh3BauXMhcR5pygNEeBHsnYXAMso/j
jnVNN7bvarcR5Td1QzMAtRfvdrrEkUd5iUI/tzxSWDvPUmSkD/t3fvsICX6DL5Jm1SSw2roHtrrX
hWOsXYqiiHC4TYjmbaR+p4P/xzGSfjOzwvcixsIK8DxeYlmmJITyUhSC/sWxf22kuSyjFZgtijdy
InDoGvTf2x+GQwShHOTefptlfL1/CWJ9ljnFKcBCbwsFz6KA6DOxFdBdABI6B7OJqonYB10ph9ya
nXsGLCUO04DcAa4nnIYEsV7GY1H4r6YsqTlBKKiYCqmVgOCtLRC+rUZjG6WhSDDmkWHwO3ZNc3CM
dZWELvLl/4IwGM4zRfD7cW4zRGF+J16KtCbswnIuhms58//gYVibMlj+PoxDs4DvotwKUx/1l666
XP6RAZPmZTBN1Mtd6gkof0YahI+/CgE0lYSQf9j2cvAyh12r0+/aEo95z+tAlt7qnMLrAd8bbDro
mtDi6gyXBv4SKhVlBmbimOa4Qm/e6A9f8zcNxt9YEtr0LjJQnezxd5mNkbvpafMoBBQtzaqMKGMw
uIF2vABGPiNy1uoEiu/ZMElv/SVC8GFIFdgAmeGHYrRimSurJnKYsGXJerutEgOeuCmvRM0rXavj
mTo9rLeD3fUlPFli3+ywsY8mBK1PY4muYywS1clNv9OJiIUczODXdWIToA39V8y3FbUCTcwgpEuk
/3uCD+yc3Nev+zCDuXsLRi/JoPJ7k2QJmfY5I3i9mjldi7kX8f5nJosHnijt5NAFBzcsl5L2f02J
MCF64Ujh65lYc+0SpGAudtBRVrjJGXSye4vVDdEbY5gEzWVfPBOqQ/gy2TxH93pA6ouFsabiqB41
KIOw/zMCwyTY/Y/uLuOHM0Kt2A1VcE2hb2vyMwMiicGTCx8CMj15AS/Qi8ZPPgxcLHgyWZVs9b8I
GjJ3Z07ml/pf55WxSDK8KGFC+SX++mRWrJ8GgwVto9sAQf0eYgptsfGFT0o32AerBb2w/tRZAxak
6jsQG2+7F59NKzSUDkDHntXeFjICah8+YRCo6nqHE+EPdbo+fcAzqP4TDEhqLXePl0pu+LMQopTU
KZ3tB/NSKWBdEPpgxDM3Fd06niuc6T7pbYVs80JXxO016/aY37fYjbVIhvAVUVq35hKFRUobF+BP
+SN44pwDhJTWh/Bsjin8PDUvoLPfE4uy9SVgO0k6FtzwyFLYXhd1hHtedxOx3q0qjQWXfAfx5JMf
GKQK4lpc/Gafhh1sXuriVSQUesRHwDKRmErE+zc6+BrS5GTtQrPNcGWuVXdsv++FT2q4RFlJOMJr
sLfL83ZsIWU132QMP5WnlQBz1dvLzYHjyIFhXv3J4bJWuXUq44xylyq0d2pwpiVGinDdEk7vl1pP
96PlInE01cg5p+AxFj6T9TfRXfZfxK5msG4+YoDwsP2evMLUaUbrcdwbjT1cT+iGi+52S2ebMKml
EF1bI2LyJ7r8ucmRQebDwdZZSDeSSHbr3HimFfMSsccDqDQCt0sA69hj6yQuacne1QiRmKqLtJOp
Td5wuu7T1Eq6iIge4/E/sxiFMlyB44OgQZ3DiM7gDhQsDSghO5sGSzA+WtSB500NnRbC2UXu4BG2
eeWerQqjssUvYsEoC+dKX4nvWRuotYuwrKlVGqYtGRfFLZEMAXCm9vCVLcl6a4O62uWAv7LKRsbx
LDsH7aRFvvBLVVJeV8WDVdAlB+SZrTpObySV3sMvZ/Arm6nDoOi5B3BnxyZYqfHoJ9NwK8sLAUPD
cSV/5yBpHzPc4w/B6AxRP6dOBTF6qdQhO8aJ3HtnNIjUPYSVTkt/wEQxM8X79TvZHXheij8X3MJh
Bb4Og/tbCPu0l3hYiofHT20h/cKj7CkajlWZwZqH3rOTjFVGc5yy0D0xWWxsDZ9Bjxx+vHoxYJTk
TGREeD0wRoBpucIiX4iQMIc6RboBOy1DYM/4oQm1vPM7xE3CYNz0JF8wcdHz3gEfBO9QJt4Vv63Z
kkwFQ+oitxBPYY3pgQatEN4Ns/NhX/LS6zIEi+OwiP03z6KkQ8JuMfDpBEnHERaHUmT/WxvjNaCR
/FNWkKEf1tHOByjqTEzWkD5eGw9c6XPSOtbhrRbaxn53+LUrEIMlpAj+9WqCHxE/zlweGCXAGpPq
Wid1SI3uOkp5AOtyJyi5gU8njMNwRk7qoFrjJRP7y0rxvS3uipNuXLpFOotXdGalzEMSyPgeEJHl
WH+wv6XIZmodstcO+1Cr0a51WT8kBsTN7+ytmJrtiAPgzSiUpwuuX9028Cy5OjDOXbLS+Mzs0C9i
jOKpdTLuhmINw8OZQKzegy7omrORXtUCxwrLkydzILMCOwenkGklagss4zizqOAt885hN4oumNbd
toMHATkffDgxkkqxsRMTC6sKSLHjLxP97g7++pdqobAgxcBxy54XyjrJT31wwddlpwzhFO1Qwfkf
KT6fvEFHb5pZKCGovzmcyTDMadGT3aojZ0uk6JE1HppWd5PSVZWCjUmIGx1vumBgun1xXVvGqLGc
Fenxy8ox7F1fBEhP1r+iRKwsK2RpV0uixxTyyC8sdc5fBwj3C0+pHYQnAAQf3IWnuETDUCjnbqTZ
GCHF1l8iPgKooJ7yhKbxIr5dHTGH0a4uRXb6+a0jVQGHE6vT/mN0rT0V7C0NWLcqOB/oaPAMQ3H4
y/SfX2sBZMqEfLeqr5pZclc8rAXKvPsRkDuKgtkZklssU+/m+wQGm56bN0s+Ffwq/6KpzJPXex2J
tgRsk82Wn5beDyHg+03nl3Bhxn9d53cVQevwf999s7ueAnV1LD3nI+gZtsRuVwFm404920Jlkz3w
QHG6GX1DgndB3lp5UiAC0UjSLvtUkpjDqfUMulqYP5UxtlNRm3R9GVYlBCgTdM+HvWcw6D/XaZ2t
O6HGqOdVsMmHS0kjBz/nEhUleuhC6e5eronM9WaVBBn8R/R3xlUuoJdFmtGNhQG+2vFEG8ZUnkFx
9VJFgSI6M/GDJEPWAV7tRmQE5ygaIsI6x/gkGy1h1iaIfLhgZykKu7X7Bk6fbuqhlbENdwTLC8iD
J5h6Wr0y9rCEKxewPF0vgklWYNCjKwpyGVs49hpHXuhFVm7OdfvCixuzEnbQZoK3iyGX7B3NdmFO
auVtMyoKqqFSgGhWcnrv2wA4vC9epDHZJneXUSuF1qnHOByG/cWdBwX9KyTXfCT4u/nAyaIXf6lW
qwqbnHVC5a4pTFAiVhPZ4FW6DtKVZwSnBvO/yRnjyqRLwog6Ho85s2rkFEH6OE970Bg5iYl/QBez
R7+okfpWdP8wXDrcZyn/aUU0UrOuWEi8yyXaGng2Y8PSooj4W9Js2Re6LBqXpf3lPUusZIbAc9D6
2eJx3nIJzVjHhR340w4NM+Z25nSaEz3O9lEfSpmf8d8FCedlhurHBi0wK5z1//csUoQ1x5TX49Up
R+mIYobKlZhUXGcrBlUGHIkb05yvxEt02VSPgIOgJJeIEoqCy/DrqIlvXYA5PxmriS9gjzZDdi2F
oAoC5bB5x9ByUME6/y/UOGshZO1jyTCh3PIEkYt+iEMgAjAiYZMJ53O0Fb9umRrEl0ncsrqCu82Y
c8Gj/QKCM8p9RA2hqzUaHFDF4MHG8FhwJFkC+0K1zstB1lsn0B/bMSG2aZD+Wn0oNcFw3MOrA+G3
Gsp/G3xfd9Twe7MmjZ3CTjnRgSpJE49bhLFVrhf5OU4n3AQ0yLsBMszp7GLe3HTdkfrpUylhmyzJ
2AJmj2VSLD61sq/b2VPFSjSZTkoLwcg2Q8oXdaGsvFCw2sp4WhWGh+R+2YAgSR3D10lfaZYasfL5
iFiJAY82Lxd3DSttI5zBmJY8MPzNI4dcc68QFZeqYor9KhUxeTf2y/+73FdthTBc5/knJFLwBzrI
BvwXqVwyvAxN7G5ogtyT7oq/UvyEPy98v4LJB7iL9OIwAcVn9u8ujgDA3vDdWFd1KBcDgnit3O8q
TZmMF9nMxd/dZ/HwYJ3ETunKUdYPd+5hfvMa1qzw+OzYpKIiWV6iXCMnA9l38gxftaBGaEvgWOan
TS9kL0KUjQML+EaxuJU0s4xtlZxVB+InzW73LTCPOEXe00k2mxNyFdCyvW9D/mKKKWYW+n/+XWsi
gSoOfOfW61qkKYrwaWzwGwkWNZiXjONfn8LuAHA3mYjZ3CevXck+3RwcPbrOfZlHlIrvKAT8u4yp
PrTbxK2hVfUpAdrhLB07+4fSM+YicetJmGyqkL6gzCkPmjJdGIS3smjxzgTebZCxo412RsaQRK9b
ITS0EJtjSbxgWLER/zjiRxpMV1btcA76dNlsTYGU+cl/SgI7ZLsm5afAsTcEGLy2ZQRSLsuAg+Oi
v5asPH+k4rmnPyFlr8ioDFXAVYmNXz+tU0vAn6dbVd23OuI/hp4s2tY3T3FL3rhzEfe4nml7lqVA
KTW9dqttZXJFzVAFUmE2HXFJ1yQNVxh2QsLGZUEC+3lmGN4w2FSAvXlNCNTAO85wEP79m16Wrcci
Q2S3LDiAZeW/pTUQIusUefU6O8mhx4uwWE1N7xveG16Uga/yZP3jTdDwkZPUVzsSWWsT+VZ2YmWh
38V9Fis7GEHs4c7xR9RovuegrBAQfcY2xhsppAA6K+3h+8fPF+eKGCBVVqnXMG17SKFLbyuX5n2I
eYRaUa7McBtjeheQYS9YCVOu7mP2d9/PZDry6mNP0rnjTMtE4m1hLvmEIVE9tX8Sgn0Zx6NRAoIu
vwiReloutOy8BnIoHakVVcqS2bNFGuvWFXtOTnrcMD3ysXO7fwBRPVQHIuvk5SaUlZBmPcm+rlIM
6t+2FO0UPPp72ZzBDb7Puc9hIktpuMGhOZJ/l4bCXuIeoOa8Q847DlbwqGVQQ3IX4u9c41nnRn+d
nY3JMxsQ+Y9Zs+RSUf1x6rHg+tp1jCeY+mE7k7OBvZTbbYviCg1okEBcME+mJCF13K1rFDknYe2I
umNENbMkVh0gKvImqY05iYZ2ENhdpQp/uq6VOi+ylKnGS06wBArRKqvZyNHk5Y4GczFKNo9aRRFB
HJGCNDwhKKrChJqfngDIQU01KuADaNDNB3PJFmjnMP4efCT9E2S6ypZ3rw+055bW0rNXXT+QyVwT
gpMrM+NXZxCdtS0YTD/pY1fWjyIb5iK44evc+g/Sl+OfkfphlJHYN21iO+zTJSE5qM6I46nf+leh
aXwRYWbJXAIWp+vq7TExE0v3s5T1v7+gtstXIfF2OjNDjL+Ak9xjtuohv//Cktu9F1bLxa3G4ibR
xn6wTEAmv/BTc4rNluaQOrfXj1v6JjASDRRk4xPwI8t/UqthkRYiP4AgBbgfutVj2A/4ry0Bp5/A
S8Rtker/fYRojWxAbNZCNjIWKRvA/T0zFK3XcpqX+dlOA51TJmceqj2nYmUEO8AYbW426p0BaHhE
/WIMGcQWC147/ChhGx6gPPdSOH/3/ylwOCOBt+jz4raWuVO9pdXRpljUdLKTuMTXhwaLvzHv1FNv
0U7vuKl3kGNY8UL1XDx6uTmH09dHzKbHstiTCE8kKlvRFmiJRHWVP9lAyvXnqR1hwBVWjBf8dBMf
hXSWy929xghBuA/ycSGV6bkYDFxKJuNzYjFwA8IULmhfNDp9kmAi3jKpHtvnCMhvSdxU6b/JyiYX
1KhtimBi2v9wJPhoAdMD31qjvGhQf9p3jbv96zAf0veu7iEeod3TuwTPI4FGklIblxoUSS9BMqtZ
meOTF92fVijryN7XygMZNrKaxsGT7G4icA5Wt7FP4DkPp92iC5mYLXtj+pg7D7Zbg9QeSACfFFyp
Kzd9mMJZZ0/jSTZEWzeJSbngHOOzuZbJ6gFgy/Czh5AAc08B81bZuatmouGzD8uorQmACJZrWyGy
0ES4Yf+UiNSjhawsJ6CW7yteN/9LqZTGm0t5zZCtkvi/OJuHOkGBWS7GUn0hX7HuI8UrQRRIQduM
sYieeP/SWrFGZjBnXz45Ct5swokmPvyyy1rCTQvsoGwqp7vPHrwhryKBPEgsr3fEbj2ckrgNzdON
DITelgV/H+HXleHXnS+cloTrOhNSjPlAgBYbaw8LtLNAszebnstYMasSdTnTkm+4mJ2Fw+1bCHxt
RY62bvPAZ3yXg/1JeNso+xuz1HlYTG5MvRtEsByGQTZdUhwafyRb6XROlmgutozJnEwZ0AAabXI+
/63YDELz2xlghfx7q3w3EcTRwNL8cLjHm7HLjfNQi3sw+I/n73sPaZsIvxUZGa199HWPIybRYkJU
5nTCsIwK5NWqo7SJtEdPMR0gHjNR+3GbR41hE8zJjgAPSI5drK+d7T0N/LQs2U98ZRek4BL9KBKH
t+W8Yv4nc82vzCQhhQJtX7J0rfH+ujD4u11XtqEJEySuB3SNd3LpgU0T/AsNna2rtDbvPl8/OFQN
u3hLsK0Qr9jttWcFDmLSZRn7/Df4hAh5dnojF0GMFSLkez3Ib7tc+fHJ23X3eimJ2JRxfDL3NGGb
X9WIjdgiX5/HLkjM0zKxtBLEkVly5d6pqW4Ekttg6Z8HbdLuyqY0iBxb7rdFy37veFGNG//pFprF
fcIc6gKoCLJinrXuymH76MBMSdEaXDDgHNBnfUbMpXWFCBkAcC95kJEEqRz3UrmlZCZ6mdudsOX0
5oHbUwMK6np6rrM+aSuNza1ku0Mb3s5q9fyu8FxMxsYhyJtkd0ukiIOv05K2EZd8clsjI/xNFs85
s3SJN0nMMV8951p0Qoe5vno9E9bR3uQthlpUa2EZlrcxxCRjm99WmrFcbNzxTpJVwCOqBVlmePtw
mC0vafgx775wX7xvCevfVE/L4e4gMJaOrKAvaLiAXVszY9S8Vp8y3k8qSVB2pd5aGCYlpn89lqut
dUfnZgCMgXr/FFmMCnJQWgr9DwIkYyL7oJodJl9sgQ+kwsDzi43BA1uuaLNd6MQmO2DrQ9oft065
u66bTcFKB+EPm4uYhFX6HM7hQkaBIO+KtUWdBqWqB1j+OEGv4f/Eb1yOmmKjkxdhDBk0H3De5IDO
tekw9P4tb/n5nmJsMnP2sYoBOSZjk+Ix1rAqVtJjMGIsiSojqMSfryKRUoHPvSI5k4LXtNSxxcat
8Serg9LOUlOXwx0dIakz5Y+fCFYPl0mGJHskf+feAoyUE6MB7668nI6IimuLQoyOstYXc9gvhC1K
7VImC5XTsKPQ2IaAEWR6gsLjIHrR67srM2f1A/jlrTwi1Wm0VwJpYPFo+LgAYb05X7hDQ83ms2ZU
rHtR51Q+qJYHcw5LayKUlBO1/COs2SOFArZbSa+mc6OIbhqPQkYsq9EocjvM/r+l+mTuAyFIjPCc
knjISZMXg9TJNxkWXdFdidKOcpoG7VSKvHgp9EgPvS5fIBOoBFwzLhuz+07/Pn32iwM9IQf1eOhS
HGFmVJ55Gyee7/M4b/OyZgRqUabqw/D4mbTic6MkRsLCCRKtED4mhjmrPYGpZRVDkLInW6QQiqda
ScMtUsXxg4Dt8hKtBpwyeeCYnbLe/iHObb/dnFovz/V8ab/50eszKmdjoSoiJtDFPYPgxX/8z1SJ
8DwEG/JKLeU6P/0NxYgmiGcOgdtY72PISMHB3clvuELNX7kXWV+wtJWmop7gMtWH6isrGp4zuc6u
L9GMhsS6yuLfT0zZdLobvxuHS3UQ4KYDSVXVM7tneVx2UmJn3EvZ++TXYh3VpO8w4MiP5knALbc5
eoQskvQiK6ydwH/aNWurBBHqR4JrPD3T9SahSs58AyLEska0jgp1nL4oYIP4IpQCwqFhzu6L3mpr
S+JNpZa9upmk9o30MT7D4siK1IFU3JNNAcLMHQ7nFLv6yH9xsHnObMf4ikZAxmvRtGqGTzd3EtrS
HwnRdNXsRpyF3p0ljiD4AmxsK38vT7sM0bMwxEmDdG667OE8xcz5WhGPMHZULaDdMEYGym1rhv6A
xNA4EmIqlHHgMpph330gFZRU7syh7IbiiIqT4dTmWzhNNrFNl2lQB6a9bcSV74C+3RzbGPEUS9yl
AS3yrsQJUytPjyxp30HciYAisOje013LW1ADQYbNHt3XWzeb+pfc9qvA2ATxfkm3N0CpXHl46ytW
1GW1YcRiK3t/j5hSFWPweAVuqZ/kRfs3aJyJAuREMc47POKjErbweoj9+vzt0LUDocLEZR/bPrGz
ms+LduUZLtsYiCxhfWUWM3AxTjdrISL+dhXDJrMijR9UBMj/NaTZEcv2qtXTc0DrJL/CGe5/NhFo
vkJox+cDPDaLB9H3b52a4UmslV8hPnLINVCiIaMDbDR4wElgFobCV1xeFbxfyrYCfEr9+90uRbsV
gUk9FlmDX4R9EQYqnJxCKebA4j/Mh4cvME5/+6E/FRi4wqewM2YHDXJyoP36L1I7wSeY45ivKkmL
T1saPh2CjGtw1ZyZXTn6e0Wp0UQi0BugnYkg+uLYVwCXz963IUxGjPdp41NpMC5j49pIcgbcEEl7
CW9kMlY514igrkC+MuL/NlSzk6or1DHwx8M9k62f8s3mwElXkQQy1URsjaUCbK8izQ5e4wDb4Req
694SsXvsCkvjq4WFVLaW5KmMM5ypH+TGqmd7QaCbyr07Wvw+/p1iUfluZjhq3fn3N+HPrfcyvLwr
pArz022ySYXfdV1WUEVAlZD6P363H5Cpfv+CQ98fXH6LFZDBaGayp9I4GpgtPhhD+Yu3JOKAqeFh
BeSfbZ0CrFZEAR9HIDjLqwAhtaXEc4hqWPEPKt3+ssyYVSQvaGWRFjVlkYIjGfWm6fGBeyHPyMgd
t4RA1IhAGoFdHVGh8t0TO21TFnF+G57q2n6a4hrPc8ov49IK3WGx5FiwnNBaI/2ZKvuQ0MnZpFs6
NhWo0Oktq38UDJCGH1NIKzy4sN9DIkVi2lyrcfvpUnxCN9uBfbwhphC3MafqoGzj65ML4Idk6tUi
P916/ScL3svrq8fShf89+XKcTVddb+oIMyA228xkLM52Hb2t2ewHZjnA4cii5vQ6EmRa5WjOe2gH
dV0xRq9MKydneIdPT6LZ6JEXed2kXgZAoIR7RdCjsHBltiMJyh0pKk148a+QDO+nWtPVxcnn6y/g
p89ukBoDJN/33qH+Km2+fTxUA5ZmSBkEJIm90QVWTzbHcK1RODfTIuvHkOyQjuvka3CUIagzr3hm
ucr7TjR6qSshvKsfkcj25Xyb9yrlkKCBL2pRNbAZr2Y7pWQIDSmiip7o9NWsg8bKr+/ug41yTQT2
s1gYmLuBwMchfrkyBI1dzQSJKkmvjwzQcuNq6wMAnagzWMjcI6jIrete2D/4bYvQSAXE/WEByb2P
z+xOw3Ur10zsU49bVVb+MC6tcNE7db56nNNynrM7YkOCvfbvCPOTO3EnTl9UQGJNrUHJqIdhXAfd
US+NSJswlyUhIg65B4DyFJxQcxgu8edVYQub4TrcszfsYe4Rv/vZlgF1ucc7IblKVXasCYLVqFjT
ugQAicwCGbKDBcr+kU4w38Sy2g/GYYW3pkpkaQ6YRJBpyKgcebPM0l+JMU20UX/d3HZFIj9h4ndS
q1BlqM99qGUedS4C+qoV1ziNNUJd5Bc670xMHB7OsUsgIiJjfPKwukpajkWo3V4v2m1JdfZwQ58C
yRIAODua/oOdFucawQiJ4HBlKYuEfqHzGsDJSxARMFKDYwS+KKjiDF3hJiwXTzqXtQk/gN2TlYwq
Q/Vp+Lqvb2WMJueU0C40OP3eUPPgkem2X4NpFDfUN3CL1dwBGFKBEIE2vPJdRyEr6MuW93vIPzAt
laounhKw6CxrGYQ8h+IK4X5x/r3Fx8SKTIVcFWauVeYRymT1Z4RpSXehGjdOpDS/sgvEBJJMYG+K
rBQTrWYCrkDOQi5czaiLgPwxa5KTmZ1Ge51eg/5P61OY0DHZWnrtoOA/2z9FZj0Og+ADu+nCm5hk
QfzdZoJlBQHjcpqwo/Te8eUjLzKqS6btHaBt0qM2O67XcQwpWWpTyTB2IgzNe00uTrX+QJfHXp92
hy44dttgpWFsbc/a8ORZ23GoRtrk1ACUHUeokXpRt2AWBwBhb860bAaAwtmTY0XuXQqJkdtpnePX
fFq/r4yf6paV18eRDhEuXzywKyTSHq09Sh8t/992uol4MQbRLy7ALvx5FnRqbNEwRWDsAdIZF0kD
z9LjvaG6bR1wH5Hq3wgUqi0CBnmAM/3ih4zUzljI87tOWhm1fEzZQuKjLBaVw6eY6rHyGcOjBF87
gktWAybZ6GhcKaULHMT4Ii9RDEUl3c4r4MrbG763FYek4etUo2zI/jrpqEJ+r0T2/a8RMMPtBAKS
NJkzk24FByDoaV8rWrNDl+a1ObLi4GbNwcI2gFrWf8UKrujQ6he+6LDYmD/GFtuQaLf2QeA36axe
ndfEnX2PKq0PgkHJRu9QjBuCqYH0UApJxmeovoIpqv5lx8n6IeXS0sgci47JejE0HDgyPyI9mEK3
fFkxK+56sui7WrErjqFyCfarq6iKpZUmNp1mqMFrX4ia6aFzPnAtKOsHnfLYz2IGNypcsaaFLQmp
gQSeHUSxPSWSuSi4RMoZ2A3HkjD6ie4xF6+dQ0IoYgBonJmDQe9cK7v1H51nfr3p/yfil2U5IOa9
YnpQGYdvkMgmvG9mI+99wA8lcgBqbOOBH1aWbbTFn+BAbRx7sAgE1udtbf128eYpAQHulqlkg5Zv
0qQ6Zo42LaVeCnmDHJF0ecP6L1UWKoUsKJVGFiQqG2i7lr+AQBxyruaMn2u/YCoA6PYDdIfO7pVr
0zfvM8o7QmPKWlmdKudiNpgtjIu+OuHUsrsLJ1aMJip/0rbnqhsnWe410CVuPSrxQhvW1lnDDhiG
sADtGhv8q6kSss8yeQZTNj0zPgg8LQfJ6nlKOCSVu6naejaoYIgrUy3nrrny31cyJv9s3aDBl2pm
Qb/47weMzFw995OTvX1gX12mXpw3OGI+kp7TiOP+B2/o6bI3y4h3zzRsC4i43ImQqYyvwGaEkGSi
LW64lFHdoEbaN/H37Q3aezq6WmXro2rYvucCw2kPvOtQWUuhSx3vkLa0dzTkowtp3/PYuI1Yr3Cn
uFyXqOJEZTbloNMywBe/E+VMzoZRSxZ7MBQo0FkYCcpbIuiQYp9/wONtL6fCWzioQSm9mofHXe2Q
O0D26yWDCSMKHI16LOEN6FEVLXhvzcUS3lTvBACFut96aG0hHv3buw9BDUSw63GBnRVse23DtxqB
y5NsHqK8ufXoMAgQkI6Wcul83I+cynl7VH0lzOmvrmw5whOrJ/Ww+gk3s/9xjj0lRGBrOaVV7eVp
bTllkkteTVRR+7Zt4kSRlLWuNcoE54anHTHBcmuQXs9LFMwYvsL33mruOjaHmim0PGU43RNGwJtI
Ucct3O8v9HriioFgtqbdh2BvQ7tBoGKHaX4b7k21/4RBmhZ7Mfg5p6YZw2dOwL4qlBykB9Jbk6dp
FPqIxBLesL5e2ciNAHGEPzzMkm4rq2MGndui7EKpjGWhOZycDxq58CXeK+vGC+burSk0Y7C1s0Bv
ZWWpcNFkJTiX2aUi+JB42xanQB1UAk+o3Taz243DjdD4HGedM39yux81P+CnzBFo5A0rLwk3RKqX
9gYV81en6/YkJp7bw/X/gZGpLZdx36PXMq3GPAtoFsQSyl1wGQmFYBnLOBdS0E85yjUQc2XrzN7D
JqZGhdbIJWYBm5jxqIXIYW84JCv0m1F+ewqj3soivzARgMpRceu7JqdCEKeWCb9CCGRbUmeSOMl3
WTn0b5wIZvVXYSweH/F9DcDSJmDOh9M6rs1U3cZKfeA1wX+yhTMzazdEyDhx2d4iNHxYk0ATRcXG
8NlR0DT7qLTJj/nJpaAOcMA+scT0CgZF6qp+XVrJDl9hOHdCjA4gjoFLxMZt31nEcXU0+hWg0YF/
/AV3eIpnx0+v1rAVetwaLbMFzwPEtqvDiXG6cOM6GaZWgOYHjsMGDt5legaEg6Iym4loZ5Kx0Aod
JBkO59kjgHaSZ67Q/CdnXPTv873WWXe/n+5We2XEKgJi+QsaPyUl87gVcRLhVz7CXGcbuOVzvzXX
yELlcfa8B4HYrof+yWCluAZ6Bh1aFnYy74f7+F3t40ezE4gBnMzHHpltY5QIe/TJS/GqexGkkcZw
bPEcsw/8Ou3pBlqJ7DC0h5oZspOM1g96yYQQH+vXaCqRzA0D1Rq04GsE7kUnc/aGu7AQVAWAmgBt
RWBvPjh3kiHsonxaLtWKuXQB4FB5SLdPgbIiqij6lnwWfH77u1dPO3PXwfBHJnHZ3YFCLAyjnPLH
Y/7hyESWEF6Aju9BFEhQefSYk+haZ7Y6NhpFShtZstLNPsWKZR2spKvy0/Dst6GoXjmsROhF7BSZ
4Gb/84zrD2l2UyDbx8/BOR4FCF4dCUbnPfN0IR/oUDQ3CL6j0IbMAbDCgHXhsg5HlBENy0Q7lctK
D3p0wtVfZp2jcmJgBAveIcSu/m8J/o47BG1O1DKJXj60KUZnu/8oEKJFZ/VunE7hkCVgxbZUvk2e
EPe4Ewijl8odhmAoeISYvHRDdJhDYHLwVV3GDJs9FZFgcib4ZtyM753lB1Ovq0i/rXyGGvH0mnh/
Jlb8kZNN/0JGHBVz9px5TNeNGpuk21M/wb+7sRhifjWE5JebuA9CrQJ0lDPmsdmaZQVz7A8sYXbE
2EwjcTZa72lViiLwQgBiPsAQ4L/WMgpq9wc2NnSEi8w246dphwNEQf63f3yZ0HN8u60INn8CsHoY
fyohouEVi8XtcghOs8DBl8tYDOHDquVmzXwh7s5hhfjEl1XF9o/bXSR6WI2sutnW9guTU+IdYDwr
IlzQ5c1L1rPDQAKxXARY99gHYtOzqxLt7Aaf5EWnuUNqOucC8d5+8e+DihaM01NmwyixLK+47sRq
pLlkpfKu6YW9rsnvxvmQWSYYc2zYRmbtG81y8JLPWCf6Sq7kpLEok0kkzn6fLdFGUzLImfMQbCUm
XGx0W3zB+rW1ltZ4eOUCexP+AYdSyJQZguPCt1GoS3mvoZj/NqnRTxg7bQgUHbD4yNujEuBnEFbE
1pZ5siECdsB2D+U3JDaGTy6n03eNsuHFO06YNWVFqwm+S57G8B5cUn0XRRDj5Yc87h3ERI+z4wpZ
NaZnP+3KkMnyI89B1CG2kQGcLEazsQfA96JWocf2bWinDU5HZl6pXHfsUqes8XptUchwA3RCM1gC
HaTe5nxLtzzjyuciuErxlv8Ejc0QWfWStir4SeOFvYByvM/gQ0iI+b30Uc7qugAQjIwOK9EiLQC7
HkPCbMb9+f+DoRpwZLNXwEXmIZHBie8+dI/c5Wzpbaij9vSNXmdY+leKXWahJ3zI96cZMQeY1Kel
pARua7NEPcTAKJDwIeFQGvm2arbKxEAnkg2u3B1EPVOuwvCiKp6rcT+x/H87EZTDRX3rgcCEMmsF
FYtcZCH7dZWYEZASt3SB7aM4CJ1+hjSbe89qjqFyDYqb7U69SBZknhP24pUjTiTUvNcc7F46tg5/
2APiL8vn/Q+3QZ4Hmy2aELLKs2VUeOb9l8XbnKrUXX2mPCfGzOmVgCaLebDzORI+y4o8pI4gW9oX
KfbtrGuUL49pSj88bAUG+K3W7GZF155dazRFg+GTFfRoHaLXCRnidqptpGTdtGkfN6AERKO4niDa
8xh+fU6fEZ5p4e5gNiact+98wy4Q1SCtm4NwMTnjZs4Iq7wsPqWipCkLRyEIMjJOkQxpUeKHINyx
HaYArNs6vN/iv+pPrNSpUF5Tkd32W+DwuhpcrMkBrk03kw415hfbdVe4uy9nR9p7TOMfFVI6IuCK
M6pOTpFdMbRfC8Gwrpys34/MVFIdbYN9ROPsFhKOIGQX8C2apmhT9dd3Mu1rJg/rKmHRI6CXxmGy
nXJj7N0VJchU7+c1ys7As73OON+iGHjcRBwABULv+gD/UjEgpUq4W4GdC5tlQLVgxCrPwA+kvLXX
U5cLve6qZw9M01d0Cv57fdqDBwKMRQSNKAXk+Pn9bdSGCsaTgjzA4EOPc2tV6zCKxOZqFMXYS1HB
c1EKWNmK0ORifNrVHfi56mCJCtZneD+a8z3t5SW6DbylvLW/04DTeyQf7FOKTiHoFbIAO2Cz/vXj
AQwQ202GFi1avnwoSw4xGh+T7Mi0fX4qN+5/2BGywrCa7ZPCOxST8KsXc32iNdJ/WOObZCSXx52A
CZSiYy8slOkiTiMFjD18LTuvz7TFPKiT1t1molNxGznxu0YrpcdIrBmGr6JfvJLoEt83ViL0+Pp+
bBGr8ZLx5bfuoY3EmJmpAURfwgKutDlNA8KnnIQB51tTMeuAYPN3yJN7+RBt0A3vq5IOLaDXS60S
PHXJUa1r+VrIAPpHgcF/T+xLFbJ1SQRKoIPFRvfRCn8zY3/FIp6vhlXRjsWZZr8yYFw4DsvOuSDw
YNtfBQVyR9Xq1YHGwl8c6kxKnMlul0K4BR8TqibihrtzONZ747AfcEGmOWIZ/nojiDuk7sBBpVdn
RamvqgYcWgK7lz/UEN6YYDdXFXw351ojqw5WGYDj2XZCgm/gbumLmT07D2zIJ1EJpc2ARBXFIudE
+2NTLoLRjTStQJNu/m6jp5jmzmrLLKL+u320Ss1q+OVN2kdhLHwj3MkeFHKNGTuBONOxNkDHFttr
FRnIQJu59Ss1lz4j6AH7xW495nX4j6tYpG/RvLjHGNJycIkLJfJ5kCAvD6D0LEbG7VJleDDzp9Hf
CVU5/Sz1RD0RUZAmqg8ikPkJ6JW4yjpmjt2U7QeGZU/lEBGxIERpgH7jZLQ5uUbGqT5/IIf85dIf
83l0mKuOhY99WARL2INd2wGgrLxvsMyZaYCMB8AjQAYFnM/qb2ag18C28Ywkmkbw6ddJsk55Valo
dE7j/ZLpHYms9tN/ItDZNcw7DctoXXK22ypfMiPtc7JpS2D1qGi2WSWvkojjTIYY/CmrioJroRaO
eT4XTHQ3DlN/kQuCQoGNrZ1qujnDxJNKSatxpWisiKMszyiqoTuE0vhaj6cmDXulPnmdyS3qvSxF
+a5Ed8bXoqWYxCHjbOOhAvTqcsiV4iJXsDAr6eM0/Gr1iX9/gnbxQeCQVn9+dxwMXpKB04rrEgCO
yFGaVm16eRQ4dba+QJG5zA4erFpCc8xTxi6xf9+xHz3WUaQ5TiKGdIjb27joETUIgSv3MtWYrLLU
YGAegoTP4iELu35fM3OBNBQSXMASUMCD9CfACZz8IRnV+BQxUSNm5myRo3FBgTlxfc2zO4ThaLpp
vNfvBDsUkKcq2ePC2+eVuK4XPZSHPSie+PWeozHSp0ksqBnh/t7CGNjhd6YjS5cgHJanWKSn72Xg
vDW0QB9IZDFSQGUlvZMb5mVbslB2hgHpYKj6dC5ydTWKRBjFBkcVVyVBiFRCCWvrBGX3hre57z69
oia63z+LhZ+xunTOExAGP+UJRNHfqakU3Q5pBcCMo+3MsREWxG4of4lQr21dNRTog67Y6+xGM4Rw
whg413TW84lKChybrtZMhb9sjn2xFEKxBmrnkFOKKE19YkmN1trUssLpE+6yHEZt1mxK0oOddG9j
/i8kWhxFCg4hPLcasBFDWnF1pGgMk37jS5eIpKMh+p8jHfhRij+/8B9oMePB6YdedExrLjw+K8eN
84u9e5oVy8WtqTkFGaESBpuf2GUQSGZ//8aE9Ak7GfP6nQDasgBWHIv5sdqGSv454fB8WbY7+U00
a2gvHkGF+U4EOM59Uihjv6tNasAfIzCSbQXecGvD1452Dw7u+J71Wyuh8blpnF6yJPKwPvJUJtrI
zi1V91K1IDyfByd74opJIVYkrkOYyTMbugYltzYRLeMkdtJsauETfhv07VYDP7+sRXMUVxqvAYzX
Jk7rZZ4ilL7YWzzrgEhfGwptvaBVFrZuEoZV2Fv6uLpyLQwjsCIuR0JEEBslVKEdq1hcTkSV3xNd
DjoJtLGFH9ra294mwfhZnIao0X0IT3/NfMsTf5wvYZhw5SbrbE+r4rBYLYmbJrHGFDKqCg3FpFjl
Eh3GZqxGR4YRnV6RS9LtX0zw8AR7v0sxX5H6cW8+R4R+axAUsNMsDfAcyyVWzWBCnmZoUuJS3LAU
kR5qPAf/NLP/9GocsGsHOMf8U4ROIpkEHMX8458eD4zPj+riYqiG4ZE3ISgKBuKqHlW0AylpdRQm
zLqCZgSmBWwzwRtigOSYM1yPF7WHvZBRVV01Hao9u1o2Dl6bgpmDsFHZ0CoUUu0wQQv2Y2kICwfV
qQ3n4Jgm7yFKkXG1GWrlG8yxifqIJsmD/WC1Rk8aeGGghpJd3h/zoMz62vk70JQ86VedD6IqrCn1
b9a069wpeNX7b2FaZaNvyjSZaC5UzrXd8NXVdd8KXKn9dSHSN24f676GbW8tX2UsSIz6SE0BCRsB
vREsWIS2dLC23G6ZgHG1ANbXj8G/CTK4aFMyUAoGW+I26gPExfwKFF6Jk1oy3ajpIOfu7jqLwFBs
TjU5NckG0KbcxNl0/jF4nXNwjA/G6yZoaaindm3Jt8GWv/MrTHpb8xAFc8suA5TLtGVxoFMtuikL
ECImc8MENg0YVf7g4bimPGaBiAYNdtL616VQmYhB6lCxWwiipnnjkMbi7ZVij+Qek/qnWzY8Ttqm
jcOJKneEy/AjeDCPTmubt6pzIe6OLgzdFxBzZQN3ykUwTtjeKaQGQB6s8PDYFXWWOoOhd/63+q1e
sEagoyRt7aA1m9MtPSIiNMFSOPOt8trj2wWDd+7wKemNLI78dvzaUjA5Y6Zmu78NFAEkDZ1BYns6
N3yPNJ2Ioq8AYD1mXJeXU8M1tC4fce2IUd5hsx1Z8w7lumVc8XsZGinNRlRgkR2fPCGeleAwAb4k
chTmDD55BqrI6aF2bgXyHPHEPIuVY3nCwLyNDY4Xp0cX9x4k3DTc9DKpz4MnLjqtfMqjMi4ion02
BqN1pqsBRPn9uNPAaMHLdmdzlGWz7cO3HO2R3ORUzvAyXpbe8Dvk17Mx41RjKiSCq13EwH+2KZDY
CDejKy2+cPzrvMslyKLEpY7s5bljCQ6cjw21qvYI7vdhtMKFAqGI1XiVPd+qnojsMIuBBZFL7+eW
pza1lsIAp6NN21I7ROYVNEr4Qzi7xqWR5Cr36zKpL7ekk2gxVAEPAyQtABwZO5dPxdHNjVPh3NTA
pMknsgT4PpWGkbrmHTU+tLb4PRCRwtVb/5nB7W+v5rRF4zvUzzTIZLQtyJ+sCSuJQT4TXjV7nLQ9
pzQhs3xPCw1ENEWqPQrM5O1/NjYZHM62S/XvMZh8oZvY+FfpDtUHIdyxIcIgFIOr66KlCtAYq6ZN
T4qBhFZZrilicxSugQekmBgQQOT+k3ESo0cx86IiEU95crDc/wyxX7FksCysYZpOPaNqy+TbzVjQ
3hkpHUV3VOTfyf1cGTCRjmYUWAqHcMPDpADj2w1FVanqsdFehFZx/kWxlGIM41c4nD66qIt2J9Yl
QAzw9vWENU3592e427CtijP/WHXw2y9Koiup1uPScKwaJVihIaP0+7k3C7B0/VMQHW5fVY5CZmxc
rZB1bdSEhDXrWkM5J4IUIg+2+VeI8qmYxI3114o0PRTS2qq+PKb82iCDZImL6vFCY4lHidwLvebz
Og9EXnZJYC+S/lrufDKVLheNskHH0gTSCw6o5zFNKqOLyhlLbJD3LAhcw2UM3hSWEk1AeaQ33zJx
L3AkAvBnQvtHxWclYVs9G1i/QfObrjoPMoohElCw4jg1VmHfhYqxU2nxddovMkb4sgT/L5rikPwQ
Gdlu6JDw/pNowI5P/GUGvqno5ZfyGnWosVdHXZIu/YLmxq+7OYxY1s/MpBg6TjtUZ6i3O7MrjMEq
B/pBHvmu7a4R9WxHwh8QUMS577//1cBPAipU2JHDx+NhjXlEeTAVxlPEYSl4xtQhloFnxLcTc2IA
NgoV7JHg1J+MpB/pwgKJ6gVV2x67fN7sk7Vf/YUFjgKxUNbOO6kutm9rPOu87dLWKIY1nCYTlys0
UgnTdU1OJKOEe2OvgApSdruVgyamDpyVUnF488c7BihS45e/9aaBV/oA74al0fl1duJwHKadrYYq
H0aK4K95U552WOP+wRhXxcGv9OzOB0dHPo4ci10fBwoHKjOknCfuuPi6H+DhbIklkR3Z59CDa8xA
68ISkKzueDO1X/UvlCy1CdHuHZqzl7tiRkpjU+YgKozmaRcpcsXXX+3wvX+Q+RLqUBtw6pnsAC8i
vSQb58aEPJjUQ9d31YDNLRxa27bylmAALd5H29CVr7gBqimOQ/uH/OXArri4repf8ttiJpZ3GJl2
m8HJ7b1J0dQDwReHFoAc4krDTFiZ46DCdF87mAoMqVJTYB7UtMSLEFTZScEkB1wgNqpP0suFzie6
bssPgwA7s+Vo6fvyqp5TrfHLYoZ9fXeT6Ay7SEEP+kHvz9UU1YwZTLx2LeQg8k0hMMddWPphqFl0
kO/K+sbazxsb01f8vO9BxRDHDwJhPfSH/f3LQjKNzsIcCaFYMy76oqTNe8wb0XuiiWvt9MAhAGt2
rE4PDD9bryToovF9VkXF+HKTTd5pJBBSkGyfYZ6nSdMZI7JWaL9ksJGDpFalm9m5Z799S48Ha1JU
2iKWClVAHj4SMlydJjLpFyfAkAgctbY3oqCe9yOyLxW5pjWfIYz526yTkXHXG1FBWrdpbeM0vDf3
5Os+Byuot1zzkl8zj+UZDeu3jx12e5Rl1t/mZ3aESHdDuEOV5vxqqM9wF2ZatbC4RGVgRBBWyqVT
az3zEt2tsGkK3a+pNRVODPRoYozFLfP3wLS4wp/LTgHIUSGFnWegj73AKgSJIhQl093pN0W1o5HP
VDVudUlBAADRAV3Uqchx6Iq98tMbmeW5H0/fouaEmo4dsJ+FzFH7wM1jAwT7JWUcUFf7r6ouQJl8
Yd/2IeX5v3jyjFyPJRN+ukv3Vjs+qf+sCyRrcEbqCeIShgGGtB5SfkJuAmdBpslL8BZnnO5ceyEU
OeGvytc7gioLJj5gyOt33mG/hsVtWQkAUC7+Ry+FQXt4pcqDpszOhPVPUamNoABQAOcbQ1yNDEan
ELt8egHV+eWcLkCLule82yjaFpWMYVCc3ODK68X+aiWHNc4nqMKBQD/YRtQeChRrUILkY10hyFuw
+PyGOCYEfAPTFA1niT4qTuTmSZYgWRrJJTDGQcILnWXWvHUZbEimpLvcMRjDP0zplOQY3HHjMcO5
4KKTkljOCjyVYy+RaRoSYqhaCJkH8jyiRAGPlJAKGRWllcB6/JVRXxInIAQ29Xp/Rf1AiOc6kzvF
8DtntJpQFMfhMRLmpCTkcyI6IKrZCl+Nq/Bmwfii+FJ7LZNzrlfOlzFeVfXT8nCCpq4VovO/7iiN
bIcY92vmJEJF+lHFyIdqGGJphU8GNFE0bWWTL1+FZiLpQj7pS7AawtqbjtVnHmJeFhI9jWm8G89s
ebNR01UjY9TwCtcChEkDj64Ufuty+CEzSH6T+O+SyJXHMyOc5u2fMcXXvbgrCQAHLAxqz/3b6plU
MatPlQLFRYyUcUtlgLC1eqnOncf5RKea5ZlTWATlljezUGzScEx1tVysSX+cpylVfOpTuxfK3DAm
BAb032E+CWiKmG+R3NKbZCVj/RVPO/AiWMQ3LD3+fuaPQDN2C2gDi5TOCzoY5Nt2OKs/KlhSD6wD
ogGgVvEicifMuAn9eA+YiVsBZTbfJ3gdXDgRm7I3nei6ndfdsT7ULgu9GqPK+tRcK41a7keUY8qQ
Hlmtu8MxZ97Bh0SpF+RNxI8guiXudPYce/ISopWI9xu/7KS8y4qqcvz1Nxgr9oAwoeNR6T/QIxpO
aDOrpMrv9QOYm5xCIUpAS9O3O0cNtYZJ/2cR7YnbGH1bP2GW2uKMTBZ07Xem4TT9XmSXZ2m7zY4D
TMN5IP4eU4IC5RTSXChZ4hOkXIWDtl80OtWGO3Q+6hdndjnmq0k6Cgllp1eWbYmZ7ZXcdMUcDvJp
gEcY1iR3Sjo75u5k9WcTjnXjPjdmt1iBfpovCD+tJzT6rtpezf8pOfss0MOX5k3ReLhasn+9fY9D
piXG5ZcDgfgqyWpHPvl5f3kMQZkH5sJf0YJHcsvUkbUhKEq4rw2YK4+FMcnsXjAxjaeNb4woJ8HA
FHksFhTO9RJRpeOBnwqO/oadkQtRa2prB/K9UO8XcxfJdZ8LJeuRevBwLQxbbOpqOOLgsr4T6qX9
MmIt2mVmB0YtK7X2Y6xfCB9Eowv+QK+ydEyqmx+LCkdYa5bKuUi7thhad2GgCmx34Dija2ffAmha
TLo89Fvym+DrMsW5y+kTs2UYwL1ujlHg7PZyJeldp5LD6tfO+em4dAFpgsXlfKrLZ0IiuYOUt8NB
Ftou1fTQUyQbYqLdqbRnGrU+JXLVUsG/R7diezIcBO/1tTlcNl23kn6tdO0iWrcwhlqeAY/kzoll
3Soo/LNDpYZMbVkF8y/HaDwbySpo1dlk5Jw5mMV6Exe7xYNm+yzKyzzf3QDn41uHK00tjM4fa4QB
qTdsSR2MRlEyF1R3nIaKHbX6IxjYA/3uzeBRwRiErU9pqPeUP4UkSvnzrckKOZELV2f9lUpXKkPd
bdUj0xP0dJQnK5z6mcmvY5XQIPu5yl4O66yDeJ3PgC2RWvV/i0sixYvOTS0Fngq8yGrx5KqIxdt6
DLIznc471U8uvx67o0ga+6ZMd3Ss2Z/R6ecIneWgNioZbpQIWfVgPK6BchEmIrrOKJAW1hftAd35
G8bjOfW5NKzGetpZkPR86tlOdfOi6Gppk10HnfOVy+YM3jIGjfpZxewhmI8eGolZ0Eh4lJXMy+/6
JnCWMT9zsXzvU1wEKqlcP1GWF7Z3zz4AA+2G8K9e0DHg4h77dmiVw9vBYIXnzFX2N01kqfbP1xoj
zlOXIf9fL9SFFuieWKfx5qiMp9o9k1V7/3xivbjOacW0w8W0PP8RJJdk0/D5GKy/rN1C2WIwbMf4
vHMlhVrcBl4BNwdrUlfaLiTNnByQVq+7GhLtyAYi5JSYvFa1ZRjtEGeqCexcq/we4HHHpSvZCdo7
/0C3g2XQvaxySs1m2mDwbeyIw+oCDBLw4IdS8jQXRMg7tVi/LmznqFbLi796ZNZtL15a4Uv7T+II
FVla5/d2oVLHjGDwWzs8/UTdzOFv5zVlTbBJKXk/1chFDrjjybDyJEuP+1S+CTXhjcm6B4tFP/y+
QV//czVmP5O4zR3Vq19ViXqNMlHDxZYDPWVsherTdwjMMzPt0gVfPDCVTue7xFf6aQ2GonfypRon
rYwnl8pJJokNgzI3IZERgZ0tASRlvPwEkUrFRd5JLLTI831Mti0cNxoV8A/msp8xWJfwiwA3OG/i
+EWWSbZZgnEJ6WR9mz0yMmvX1fUkoeVbU76XVdnlm+LdXfWSYvHcgWuChWqT2AaQgqRA/lTozcQ2
VtuF/FDjQrT69wibMHZWtMe2lXBLTBB1b+yd3/xBr7gdJxT+VdTNtFABHQ7FSBZwwZ02TlBs+moU
GSdQDCP3PtepvfQc2PJx0nNfgUhOK72RJwQcdEW3hs96ftseVi0r7jU5JiDLfNOm01d9J6+Mkczs
mosSRMFqROwhNRjtOUqh/ebwpjuXclF1uzsIP0D2Geuw7qd/SXskGiQscH5UUbdbMrqSVh/KZU9O
wHOG2toBgzXx16PLHQuviPNREsm79885kkNLUdsq/4F+7bCwyimM8yKP2UVKLkHZjflxak/M10Fd
8ySUZrpDaQ8HzNhmYb5jghfDEJJxSuwdP43fcVR4ZZBkWIS+FBLDSyufocOJabvFA7WUYJkzvYZj
R4y41uPQmD33SMviG3brAJniaGytsjY7rXXdd+XtHYIGe3nJHOwPZnyJlnfE65fXsUsbkKqmvqP2
HJ1KHnFO3E03pznyDimeOgxtn9MSxjH9NEIpVmYbdA1yA7Jws3io91maNxMdhWZPe24aFx/y5rpf
FYfQiLfzJLFWUiiekCPeIxKMPEzUUp84gPXVG84qAsXUjcD5QbMB+TGZC4cJCk40hQ99vxiGmQqd
otQF3Qw0ecRvhqjJJGSWkh0lRrILpW9qUQVWLJh+4N8hRB8U9aEwUAfBVuVr7oIo8Rv5drtq24gw
itjSr8KWUD/65//magffBSdoLbAXZ9/RIjV6G6Xb3k4fbTlwmUALyVTOBI7QvQ0Uc/pPVpl+Kuhg
FkQki2az20Bz4bWJoP8QwgGPP23qRX/d1WukxR4G0YtfexgQHfDdDdhYAJ8cG7qjx88W2qMJUsd2
50cFKD7roZoJ48AHZsKVzyj/jHe7xRU6wLBobLOTmBglJM7A0J17WOffGsG71eir3m2oLJ6K0Mne
DTrFdPgC78n5CMraJw7z3NryFvXFVHi2CGBcrNCEik6mOQ5Pv6vRoemf1lg+svMld2NBNlbn3U5B
TT2VMzl8bme5rgeO8FFY/EOK/vijcG5qvKSADr1LwGIqdUflzJiZM7RNISAmlcfzx2LygtA11YuW
lyzdocc9PSjGKlF8pg7LysPoCV776QqQmYoqfUeEVphiy9uSPL4ecX3thOLJRtS0F+EQ/KIl8eAA
C03hFud/gMmtHdJ5PgWDPHb856R88uYFsenJlXW6mVvUpXXLKrzVTQnlL8CGfVr/nI0Q3iuRl2dF
6jUnIdgeg7wdNZjT+Y4fSQaC/LFW2f+ibSjH1/RphzTuXQuyXM5gQeXYJnWEOB5DyZLoV2mu2Zzk
TOapHgpkzJ7oQgw8eTu4hWx0GRn2hPh/52E+J9D8/k5E1ax4+y7hBM/KB080/1ulGgBVv8FZaaXT
HLNQfyeRGMnOEjLogKr/OHsdCLaQHfSWHRay6PyjZEnvJccAQJ7YpV1l38tF9MTcKjF2QQdbcBGm
/+P1ei8Dv0MjlESB/2lCvLcue68EPoZfqc5IVkwBaf9ZqS7aYJxkxAcxD3bVRHa19Dh9GC9gPxdn
d5I2+4mhAvfhllpxTKB1sPLa7yNWA39TgNxUyiOZFzCgT9neT2RRHq26gyAXVWzWBBjjWBwNkUPy
Pi2Zq73sslVc1b6gmM6S98IC5NZO1fwNoMtptq3ZQ5QxHcGGHXhbLmSDFK135IuWyjp5Vov4nJou
8Od/T+8kDa6w4P08YXv2S7R6mvH3t7AQGgc8gmZWiBBTOZHVEgA2csbzneica+yYo90cHouljwgQ
VE+WmsyontIryCDbyCOp+QFD4etxEhJy43HsqFd17JZ4CcCkyWP4wzJIsZicE6StBLEuP0VTMrRt
zfYaievqEtkzoeuVoKwf9Gx+Qro5VcCQ2GNkrvAPpQgrkBt/hzUXdEUtXCIxYUELh8VkenuscBA0
5wX1MKe1QPKowAn9kRFGGKv5aaZtEOixl+1RF1sq6T9GMWn+XFFwET/YP1s+TRFRWGbBlvvOm+qM
wUiZX+KnJ65vr+LWxpS1Nu9+91YRHnXoTpJUJBH2kJD6+nmmEwhxiERYaIC2k1H4baMn38zjM04W
oxh3kjhRd1XPoJ3lihH12AHjN4rW5BaQSZInSTrBSKA71Sfg9NoajiaefULbXQPTMln+Tm5ZWVQQ
a4JmFed+jVh2GUd3qq417iXEw1zRaS+3yagSNQJ41ToeaZ9NKCmROkEKiNyTY0pOu9MSJq00jd9d
Ka47uUVLZIMTCduC8ZYBTwQQWmYg1dOW5TLttY9Sx24DTj4gov7qZRghizZFs7vA1CRY5ElCZsb6
mPaWniSZG6/j8BX0LxeZmPDjWMXtV0nGvpdK+xW+PFCkoJIrYw60JMHswo0p+/CwgLR+h5iXNxbO
zcxft4s7cxGhR95Xjj3xXNy5h/LzD6kvg/8LwXKXnclIX5FY3tnM3FD0Zr/YA7K/jFRrGJDaauAz
6wiENX1NwuET4Vl5kFHeR8mRJbdCDIyi86U0NREemJvV5rZDQO5Msqp+fyk1pPK2YbKVWiZb6c8r
Asdh5KKwrmq60sIA328UhCixgOnd5A9H0bzVD5hDZgofQq9kljf7JUUhCWPzKDM+qsi+6yiHDnEK
5c1F0po5DeVF4CWrv/uJZqNQBVsjGaxhPSS5zRCXxdsC1wbs4ZB4iApAuEh31eXQZyHC8Oyc7HYF
lDGIGhn685jdQ4qmdz7rwjTRVk4ha6vJme8uCk2nMXennQ7quHEgkW30gT/IU40qxOH03eKBKtf0
mq1mTjAZgTXdxWR7YI1/vMGzGBK3xfflhW6j5HyDU0ZKsFz7Ha6CB5E5Abk1S2bpY2LpCEfSiP0d
1UsOCoKK6hzCA2LQtuoYEfBbkZhh/1jZHxm/fdaHv+PWVdgcME0kDyIuNWa0mAmy0Fp/VUiDlS3A
Stp3egJpvkSyDaEx2rhI3zsfqbp6PXM0W1JpBlIl1G1GkwoVF8gQUXPkCleJQofAclTN7DR3wM3Y
lejXvWmC9k82Bgi8FfkmLpOXFjqMfy9TrZfp/Rw2nsM6TL/e3bsgpXCFQGNvPxrD22O2sp0rVIn0
VwN/1GkI49eM/l6Z0dMawG4ta4dpzuI1dBt6AEXe/mn0/4XpUJ2U0w8H60gDvinKHU9vCsIhwltQ
lUVdYap+9E5CFvJsZo5Tbw9hXCXB5aqUs7hkhAaGvNeaA37td+xHxR3eafOA/NyVTYDoOz9ToUtx
H3J4mcq+9GebAAhm9wWd+5xvLjPxuCSqsCw53atM2ZcNId2yOxlI4sVyYawUehYxp0DeG5CTth3K
Hsi1tFD82WdVfUzdgkVVzWrJ9LAKdhR45dnWIA7O+gPxIUWXNIfuB0jtjDAjT6uJlJXKbAd64b8y
1AusdXMRx7UFyIEJW72CmzF7HRDEZlncP4mKMmNx7jNtl9up7MEoJ+wG13MGStmZGfwww0phnO28
NCKgkd7J6Y+hLBLp/Zfy5wloBiduv/646Vv8dzc3exoeIiuzvvE2WNauN+o6p4cqTv3deLTukN7o
CLZ3JC+QSlxMosqs2PLSLMdSU+qDJESCf3j9r8RpXk8+Trjkio6KG4Muw8uryOdrRcJLXRovlKae
j2MuX8Cc4/Ng+8Bf2CJZBR5r6v4BRiJGihvQRP5mfArrTNeHt1jPWcldxTKisSd5qMSFggQVypYk
xASi48gip351/F2hMGw1LbLVXfPxAVLt5H7WZAGcfmprjIle0bzy+qMl0rEVW1sViidOncbtyy37
3KufoHye96VCWtiKf5FOQEhVyK2tpf31KtcmmXXmtOGW4ik+VmVX759Ln1LK35I/9/WQ46PIOeu7
IwGGlCho5LQpFaamsiheMj5YnVuQqFN4A51DB2KyNqHvrLdCMfc4E14ds3/WqKlcRoDhIGf8NewG
P39AzEVKxoaFYzWVSjJtHn/VoGygE3KxZhcrKK7ZAk8EU+Z8iIpMTUd3DXNs1+5HgCNYlv6FRR+C
uc0pZqX+NMFMF6o72WNc8zeiZJaUfYasZNfbBdHma6Zaa7qEl9Bxkx/NqC4JqyXaVQ3ORpvdjMJO
jDrRkpk2zIK/0ehucMegMG1LHBVb4AtpkG8u3zI0g3rViyMVWZL9HugIflcmudPKBhO5quMxPuve
YUs93tS4Bge6ziAHF079+vFP6fxODYWM+5xLbTHt5K5kEM1CY7nzFqe2BRMqeEYs976DWX7Bnm7L
2dQgbs3oR6CerS2gAEQKES51hBuN0VJuU7X1fZ0N/YAETRu5IFLEe96LmZnqD0bpoSlbiCE9CKI4
7+aonz5fjGiZH714FLUrDf+Y3Vfy64W0DxUpLuoDQjlqJlw7H3T4JoKD+0FjeAX5XoWdaQqbL37P
PTk0aALR45EmD9sXe6a1V3RHv2Gm5AXjsWFfLf1VirFsLSKx5W8WLl3SoAIYwPZdWATkDTtZGTJg
nNg0TybTTHLjmgnKm2HhfliwfwkYqolXfGJBef2MxhrvcdBvnfBcXQu3mPGsqgHZrPEGEU/JyXbo
32WDv6fE/Z9uCNfLqJPv24XuyJ1q5wruzSHTdDhbS+Jy2cuSnNtNUDk3by0jjaYOOYumbg0L1mLQ
9fZPEdiRozcWFwgZb86ijfgIw2qpEUJtOHBCp2EzTabSd8qK9H73B255eduJnkpLgtEpk1Mq9RM8
r0tM68Wae2ktFodbIofMYB/6R5/eSe6r2sc/fnxaiRxEY3jqo1qfVwP+qlejd/ooRkuAPKyj10ud
OnN27KrErhndDDsNIVERU6e6vjEpWblv7l5D7SpdxIeRjmk1TzrrwN7h5ezFffZtmEVJqZteLk0m
w2GorZkBJrzI1Sg270s90CHOkqUQj3O+Mi3yQgdCZU9NaCGGUC9ff5e5FZ6KbVrCayXV3WXmf5HM
zyP+AAn2y9dR/O1bNkTGh/LCfhFsYRZvfCfF0QT3GsSUaPxFWlW1bnNwhQEA0a7REcQ8L0Pla4ZV
j0sRSX8EotVMIBrGEXEd7Y1Uvt200enxDz3on4QfuLALU+JGtyZM86OI0k0JcbJ8UMn7A3gfs7Mc
x7PBzDZfmseZatrH3inu5UbG3CVaGDU3HV3r8J+Zpajg268Wi+txno9ShLa/SDNvUwTBnfrZzIxu
zCMMUuCCz9OOzpgHANYbxKym64mBe32Sh2zskJhlZYVh+tTsLwQgmDdAb3omZeaf4ChVuPObHM70
g4ZoUvCmzApck5s7CJEY1jSRGQQZ+juo8UdpRsSQNhM7R64laBupyIspZOXFY4MTMURgsyM9tVsF
MqXmloMLWlhSW4vWnkgYrvlmr3W9y9idyX/9yNoqxmuaOuP39cnNF6GNyZExNiPslnhgu96es7Rg
eFkPZElCQcJ85TyAGbiKrWKdhdbgiGi2545LMM3z6/0usjnAX11JlWgu7BkJaF2n2O5Xgg8Ra2NW
k343oEBxG1jOvLBu6s1ggURFxhNExd3e8HpTaTcfDffSWdOBpgG6wyc2CNjBaITaVDzKQIJS+Ds3
pry0d+EldwzagEWy3vjyBoOJvNJNW0OlVU1SSjT136fCb9vrFDun1GdAeb2A9DjCSGdbZiC6zjQH
Nn/saVcH5CC1WeN0NpihkCN3dnsypXnNEIILVO3//xbtmLjJ5O/5oU3pdYE5sy1Iz4vNmhE3AaCe
OLlRVuwL3z3//gKs7i6JXzLO+1XQH03dc2ShCC+ZF/wtVAd3UzwSBAQBGH7FP8ArflvJoXgIK2hJ
kCdi/f1dcJMOhOkKGq05AZGfJzx4XcwJjRlKSrz8sDvS5CktNwXnerPasoT4OFOOZeh09iC3i2mR
zj+G3+KEKv45I0x4hSgIKDP6Fw8ZGBUtIAy5FtKTSh6sW+i7fapluvMyYfuMXbzC5nV9BF7Vc6BS
x/mZCL/rw0kumpj66FRDOUVOImcryPjdFAIIIiqoth6TL41vSUlq5ohITf4dLk31wkhoCaFvOs8p
c94Z7G6Yl4u9/wzggiufa90mhjNScEUAHZS26TcoWmdftzxgs535iRK91icNkbuWvM/Hzmcp2F/J
ODFCTDjAj5d6omj8Inu5SsFoYzQODVhENfY8oPdUxgzD5qPqUr5cork5xOoFP8ALJcEZE6h30hWN
x8s1sqfYsSJp/TKi4OF05zAK4Y2hIFrMFD8DvS95/V3bonz+6EOauIjgUpgyrSu2u7zsoEAtk9A5
5FGCs8OdtmYeDZNEFElyCij+tL2OkQv9avvJFBbCACboC9R4V0YjLzydfAiwA9RqBwYSIv3cBhUL
tZ7X0WnBrg2NnOdzepuoeoM1etb6CdmqkcrQDJ2ERwXg5k1h/PP2Yj8N+T2kQNnG38fTUdO+ri1A
sk8LFrh58lwSyJdWUHqOiljvNuTeuUYJ87it8nAmrYUWUJXmMO+ix2O+V1CP3JBcihCgjiK4gYTS
wQ3DTiuq0nsSpIv0DZw3LRcC12yxloOL71X9OaVeKkKNlb54s7Dbh4jxtphEZaDqjiLeh3DdSOAw
0kUjzBcAFmIAG0vF/C1+wdVOkh0w/aF+5f/llEG6grRxvxN+Yt5YUiW3fkqPV+Yo61p2XCk/ZwX+
VN+hrvNLVb+adQBABXQPoytSWscuXSms/4OG6SHl7p6EamidobrG8HERpGZ0cx8+mY4xZ6PmyXLg
fJ0UdoYQQKjQscy+YoxwhyxXoJAP+qrYcJrvsfb5asgcoY/u30CcGD7JMqSyvg6Gt6m+ax/0q548
a6/zXoDNphg12np2yWOCjnn5f9QD1s+f2SYlU9DjWMmNp3SPcv+Z0xvTqriGaeUL4BJkXCE878H7
llxUFGNHXkTE0UhLFpu6UXQW6MVBMRFRpcSDBUTyzoWZR0TmzFz9+b6bB6NJixPA6ECUq8CzgdPF
FdMlB4chYfedijmUqesTWueC5/Pt5fHgvINE5zasyYJKJcE3sNE8pviSxbMt4p/MMCjeKDrQl8ty
PMf/p9HLTDw8B56X7ZqHfN25obD/nTyvHzTacv01BO6eB22AXDwQqSMO3Q896nFMudW7UcRqp9Xm
qHbcbTVJ2bGC2V+aLrYMFmMtcIh1avtwy38HW7oS5dUon9oQWPtdjNE+EiS0GLoPmkr5aTemNsM1
rjAHNvCTlqKyVS/BLtmhZ3YCOcg+xAzrvjROMxGrtsuPkddU7Zy8nVjKq8uRKLkbq4lkWNoE5Bn+
eIZrp6h8w0bCJwc+bG7b+QYKK+1EXv5NW7CHz7IZKkAgWPMTKyYbnVHSCSL+RHswkCnjUiECSrMl
a4uxqxRgv5S4sxB7xFdbYBGC1NK6KTogJ7ToMZnwuC6KFRMdfjzhU6ynwDjfzw5mxvPrOqbnZRmI
gSBTB7e9/o2zBSK6gTR+lxvDOCH5iRlf++r/P1vwAeMeSs3EGGILJBis8rN65v1+6Ey1r/6jNycE
rSgNsa7IdJIGCToqKxofjlh183MXR6BsIC5iB5PPz/4mHG4D/Ys0m+bMdZv+/WHQ9XIbtwl4vr3B
Af3aqNPgtGND63zbSGRPOTwThxdDmO0qgNM7+zVwFXisbZUPOEXBThIlVRPOYtc+Cy4vDswiejGR
Z4O7gu7NDTbKxTBk/ki66J/x5MaoQgyQq6ePJOj3JwW2dGZOHtmcOJFsV/gPbn4McdZdkwj9hMfJ
F38d+6Z97NbxyWEtaCR9RlSVrh0Bc5DdD9tQv3PjvJFxBOz3qir8zLy2IcOUZCimSVw3n5+Qc9D7
OjrrnCIsOuK7JHNNaTJnlP0AKOCHR19rFx5PtoqfKQX/xDowoRg6UjaiLVJPjkFVex41QcOu8NrT
7aIOy3h49SvxdHB8hpcSOSlrfhnPR33wU0LxQ6cHtaykaxHEDxaFjHptxD/G5aKz654tZLwkaUyf
/AwHB3vDyJUNmL6ax+JAHZsXbaJUsKTn6OeLCLzs/81n6PQRN4gdJbqpU357wkW9jhr5g6btLRrv
vh75E01fgJdQRE4hf0XuUjcEiNKQLQcfrmcNsDShDTB3Be0ySHqsHePk7FudzCqsIwlFIZ4a6TVW
N9z8jA2tLyky1zE2XTllKESsowSzbYbUkWDg6iXLzN3mwgXAlFT5VRHVfIiWr/y++KNohcq/TEBx
+r9i5IUocUGjRClsrBorJBRK/O22gVu0pIyVXI4df15untCI2uONyzYhot1No//YP6/+0QDzuBoo
QVIJ50ImbuwV13+Mtl/hqras6Ncfm36+8UxDL9lH+4JrGYwMoZv96ADCvMvT5AoD/m1gbobCvnX6
mH+xZojJp+zB1GiUKsrhQ5B1x0nmjXjCyxwHRRwkTMAqs+1ODARgl/T2caLAoB1j3UJdpbIkEeo4
DyLp/qEb4EdLu8JkcKw/J89qMXh9MxrZaZ1lz+F0gHFph5p670FQF8oohyAefoyL2N2KNGnWEIQR
8yCjMDFcdcnvzNXzUBNbWJ0GNDw/Tcj9K61NigDmM2pTw0Vmr8f2ly3Ew8lGtuI1oIeSzOFB5QAZ
rpCANQa7JHHaTAqtV8nb2mZj0ov+xfwE/k0Fc9xIYlK4znXbrIzfHd+r4fb+p8Ym7qKdrrgcrYWi
jZ4LmQRm0evD7npJb6X3JQpPafqZVzoO3NCHnMGYyGQIxxNDVGoChBdpMDM6vPCfwujonNFFGDbm
xo/aTiK/qSkpBgMpY74FLTmTXdeLmDsxU0a/3BTD1crz+L7c7WPYc7UIAFCr9WfXULCTNmmmQzp8
am/t6XglyWC7SupHxgnYiYt2XgelxbqLglMGcnr1+IwsWf59+TQeBkdzUlyo+D7YWxGrfb+LlngD
wzuiRZBAbq4pwsTh66jH8Uz1X0uGrV1w2N8xap7EqK8M2iTQ+R4ZLoxvV1kfMa17u8IRiwKGNKM5
vkivxAfIMLQIT1Gjo6qNoh1DKfV8GRs1De1JlpzHavfxrQR6rDHlePBpwxctw76WW4fmx+BQHdkG
ZuuxEe2fSXysfmwnaSTZ9zOZPc8Szl8NHwwr0CVlCpYxaghOjx9QePhBeJOKmIzizFJhzp9U4ORA
C9rr8E1IEytr7Am7V8OWaHjCQ5ng2A3lw5h4pqrL1qzrxGo+xsRv9WtWh2mgBmHuMPB2tea9GnvR
Lzrdbb5D0Y6ymHDNSeyigaly4SQ0dby6ly6NEQn6dg+0Bto4SNEpW+9a0A4WrHb5JVFHvkR48sKS
uamkXVJqyCNpCXM6iNWrnrCF2Nz5mOGcUJBHgatrHQX+j28ojwUa9x+CvHL6WBdAyK/S/d+X1Oaa
zyPZ+Run6mnZAQuZzaxjeN82Kxov/PpGI5A6/OhmyMMJXS5/Yp8CFB98mx+gsHNei3PHCU9bSOqE
mA1AmVcoIwTv8ewZJWM0AuERRGd7HdYjs4ZRSqFZBH921BJMq1f1K5ZTWBj1YzMogxeG70HyQMHn
rGtRTm8Ahy/sLh7vU1HIEyY1SBwSpzg66plodYbnpotVN0Hx3EyGy+vnxoGf3q87F2jXUPY9jRLP
yXQhJRjSBnx9+sIcEyLDjg2dbvhAGK1lcLY4DGvz8X9ebECv9OKD+l+9zafA9HyDsopMOhxAozzb
Te+wP6r70uMb7VixnTVt8KDCLeDIb6kDY8/UcgXf/LVQ/h93mxVpL7DNqIgSAspxmZ1m1ey2fiGP
Rc1+TZH8Piyo1SIG17iOnyRWrPyWFU9IZlGBQ2qQbyBUeB/ft+R12ab8d679uwIEG24jGzz9qtf4
EEoDAxGlJ/gDxvtpLKz4HMiyoDMnKdMAssDDaSlQ4R2S3S+6KQQRwVXk7LmWWf0a+yFbMV89VrsO
JYpHBgT0gbFEAgdQiqVh4q2SNpTcbjBsg+E32ZKlAZHxjPVRK50xA5xNksPrtNU40SJp/z6l1sUN
5YiiBeb2UqwKwvst8f4lZAz2MMZT8vxG4I4PKz8SvocVAcHMxnZUVv4a8azRH34GJ8I6uRl0m1Sf
rxkHnP0rmSkunGmw3sOsKrdzn4KUfFhwKZ1ohZqCWf+MAQdJBsOaleLd+jG78pSBTWJRx/zFyY2G
Ab47O/dFO5RFcCkT9yAZC2UfiJ+/93laiRmrWKIbvYxtlPjWIspRKU6QJFSkaX7AlKLs9WoeLyzz
6W4DJjuJ+N7qbHz5VJjd962L6xxkahSUVTmj48OaFBjlztZMVbcunhRdEHgsqAaAfruRgaNoPFNw
t9ZZA2kT5c6y8vbBJmqJHI1QEUqNq7mbQ1eVbnlX6vdM1pMaxwhRJNvbsuqLZrGgb3x6RUj3m9Aa
1BDZ1sZqvXLcapbQoAM3Xt6dQTYvTgeeIhAtt3tnTkF42lkOlcyJKUK2bVUoncrnpQnlT5JdMjvy
sjKYI3muvsgow/CZaWM002ihMCfkHvxVNgMQHn9bECgW18JdZrafwCj/zpixftEnRBdA9dyZR6ZZ
P4o0CbYFrVNXeIF6PdLK+12mXw2BCtHXy3w5h+W4m9aylmwTVCG14+GBMb3CYGG8GvAKjRfwCLUt
XQV0Wo2va4K3ZTVukvZeZz4QgjReN8L8xtdhnbmkIr0mJyD/RN5+BDqvAVTeo4btv+V38FibK95U
SjlUsQdCkKBXxYiWxEyDCf2AhLF5YUI4hJFgLG+wKH3Zgc/a7Y0CuaZGa47zTcko4IF/AZpD4Osx
FkFF0MSC8YClJMbmLQ6KdNXW/nFuS9wNYTcoc5NFlPb9Ik2GDdaP8sfXsfTeho93hIgN/jI5ohWs
g+pYbe0BT0S3ZSw/GTn19p8z/NDMna1MXqCpcjk6+gUYSNiAbXlKKEQp7FX5+CYn0zl5zuqOdqIk
YAb0Dz0PK+/TT5r97iODGdLBbyx1s0kuUulhwImHidQYqZkpTh4xrc5joE9z+FxEgQ4icUDu50x5
L3pC/AL99tQACjgtCA37sDmiFgqbKP32wqekKzq28BBJ3W0sEqv6oALOmO86sP6SN3vWVlJaTB2L
WxrMReDkH7lRd748YOpclazJzPWGtBTLGPBGZ/7JumwudJK6L6I2WoumMnjZAG8LvA5jcpoig6NT
QVqY74JA1x+cawri6np0YZIXwIbggr+8+34/eIPOgxGszdXAn4Z/V4l5/Q/LfRmaf2FN3DXr5j8j
SF+SfrIb1xjwsx7oBcpUh25Th4A1bhZ0rvStgd6QLMoKwVdlWn0MoCKzQkldgv6xVL+PiisnAhhc
0B9hCITSRbLr44Oje8ZVWJvIUeEfS+fisctkLZPlKBjpVJ5gbPHIAf4vl0/4Ir/RYd12BQNYa7VP
V2m0Tagl4aJo1wroW3913Ybxtt/KDn20qlPnEKNEHqplPloJxF6/RKSdVMDaF6rggpZMZIr502vd
ernf/HrwXs+X6rqNx/8Ud5jK72u6aLBxzfd4Uen6C5EklTUogQNZJ9tj9W8GjTUPaSB3q+641xGF
BpDl5H+crDhKO+N/P0RMkTiS4oWhjywgw5VxSALLtROeeZ2hyXNGrmHTlLumMGP2HjurSmYqO/Gb
Z0s2t6nwAYMQGwHyiZsNl9OQYUtiNuzopPuXYm9UxLhVADN3qxKPFB4oli7HHFbabnk4cTRQCaqt
V5Fvdkluf18PQjoFPMI3FoxN80KPx9MshcnE/E553aZsGWScem4kggq9p3w9d8z80B25APtMb0r/
BEtAAS5MQAzgRpEpbAArwgFseZnjNTvSgHGtOKeTRE7Naaqz8nC3AgQZRJTxW+6pgp7X6sNwGFI7
528PVHN7Kn+fmdhknFBi9OvfCSsIFwSKRKMlHvQinGI3qZAQJ4dKyOu67YREHis5vHDk9ErB0P8V
Je1c8Ca8ILBbRSbQyDZvny5Jp/WAlobvmCTjk6MSKBegsk9JTIGTrLPzd8L6e1ojSXcVdSDLuMxR
RVy1H6IHCs2zzNwAvD48MfUp3+heLemLyXvwBwVaW6NE48Nlg+fwTb7dhh6mdDTjIJsVLig8QRPy
iBJzkPWwZqgDQJbvmC0iAtstUqDeEQEMV5CRjDxwVMD+YIza+SZjV2JBjFYnRPyYvOsFm8wadXcS
DhwklZS0QQWtX5iwEyexitV82z9M+XtEQL6zua8o1jQTBD2crnK0s7QvXkhwwTAdIIWHd1SBjuoL
20vCfWcPLbRyC0eO0EqY6A38RM7goB7glHWuWxnvaSk+xBUcYXYkPerVACI1hIKEwWxbdjR/fmOS
orgy/Ss7JmJqOm5drSg39WzkpLZ4MByZH+JRflR1+JekMT2UjAG80CUXxLoYYp93koLlfMHcybXO
rdtqqkFP+cF5VCq07/lXXjClWVUdmU0m92ETuU/Jv6dOk4wcjVbzihx5BVbOTI8Jji5ygzBk/Ouc
U8bJ7fCxZIwNReDmcl0Rk9E+dqcABLdXSiL23YC9gKQp2cadA1O13OtvdLI8Xnh4KLhEjLmDH14c
chIcLGV5RaMy5CAIZOzo/HoIckAvyHXxSyDyBhbM9+3g+WgWbO6jZ+mCiuPNfYZTPdEms2FSiScG
hPd6iaO46UvR3RLwo6qfnAXhXBCfZ3+q+cuPt3DuqvTUKlSOFYgRuZHDev8flffTGemTzuSE6egb
pJu30zJ52LyglU2jsfZXUielQJLsnK+M6xfeamoDafdqihD/P+9hFmt69lNO7T6UBmVPX2aNVVd9
wNR/La4qE/0BTN87RYcyXwRD+qgFzAz/lRcQpq5vA3FCFTzzbZJlyMzN10VV2pSpbOy4SWGNkc0g
4XbU2egmJzcwlyuDgridMf5W/U0+Zpkv4XXophMp5E2Jx/Z3HiaiO1T2UAAycpz+AvtdaETIPU7V
yIz7lIBSfJyDE554NM7SMsBa/breB4Uufxwz1bYEsRqTN+PakHOMv8Eqknevpgau99zLh2Z35GNB
ah8dN/qRi6ArsMj9B+q3srgPXSang8zCL2KbB09Mrj7Pl+6RSeog8FgZ9pJ0iLew+XwZo+1YTZIX
uBQakZZCpwtzYHREDqHo+pSiPVR9Mfwu1vC8Z4MC1JF5SiBnEpmucwNqTReDg2sXiit0Nytb3GUJ
ITQAm1/nEDoY1EggdRwI6Q4NmeL2cYlwTTCOSuM5wDu6fyvwdCBEjnOCi9wXZ9nu++5lvJ9oCycn
sAFw56iqY8yKVywhk/X6um2p4MHT34nPbl31tfwjHPjmSVW3gaWLP9HYbzMiVWK7nBS5FFaof84+
SemlXsaU7FRYgD4jo5g2s2eGYOgvzbRyyRAh+TO1osRwqcpGuL6aoJc1ajIaiGDdeCagM4Dh07gx
n5T6s5QgMuDLHwlWg+facJ45RQsdrNINjyJ+okU4EkCEGlPKBXKvkPJNEI+XhYL7ieBtzzpizFgH
m5zdJQTKX1tM5eydLOUeFpDei75ryDSN8QTvt/mZZJRxs6Vq7iFV4p4Ky+a+BfKT8dvKZnsxQjSW
zKemw5e2ynZxWmhXo3N9AeNkrgFukHvQEH9dwZ4UPDFfoAjAOgxYM0vju6WC/v5X7G93GGmofMLY
22vZ7zpoz9W/JvONMSAdyRRnrNOp9FsXBPkNAKxQ70ZOkp+BbFw8OKCkqJ3G0VuSaZGHilLPNT16
ONlMoWeZV6I+yGXnOWdSDmKiEcJqiZ6mpjNVuP/TJDu7tTWquKPkbOYmdmsUZOI64S2e23WYQ4fP
yb5MNBDR1E0QgKGHh77YoN0HI0amgIFFas2HJVcjSUGD8RLMwtVRPSgRZkxAznZxXcXXwCvq8sCF
BuWAmvjGPH4eQJ2i1Iy/Qohr8Y42iR96OO86bZOKACwQeXBvRmxIQzaGEabM1gZA+YYmep8fA5I4
HMBSjDUv55OlhsnrOPgxzspnjPsn7XTceDz3SPi6AOZq2U9xH/689vhmDSX1WNm4jRfBx4qrjbcm
lTTZLLAki6nymU2wwAZOuNupfbazvtQzSHvpZXolRNh4lW/+D0hkUMd3b2H/heungKo+Cl7uCeb6
bbG/0wh+aUoHYId5AyStkSfvYJ1K5Zn7HXVsYRc2Vi0g6OMxonJhNgiwgVBueFVKk6anfOwDlowA
gkEJmy19iqAU2AerFbjRNkHS8PssKwgNsUfF6TAVPFUb3YgdLJgOuSQXd9u8erEyGXUXzLSOGCCb
HWzGEK81cumyfVclVwaIKbTBhhv2j//TYZW7hPEvCVH74FUmLtfIQvoaxyT9HP0FvpEkSFwFN/bA
dzU5pPm09cvdSpSejCFMHoehRVmUk7mZWWzXBGJrlho8GTFxvRTP33bBHJkKcgw3OR0XSvVh5f9v
/exKl3CCfz0aes0ytt2LSEm+z4sQLROtl+ppdwHetEkc8iH8DykjnJOpuW7Ct8qj/jkr8CuJ1CSJ
fiRkbARTgNFUXTlFph1pt05zCVr8NSirdgLpALhLTxeDmzL6mlG/b2hO2vZGY9AZVfy3SPOn/2a9
hB2ITDKR6TMsDOimez7qhiB02khxDfeN6zMkfaKpV6sZYh+m7A2sAtzrIag7xV00gfcI2JnjVKcC
y1EOvOTTJM8UXR85Pvs6LfIH3/0RXeU/JCsuyaAgpZirjftIHPYGRbXdkASYp9O0xr8c2MlcP0fe
8BkBq4PXYgylNMPFwJ8DrU/hoyB+J79P3wsNZDx5dhHVd92AhJ792g0DbchCJpvYQJWCmBO0HOuN
UGoRjJ41D1/JqeSqiG1KKfVxMfig9p5oHnSgRwNwUYemBfUmKn7uXvN6aqEmiXv/J7W/Y5Aw0DDI
dDxuWACD66ZNnX1eZaaqWewWBWobwRRf7vnwXdUsXciRqMLhizSyhMA+9ORpkXmYaeZTEPiWPCnY
Yd0qaF8mdsYueck8kG6ZKFyT1FrGiFemrh4GGIshehr9WR1ajV/nt5N0Yvcq0VbfrhZzYsTHcH9Z
XXU9JxZjeymf6Kdj7fm86xErYt0Bj+eQrfw6ybcEiIpO7xzHT8oteRQYehM32ikdTNqJByEbyT8Z
ck3aLLc1/qLEFsm1FCMIJcImsWjfGKSJPVetAEHgBfdeIGgmeruYmaQIP3iQfAzt/TwX1OrXWst8
K9V1SUIJ4JOajNcHT6a8zoOjYyjffBBcLRAT8kqRwGaVPm4isdpwiDyUvnKf9JJTVJatVJartLLh
slZs9ZNHtbMLKWdzk3c4HH/IH8k9WZEGT+ePKwdsnsuzcud0HL6Yt1KzNy8NhLDOKdAckq3RZPwB
C21Ji1WXCdKDEWOkxl3cxOZBHnAlfn8nmujbMzJdusMLpYIPN8ztE1R9aNuc/bcbkkJiOz109Sc0
86MnQh14zHgRxvsNggAL7T3wgoYcU6zqO3y/iLyZXGBk7/b0XSJpleQuMLuQFyMXp+6cK+auQfR9
7VYhMi/uqg/qCDTxMrBudk1qrOjjavhNYO73g+DZKWUWZbtK4szTGPdL5jJ9L8qJcb3G2PLaCWVe
2r14fuFNWf9K4X8RYfzjCAz8kpQia3hNu7LugHauVsz10oYArNVJdbV9Cji1Azygc0K7feQBIc68
1Y+Yv4qwp7KMlqYtKQeIrbALqd9kFPgz0ZIdlL6GFqjsTQ+vDwrB4M2yOT94ia0i9bU67Ml/MxK8
XXV5iiT6dBP/bowahvjeIRDWnEGEHOTcm5G1yPnVtXsX2uNhCxLcdC9rpS1fdyic3uSxgyrUNbF7
4ol60/bKH3Q7tAdqzAAXOTprV7jXUdwDjGVUbGyeDjtZw6sYJBmfbBvs5UVpuAvZR+MhuRej87JP
gIZu5Qy++MvIDNEO6Yj9xaLJNGRTNSgBA5xkS4eloAVBS3MzGcgacI2wPb3fpbN4H1NUjBlaQqVs
kjI5EtZkI0p82VrVtpt2kASNxpQxO1dMXMuHe8gWTR7PdV90jYXL+clcSg/T5TsW1/5TaOodYCYI
mmIvfK8O8tu0CogPWmvrgVBRy10db1GKx7CD0Sb/rWhMAIq2k1pkZZIyengcBo2OVYj9KSYWpJ42
Mwq9RSpxtteIMfDwnuOf+P6bCaYAXLvmwbI7Zh8caND3t7hK6Mdam0DRbUL9nmbRqJ8wextW/9Pq
axF15buHvCOnu2O+UOMgYjiDAeoAj/vvDMmtvDtwrhnqXFIfUXlg9MI/pItQ92+Y8i2xIvNs3teZ
6VltAqnLDK5S6Bnp8vkkbM/C6hbm4hJ2YwjfrCQ2/aJHA8pPfq6nQgZDvRNjbUmA0HhctnmN0hog
28ZuzOy+ZDtMxbU6Nll9eCLy5sifLFcT9An9qshNd2GnZG4FMM66QCYLgQnSJsWFLsGWchVgKj3o
dXJaxTpHjYc6uTewAzkYPOC+uPPWvup7/8B/2Pc2V3VfnhfFwfT6NuHNykf9ykVIPK+0DR6b4GKP
A58bH0pmQ1kqQm5M/PggH+aBDDFCU+Bz1K/a/s7Z2GangInjdNgkqe4ZRfUA6jd73QSa7PKICtXe
Cugp7YT5A3hS8pbmN0MuNbaXCM65OybFGokNf9vpGSi4cYNyTAHqmecxR8T5kJsMqw+8J4hfGqh6
IIqMBwNdbYusWJBr2XMzGzBUk/GomsjH2EEBt4xkTIZxVOSmA6h5E+peK4Sv24+q8iR9jbHah/VH
vrMx6IcESGhBh6Jz5OFwlfrRLYV0N1/cfykerM98h9sEbNG5G6j9UE72bRxTWnw69zsQ3Lc1c8vV
6e83ImqzyON2KiEpUmoahEQpSL+EOPrg7hMsx0iVKS/1oqvh87i8nZRV7iKDy1qnAfw4ayKA65of
lcx98C5e9eMhVUCpqu2L5csUedwLh89iRFAvN1kjmTroDLnYDHdINFdrMlnS94G2Akh5RbAVdR/v
euj+rkSNC3GYOrpbbMZZ+1QzsX9I5EmAtD3UyPmGlgN/tp+Xr8rFXJ/H9uHbuMPbTGxvIvZh8ZPA
mjFiBkhnzhdJeXGQBTDcXcHWS0iVfSYkKsi11h2zqVcd4pd9AkKiTHrYoQaG8JIBOTWJhi4dZB6L
Tsq0M0Sk8TB9heN5zXMiHBlqhQn0kmM0jcyNHPB6pR1YAmVL57cQPxzlIZ0BoRMxEKEjtCpV1r3o
gw5id8z3oBsx6copuyHoKFN8/v1+TUhPzIIicd9iPKbvGeqkThzVFLG1bXIz4rgZZI7mf/TrIrjT
rppwlnmNOjJXX64OTtgsTsgWAisk5UX6pmuAXZX67L3h62iKjQjUFNVZDuoJBRKCPbojh06NlL0X
w59rNE+2NMPFTAxTELq4vYR6/OYG9NTOUlGcO1MdN3mrTiPkQA3sKYiNSwvyJVRpf9kMc1HCn1Nh
rkom3CQw1KRm0mtOau2NM+yMFNNVHGgKSQY8Nggxb6uHtRYd+X80jJruhrcSLrpRqAoQUV3nTjhc
+wAaLK+aIaCsVXMZ2SkBv7q8sU7D0Nxvdz4gnqVVOyKxP41sRjNsbDaVnt7B6cfzswOac4ChQtI0
dDsNI8MmFS5f+Er7jDtvcrmkb/eSiivQpvyJaUqwslfHCdCyChEfTrFyvo0pskgr9zn5Jk4TacrK
mHOMdAGB0C/yyEqiqMFQbnDFvKGJk5BValg7O5cxEYZkBN3O4v0qqbeVwqnZ43gwjK553kFDQtwk
9LI8xw0hz7egtdzX3VaIEM8SvW5PYw5YuSPuRwjZyx1ooVA7Wo4wH+RCIMGEpdmi4zSv6FwPdphV
2aOpaW+oRaCNnMNpQoRPY6Ww2oeSxUQxbgZfMv+YF7r8tr8m4YIldR64bvPdWTDrhNxytkSRJM/Y
mZBzPG5vIB+PY8yY1/0DZssaOuDz2z6UOzAz+EQpb52JU0j7R4obgP9hJgpqlhFvSZLE4AYrbLa9
kUE621X+nyzVFLWNl8QP9X2bBaugntUMx8imkYDcAb7JFbA4lR+mgDtWO9/Lf7uc26+1rkyW3WGS
CLMggrRgdV6K64UuyWLtHzeeYrNgjmZ94HV4rTG0Gli3C1RK8JZd00M5ZE3h322yWCgTUc+pObLA
9H0UXDNTFWigtMkuUlE0n8MxgeSwfCzpY1WlxcTv0DJ08XDxTLkYOhiu2SE0KX1qbGVSYIdtpsBB
QUe4hnhnq1gnQQz9CxtNsz/GSkDUuT1N4BiWtVA1BvJgxQcWaqJWYvZIfoX58wqPPgcwyf8AB2us
uZX76449hWt7q6WjbTfKTzeZ/Z3FEjU+xQ6OquwomQRGCH1iQ4lCKUzgSiduW8uIW3DJgMJQk5LR
p3iqIZE0IcRYiJyUg15qjWem088yFZohwkJk4RF3IjwIybSuegJux0IJIq3JNhwbDaWZD9Fu7wh4
xc3WF4hexeExWObV/HENCTVu7si4FZAq73QJwBVrDET4spoQDDQHrIXOOLZCWZa0BVOnWbDMX/rK
0b2je7QBvZaUjG6P3YY6pIeqryu4YIk/tGQVxLh/THda+VYSkV++lYAb02h76Vc8kXrF3a+UEhpP
hjS83h83zZKqiNWVEbQvZmt/ro72QmpuRJ5DmDlUbLrh5whWrMN7ANqEkm9Uqrp1amKJpSDr9oJK
kbRjMsmLzLhsh13znMj200f7pOc+6AQ8pOS9PSKz23uOVHct1+QcoXbQVXwjAncIcpvcYePTomdI
DYKLPNDSO9K0BJQWu6jUzReyAWfOwcgSgKHChTpkuCWUZtI1eEjBLlyp5sgJ1MFhoBYeaadgggEw
wOJhTIHBlA12r4gJFANe/jJuuXUBI0agtkk5ZaPahMw8HeXqtnAJEkz3XO7to7JPY3oebTGB4vpx
FoFK/0Vp8/ezaUl9ZKBQ5ukLFNcrtMRxVxttCDVJYutY0YAMG9NDnc3pMZRhkEz6in2WcLzo40GW
mDLPyRKKbGuP9wFWWe32r2iWyG4uL3aEjenzxKyBVenFTiLc5X34kEKVb+Wn6EH3ZMV7HHuhT5Cu
2dwixCudx6xIAkyyXIkfa8cyrFlj1TQiNjh8DtfXW9G9KNyBUM7EuK/TvYK09GVdcJU96SbCopF9
1/NIgcjsb+5COWiB55CVc42tN5C2gvg2boO83fPLeDCxrnF8LNoN8uvV3/sZqiBOOZ4ZhEgvByGh
YXqu7ShDvEtj5xeLOD/LGKe+BnbWQ7LmfXplsA4PDrj0fRs+a6tJL5Bc0uj3TwAmJma5LqEIaf8S
JQG3wen6vZlpNVYp3ObWpe0loTMTKaUB3pkkJ8pcI93Y68oUiKDkITMWbZgwduyRz63czyiSQV27
wOl9iiUAw1ndzID3Y+19PSNGJnk30EaXWhL8wZSiOHn67gRXZIs1H+W+u++jKfPRFxTUi5iIoWlv
zWddbM+xfD5sooVecGmTsoqn/SE22k/IZp5DtopZy/ikhlQ5EvExQhBSfV19nZDLn82hGW7Nqt1s
qkKnu//2kWbUnmjvyryIc21PjItviFcGBwhXTqvO46IDihxb3gen/pErk08XpRN7TTsHqnTMEy/W
+K9cWI4g96vjE3Z9dxluhcMW/y5IC1VLucyoAAmDvAdkCzO60XumlLhZTVeHlDsqsOSTt0upYG8m
YNgTFxMDLTB669yzbUlktStnjyqJM/1Ki3tjY+YIkrlvyPvla2xKMGrF8uCZFhSlFM+f4cx81Ojn
4r5m8a2p6P6PVVBK/kFzjZczLtjSalK0X7GZowzkDtBH3EyOMGE9hQTK+70nwPTw9xmQHOzYXCMV
KC570TUIgfX9glGABtItWnL9Ha8ZLI26VjkpRPeAw1sCBDw68pidJi+LC3Tr0ctubGP0DIrDEMk3
9iZdKw1mDVPvdfh45cpY+YsEgcL58V2JzWHNLcUd/uHSuD8HWoMBTMVNNei+VZidRR8gF68gdIg3
43uk0cldNfepwskkYRm9haatab1V04C09B0qtovhHBTT46sGz6wCLuKWCS+NHExi+JBtyQf6/quM
aWcHhKKHfiCy/BfGnJcjtMDXEaeCPmzSt5PCnJbY14HwD912Oi2iwywoZIdZGMjuc/LOroqCO8fh
Ft2B+/1OkZZFkfULanc71m5Xl2oV3Ut+ViiYm9fHXFCSTr5Jv7et10NpJ+OE4H34LerDc4JO98na
uXXi2Ow8RQli0kaAwJb3I/TXIzo9Rl5HduYWjeSrkpIRNvcrUrJgH468OSevPIkW8mk5dwOjA6ge
YK8pc+OFMaht0xI6A5t2qhBVXeb45khuha7vp8bhOBiTcRQBNEnKc4BE5dN5HTDUyYpUx8rJcaT6
sB2vvrG8dZdzhSrOhLVlifcu9hiS3S/IW5vVDLIR3lJpG1ECClqr4pa0sXYSMIJdIn5Yv1J95pis
4izCE/12SwRZCtY0H/7+04izsMPnAmLrUDw5MO7Wg6nq8XWZp+h5hn9G0bQW0acTZ5iUmCYHtP6R
LGFapmWb+LvCf+cgMAvmtjdnG2qACpDJ11U3g31KGKtY5L79MF07JIlErzCFOQkk6IoyWBuVh2kM
OiZYOv/L6BFl1EghYDl7P/q/5rUQrRTlYE3xOr8nhSuuqJjw9G5Ino4Rtn86k5tX9Jy3PIRGzs3+
G1xG2ZSDVZ7IVKADm1VRVePvRLtaw8cPDmS4BsxZKnjcz6F/N1iejK7gYrzxC4vgqjIAsqMdtqtU
81O3kWKL1miNAivzLAv4QgvQIKePuVD3bQHMJU4psWvub6DaqBO4gXV/suXNRxyFGu1SgtGOnbDe
h0oemeXtPBuxLCHZ3/oKumUy8xt7PgiQuqjoc9pY/y2C6VR2euo+RARWVNopfHUrDiHicFJvDHwj
bOjRqOOOm775wnjpf25PGPkDyz0qBmwnX/bqeoO+IO6hL2nY0/DvGuW+tlCXceY+4nZZdZhYjKqp
CVDHgGQ1zoVky65C0gzW8rvnLbzQs1I+GIIz5i4YSc21F0j7K/7DfHK/t6AqDUeXl4BqnDa16G0Y
ryEHfKZ1KZMZAHTKzAATgbMTZGHSJ4bcLIGkDjaIi0uoytu6kvc/Cr735hxiDsAbPvXj4iomoFOg
aVk9tVEseSpJLU2ijGVnmr9YiY9MF4z5bb5eoF0VF+8AI5jgWhGCzqdmpl6jBlOIPaDZjgTVKrsO
e1KgtKNuo/AAQ/nX9TmHwaYYfkh5qlyURqzId7lg0tqfyAy1SoVmI+NtIp03pugLmZs65YxOXMU7
3SNHB6fUJ3yXVlupck5+dI82ZGy/qnxxx8840imLZUkh7b2hp3J+iPCoZeQMlzQo0BJPa+5yfc3q
9gXUeZJWx6ZRMd4QK9bd6ahUBP6TEU+fGCFME4UVf7eOW4ROfwfdjoyYmRMdXUhit8js+UuRk8E2
fyoqTx/l/l2RBGngRsVggu4q/QOdOL7W719Sj1iGsuNql2k2syWtMYmc+0fEbmT2j7MxIsq7aOtr
O+EPeiWRYIAAT1oeUZSbHO9Hj3OdJCyd9jumPgqAKrOOUtSAK01UfAbJdwm5Mci2ANcdi/JzV6jH
l84KqWae+//ghJYknmez8W4DEqnmR829vTROuW0kW8ILPi0KI84OdpHM32HC9VPR1Be0vHG1ky9X
94dT9o3qf6k/ryr7Abb3OQpzoq6SfVAbdPA8y317l6zoPo++ddhyekO5issw1Jb+qBAWE6/vJvzE
cwVSZ9JuitC3XXw4JEx7otWff4ob+XzmYCqEiYx3WaBF5QKnBt+CMpGLnBaEgG6gXa3gacNeOnDo
Dh338fKxFOWTGMbEs/vfm9Qgbu+yJ9gMdkjUR1XbVlc6hfmNxjHyW/8p+a6krbTuNwv+c5fih1fn
tBgNNs7BerdeAaPaD4R1sWnK2UlLXdaNY1wNojp0f7HaG+g4yKjPE09m0DR7Dbx1axgamS4DbmGA
5wTHzOgdw/zogYPiijBmAyupRd8jMITL8g9DkB9uyzE3FQvZmQcdaQRQOG9vI7yKJzT3fWGL4Hz/
/kQ/dzb77etFT/0jaPddabDdFpQVqYK16dRRG/NfX7P6zTVmAFIm665AtnY9Z43a3Wen6sr//o92
UnUDF6AWocbUu3nmscdTFErwjzOJANZZv5FbNqM15mXycYV/+1i6CvyYDrLzUgbNrMVR3tgTBL6M
0vJjUElSFFPzui8DulczwJOUBkanc5wZeR/gT9VDkzHQOGKx57X7X2RcJptj5V6IitoUlxqWitN4
AxqNDhODdhracWLmtjqgfTMiLusUDTzJB+lelsZ0JP3hHcL5EE1TUyRA43xJc91E0g3gWT5UKfgw
clYwPBd9SZqWA6zRHsp2Od10PRQkTO6okWyE/yv39d54yOKe/i0ccbLfcuvNezA6lvGCVmFnFWX3
vvo0TQeZ/rRW4YkXsoAkAHcSMvrT6Cp5KgpDi0zMnpLl+Ju8SaPFmvwOrStoSskbt8DR49Qi1EMI
NZoC7pOKCLR49t8KkfBo115LfQjakF7pSTq+1ZfTnHLxr29AE1FauAPfQnvTnmXJo9Re52WtzevE
6T9FT4pMaHgjQzwrXUcDzNPRxXr5uUftci5NY3pVY2MNyIztqh8WRwkRzBveXzgqKfMxPKU7sKf/
XZo5V2+mpqT4jFtxzf3HXlZqOii8eApNQovpHfZh8rfwlGDi5AA/PnBN3F9U5oUH2rvbZli+o8hK
10KJ1dqUeG/Qj0YRARxKQUw6//yP2WsnNHfXqaAr3YLmm2/kUV1tZRvzkLJfReI8wWLSVee8pp8Y
UgG7f5wo0WUx73AlYBZAVewo4DzAGmg/A4HKkGcp2qyY+tF59LeI5hGYa5oHMStY2M9Ghg0MQrs9
LFnmKzN18lL3QXUxFK3ErvFNQZ+RhN9PqFjWMy3I4sma1sH4O1eGBZI6RIk7p9UFkFNZtqbR6wTN
1TaNfViQNBXGoVODjhRUbTrik3bbhgcTCPu7M8R18CB5rb3J2CSaDrukSwCCs8y2bhkmFPizc5XS
OzvwLOYENS31tKpmZ4NeEIThNYRMFFl/zXRWZhJy/sG0llffbZyt0AQbeUCm4p5oVLZFkQUE0Zq3
cBouOWl32zH1cHgSE9x7BSxEJN2eOCE2wQpqDetVqYyR0oGkb9CJ9XQknMK2nJyk7Wm/K5MF/FwF
Dd7wQHsR4B/qh7iX5s8xdpcpfS63n+PyGVg/fxlE+cRhUZ9QQl8C1I8CuwZ8zdPywEp8mxMjjBef
gjtHI8YgIZaFVuwhd//blYXt2lKc5nIh86omCGYqGj8ilmPZqFnhchYVygTC66d5dtNIe4AkiB2i
gjdM+z1/RaB1VBXQVP19V9yq6jfJotdC2eUlfU4nfrFhq9RVBBLdpE9HrjGSsWTrgNJn5ExjMQ/P
E99flKnaPkK7y0QFhmkmjEAYV1c9Qxm4aNQs6EPz2XvJn+8IXudZQaR6BMVWy4UUZ7BQKpe+71aW
kCPhQL8mS77laVCELgZdnfuLtjmD/wYzxci8ofTowC30+tGX0X1GHuXAXZvvfMpsrk0gz64vr6H7
rjEQw9Iy6Pv/ER52wVWNAt1obWnItl4Nn86SY7/fV1mA6BWExy4yU8/vmgKMO+aGwWyVkSYDen2j
HBq6tc0XleelEksjAzH05T3a/X4qsUWzzhbcca0+RPnk8SZaDTMMd5ZK/78m3tEzLSGesfy1QBZx
/S+Z/QOZaxf3kxsBBrWR5pvkk/1jhngSJbKR3u9V4Ae+P5PpWnLDZ8DZ9tr8YxJdA/MoNG6OVjZn
/YqWYK4btQxMTfmRb/J3p46Ur2wHQV+bDittMKynL5FSVkEAFtGKCEyGW3d7n4xi7U9v7Q+zycgy
PJCtJ/p3MM9mGHv6BMBkgdGkDTzsIFd2a+DU6TWD1YZRPwqb8w3U5ymAjwHHNm3pMI7d7PfcwnM/
JvTA0h5iirPhegqWlPsoQe4Q6Zx3AcO5KEmP/c5mOzhXskjIY0yKoVuiYYaHchTH4V6wrBIdxiO1
ZejdxI8GRItB3qm3Xm+EbafMbO9gAFB6L8oI2EJoxcQqaACA9kySsL6pzz8GM0Ke8TWAt3V0sgwr
Gu2QFcj1G7Dk5QF/pUSKvNBLMqoYZsFfZTLneBs2hQNp1reP2HpvfMlyXUdhImbyYCcqk6Aothmz
7ajk1ZFIzwuAPmB83vNOwGkSqaO0Syn2b7REyVQm/rz7IdqM9U6PxMbNEc48J1ACjh590QSm8YI2
sQu5Q9wsjTDj5enTnX7cCajuA4bNpU5glALffKPjs9s09C4D6JabBu1SKxrnd8VLdx1jHhq/zWf6
WhulDpV0ra6uB5J0JFbANRVrzh8seqUG2+P2TZm7os8CahkDI2tOGASBpwq+/uyJ+gNKFDoDGCQ3
WCKs5+xezXqqPC+v1ga5j2WKuxbz8cxbJCdU9tW1ZGOK4iMwvrucGO/J2DZ7ERdVbnIBeKtrj+xZ
sIqauqTurX/EvJryzuqt8+tbdB4D6p7lDX7lvEjTqaIE3WMFqjmn+IAQvD6QWMk+emvOEAxkmHDH
f+c/nZvAYbh0SQJs9LgQ9iCedX0moz66/VxrVGMpIzoB91R4p9q95Evc0q47ZQxIz+3f4Yps3Jmz
8NQQiGjXmsh2Zkb54JNjilDLgzh2VPA5SwZOdbcMsD3wJcm1gT44Z6JO7zwErPtavxlhci2XuCfx
qqVtZKQj486JiILGFNW+fDY/AsYI8x5FOebCSRiHAORSySppH3fCCsAApvFWAQNnP8IrDfABk81+
Ag61AsRajZ7Wc9mDOm/45Qjv0Q4RL2CKvzbxsi/R8nQMbYMj1PfpCftoW6/CE5QGsShLHp+Fj4r3
MDLYAs2cRgaZyesERdHmCzVZMDpxXZUnpQYvUkn4Erbv+OpxUW1mIzzS9XUXEKMuwrz65Gfkj4ju
j2EwRstRxuF3o6erp954+wN+63iZ4urAZqztpQ9wIXeBCkjSvjbOyS5+ZqInS6pETJw0FNErWBRb
PYeb6uT9aYLtPDZa+MVQ2DvGMj4cI0hUdmzDaIF3WZEUzby8ZGWfQiS8ORKLvDL+8SZL/w27ajqe
/zAHmmBogcBfL4nEfTXDduRtPm2efRAjvs8nGxpk+dHuxl6GdK+GqLv4sVhvszZtJGMNMLS5nzPG
eeZLLLp7RsrpI1lT60mTw8xLzV2szQN9AIpPxWZJsiguSJ5VepDv2oE6YwrBFCwvtuEmefYvutHv
iJHDaTbubFWhB+mdZ5eplhZRHG7UrDdWJYbgKRJg+V9ATqakg2+C36npiZgBuFgY5WYKocP1jsrd
6CdAPzbiRFW2/ahUcULRB23FPbo6KBEuiLqdGm4GoK/VfUJuUhd1v3aVsRQR145+Z+cXrU/T70sY
qgxMpj5k2Qs8OUieRV7dmlAMG6gjnJD3OxzLWgSmGLBgUrR2pnCK/cSedrNKiGa/rxjGesQXC5Ah
yoXpnJpRRToYPFJOTLJdGgvD/w6SUxftlPt3JoV1Q1jZXkmyanXVnybO4KE38xnuZFo74p2nUBWf
2AxDqm0nPDd3nL+MztTjRwq8qTeoZJXAh96fpEhYUOIlOWpHVkq6d70cSdPLb7sMe5cdDD7Uyjc/
58XgfTq85IEIXQ+grGaE+r8g7t90dgqepTG2OSLFkMk7N8Ey+lDldu/ZE3dYh8b13mEB7VmXJ0mY
tF5kldfM3bYgRzHIF4AkanVTwXRviSJHMhI5jeMtR8OJcxNPgbrxXJpTqObrBOP0bdlGzwVhHZem
BIBjVqiMXrGhkwWCigvMEn/LzUD/0JeffS8hmA7RuQM80NRcJA6U6omw3zKBADB2fDjaZ/1vsAc1
5AmMWIi4qJ9w5eZ1U+9Sz+W8ojPfJ3CtQoxMt8q3KEbqoohkYUq7/M36XA+TP/br4zlp59Z5VUK5
RcpC+DULdZ65K8on/xgBOKQRMe10MN0M7DeGosvrpBkw6KE3vjsunWPgDQHk8eMEGS374JKeGPdh
+b3L9czd5Y8XL9lNAAl25kuM2T/LrLT+duUtiuo+xu73ieqzhHl+9dpl2VsE+bD2WIplRE8lXkom
grAOdsed2HBR9Xf3KTA5vZvQG9fhTfgWFKQ5xRCmQDMMjYYVjlDBTjfNI9HCx7aditjD/ZhGGiHd
CUUAaKbDn2u8ul9J5xviq+MCc8En26I0wNe3uayPZYrO3XzP/0YTVtsQJNLFt6oJhuQTiPlGV4g7
35mk44OicbnIYvWuB9iePkqGEI8ZP7vMm/1dLShwKZCt663rg+75UUNncjiVH+8tSk+MMVyDtqlz
nUE65PrwTEcpq55Crd+/boJ3lkGAUxU0Yrt8GgFkFpUR39J20q4J+KqAygYAxYj43SysBSy7pBKt
I3iYWVywCUyKRIGbdZ7ymgXgxAtvlxnMSJp51StXsnUrIl5PN8pGUs+SLM5LjzS2IqM+m8Mzumho
biuXsFz5jfIfERI1X5y8EwkZ5O4iUfe3+vsQiMie+G/J2SII+F4NygnNB+XITW0FaYFAP+r4jos6
CJ/HNZv3U+34WZufg062bz9IRNuCjqG/M0Wbvg1TeogU3PQpcIBRYB5UYm3H8XzaqizhiOKBLIvr
ZKI9NYkmeacgoL9KAUGG/ukKq9WBddYjwGen7MUC994DgihuLbY6Lw5uavpnHg7V6hiGfM5LmG3z
bSVrlMH1YcxLCR+zKsnwXBKBpMj5R7wXAmlze2/6gWcT6MhjcObONB20IJk2n+X/CEVenc98RE3s
Yi6zoEfzMXUBYZD+PmG/4fCABObdgEnLHg1YeYz78PEYOIRkhXXmEpf/7n82qjxhUvPKF96DfOb0
gaToGmzbgF9P0IW+95bT/sWdoAy+9luTlFyb4nsanZ0cZgbuZHoeLNP0FnBjH5TgAa8AE0o6R0ge
FYC0ckTsLuMJg29+O+XLr74SQtWjrVeLVBjIDbXidw+RClXlMqcwka/sWECJiDlE3SJRJkQUItz5
EPHtkXBYOIND530PJmcMHPJyhSut5ZDFJHl6eZbOpRhmNlriUyevYlXotQ+YPHfEHlYOOWBk+4bY
vBU6ECYbDgqCPwWy5FGNYb6dg53rTKs6ZxDLPqaeoDLHxsnoIblzh8F6Ksm2I2K2nl22zYgbHalv
dZbO3xD5jgr8DegHY2NLEdZ0LOI8zgh/jYDj1BzcpnI1t1MZ5F+vzQOwML9U+ZdOeNVsoZ19aq8y
f0QezLov9DC+FdHqWQdnUZYLT0xir0LVvdnkflAOVC31IPbVoukbCLr7JDpGSp9TztnIqtZKGrXg
MqJri0G2z3CJGtWuHelIHZSlnDq2mPN8FrThsGSGf/VCjV06lpJBRFeEEznUlbqd23zs/jBuyr3U
ljLvCROFnHi+kCRpIF1Ux2xwjMuNn5lcSypVRA2+iu/swbFLgkH+Q0mdECdXyqR5dXuRJryKoopm
sFsWFQtmNxL8jee6Q6/wIVi6EW8ZNLdWJ3uJdrVyi3YBGwLG4CZ5t69pItFSLRLUlEaNdXQzZb0f
rbUKByQq6fqxBpLtkVZLXcggEmoYm/YNJ4kUajg3R08Bgh4J3Nh4nO+0LxTPMc7yEpPyX6N/G5HW
SZNaIhsrgOeyQ10m+fC+1bvZlV07X0pjGiztErje4x8IBQ1jnvzuYKLakDoWDz5syBPM6hCMo3aM
O5zNxR4LB9wrnUzfB3J3JseNfq5x4C3w3bSCqb8w+JXugZSzZiSaSrzHHIrtkBkePDsFTxHAtJNn
3y4EH+LaFSOdEDvq+KRSCbPGXYKPzAdUL7azeGFdKJUUw2K7LAiNG94KvML5ST2jJIRBC8Rw1Rsu
AhMvZXjbJ3g2TbtvR8A09hGurcpLxXSmTTWlXYLzo8TCpnEcd9GuE8t/kd7lOhip9FtVx5l+MT7I
D4JklYZ+StnKih5fxDrm7qovYz/rhFm2Eb9vjGhRLyTDHdIY7bdvDDotivMcCotk54cYYWyMuRJI
abVJvLPA32OHotYWdpkDnGzsKCcIBy2IVp0nOBUFJW/zmRgyCPdnpetTEt87ITnWznzBc8jF0i+P
vXUrc/lvEmryEKn0XvJIzNiHDoOFKYtATaW1etrDKy0CzCRT8GRwggQdT2XU7awEATep9bfHSeSh
V1iz+/ZYoAfvoMvpJkeOlwI1P4C/TE2W0eEy6Mc++S8L+McU9qtsguimstfg7xEU5tQ6FiXUUBu+
sm3CKoLEAPAjlbZNRfrJuaTbBxzAujvZl6nRjqC1W+ayWp9AVjJXxoYZR/Nx1VEeQSJ7anUVF3Qo
L0pP1MlRhjZLM6glqKF2T9r3ZcxyIuQmKfvt6hVVDnoLVZL0j1RYpRl8bALdJ9kOb88O1v/rqAKl
ihk+jfQbiHfXLS4U8wuqZsMdc6xhRVn/uFBqBM7KmcTH1qAyo61vD2EnVC3kY626AItdOpu79R/d
XtjxedQAW6CeWBcenpO+lR4gf6MH9/HHFr/V7DDMbchjhqKztos95QCcpAOQIJ4L8G60XSV3z6xu
wLnjIVogvpvS4swIcuXhd/Qe3rZ7HbKPIWBbj38Og0XQiN/8XBINUzpcS49OcoWJnLXyZFQg1n8Y
tsrVBHDjB4/q5LCOqYsMPq53tVCgFXmamsDVj29zByd+jDCbmwcT0ypm/4WKPqUxivzlSL+7i5uo
Hn7zQNcRuiFlc98isvLGY6pemW/EV/nIt1JpLexxOgjeEKZDGLlxoVFsHdSp1jD6mPT2V8fFX6py
/lzOtXTmEaJUnDnYhP+dbXhuNXs/OWcd8JtdgE1cwMJUx227BJ4uA6wZUljmgjH6wtM+dWdgXncA
WkRmSBVgL1MnJ551I1XZDFtv4uZ45V5TuCr1y/uyPMnSIKocb83gh35N2zJve8l+MuyYM2mgZJtc
eueT9307oWoCNB4IPc+5QKn3G/xbFttXrbCUXMEbnfFGMwEVqwekQ+w1+1+KEaD6CF8Ivltf4Jv2
Amxvj6LFJrx7lGWlfDRt+BdPc+xOPPObv3s2YtPOcOdOf93hucXMgxGkNMG5eVHgDr4i6Rtw27g8
2y6AFna4v7JmIi1mRFGOtgHBW4wDt5NsKp8/vG/soP5Ew3ilaR2LwmY9WM/Xigu0iE4jurSN18HU
9wbQrL+8zKUoGODGfz+WFycDBb9Lgt41Il/Mu1D7SEK4D60Eo3EBk4/zR/IOwBxZ1adaU3L/iq0/
OUApnvMjgvn0e5z+AybPo8jC83vVP7iI3wonrwJpMTL7TeVtEarHCd6YMURfimvTNr108BsvLHsj
mWf7CBT5nDe2IANdqIm2vHiMumDnfOJEN6pIsdWDKYrxA2VZLQqbr7VwjRNynkP5cudmfO82XI5n
s3iz6tgEggFOTAn6RLsZl+fLzax2LKsXZTIaBZC25NChclcH+Hru4p8fSsfPXhrDjTTRFI7jNeZz
oeg+JjvIFaGBQPrIIX5JFgmV/m4j8dF6wQOLIh4p4DUO67D150aCsW58w7iQSG/DNbSQ+JhY2QTU
T2i9GjYYheYK8TotH3nerzP+byHzCzf+adLS1xF5D03Lin/A5vYO2mQHi7h+3eeKVzHeEtkqGQWT
78AxaBa6Lu3zDNl1lrSgMUszNFGpJiM9GSG2Bq1T6nvWaOcAQm3yE++lcKF9z7v8IPTJY4xiEdZ/
4Yyz1qz5jyAISQt13MF4/CUe8kRnCfBSQTlqyDZUjlIomOaSJtN95z9aeWDRxY8SuYwEXztUs554
FLJ+RL86ots20C3p2p6p58nm19QT+hyTm0m6c1eWJhSYouitCXz2FUUdS35Nke2hEnqbt0Xux5ye
zN6VT5ODv87QIlljZB5/Bobu+S4KJi3IFRRP7XvU3XSoby4wbjNyOk/MdN4BO+lZ3W2QS4ENZLcB
6UKPJstkAqtJ3V9jO3CB2bRYBRH2Rv5RsJSXJeZwCpO3GsY73xExYXHXsZJAwH0lu44BT6NvGCUt
9o/FzhNEKFNWz6ssG33WWHJdTV6oLi6Kpmfzuz4BqkA/LOKYDjiEy0g0Eiif4v/emF1UjzqroLiw
mpG6pyFirWjo6QhFlVKuJA9oeYGySapH4tz16z1NBgKHIi4Y6zqaHz0T+h/nenw1Zy1nQert7HDY
jd7vhdnjeLnNbKAGmVTCGkjzbwkZcEjGyGZyrYN5PP0pAR6MSV81VWgkshLEprX/Vgx8FdlVyxAv
tmM6NlUZ0OsoVAvvvwkuyEal8xfmIDmeoIHCAQHXmFGy3XnIN36zBnz0LVnjXpKCd/XNsntLj2IK
0xG3lDM9MJe9pnM6pcqWkMqkz9ylO1NlkxS/Fdku6hX0pKJp55yaASj7r5b00lSZUjfkEtrJ4f4G
jGtl3bvnWamxN0xSNMKNhELRfilZQQINLCx5ryf9hyn/Zyy8doz3jGriMn4jslnzSTVwllo7JuTZ
T2TpSq3sU+L63c3fQLtOpL+ITNmyrE652KURnoGm4jXsk4mXvh7f6KJOD9cyUIOmkp5x4CCYltT1
sIVfcMAAv81RwkOOnA0HuNoaB12SgfMO2n4zCzwBtTBCqqg8BE03InmVcqrZeS7bz9KvfiOPHHGn
fTB5FLTtiE1Pxrnf/8xjz7GusmQvuqX+Q4Yblh3myicAqp/z7xIUOk98HyZJYtO2SDTF9MWax5l4
q/h3HesRxlpMTUtoJFPE0zCaHlOo54LeFhdK4TqfKsY2v1fnhK5K0KdMjRjgmsZzNMPRTSdr3rfK
U4ol04cPH2AsRJjuPIII9T5QohfbsHJkTbDKp6Qx6yLI2PCXmTYQIdUXPAMJ/yjDSIzQWuASZufj
0D9InBwFwDUqqPdQT2UftHOpss5JGhUdNzEqRyMqTxMgnwaDPkyDyBoRsB5u1R/sqpDx9D1ALkfS
OfRnCUJLQFNBqBQrbTMk9HsM/8nXnYDKdT3wJiBAZ2C5me7V8dkHTuk5I2g9gYmuGASfkxtfOgUv
ImfF4oYEZgd7qaFG6RmWrpFSVkVdwAPSiLIgz4X6jJxaZBt6hwCZbq9qTg2LfjENFCEBHhrQ5tJI
FKYH4pm+Z8AfLX22HeT0uzQfJ2a/6Cp64P/gE7qWmQnQIEejnp/kPST+QO5MhjFyTau5jBHheymC
at0jWLKdGlLBv7PGFy3fLCTuDR3Jhl+Gg8bZ2DsnR2Af8xqgpTd9L/80YsJ7EZsKiH1hImXFZjgY
dSEWQ89jhF4hclO7AMqbUvwCQQOwcsJGOB037//wbJnzWxGti73MI1YzS/qGLyb5i9icnHckx0xb
DsSMGgpg1gvxieZwlHzTOOtne4WXKKGFpdWHNrIRHS4IB680vtL1JVsSshBNTfcOiDKUFM1aJEl6
hzEYb1zynC7V5veq1HN6BuNcJVyHjTi1Z4LtxpnvKfj7BzaWJ4zUyNdFwc2jY93vgzR9kSwRpV2Q
qjunx8PsHY85N1/5kx8/vDZFj0MOnw5903RFlB4ZdnduzZIiQZ4MsjtI7xcWenum3/J7wd8L+qGp
ZgxceDaYfEZ7naMT22Y8bi/TD5cM3Xy2midDo9PxyCU+kYDtaG0W4dCwLvc2icCXtjQvfY+PgDvJ
ywjSfHEdGxYF/BP8YjcmIJ97+gxnTWod78ZybkR9v+niTeGUHWiW40DhJFCYt4W03mkQ/tVkEmTB
jOjdBAwB5tQRr2SRPPqyPMkhKEIJFzoj98ntthzaVIimJfVYhBT6lVnFEtQW/7PdOyai/bBaMO+q
T3tqg3iKUu5LbSLFg1KO1e9QuxFGEBHN5aWn+jwxXIXEW56g+k7k7y9s11zJ2BKmbn8FcSaA5A8R
WRCyZZwYjQ3TdmCrJriym66TA5cUgx/G0cKQ4eNBM4zjFFxbLkpY7IoCcbGSXhKg+buV6UWmtIh0
+9lbt52/OvI/9tbx3h2YVgjRN9mW1G1kpwOS1br74Ovrbpv/SaBXwY59M4HBGFnZhh/QT7tpZRkM
8fHaxf7LWQRxm6Nrs4MMr8KgnHSSEd14zeLqVSHpX4xz5a9UgXqwCTukxl+/sDn6LDlyClBHX/Wz
e1Qib0pjjQOKHe7/P6gr/cdHnAyLn4A+ThL0SBIIkvklZFh7k/U3/QNygrX3Z9mkIiro/kuVLJh2
5AL/KtAqEQ/1RfiFnCnHgyVWqx3hWdhqyEhgs/1nLibEe0j76gPGzooWLSNzwsJPFBsVALcPHIJ6
Mj9wMxE9hKzZ1aQdePTRAijpX3ESudiklq/yCz6vdwBFUHdqsJgMR3xPdUTas9swMagv7VPt5Toe
DUIDZitrLbJn7rXcvz6pIstq7uLh8Jf80z8fxWlhmpb2NrcrN5Ya5nZCz8bSL+68PvlvW3O/KGj1
1xW8ATk9Ze96XhgyQBXGhGBZ7PXwk9Tb/7OZ5PtDEfcWaHe22uOpYo2jSjk4nxVq3pLbgYsIMZou
r0dbLDI235tJCC0LxlpBwGfdfNmna5OVRuao4C5J/hqFZ9cWjMbIB/foS0QZpMZCEEzdEpG0nEuv
RYJ9jb3udBBfRisXsTbDjQ6QwuOmbXfR8CjIAgVI6bpw+7iZhoHM/aKurjEhyPANkgOXvIdmV4KF
N6h/icI7wEiIHRFzNdI0F7A5cWI5HBUgGcMcOzrc0eCGJcMh5Xr5sAoFjrkayPpGiRrEi/MAUlO0
EqzLFmAvPxS31zyhvuiPlVMThwl15cv//pH1Lv2CzZngbET5l/UsN7D3SKH0l3asRBSIKJ3AAv51
eTmXcyui9bTXJu/lQVbPA+gJnzYnNqbB4t/nwydJC7K0hX5PdOdYt4dRMbsR84wRYY12I6AXBEsO
vek57wlkKL8d8trtCPDQma9G/6Sx0iHeG5pEZMruEEcXA8Fdc7x1Sev4SWwkg4OGtZO8pYULM88z
KxwSh5HiN/tIP3yyfxU16QmdU1Rn16w9kVAqlhru/TtLteIrWwuzhIPryxp1K9nXBY8CAxE1z63T
kt4EuGWoUiwx1ZwGw88s5frpT5saB2BH6Ocz3TW31d0+uI77IZZcHzlSpTWgx+3YYs9OOgqi2oaE
dgHg8TDl1CG4L880/CzIfqbdRm6SwkqOVsENoJ7tjThFbKTWnxrRMzpgc0j0HNfVrXb+X+UqeZl9
S+Zgk1xCP6tkh0Yo/xFk6QfP55U5OjLOKMuhO4ewkdpErx6rYVPyJLkoSAsidFKTtJEf8LKO+U/+
lbqrhzjBtseFXVR6D9ARu0j12J9Gvq9elRaK/2V7Yf44iAQiSnNX6c9Yr3lhglR0IEdEJhRfB7R8
aZ54Fh3tQoKxgyK/jbj1ULVRHeb+Z81v8cwiZyChafx8m+SqlXgmwO5rfYqH+U2Lch0UZuXnxu9P
MHE6Cy1Xw/l8VEFB9/s/ZGvZBJgnONeNLOJkuTB5jN3VZxmA3mTq+aVfQcnKzoMemAdgusHrezgl
WYLqIs54xOF0ogWNFJvBUTyHkdLRsfV1T+Sf2EHe40MkJA0Ln8K0aNL0an9fagOi2/qJ/AFDEH1w
bbPMgBuK1PAuhEaGSY5F1O0K2hRWaCd+D+H36MliBZkC6LW1zsC6xaWpEvHfISr5SYEw/qDPJIqC
PG9lk6glc5g/l0c/yHohpGnxh4OeBmUqHveSZJxPkrJ49zcjUFYwoYs3ZPAhnmCsefWqb4Nse6Ru
vzNKHOrrwDU4O94aoNQTzj11kMEp3v/EW+qeITolAKRs/l5DgLrENeJY/U8Q6S647sboK9MxmENj
X7/6O2/vXjU9CTft376EijCGdskunPMJscOEQhWRZ+Yx7d/Xoq1ZyqgEvDFm9nW1LFIYAGdkCQZa
Zmpvcy7oI7mgWrSFkoS2MbsZPMR3d4hIErddYXPJ1+slVeJ3zGDp7MQFMQ8bcvhYSC5T/Hod4EU/
/R5YV8gF+stq85SwLywBOqCTj+BMMeGyYDNRR4INv5KxF4bM9BH6FjF/J6Iris9+y0q5qORRvH2y
HgrjVfSM+++mBh9N3vffRHI0E6UTeaRX299xD1bshsRApSEJtjekIOOMQIOXf6g2QRcmiYNh/QWd
+NzOaoT5bwvhwm/ZB/3afDAEbXYMg6CSc1ugmFa/qJp23Hqar1gx20W7EfllMQFYhZR48/iFwJVK
FsS1M1PGlGK9rHnOY8cAh7FGJb8P56ykzOsVM+IsQ+iABIZ09+ib7MvisMKEUnXcHOJaAnV/eczd
ia5NXTd4cHqnNS90cwlt6tZsixZLVlMaggw2uM3uhgYIa8d/OhabMWQ7uJlKPTk+Bo65vnBxiyqi
T8T0KvcZFbd/1pGNR9EY+77OZygadJFWumYJVSwZHJjOqtv2CamV8dIAWRCexTJqt092CtU2glcH
1wG7W4SZwKjD6Ladzt1X5dHqR5bBPWePgWsPLz+CnAelDtGG4109ToNvB59QRZsyRrbaMN7tkO2e
Wh8JUpzKD3GxOhcI/q8zUPDmuJGQITB2OcIQDUZ418KwL9UROW387Gw2OpBkOtQC2WmR+4O4wTlu
71LBGZKgB5VIfXFDqHjhKi5phX2aCAYUpVM2HhLtnWayofBznxaEn35iUNQJhYn4FXf+RAGhruCS
QDuRBrDQsVyUwlOZ+VmdHkVd6waYb1bk+/lDDMBMJlGIFgOwz5AHzQPzn5iCPwC76sWp3C1gB3/Y
0smFdnvOwh8QjhUDL5EfOP1pqw8maMsyMny4tuVesL93YhKy+yPnYNsAnfV4k+AaQr1neYeM8DWW
QoTMwZKVjN3Mgzwgu6D3WJY7slgem0UWIQl9AKygdPXRkJ2SXlikeEhGLlmxlEcGdb0zFgGnj6Bq
r8i1EDlvHlvWLPC0tAjrkRBgVOTGBydXt1VqWFApDVe4JY2cUlNkmhkkdmcuCVdM1FxFcmZprf6a
gjweDaGX8+RXfabkXiLQK7YRcdPqt+Hl9mrQpT6iYwxJYtOqJ/Wh1eV/fFgXp7kEF0MqkJI4rLTu
16Vr7ltqXQZDgdCcmm2ijoC+47gS08Z9b1IF9XGqXXjrYQiqO2+BPp6q/WFm5ZXglu/2XjAxY9I8
FbVsEZrHrGp9CdWS9YaTwGpFjrBSOOnLuoXhqsDf5dyTvVEB1BlR6RChp6KGMHc11kfY1TgKiNpu
gpNrbx6+sX276uEATIlX+burVM6hWSn1Q3z4Yi8s36H8ZmNiWPx6qsPEbL0rvHZhi2m0i587uRfw
S27wi4mCfi+BVKmg38jFCLAkZIHqsCkK4Te3PlCrgUIKfAHsudLTSI2HWVeN3FQ8ZWSa+6kwgEvF
Y4l+sWAY+RWfn38RFIgWxB9w3ZJjVanyiAiOnS70dJOChPUwv4tpyyZZsTypM+haEGmL7JeQN1nY
lHbUeE81Rtq393OHYWNWfVQvwhkRXhcB5XSrTYQ8QXFYQDppiPRVOB9zl7b5HEndvNpntlOsnmpq
YOVhmD+fR8uF+O96ZCCU6m+RlDImN/zTS0SQ2Hhclo2jRtnX1XxLew82TLHS8AtmnOGTE94ePgeh
9EFBum7rbi3WBXEcLN0L1GT1a20KzUlTSjkYfR1U7Z9ggIEdZeqxNr4Q31391W64mW1TzieKzAxJ
FaPD5j5Ncybic6xVEdKggcryz3PNfyrHtIotHd1HuPTRS/Wq2I82372+AiC6MW7KcRpPdjoHwpdp
RYdcQ6QgnYDDqxS1rvP0si3SknDHEZ5y6VBDKV4RrTZY+e3RA9z4a5IXPW9lTDOK2wGES3nQ9nh9
CYO6LIjWkc/GE548mNHXIiYlM1hJCjZoBjb82/H64MRaOpXWTPBHxXuhkXemNYTlHBXJGlNingpQ
3cYUYWCWe0mAwVU+KwwDAbRP0/fZJwjbtTNar2CiBR0hxVfHx3Gb1nj7TBBELABemNcF9U8wCSXz
bJ/2jXV9GDikzXLnSM6hYMTiJUfHEkSSw/VyfLxJsD3GIp+aF5VXLB39W9l8cueuW9ohin96WN2u
qGDzuveI97BT6sxA/GJih3sibYSPgtRkr/YXH773lCODOdKFoESSzAdeQv3cspmX4srAa6WY+VnP
mKF5wZNDx8rW/MprHMYrhQcQgfXj6vAm7dZgVtlx9sbd70cOpgYwRFTI5mAJIgrEg7fa8RiFCnJ0
JpCf5B0v2nF03lkKpwp/RMDeBRlB4+am8k6mAIGNkNg+Ff00dzssVpbrRk+Od7DRgcS5KM6qG2+w
yem2llGrUbvWnv/D4HP2bCFCZ4h7JFFCEQQ6jPpHd/2TO1/ZTU/bWZ6kH9+MX/rAe8PGfcwZzbbL
tbiR2wdO+ye9ByZZ+ZPT/sdpNQVnQxq2UdwltAiubTYY2N6qo783y8+1/daTYTvn54HIcOSgY1p/
FORR/kECV9GehwTrvoMCQ4+j/WbGmI/BjIRaVXLTaHWfhUFA6ipNZzhBr3kSY844N+VyrFhcau0M
k4u6tZG60kf5daUkaJoKW++IU7zHaHI3DJfHtBbyfCyGRbN84VPBqVqGPz6x5tFyJf/a6o+a0UFG
IuRdJyj8xbZ9YqsPblnNxbfVCNu6o85gWT122TVv4soPj3ZSWlSUQdiSGOunS+pAzheifFLM1x6E
oMjEh5bvMdI4UWGzWHObpN/IP4OTi6+TZPrzCE938kYNsQKgRXfUyBFeavrkR/b24IRvvGgOo6zb
xLUcwixuTi7p+0bW4UgDSfTexJF6cUydBWNFSCPg65tMt8uHRK7p8FPQOr4x+wIFY4i8suT5Qiap
eLWZpODliAZKTR8Jklt7vjHsatlRVOWbjh7YEs1LRVOZsOEsg2eCt9Ca7Dxcdgym6a+YA7JwPV8R
tv1T/8smKrAilNSsMsf3ukXW5ytEZIa2Voi3pnoBXnuaP6bLeksfM+pyagOn3vkBm8FDXj75ZN01
4XrLrG3LZPZQ0Ehl+UUWbs2nJuOxz3I6f0GLZr/RyVko/qTU31ONXtIBXJwPg16RBJfRp16eh/LG
tMtfcaFPL/rPv/NoB78dWRPTn/xVy0iLo6I9FR7YJSyia3anj4u6WpAkqQppokC7Jy4bbc91N9pH
zYANHg9/cCY/VW6Vnuub6shxdadostaxa4DsDh1dLUTxd3TNVW6FhvkPlCFInGFDVA2YpW9iSlTf
Sp+w7aruvy8bbOfvd04l1N5KPSL5DHP2L4ook9GupuexLqXkU1Y67rFOkkhmpPfxduQ5zcYhLLrW
1rI0WqW44iyYydnHURn6LDonXJRWGT92gJkqTP1JRpSM6qWsVvgIMErHNp+P0ftZSTTIZ7K2ytfL
MGkSJD5IdsBv8H3iujvagIlFh7dGYQgs61mvpc6VJEFljEHdqWWbhm1YBfHp6MVJ+yuTv/9LXDCF
p5GsR3qO6aA67F08TDJd2yuL9W9vNV3/KdMinSzmfvgBgJ8DRPQBadvUa3nHIt1v7roN2aaJGb6J
sBSC3e1nit8pvoKIc3bUJ1TiH++e/9sT4iM4qEHNDoUE0Tai0hnBRalAOAIKja/b2D4AjLLbHsJV
WG4IAa2tXq+vDI5K4oQXDEndgewVwHVU55AZuhHxALuxN5jbPNzeYcmBE3eP3dAzBRdcpgWsG3TR
592gOpKeCdAYwhCh60C+JrLHLJh5tel81nFg6+PoGtgMAAkNpG+Ozt/cYfFhi1+RuB0ItB4aDTES
M/m8z8F2b8YjYR6gaBsjmUXwDwluLjrsvsZrlx9IojelRqOBBCtdZ5so34TpkWQ8kJpKR67mnpbk
DDhLbQqiKAvriZOfVPDlpvluiBhafI5F/CeCV0hiutE7SpsW9wT9iIGvRvavCXF90DcO0EwVRlAW
RagKbRAAPXcG1/IriJApSnPYt+EZ/GAmwXCEmC55eWCXl2f4LMuBhSkagcx+2dmJy8Id0+QEVOC2
kYTEdVmC3Mvhf5TW2SRdOuvWZiutQu6+RAc/euxCimID17nEerxvV4cWn/pR/crJvKrqRqVtCWr4
MrGF9jevomprexqib+24mEQZhrxLAd0geefsoLAo4HK9Om35f2ey7Ha/3vzhKGxTi//XffKf7Y8V
ljL0x4nnsL913Nw5jtQdHBzp1uoLNqJXucm9830pUsyLaehte62YVwJ5e4ykNQheu3fhoL4H0gSA
gU3rHwBA5yYlBTSU9zVCP+jVdE37y/kQMHP8ATFv97OGmwN+GjvK0PFwWOZazerBcT8WFxOKvE+L
W6iSNttnnfFP8oBq93RDTsuXnvmXDKGbSp86A8jzIQizUT+lclU9HzpflxHwmfgKO3JQLNKgs8sv
SLt0j04Z/Kg3Jjg8yq8m9sV4ZW+fNOQrjWrpNcBH68JOj71XylGT/uX7XwvnTqdVplsdeujq/QPi
pvllA5LTYPQMZ1VQC9zSAIxCg1wHPFFOZGXZQPv4Zfjz8pMYjmspyzxH8hePma9GxQfY27uH3q7H
J0nHa9kiSPjg2E1sqpuLKbCqHQkBGRMta0hMC6z9M27r/N0AB2Jq8rnmcjElJ3enlt2sSvt9IER/
9HnNj3neD+yuP8vijW+Zo+W0VWMtU3NLS12JjqfsvdP5GHdzV+7sj3knfmMm9Y0ldYuGJiGd63yX
XEMyv0Z2EcqVeNlbeJmKiTqSqtXPQl9lAknXM+k5NjPYLebxCVsIP2Y/fMA6ZAGXA2ucmhr6jFaN
sq5E0wLY0qSblmwmFA/f0VTgnae13rY/3m4bWj/J06JJh6ODnn3ZwBL92ZiGEqltRQcXUGQoHVvx
RrIbuU4heQtX93uJ8xbB6QkMyyEurKORuVpbiGpKBHzEIncsie5gqM/pdRxnjO3g9u424FvaJsCi
WLSUwsbK/EKxDetr9ODtmRNxWsbQ3JL7yCegK0q0a0Ho27N8SCDZ9tnJaWHRlA68zLJghu0H+b8E
MLUBNvjrzx+nzn8IRHtBdtnJ+a8yklkNGTOGu4Mn8hcabBNgiQIc1KL5qKQiKDgjVsokxFP/OBBo
qlcpkiOh4GsXgu2bgD9SvInRLjySF16Qip61pkDzZpXruuE3r6PphYr4Qqj2Btt47l1TJeWe34HF
kI23qkC6gZXdBq0nwpJHfuwweywmXNq+oJFUn7kO0BymTI53TN/I5KYtkqzJKljZTmOpVKj9TSI9
WENZXkdlR1r18FK0Xaikb1UycQuVBxHkNTUQ4QWvgXApcorT9DKcicA+oIPdcbn0LlX4PychcTpy
QR9J7i2cY+BT9JyWW3aBLb50WKEHQ9iXay6jcxFe8wA13XnH+pkMKDENZOJf60mWjmNtYWuEFqjL
icHg45/gkOhc9XUy4izpqnVZWWIsOePqFSeBVVSxB3q91RJ+nFwV8UXi1Jbw7M9OEDsJg6ekY8uj
r9exdtD7gzHhe+MXu9VvjhB0RvYsBph36/ThqK9jK7BnaWbA4XEYOLm2enEZMzHLHgGQMaANQH+y
qxoon2kb0HKlMIYJiWOy4Z2is3+c2fKOv0IK3We/XBf8Ea+uFUozzTKx5b3qkBGo4l1WERFUsQk0
spbKvRNXtflldbGMDviFBlLT6WyI6mDvwQ/NZOBOVMUzTceVM1EVgQJahaYnt5lr8SjVjVF9z7ul
G20okaZffxkjNqH9OlQsEzH3hvwk6IietyIPbVh24zc9nXOqvVQeQ6T9pYRuR0+RvLfdc3olgnlV
edRjUzJ57SxfGpzzOKOhm30RlRGwo2nmMVRll/lQ6pfGAyrHLug6gx4JdxlPKt67dwjtHWvHRdC7
P7TWjmEWNfd0YMh8MA0y3zWGfRT8ZSrdD6/TMjCyC84isHzTnyxxtvN+7cMHutvqkca7UUHPkPoq
7UH+Q4IARN/PNrol85YkvuDPmmUvwt0qU4MSW8jciqiul4JlP4WNbNFm/yDL6zP7uo9qRJgUaTT5
80LBLRQ7eWrJ22fA2TMaYEleCQSSD+7F6sKq0fau1k5DqvT0RSPV2avRefwpd6F21zKFZ0QvTOvi
bz9CwsptYnscrqFJIMKly6Pj9GlxEUm9ZvGtjkHtK2bQohVkl0RYmK58Ffd8w0+KD6PFR4oUjU+F
eL991++LfGmeHQUQD58CjlRZDfj36ckIwJjy0bZb8rVVXm+zHYPoN4YRroqI5jI7EBKEOV+GBtPz
WGNoJ5jr7gRuLXVFD3QNOCK0XoX3IP9V/BZR6cEomAOhZJLhI5r1JI/nZ86qXKrntTiBkwYu/Rvr
0witrE65qZX/ZqK0BRJhkREF4bjg9jq8SRpXD3/epxyPa62gcBGlrsVBQVQRMAsRIMsl34WYmhfi
pfqsxRA1d92Wxqk3KP3J/Q+T4dXsE//B380bV73o2BKQglJaiijusQ2EgNLMyOuD7UPFwkmF0a9A
R+6dRA6GTZc5Pe3MHWqZfvOvDJfF8tSckoyFHLkuAuke4yOEITCQKdinZxgqb68sJzLMPtby3ZM/
oT5FIgdlF2H8aswhmzhi7EWVTrRocXU+oKcvHSHxPyKSm8wW+Sn2w4rdvSiU5E8qCg7qhRxvGnBy
0iiZFGpVvmMR8CY9xli2VEi4C+6PnHj/F4rrmPdzZq8QB3IXXN+iT1M7qSKcj9KJ994hCoDx8Qcq
5twXpVSOsQfIo6QBZSLhsLPlXL02JO8XG5PbTnyH6VPu8o/YPI9CUpks4orw8P0GOF2z8pGhtoFM
xN4E6iNO1xlvFtYs4jBgnEQZ0byn1nqR/6B+yt290ThJaU24oCEFdFYxu5bxl8lh4pUM/t5KBoCg
tiIp4fTIfyXPoQH85QAtz8M+DGMSXYsgdwL2LWZkiczdl/xtv47yffPIWtkzmWn0tZSumFQKiGVz
G2ZxxGEhCTlO2e4Qeix1/iV+8anB3ZcqETDru+5r8QirNWvht3JFTwysPPecB4iuq+0HwZ2WODpv
7/mndK8TCi3fbyLhaMxk2ljv26RJKXZjSGkTCB7Q/MYbtmba+JF8q3Ox1WJ1Fak2hijo/5xBESks
yKImxAmjv9tys3EJv241zj4XFvueS6wsem3NL4OFwStikwwnHzoLHfKalcIyM4exQUc3otBUdXjZ
qV9tSumW5c8OPSsQer8lZw/9nyMwNO1UcTrzyNFDQ/JxIbvHI69qrz6rcTp07pi/rfSLpWAVqEfj
zJBqMTEJWiD73Q8AGCX7ml4qQmEOcnptrhHKDlHhH/XN2+Xqh7pdxYGZAgEetpvbtxfgFIeJWY7G
Ge0kW9kw1ItPLVpyWQx0iIbdd1/zjKo7Bu+NMlaoNRaw3fd0Wa3N9PC97pfv1tEY9vKNZrggc6tP
XC45vgQDNBYjMFPOOkS6mRB2BY0wdjhSlpkGQspfUtJyHA7ZnDDQATaDfv+Vdh877OexBMkG9tsP
uOGRrcb61Y9DwnDMf0fLn59MZnNSDzfPbwJFhvR5Fz8zYoORAXnXbojALygCcKe32GLk9BLyNO0x
ezOIq2gH11nwdtRV3cuFWN58wnMRdNouBqNYUnLG67ulYU3OrcPOypt83++s+NAPk72/KBSsnevM
i04O1ozLWdP8Y0zPl10wp093GpNyp4LkV1dDz4mT2jAN0vbGX3Pfdm3vOPYhjlPtikaUErgfhZjf
WwEHdb5TnydyKoHR46+pyIJ3JA46gbT+6TA7DN29hUU8faHKIWUW02NdzFfuHJHeWEz1aWxUdYyA
vjP070PtjGvyzIFrtAxXCS8badDKHZqOD6NKk3LFfovk1KQF6nHKSmpaWklhE8k8Yhva/ODHS7z4
GbRYc++nvDKXGe4EaLovMnDDJ03kQ4RCSQ1osnKaDeT9n+N1yRV846pKwL3FLc19Tj8eiGWlBGjR
QSeg0v7LfMK5HER5MLHqYqK58eXnavV6XqscIaNHjLV+oc58Y5gNSXI9fWQ02kuVzJuGpoj/7URw
hrCkAkEqqZwl90SrsCUcwYwyp2xHmfDPL9QHhxaDF7eukRDYbkmvNZ3zXj66Yz1lOAfo2ogbRPvK
HFchQyFhgexag2tO5Dm/K51K1YcJJCRkGomEzFe2v0mgEh/GqdNbnjO1MFEX9NZZtPi2/qLIh+eg
/D6lP4K4RigDNyCmhrLkfM/biCk3MwlUu+t0Eq5yLLEzbLzEromvd4AVPhmYnwWbsxxVlOD0cJx0
B9YdniLLjSake3eviRoG97Up1r4PhM4341ZbgMU2TTIg6H6WM4VYtAfudtYflbtkw8KdIAYOmj76
gKiCrfwA1vqv1KIBmYASX/N7640ksb3YspzY1T5JVysYEb1Er8h9inIf9oMC4fvtpf2jE2TkzxwJ
C3DIfbO3T80MpZvoEvEA+Kr1OqD1OcC17DaBQOZKhkf7nEMXRiARNIMrBSQf0EAxKQqHtk5HiclO
vsclWmcIqUbKNFyAnra1FlYpDhU3YmarpUH5U00Bc6+58+rnm/XQstTICAGWsELgsVEdQW+6z9vY
sfuKgFW0WNMeopeuoc5NcapDzQOThFzKA+SWOZQAMFWotSFsNZe4t8UFd5kIoTJJ1OIam53s9lEV
zMjZu36rUsdQiyaNkmzBvVFL6GwdrmpIQGAIZHfc6pJnzdYm9f0XBkfglHbgd6uxJQVxI9yERODb
WSqBueOcMovokzUEnvrp/nUNSumbG+aOx8bQFh0AEGEKSGhIZvwJPIwM1rKNADgBdKxvbWIUJKWj
GUmH3Qw59zaDCKWo+IKeGMfPjRIqNj/McIgruavk/owJVt3Fdmx91yElmQDyYsfpev8pAWiV8iNV
ZpaXjgFeFXEpYk9XfRA6NugDdIPmuxFc7MD9qQZ2Z4536njmgbQhQFIb1ch+tfSwvxzRQiI51ZPn
xsIoc8ySdS+XS3ILjojsjumYVIgkmUONmJa/ey2jv6xs8zlIux6JwLhK1eplKLb2U+/x9WuXveW2
Lob3DK18yzvIH/KuyrdKAcwr1pF5cNu3cZx4X/zOZInJC5tHZIWn7DDqf5DfpH0oTXsQjrXT4xRl
1BxaYobWwIXrJKzWJpuHT4tvOYpIXjyUJjUtVlaVvFrdE0iq/rDxACmw0nYRswS38w8gzun90OSJ
E6V9KGFyOrmMeC7nqKWkoLsmemIGRY9yN9cw0x/b4jLptAaAlrAfGte8xAmhozKqUxOng8vn3JqB
4oSNkw4J+vl7Tl4xPYTpjWKYDi3EGljQ/wjEbe9/5HSDaFjIjM7/P8NkM2HD5il3O1Y5Pnqy44Nb
+sBtGnpm9uSB36cUAFM6qqBFxGcOi0wqjSeUMv/TW3xm7s+f0/fVNNwJn1MygGMtEck33LrmM0Gc
VAhgW3wGUjvoJD3ClGUP6fzhvLY4lvQYKfvGQwI1CekHT4PR/e3sijNmKuUtw6lTUIEYCuonxcET
d5/Kxkf3jc/lKh91R59ohb9y9ejRU77Oy4CUOqJiccMsQzwLahYH4bdKCuAcNoMZa08J9qwJsVRw
J+1vWM4JNk6hC02U9EL8CDj0HGS1bNOyN7fyfTSqUGochuCA16hbgJZwFnmhurZDvZ+rhHHvc6I0
EGuhs3EPtRzswXzlXwDl8MIOR8isy5Aghiqf5IFZXGUwUeYlOW5g8DTYwzNVxlK8jEuUZsDnq+Bv
KZAhB3s5p77MYnyyH7QzTwaasALodyt1vagF04uRtu05b6Mrc/L3klriNVlyB2uoMNCFm7OkGSom
2NZqzsCCqZXgTLACK2n1dFEDQInKQaIRg7SrOYChVKyOyeT3aENHpsQplcUU/PLKWdYGsqfW6g+W
w7vLPJm9/3KaU6SVL/bn4+NxaRS6XoNu1BRwvHR18rhnZO1QXtCHTdnysz9hxAK5aEQW+lW6YFqD
4gQw6Ta1vZxzQYM+3gXIJ+Sk8n+vIiYhwiYY/KCXpVDXchH8mIatI2wPc5miZdSGDiasL6h8F26A
CkBe2HlOf0+5gBSjQuKSAEL3tf1D5Ig8GbguryHdn+NldM7w6Capd2TIEy3j0bpDRY8w3IW08iYk
XHFX/N6AmsZSuDKth/+IRsHUT3g68jpDDQ2D7QHja7rCjFGy30FIQGXg6CU6sgC1FZrTKxRvN4St
fV6NucdJ/eYnuTHCa3t00pQd6/Sn08wGKdcORy5BhGJlN10pst89+YF8y4ulB3DWD76/v7qj43hG
Jo2dhf06rAAuCCWoAEeG3m0K2BFORVNG5zKY2rh485XcocyYn3yP6EP2nG4hoM8AvdLY55RdLYfU
tknfDtak/JUimBHGDO490G6Oyjl+P7XwCLbENuJafD43jbMh2SjmeBfJLj/v+UXZGY7CzfVUD/ZF
EzHv3F1TfJfKRzGC0lbpiax/QV6TFKVs4mGyupRodXYTLe/emjodfk53xV6TTqYHtZMeLYjg+ols
8M2FvW1QzqCp9uFp8SnKlDFLHNGNSvhG4RuF4HQhoNkuGX6CDwQaEBquYdQyyVhknaVjUIdcMSkN
9tLE7yLrLbtf9jbl849dZLE91mqOx8ttYyK8DAvM//dI8o02GSCDyTT05sZR2ITbv8o4CKk9EwwQ
dGYI6FByC8OsTZBo0mboC38Mu0SX4O+veyAefagCpScL3UfP5DBnGFz9HGvTu7JzO0+0R4v9aVC8
rJztWId4orhce87ZUIwXY8I3mbl2dqpVqmEBS5Sm/qfU/dTpcerxqJc8TOPOTxOaJuckiDV4abCV
qBOS+lwgzQNEQ7rVD4u8lOXyUyQrLyvnCBvhqFz2q1ZrVO7snx86vsGyY8rUibO75pzA63gBpwSf
+DVVYf+uyiZjCpxwk2bTfxOPY2/UjM1DYl1vAHGzV5H9W0kejziEA2hPTIeZ6Xe84Jl7vaNvb3lv
LYNbmSnDdrFGP8ws1nXobgiKJcesrZiMVzvv1vjVl/pCOMa1iX4TqVN7baSUHpHhvLku0PFkmZlD
mZzILmXrtlN5YuQxrqOacet0ipgtpXCGZXZEQcSHA1cs7pJ3M2b3BHxr9QANGFPpP1ChW65PHeku
iWl1AcGoiJGE3t2vg0TAS/Uswp2FLn7hQ9YxLkJNG3yIlmT+yLOQVDrQKj9/DNKWKMn6dQWhWg+A
DkBRo6NxtVMNr2ZGS3StZeiQ4NpZaDHQzs5UbypxEUholafGhjxMLIxdIMEqZF1M836R7QyFO4Pn
BoSzFBu1XYHvyTIwRhIDwydDBKoAxs65yX2tyyi+hFW/IG8AmPuLUcMq9bLWGTzLiKOOPecgP8jy
cTmHWlopPbkUj0nKsu7W0sgGd+QI+vC7sgkmezCSUxbIIrQ5gsa85groR38E2g34WCTp2fWrJ7NI
SW07OmMXCvgUzjaJpGoIGGLyYlAf3HNuvwEH1/I5xxBcZmSSJpHV0+Wc9zg4FpPWXg4/MbbGygzM
CZfFucsggt+j9X64T95WmXFeleB7ZGDPsaMrTDf/r+DmMNP5s9PeYDZAtcMVyBYKli2T07zuXp88
nVFCtczZP6AK5TnzMCYGAgQ2hYVHzMXlsw6uXQBRjlUldlr0BiJFaY2SrR5jTWiIOugVYdozYOCB
Tbv2ARwpJ08XejCUVH0Yb0ymrGAuuO+BNhUHLJe+yFo3V51QDLr0eLOqXlYeaF9qnKDGrv4yB2Ay
5lQ/2lcCMAbafpx0fKmELD7umcEHvfiiSM7hZboJCSZnHKWmzW8t/R3ErhHbOaUQFs1cNDAhYR56
fbkRWi570xRRlI/n6mHCsDY5muvx2NIlblj1hP3SQCoy3leAkrvWXnEsoN7S8rXY6dl1p4eDrL+o
8KTyC6z8dXSV7HIZ1OmyufVEjUHFQFzMdubR2/3OuYGkuvVnovYv34wNEeN6HsFHABpco41vh67K
CluvdEAA5NWlSefchBPJ4UaOHFv4nZOe/9nbtMM3iazUEaHhBGKhADVqWIFu2qyEfLVoiBAEwWAw
dgi/F+0BuiEH3xrwbY+BLHycObb+W0Uox5eG7r4TVyjTwiLCsWNHU0RqpzlAF2PAjn6c4rastx9s
k1QSp4uDgKxA2xnd98pIIX87JL5VDegZRjyli/m2dvUr5ONq4sOu6k0iA6yTFn+FT6bbvszuzmS5
HEtFpdaU2IiDoR6VLmja31lkp5rRUCDqJYJXeU9opp6yBf6GGV9VFfVGXV3VFoCTvaxyzRK0/CGJ
F6lDmx5vopxcBusBMEYnEUU152lSzI4JBo+esHI+O3nBa41luRmiQ2PY78DMEglWEac2QbZlvp61
L9C2d9knL2cJyKofOiCDyd2kjkwogE/hZmf6O5UkyGosqpSqvXx1kE+FrLz7SKV6KbYHkmfYE+k5
FGCSYQ0QOrAT5byP1/OsDYuvOeUCIA2ICtie6dDVK4OQ8kcNJr/IZOeM3P1P7QieDJW63f63YwE3
+bCSsGAzi6lAfoGGiWToYAMkb2+IaRc8sLFlh6VlvrZ4O96vegyFkQ2MKEy9tmD7cKDIz520nsV9
H2R/eV8zinf9U897pjaAgdC5FGTTfkpM9h5SYhZjbEBYrvlR+x+z/BYmI5A4wICGcbWA7yqP/fBe
q7UIJzuu1smKKql8h6qn8CVjHDaCP10b0GB8/xCxwhixzVonfiClho70JBmYjfQxERr96Z5a72Ua
Q6Q12TnUdq/5gEcBMJGGvTopt+S5fA6OD7l8LwQpgo0lzVyKdBce5aJOuopsTfbXP2I9P8F9lmZb
SW0yKMxwA/op7Z0JtzQu4J6LEff+331MJS43hnq3RmIwGnDke8tsYk+GbY5dD3tOYIMBs1vgBSdB
zFMmYwdcSEdPfr3h8yqFQ//hqVg8LGkcaItPMXCIur2fQKkJ+Rtd9neLeUna68Xs1rbnCCO2FbTY
rIq/PkwpUDcS1w0+lRpgxYkhIasgTpwXZ91P0mC3G4iwpzzcop/KmJv9Xw5IJR/2e9VLnCOXP0hK
CP1p2VAHmDS96uN1MXKO2llXTWvCu+DjFLpjbG+G8ptzYC9cbXb6ylfmNMySIEzF8u5SUlaBoc5R
KYqx86T0fZ5DXxNuh/YFDe5h17UkRoteC3A9HHfFAIm4GxLM/A8pXjybri9XaaZtHRUTGmDlQnQa
wc4sBkGy0n1JxtI22AJKotDj8GT9wjuR0t+yuRYJGozkTigjM2zLgB4n3eWc7qezm2SQJdeuljrT
fpyGN7xTBAyVMQfl406x3dp69yjibCV8SxA0bTxhm3NlQ9koMUlO+kO0DVL+Qxj5+VclLGA+3Zc0
kRHNPOqs4H4MphhNMYGah/vEd0Q89Qc+B6Kx0pfSokxlo/ZNachxRK8Vj3FXlK9fvrPwgZgobd1N
Z7jC3qZUMm+QRQS01+9rKMQhg7tVEYkZwGHdIfifxuh6ObmVgo71ZYpTBM5WFHTIZNPcLilPHdSa
//me8q0dehnwAMbaW307uvwzRN0IlS0KJHa148KWIQ9Zn0H10GQ1GWMP7bGg1T6Du6Y7EPn8Lakc
gFi3/EjjKeJng0g+NgNaBIPE+V5iER9i06El9YgXrCcNVn6eJLYiMzwpxe4zfOK+pgDK3CBVxQJp
FadSZYM8lFrmVHD41PzgYPqpInx8JCdpdzmkFTaEUfQ9C1VrpiDPv8Im4NlDH443G5atCHW2t6/m
EDwSKgwIHYT1uC65OJINKkGm1C2CCcF/y31MZBeFOj+DndmRmjr5VweFq74G9nqrZVDDUzXtxjxt
NBCv6nN/aX4iDbiICHdw3ZmisFCwnsqwd7LmNYhU/ITa4Q+HlaekKsJ9OzWnE7P7nTQdpldYHjBB
F5CaiLRsEDdNcWpsYMHoKr385RgxE7ylaxlDkV78JHaTtjaBnwxK4W/xb01LB8I11J6blDKJpxom
81yqbkJrgNIjaMb4Us8rLHsVRbLZH90tA+9rDEhHA7+0aHgbGx41SaNskBOFTmvxKVm5zI/MTz3s
rH8oMqswP8Xq49z0cpZxUwb3AjBeCWOcQ4J5IHSepbU73xmQzhVFyWanfHZB+hsjASKh9fof6N6a
D0cDBbpsWEQetsc/rrugPa6u4c3iPgAYhtIqEmHqfTCryVU2IgqZ9e1SNdJedasN3T5R4otpbsRq
p9TOrAW8pUuix4vQLD2Q34B6xlUFMGgaAkM4tuLF3yEoXREXwzvw48ZZ2vy7Ltvvhch45eIuDhLK
FTZKjb8qpGfW3V2akpzKjolqMCFAA2WSlof2qC3jf/v+MxZxAGz+RRu5LyfXfeUWGMrF0eSKXAK/
xAnbApzDlcRKCWIZb4D7fbBkXWZh4dhW9x9Y18LcCQ0Eux4vro0EksWTnxspj5yTgiczQuHUCwYs
6KPQ3/C4A+LC6xfQQnJPJYUYNoYi0WjLO87uqbsggvfJLBhgYOHuT1O3/Ca6v7PqhdgY9b4+KIS9
EauaGMxwAIxvB5AEeYfaFVFMsw8ovYSrZjrwtfGs3dw7NdRO+Y5Kk2MhGZ1NNiLxivHO/X4ShYao
Qjl1734VhcZTplRJ8PkNkVYFCq50EPYbIsPgC9PSpsJ83gcTc3aAUoXITlFSMGEiNxvA6/93YOtK
Q+QPjzLtvkKrtEFqlEkqTVvxaTsiDLck1NDL8fWNkO8PQ+AQypu6JkBnQh6xEUQIW57Z1AXvMnbY
r3/0WXfwfieZi0tIIn0769rOkaWPB9Iw2W3oo/jmgry0sM2mpv8sb1fS4HPMcNFscTqNoGmPYZMl
61DFmigKSZNInonMX1/+EHOQNom750nQmO769wUOHBpdYuO/otBlDSZP0YXbL8EWjj0W14HRlabz
iUljFKUWTzAsTNFp8BVmiYiA9xJIDmaGuYzHXPuiJfxECugW1HyVlxUCB33wn/sZKIUc1ksvv6bd
pVhXr5Gw7XqfoeyOjxWgMPPl12kM4MqtlMUq0wZPmb+mBZjevI/R3VMEUo8cFddFRQd+yzbT8NUZ
MoHTZYcUn/wzu10aZpdUAefRamugRvpNJRFQw+rXhN7ccvXeKMm+ZfuAD3BMX0i+QRbSLWfniZnL
2qQ6LK8KSkdwYYX9ZiOcV3r1XPWd/FN1LkSqbcfHlHcVN5vobU7AfQgfqvIwJd7E2inPXCdWzgJk
+vQo4dcPWJdm+fKvy0Yj97cVK3onve77WQhCoaw0u880avXiSqm2g10AlY6wDqsZVgQ+rdAmAPi+
MAiBqUUU9InLJe5uyuqKs65k5sT+Kurt8E1a7rpmAJ/gLJT1b3fDZr+TpYOZ/aJjh6mUYhCR78JR
6xao5szen/su1L4JRLNlC4k1TBUCg7oX5eqIdGteHKFNZumptLJg/OWy18RHXDUriKjQAd8aWn7V
L4gTAhjvPjbepwE1hSkxnld3iRte5pQ+J0uIO1Cosy2rG4tDeZxkPSQmeNAPSwzd9/T9n39auZJB
dSP9CBPOPDoteS8i4BbYKlU+aDf/1GCbSeTcnHR10u7ol9jeXSCZSRyGZaxleBpWo63gtLqFHq1A
ab4H69LQZWjYPQqRTtZgpa+YLQ1TAuGy7zC/RMQLCjf7dxKz3dHwWLc9Qdo2PWQh2m2XC1J/c5AK
9JM3GyRR/QV00pOwvBe8IeaukAIXYIK+E/VReYLjdzNT4E/8bpkTpZ+D9duaoaKh3M5dv2iiFtTO
aFvi/3ReI1eZPh6vIoH40OPt5ciCbaC2wyzD65JltDt9KKIDMv+sB9aoPnlWW7/zmPMOZD+DSoQh
VtadTmME8jJwmMFZ6y2GtrYc3vT3rYIXq5f+PPiQnvvMg5CZvuZSM2aFHUc9+JEaRVr8G75pKzgs
zlLZaeKsvpmKpw0L6ayjvPIggFdxhS7QRhGlyyj94QRgGdt/dsD09pndbG8jYzkIGl8O+k6PvlYw
fO+4r7CTOfT7XumP5Tlad1zwfzvQ8dd7Ae6AzVU2wo75ZX95RSR9vYjm0u4zdLw56rjpHhBixo/L
UNjtkhdJibnCNULQmQrrW1Ok+RJZECTIqMhAs91UfLf3sjUgEbrStNWbUWvdm5LN8xjUH+INJcEX
zu6PNXQNjIoG1iG9Cp+gR7hSz8JQVAs7cY62vbjteahs589LyfgPWUZbP88JtcCIU0dFHc9JxzdE
2DLKl0B8/2S/IZBQSk4/gEODBbqaFXRLOmKFY0Ccj8UqYM2Gi1B7cVUYrdZX9nz5eHCHomsHoSAa
PJ7dpxmYkJgKowF3okNTCgqSIaHRg1rA1Tc1CNDOLNMXM9yLph0qoIG5+GLs68hwCQOT33APmAAc
FPDBr1SddYfshJCppyJgYhbKRe/Vd4U4Ywlax/3rdYzz0+2mjMq1WVjZY7P+v+KprJ9NQDGbO/rV
SNSHk/2wGxlIe3PZewrffchjM8fa8JLxRPJQbtxwHBlxFF18b62Ocuj6IgIY7+qP1Lw4KXM0fNwr
54of/p/Y8Bpo6IUs4IxkbtMafDGI8xb6q7/e+wDq75W0fMu2116SJ8EJF1AnrQvqRUCS+KyS059/
B3Jl/c2pyPRab0b/LlepN8dF6Uc7j3eId6d8ogxvgaKiZvUOUgxubEpy+vygwG6HKAgG9LSdLaCg
53ZU6qvCe/ts+7en5773gi2jY9B8ek9us6+MAVMX9dGPQ/+0S7yr3RvKPzM6HTODpKESAAzZjY1t
Q3gzSKVsf7lJ4PbdL5D7raWFkqzv0Q2nsj6AuFYqAO3GV/V9tJ4/p5b5SEnU2fnVCzCCsxZ/BtTA
dECnANJ8LCGHRVpQWogR8yM4b3q9w6a6H7tp456kJ72NxiBn8aEmf/fSS/J2UmBqGUoD4ZrVORkP
5Rmg/ulhYbtrF4wxhAzZE7ATqQ9oPyhS7TlNmAZFXSVL7QVDzCZKxoNbLZXRBm0a3xRQgRry5S3E
Ht5wLnkSzHBw43+N3SoDAl1QHR5GlERnc3ec9CBOb99x7xUrMr2eAxTtAwvq70y+oHrDxXKQuegy
u8T6DxaqdP7pJVcMkOQbSxhnaRMzlRCXqgcGeLw/CfNTMXWpKEzGRaCRHnrIeZwbnOdIWU3rIWdm
mb+wj+vrz/esHW4TsBUpLHrwO3FJvo3+dU4Rgdn8Arr28dN27/3IU9szCSKECr9qWvO5eHvb7r5f
Nb5DddEeNEDUgM3zFiGaHFDP3h/QDTphlYzGHbo+qM5n39KicRKGdUT7T4QZm/aE84Q7ruB9U/Pt
TqdHGAupXgsWlTk3CRWnNzgIitqwMa1j4+TmxT+T5UtGalliWfzu4c7agcDWziWnPSWwDwUVLVe1
0z7pY+l7wbnJzdFaKJR8yBzJZY+50sFK5mxkYD2OCdO5goljHCwVMBkpNoUgl1T5nZB8DAbxlgh+
yV2OkfBJxX5LLB9dksaBFmRBSXfZ0QnRb8TsDN8WEj0HRXOiv8Jkgbb64vHLXTR5G/srGtlahgAp
V4iFIZMRangCM0ZCYWeLKjymudHRg/6zW94LAYoJyqed3x/62uLQo/PS/fF0Jlk5+70zq+RC+rGX
MYkSQ1aW1PBIG/de9q9F4F0uDEXrr0iYKXfOXcBC6XBRWE3kh3WlE3eJ4bqks0u2SJ776GGYD5iu
ZAb9V0rsQ5rO123zysluu/9cHXTctAJaXHJdyqHiNjk9vWoFo/yFGemyPZpsINrYpxS8QQUkSIzw
QFAExPDxq+/uGMqKy9pjhP7VQvaVcwTCJo19w1AYlMsQkwRD5Fi2IbLVotuhR4gWbCZvdg9Avymq
P2zzSxqrTYrTfKk4Y804tBCnmKxFXrod1UCKqyVF8o+j0k7CJcG0y3l4RID1dMS3iMn/xA2/spIG
3K5uQIJCbNzCy4fy9jcAqCiXsjy6Q4CL7f7quZhQMmNs75iNyW4I95G3KoFGTSKgyaNZ85r70kt5
3SGZn1YbFf5D7RO0c3K2j5863lsJAFYkktO9iZV2uY1jM+2SdkSvuWmyC78279JJkxh1X79+4Hou
OYcd4SHynesrSKB8P7beXba7btladr4aQ7gkrh0vweDoWpdUV3cXI1yFjS4OqV/9HGDDHAeVpYWU
ny/8e4BAH1lLpu0lbLO/V7LTyisUNXSi2NHJ4VBVI4s4mZpytoga6X0StPdEUknbXuYhtsKtpd9f
aKL+4VgSS8EhTOinIqHB54kUjdxIZFOa1CPKcaq5O4TM84pHpr7ghjfHm0FbFdHNg2MV5QCBbpw7
R0kvSYp9o/GCDqrFzKk/6JJbvd8rO7J/5q/P4LxlrcEV2pGJaf42V6sDubZcntYwxCDKDXoCsRAd
yDGyqbhm2cxFiWqV2A0dmhJ8Ub3aXhXafR+a033T1o3wJ+AwId8dbX+AXYA5m/PPa0XZNhjy0VfU
+E5+AY9PqCphZ2imxgjJYyNefJUP3NkfRHg+CBAKg4xxnMGwL3kyI0NMkGSJK+NNsgzeISkOnlRu
hVFKzaCZ4WnYuUdRbvoGX2gvCs5HxkVai5LETdqj3dvFUAxgsaQMIXpcJezF21pVjMstJTNTFk8m
SiDkQ76UDl1tDCyLDHEjWZrE6KWB9Z/GCaJDaGzZ90+2/kQkexALQmzZALAqnn7PUW8kSs37+JZd
FghlYSfGlV5A4h3Ume4yILLSbDfbnHMY1A3uTd/ds9h55wZQ8kYPpa0X/CDqCFt2hgMUfzbsGw1o
VtyS+I5N3+FGqg8Fg3YV8pk1RLDTjvdOwnIrOBstkJNRRq8/fWhTKNQI8h0YrCsKBgTgGbZxxoaz
+AodX1MevYXc7nIWzr4EvK3au03aXN2O/17NoRACEuJgiUEh9D0k2CyT369dtLPb3Gb3qc7ADWeq
LCZt0gA41fwJXzVdnkLs/WBZX1wFo1NV7C8OlfyGkePfCOjRJXEy4IjgasJP3yAoizwLAUqpAArf
qZ6Z/uPjoNhJzGPJMpbk1uMQ9s7OTtveLEJJFIYCYS0D4NTguEMrV0KZzU+pJYPFnb2K8rCQCDIa
wY540q/2F5MjWZ6vRqVyVRm69W9oWXunqPcUy7BSIrqOlfp3zJnZY6ZFsT7K5imUNDDa90thoDT2
ft5hKLkxWYzEclpIObjUQLHqo4f+B3dsizjUb+5Mj1cigFigRP3/2PbJllj75pJdAd4h5MscFNlc
3hZWZSStaZr5+1x8/MFNsdkKj0jjQjqDgp1A5TokqpiLX3wRfy8AIiWpsQQ9c0clf7I0XWAsAUQr
Prs5t+m3l5h44T4j5SgffErSJCxYDJgz/024NBXqWAdYr6u6rKzONtxJCaJdmXjlbdV39oLbGjcs
H3ABsk/Q2lyY2QkMO5hs+OQEGOPyJe/W7W37RMxUUzohvrUOTfeiS3tY007Ep74eLfPegGAYqz+Y
OswrBm40lFnocCDsAsQ2UhXHOf94PtAmnP4ggL+dG7mAoHuejqsC7zfPoZmj+dF35OYV9s9P/0hZ
2lfDm1aU4u2x2NlWFwcJ/5QA/m53swCS5zj3gEhnosgQHrMvLUZeMErVorusVBB50rYVXhCpf28F
5Pib37hQJBsLfhiuQ92tV3I4ktx/h/ZO8nFNXgSxP86KwhZCDMxL10/Le7BENRk7gJP5c/qNzX1l
phavlVgi3TrgGvFCgqVbtxse8Wt+Fu8P3TIj4mMrbR+FNUCXXBjfyz4uw2+zt+QpD4XX/1wd2KIJ
AFZi8nMx8lqU1nn/5wckGKDpWakwjT0pqD7v4P76n6xZin1ethZntfpJEGSoLADbSL/xkyYRR43F
BRcT5yA0Rte7VEMbSONIdSD6DsjyZb03qdN+vZgNOrgs+x51+9n8bvh35KQ90JVqyiBVHl/rJMPq
QTgaUVFvV8TWJVRWMEq8l2/TgtixSSLshQlnKNS3J1/dl1KCfG79QoFwOnSFNt/iEDQyQgYUJJXz
PiE1nXAyCkHyJsGGAFMarxobn50Us3YXbAHSdv/zOKUSYmqg7LcwBvI7IZ7+QPmtM3YT5DJzWXqJ
Luixn9k5qcV4rv3ABgCAEYa+ViQZKpfq8/xH7rwLx3qUbozcNtUp8XCejggachvOvttb2obgzCa5
7Ub2m1RTl/0+B9qNkzWMuKB+MQ4dlhKyDiPgLDkU+q0dL+1QalV44zBar3lwwTJxmCZkqyjZklTr
xBw6MTEb2IS79Uy829DiKi4cBxtU2Vee4a2+fkesCLvcDQbwwyKK3aSM66ki9VsaNkP6qFduAQsT
xH6JGjdQH9s1mEIKh0+DqzgRojGEmbq/r7EU6d5BsFyl0a8vYg6QqGc1KAYwC0EJGUvxufK9HfXc
4OU01gsUEOJllySNwFj3X4VPFbYBgnNBprtIzAB/MQVBZo/n7APDameNjMhq3e2IomvUK+45hrNa
PJAoT4ULVWSFEbxAm3ySAkHtCSeWya8033B+0xpuej8TLbfnpHyIjVPtIytfrh3G4mqtSydJTBJm
FXs1WENtVR3eJpqmxu2WrxelYfQN3Kpw2+dNpg+1Sl343lB1LsabFFNIjkNN7d3QZzNjOh/Au3aK
c3GVu68MMz3JAmAapdsZDBFvzwTwtC9JPVOIxFyFBZGYCnmh9tP2h/LnEr7GfjbtJlpIKoU5Ze75
1/GDtpaSXieLbLiYpJewFhtABaO1p3JXAbw25IOdnoG6yAh/K0AvH1cZPX8U6S2MVWZ0FI7Wd0k6
lRapbrbpDv6IlAqCkjhAD4hSn5D/xGmugTxCEuGshYmdzKv90EKCrWSdBHxEuqZ6u+i3f+Z7/qGo
CefsmkuWIkjmRvl4ZEUGSqkd0GpxnN0rZWpgntIbu7dT+6NQZFpkvePOe9DrvPikRusx9e7LHPev
XPWd+FWcsZwqVK5sDnRoG9N9A83A5mVIApxAEkdlHyKzwxRUtd5/V6Yy6XfpkH2lpkgN8sA5NUV1
Eao2GGtH16TrVklecdGCrVS2QjJyJI9ZUxuOKFQjMS6Gz8oSiTuMtPd13Xi+AJrH8HEp3TNBsqh1
jYqtpeeUuu4lhecEMagrDkGTQge3Wh4vzzr6FqcQQ5S+/T0tmsD+HfJrh4aqYoK0xk+mTsp3LVyO
7PRtky+NwOYLOgZcUB2TnBTGcP7HcXsvJ4B4MCpKPpU5wHfwnXRsUYHDfniG56G28jtpAreDuUmf
TfkN+htjybw1sC1jnsIqAZ8RZeLNutTRmnW6UXdrCtzFbYlwSszo1/B+ldFwyMF8QdDAyeSJuzjk
gi76TMIEokXA038UDTE2edLeCW63UvdAXO5lwE06WbWR+YG6fQnpeyw9IK2cnZbo/RAnshJlSBxW
nDtG8FRiHG3gMQHhg/OSCBSvL/EfQbZOkf+f+tvZr/+M8aKeb1RTZQ6Wld0bhXibDFPQhL8hRHa7
Rpupk1zuA7IHUEdRAu7DjT7/Y1vemVRb1LaX/IGpwus/5Z2JGSsc2SurEsSt62Ovwuy7OlaxoS2C
+oSnMQoT3VBpMaZrzQnS6eCH4MYZvvWSkl18ODNkSLolAoJYgElbS7F6ZD5b3bsr0Zu2oHZLgEIV
prOt560xCU27AQ40uoZ6ZrZYCpEy0qTXZ+Kw3a8QmKa0OmCCx6+SymjlKT3nxaoezfKVNke+rUQy
uJzz5IzmQ2pcx/sp8BUOhiWPlxtgruqD873/7jbyWy8ZOh20/8RxX/JUg7kpHovlNyiNkJWaYJMd
IJQqzvTu7lqkUNTuvZfyeVNbt4+lTJw/A5FaGr0LC0AjtO9ElYb73QV/gbbtC2m415bBF1HdLPwG
JyUJYLJC2QxlClDktSAK5b0irofHFGjP9ZQ5sGWyMlBI2lUXY2TIwxmqRl2buwWwM71Bt+Cvx1zM
8kacEqF30FyekgQ0JSWcsO/hiByoSnA/CtKlL1bKuB/nK4yq2o+HAaT8I0xCIjSwzPRhhPtK1QYH
WH18diMtfliiysycIpjNpZWwMbpH9BBzPCWHDuxay3l4sv5EmQ7sVGc7+Yscn4bdpRLKgzT2duWs
/qjtcoQcT/ead8W47frQ4Ewn3iNvlgrOZ4957g2ISWjMw+Ehkyn2pvK1lYA/hsMexxGT0wIcoxij
tsS5xPXSUL5qkTLDFAQUFsRVW3DSIyFo9nqxBMfFewVE+9EpzILAtOAw/vmEot4HwkM//Iu3DfY5
lGD2fqlT4zZywnNesLm+XUkLbOSz3YAhXr+SoDe9wJmNrptq4IYbcjwcZlpi2uhaphBz3heejr0u
aScq5bw4V2yQTCjwE0NNEGXTh62lpWCpJtoJqeNdAwk/rnuh2il0RihCOsMIHM1R9mtvf125un2k
5a4haqvybSx+DR/NL0AnzKugsWx1VHXbtiznCR9yVgbwQyTNcPtkzFluFCmdIEDCsx/1OTfuH0rC
9qPgEWDTphEE0cLtuccUQi02t1Td1YV4i4BsP6ftQZREUgNH4kPGdx/OQjFVuYFw/mILN3eH7bKt
ZOMbGl555nvRt2wjbRuhoSKzFc3fCjZQKwFpkBKcBBOC7WZqnehGr8ZaHFrbwHtQHgGGlployNDP
M+6sUD8IKR8MUCqxIFckYAtffqqRTFHEI8m6+iUEL4lP02BUK+n+75XJZbRlZC1bS/SbRp4wH40n
lVQo7X8nmOPLzwvPUZgWAx5Lqfp74bLnH4W9t3/X1s+Vc0jrSXPwnWqzG5CQ/IQhaTl7CX6/mEzU
qQJSJQYjECnkJIWL0DrAFDDGlAfDdJWBb6s9iJRFI1K/e97ZEvld13C3GoRSjnRTePIM0hBNT4AZ
ztfBVl5dr2MWkYGEd5svSqzjN/gjnX2zAz7fi6cNnhS9X63O0ddI7loVEoGq2rJpO0s2G5MOM6Le
CUXhcjHb/UzDV5CUG+FrS++es7NDMcFnIxyhPz8/t+jPlFwDKsaIqpmYS9CF6xzql5VmHa8Sx3KY
VSnSCDUovcLwEuXM1b+ikd3qktdLJHwZ5QB8A5puxeSITjVC4f9qegMQtj9+lD/OvMzS3+pc+NH6
e/Hx1km1Xp9lthQdRFTEab9MqQSWC91JoiWeGBC4gkPDHE+YWRFntq3PquWnqClPSg71nysRpLTu
cfXf3kXVu4uv48nZMlG3ob2jHwD/qmv6Cy/nae9vOrALoR/LMLsdbkbxfnz+2nuQsQU+JDEGH92F
wzQQxIct9IGpWItZcFGb68NcjRO6J0s1U/X36JBHHZJm7jAYcM8g75RAlytOul33oZvFd9EJqVaa
1cTkk1DEHZJBSkuuUVVsQjZ5m75BF4dSKwV0m2crm9h5WOeR2Jeuu/a2XRe7D8+rkex40P/qdrWf
I3utRyX1IGBrUbfWaw4aMx0jr2eUFNwWzkTK3/fvllcsXhLIMwRsuIUy62qNx091uQFs5pDNLYg7
wfdApQWF+Zi2QC9rvzZejv3eNbgaQJnnRkcnRfUJiK2WdBU5UF0LOhlPSvAKpkHpj60S3ZqAkoCu
Pq7kjYHf1o03t6r/Kww0c+OfLGGAIgFt0YxDAKWMXqM9w95xkj1vVQKNgxjrt4NRR76/vH4ce0Iz
lboMzDUpNTFF4BgCmk0iJClmWsqjy/eXDV5S7owFHYPN4DXvne7HgDKHpOIm0kwRoC33lowqjwHw
YPDKjW81H40qHhx5N/oH0KAZnpoqMjuOvCKTgtg69Lx48SQ8HdHE3rspcdSiGcX0pQT/DB72gdnQ
42wzq8hbZ+ApovaXsOIF+e+DHInpOdVd6C8ysDYr+yu4yL/T3dC9C4f/hnq2h6TYdU2+46pcXBXp
yjxbwq3OWY++Om4ztyu3ajrXZtSYMXSZWE1ae4sBgeEJd7U2czE9Q4jsi/vnflw/QhESET9vwm+4
Es5BHmHmA+OM2V4N3208hT5SdM0hD1azOXyyuQMVlqy3pGjvkH7Q3Wby+ZyiLLdx1zm+SiF/Wu43
pzk98VipL4HufmtOKja/iBAZyiUq1Rq6BP9QiFk14rTAmM/tgAygCXa9SAhxZF4P2o6/WOL9TWWa
uQJlzH8ygvrKmghTzeNPUmKhpR9oLGjDTB1f3r84i2viaFkApK8CLEQCx1Mo5JY22R4BeM5zxZY1
bNlvja/kpvMrRysaJ+V9Fyt7lPkSH1omfZ2QPlAHqoPk7VVa/r4MxfE/bz+UwhYb1501iRgXBzzI
hhiYk4X2e8lt447qV9ByxRSVLNq3RZ6duDJsZ/117ucXADGvDh3oAZ7od79D5deWy94Nm5jy+w+j
oBqx14rl7uSYhK5QAIzw/TQQ90s/rRHBvg+Wi54QXOYOydZeHuxVxh6muDI3LmXT6g6QUOCyNhgO
SQYviiUq1IxDCYtKODUia25bNmYsIy5PEEMf42Jcz4ktnfROY3vXlx8fSTZikTzywRGZtSMfBRHA
lk/lfDK8cbO2cjoIe1r8GWR4zZT/i9N8vrp9qfgh3+DLpOejU8ipiFVc/qB1H3LBQJSk2JuL8T2P
55l7+dViMz1uITUnLcg9RM8g7Lw1Ls+8+1x16LF6qQwtI00yH4+3bqm2Ky/cKJnp17ZH6LFQRSN1
x1+TX1kwsFw/N2c2MAMZsZxvEahNevPzptfSTS1DdW66QWJS+yyDCfT0KBW9N29BP3881xuFP/Nk
YtQfU2wrD5nLDoHvw110JtCHRIkArwhgyKn9Fsdk/D6HR+35zoNsO0Mx66d5RLlXxU1uqZtlA5sf
Wcd2QaDG9ukT4O+vhpkN3fP4/LzK4E8Y0ALbDLhnKuHSuMap1OkBPePtllUCBGkUwWP4R4wH5X/N
K+CsNlbDmx+bhoVWwBtsc3MUYXS+yydJh/jC5igdBx152pXX/OmBUL8az7kR85Bajl1rJWpOOS0a
AJlTDWZUr3LQ3anBvqRgMhhSu7rWcl1aDjVK9dX855VujIz+oX7A+rfJiYmHWztbusZKwow9a5Q4
fXMRO99sVIm+pnfrWe7Lr63b0CMMUR7hOQoXy35PqDBOXhEPyNbsaSocaAe4gbufVIa0oJAPeG52
bQEsTOK33aVFNyKoouS5yajH/GDf04jLnXLe5hMqSEh16lY/pJL5ZBGdxwDJl8ordSevxqthVgFC
cGnw7d0y/QS6W1oNPhgaMKs2bGhUB98EgxeGfWLaliS4itJskFhrq1aLxMYiDauqN472C7DYknsh
RacA+342Ph+Qw2VeLIfuArlRYzUVE3Z1xw7skMLobXhTEWV8nybdkWRPtJqufux7DMctMhGPtGop
ndvtLrFejTx8dmvGO0ZA6edAtXDZs4HUQEsguKs0mr++P8qJ1uAkZXNl6/2Vsnq8hhv/W+j1zOP7
wrDtuMtx6GqFO0g9icGLrceJZxRKIK3erwVipAQvhduI3U07AKT55Zi3lRbIcIRhXLmGJWqgHc7N
WOuMPg+al+adRSTxul/2Cdn3r8RwIoc0b/4759fanTJV36UBeX3i3RLrM6UHnMnGYHuvD/Q2XvpG
vNMky9Nw0BqBN/OBqclkpbGiI9Dic54EXr/XxvvG5zpAOAck6chTie1yiTYdL6Na9bHEaD3spS/j
nRmQi4F1fMdNxukPGyVwXbo/8h6t3xaMPbd0lU3SwAHqLRopaewZVNjeHlLLC2+NPwKSHvVvLBMv
cxDw0SPK/9HL8Z+Eny1HekA0KpRAEvMd2o2aOQy3s2dpJd6NYbtePCCT0DA3e7xi8k0FhTc88Dkd
bMA8vUCk3vNcGiiPwogglv4F485dnIVLR5iBS0paUfuc46JMhjWvsXPXzhCpJZgkMNxICaZrZ/QC
+AJ2Xrq5wlECxHJdgvvu3ok+SgXSIKdHK0RQOdL/yg65nxrzy1cZ1o56EZcWCVXunRl/Zb4tix+t
Vdy3s+TFPWsjXToGhB/FZ3JER6ZE69wmAz8Vi99q0Izq6H/VRn42Z37dODwhiQHUfvS5k28O67+1
TkUjTjELRj4F1AVGA9IZ4N2lVtjAogUeJyNXmpm54dSRDeDqTnUUmyXeyAvz5+AEx14nund22ByR
J/4s4OGkUnnM/1id+k7DQLdiPtMjHfZeYB0EsyDn8aubmYykxMr/MBw+aFSMJdG6/k3yAIc/ea8J
qicI6ax+mBX29xMT00ohtyFJOC8Ms79MhXdPk/vHxW+kA2dRh9NABbEaOjlWilxsKqkKumoo5hIG
MuwOFCxLbIbqpIWkvOcxAzgYBarHK0FK9U+Ey1wWiWneD1+nyiefkYCYoMJx+NCSC4n6TrZ68VWk
atdO41SH+BZvvr6Thm6z+Kpw9F9KpXTuSLFGj2GTl3iDyycNxaMaKQXP/AAUlfcuNJzo1sTVSSAQ
zsrXGp0bXpXUt0Icww1ZNMPoFixeVHHYWScQ5uX8de8gFO4iEHm63wdpAQ7bHduj6rLRq+f6KPoI
O8/dpQuwaqbshNOxNnVLkWHp8BkBoE8zZIO6p/aY0FGK46cZPeLws6kfw+jpGmQdoncyB7tNjHc2
rY+HWrrubtBAHj+7W1VECy1x0oKDQ7tUQpj4ns68o/Hu9EmwL3Yx+jv7GUTuUS2LWugDNP1Ff6Rl
/RTz9tcLUadfc6EsLPNt0u0/4jVwZvz6lmQq11nEWhsocbQhbDVlnUJOIhr4cJ/SvnhW+WVA6pJc
N29/0bEWWNZk4ml8nCUGDFqsxPgLm/YpWCDH+RVZYRUh0DBS2PzPYvyBdbAk4k6sjWbQggGf1brP
K0Ii5dbj2aDf5tLT9qSL9GqV1WdpkMSkie7/2OoTZvRAPyRLe9N0AgIUL9ByFDwFXHQGbRKsbfhj
DdaKn1D9nuqszRCJq1L0bl0PbAcO0H/rNXD4gl4Odl4VQPBpjexXP6T/R1Ow9hgTiq9/Nzj3t/Ym
SgmT90rC/ub8Ap6aI3GrObl5+grfVoxOG7atXUAcHBQuKVxVQkXMmgG6s7uR1ob1vwW0m1pP5Y3c
kbPyn9O/38ero9Ht86OB6d8cg7psQKWfh/ItUTwuNr8lMUKH1oLoRQzjzfIE3492iD9PaI4AGz8G
iCR5pCu3yeD0mKBOt0aM72YiTr/O8ESD8XvWhul1bazROuNrssdtiylzaJyGyzR9FJhRoJy5uRWs
guRgs3uEoYgXhmwszsb5Cxl8WogweTiavtbIvSIlev7291L3FyB4j95Y5kSYGlYiMjc70aXeMPdJ
txnSxYdAe0ruSJ7l+9GKyBcpuUPBNjffPu/aykgNsL9Y+i0b4IhGTm/yvngnA5beh341legtYIfR
prijr+9WivMGBi0PWyK3DUnHeRBCJuqZJkvl21NOQoi7HXFWZdx4hid5YMRzT+bN6F533KlKi0Jn
vOaLib0guu4dIsYLib+Jzw+BcGjW+m/gcldUe2QCV5GtJN2nCwB2aQZ/jxSOqp8er1XUerrxD4Ji
5+YeV8nEGz1uy6BMEpgNZHw/GASbB6FCz/Kg7Lsm3M630KKcjF+8v28vNMwIYO5uF5J2+tk2UBU3
fyT7iskqOt6mlHq2Oiv482qxghkLg2RUNzjjLFTggO02UA0zcr/H1xPIgRI+f+orf5FyYHoAeh+W
BVHB/kKDMNIM0ZRa9d+5SKPz/6hg3tDYWUeX8DWomBpLi7YHGFaCDCifu6m/vm+reIhpVbzFMg6A
/XDyItocG5ts9Di+zXqAml83jRfFA1MSjvrD8vOiQZiEEugCiT+goEIt8clYTVLGAka1XqzYCtFs
CgVI5GMpznPx2ETO4DVPruQhZ68kUZ5OuhO0nAfbqg3rH97HuIDPAZQfplarXKSbbHr8NE0aRGsQ
wASt0I7389+pnqIrq7/9roNOenBZmb+TbYSe5oo3m+xC7MPfxWAHHJWLpK+5HKIqNvge6PmuWLiH
8hggyTpu/O9EsmLD+9SUfIiVSLyFYYWCqfsxypKaIYKRt2Yivxw3gMsSu1F9I28RCrzpDHxAcQxs
BwkBjbWJcGcc6JRIRDYaB4HV/TLBppQs4pA1D8HtzZRFjl1oN0rM4xMcAjEY1fb685JVfLCSOy+1
4vr7q7GuP3my+z8epBFEnCbF8dtJfTddhabZNHThBWFgg+eopnWw5UnGcyVCI9yGueW0uwetYW0/
DNcSrgAGJPbydF73RLF2xujbgMEVhp+PhTqMvWisBnuZ8ggWi0zmSTEfFrjo5P2y17DZziPjzQoI
NvoK7YD6e27J14jtRVP4GppOF5yXzRLRBMC97Aob0V5+ptnSeYsiUf6RdO8KqkqnkFTBE07Z68vc
gnwGHocFKyxaBS2gjv4NtzXuIRYR0h1Lt5A1WE8E0kVf0MgHPIRBxJd+CNoUvgSvqx6yQ6MpPIny
Dzh4qiTDqDl2JvXzOqY7FGs/FYOYVtBpGvNWrztU14GyS82sS7mWqejRe8ITIND669r8nl+nkULP
KxPD+wrkV8TwkZ84cse81O4AAveeHiZOMC7fQAaK4vNRWTTuVywj1n/3YM+Z0hG0udviqRKHz1Id
Y53Yyvr5VKFUG+F4x7P7BirWZKNqG5EWxCE+9smuQzNCKD/JYrHXUTCi9jR2ojoJy40TpLSqrJPv
yPLM0dQY4qEylofyovw3Hw6h87SBVh3ghUjRewtxVACJiGti96xPCdSgL8H+Hwm+OYvHjMztYM+y
voBP+cmNarcN0OeMyy360LLTlEPovzDnaCA0FAUEUuXS9WDSOa+nJhpfYn9WKdIrMvYbxOmlSJsp
HH1yiWPY4UXKN90RxdIs6HOJESj0e6phY3IxXBSjwuR1c+zP/J2HM0DCFHQM1Eyi3nDZvA/E6eQs
HwR9C79hEp9I8+WgYSrXr9aW8yP5f+2Xr+gJSu1XFeN/FGtcqdGz/SyZ0hXw3Xoe6uqFXIvEcMcL
T4FxHfg8G5vNYG0WvC66VNdoW734F4MlYv+J2jigk4XMLjUQO+oj9Wv2cZx0GV5bMUZoXnZIJyfW
iOoV9wqW5CTmVd55OEj9/0jtqdJS640GnMj0G3VIcmlqRB4kn3fwTF2NsO19s4G/ZplIEJK7hGAH
Kqcn22XlbkTh9r683oefqK/P3uaV73IaM8lgipgW0hMhQRfkCpKN9lxx+j9StbWBveXoGx5gp2oS
RSgjlWUPwXlChGxiv8Sp0jlJbCPUD/9oZE7sOCAFKsjhgdTS6flCd2rM2U678Ga3pp3hpM5bX0nI
yFol8LkEhiMzyIXJpNbi8iCNJGqzhAN/YpDSLGNpJmmC2yrbCaddMeoY2mmqI2xda7Qrjd3i1BoJ
+kJZXuLVEhlMtTwlGCH3/SpLsIdv9zR+aWR0QS2lon4KnCchL2BYBeboDSPFxUH3LtzFebXdE0NQ
6i4J+EA+a/5aWEFAjEFP1mt+kNbskZmMxXHXt1W9HJL/F8FBNKO7tqFe6cr+F9P0GrbuRnWvnHI6
juFS4znIzC/JR/G45Ftn+wHuakd0lUq5UsaVvIZRtGnRQKfSUw4ej3zpjqlfzrdjru44Lsl+qlZO
yqt1KGjZcPBrKfDhmQRI9IsIs3b5rhMP5Ve34wD/ZPVfOwy3x9ag2iQYx3Gi4djqc7VxNTfZY2tJ
8agBuGkZAYG3bNdTtGERv5m9115FVgwwxq4U8D/jkvkKW3oheiGrwsuGJtXafBS6VgnL7Z9OFPzB
owAJqjEudWS9kBzw0cRDqyPd4DHalWpdEH/7+ISNLIEwwzHepn+WZ0+8S7AwGreg4RDmafUqFptm
/MeS6/Tg3kVunLlDiNklNrmDp/rvGzWDAH2GWQxxFatkO/jXoNeoH9H+CPLKU/Yv329jiGCziA1R
aFok6V3Eexd0oxwqSm6YFpamSktwNIcqE3sC+K2jHninURMaua+Nbs9kdGHcLSRVprGspNC9i+HK
TA6oh+yi3KAvGUcJLUftpxEwSC3jFZZyNstDdmYJmloYA3+FKTKYZvuO2eiBN88klzb5VwPK5NX6
Nd3zSFE+nocRxqz3S6LCA41zn0jz61wwUAg8UDAgEewxEEnZYcYGZS89gqDNnESGRvnwBc05RbdC
Ad03VtnOiMX1xuUa6ih6dxz5Sm9up+lh7jR/O40QhfHidHJvGh5C8L6fhPhmH9S5CuDmsQbdfoNC
9fdcB826WbkqLKMXrJE/PIJEqRSoHOezHZyH5h5h1sL5sBH2i0M8enypjFVyZi4HiiGQOc+EiSLq
AdXj6ob/KLqhGmRGB5Km+kAhdvNV8VrGoKnVlU2Do66TEDIy5nYvMynUbKA8kHucvTwycw7VfsTR
Z8fdOoYq0l46BUdj2TN6QVVKBwPJTlLTYEtSq6TBMzLEC3V73jvddfHwY1yHJtwFGywshfVS16a4
Rzvi+9DgYKjOUWETgt8W6wc1aqWIdKFGfUY7P1pVaLUtWmvUTthyRjPPCO1dg40UXj/XoBUA/Ltl
grp+aC1WOR97M/HmOrB7yIZY7XcCWB5/ikqXuQ8BMCKQ1Wl+HWz5mFduInJhWFbG4dWO+7YBPcf4
damhovvTwpGroSePY/s7uSuiGgz7Qt6LCmxehLRCkXkPAUw75frATn7awwgO8u1tf/tMsun8uFTh
rX3MFrFSAj0c8vepiJJAAPoIBPII3KtNo2ZO+DKByNN7KWfaAljSloAH2INdZDt6xtaCz880viqq
pE8hIlDnEdwf0ZPZoSTmVYX46vYsuaSFlf6cisieh5rHjL1JDMkemsN5A7ICnITB9+l5p3xDt5Z2
0d4GJ1bBb7dN7J2j7vWgRWcannPhGN7l5SCXYP+9xvm+Gc25eCMe3FmVu3EFdZ0xBN/t7Un1NVGQ
1E/SHL1WLfvvzCETEJEBDK0yGaVwA/flrDuUh4CTqHdzAh7zGIpbls5ft7pjh3IHGtSesPD91ops
6kAjG6tK4ilumYOooK77Rv7N0KMGwHLrmBQzWrT3mnCaiYmXiK5IK+FZqZ1+f+WUWn0rwdsT3I+g
VA5MmUcGiCGD3eOeYCUx9ysIYYU1uOcj/T40s7+dl8u/9e9GPgOVJj8XGEdWGyyWsGCxWGjwjjp9
72Cd0XgS+UM9A271j+pepfL7sokCPFEMk5DmQMUc7i8mf2OrQHIgnGpYPCtxwnSLtG6tgmfctGxv
8uOKqdL+gI3BW8YGytzt4Pq1ay2kMo1ti753mJZngCjc9kgJoBIk84boUZL7+kfGrCpjHzdDiIKJ
tKp+DthvdKKuEnPsTZWwLxswpXw7R9/PS25xJgsZqqj4d8o8nvJjC5Ko2HdWO5fIBmLVsIdmV5xM
Gtj37vRfCmV21mY2BC/KLWCEvS/FBiokpLPrrSa+o60xyqt9+oc7/AgPQtrmcVPAKdTEqJu5WH7W
PF8ORsh2nVuDO+tXcqev2LB+C2tppIzPxwW8jG5HmJfgeQkqoEuIGki+ULDhW/hqIg2tUxD9PvW2
vNQQk7GGvY5m18zAnyR4yYkRCYSrt6P8Nqn3TthSSp4b4eBGtBwXMPut4HLqvnZ6hR7Dv6HoAebq
3FTe4ZIuFCrUbbc4V3jf+haYM4g7WY0ypRx+NMc4p0jd3AYVndghHbXkFCxqN6Dtuv55K8GiQck6
wWTULR9mfwPdXub1guY6EYWu3CWyEnrtIpKVmVPfkhi9RSC/DoavO80Zx+QnORiN+0VM2JOWsrIR
updQm5Kk3fk5vj8pdWRgIV9bTHiAdk+QGcKxm5zh+ySgfo5vbBTe/veT+D9GBiIjvURER8jSw3PJ
AWgo94MdHpdBIiFkh5pahWjUiLuuPlSSEYgGoDFVsyrcTbDIGCYAmRH6/2hiGY5WCIyqDgy3q6jU
EGN0KlLNYvdybAmIsNhbsF1tw/k+ardHRB1zjQdoVAWXEJILfbq9ZIvcUnXB4gXgE6TdDfDH5NLp
2vsBgAVS/SHJqr+K6Gkuxs0pFD75rwFbp5gNtBrbdQ2o3KCd+MaOuRSx1uQUgJpVLUP8mqoUREml
pX70bFBLkgFcFVqJQrvqoHpL+KeDOqn1HrW47KKnAU1mxBkdyAhbghf5jB3ZRE5VTVWjB5SYDnJG
JGfkxQwPV/xC5kv6v9dNZyroe5H5N1ibX0ThjqakZwd/lai3fsfMb9o8SKF15YcbLTEwNJ7IrUL5
rIsJ1X77+/Cck8iqFHGVapQ9r0gHhuFbTKDrUM9lJJYLdrHl2kSDv4zjg/+n++c+c/LAQqzy1leF
EKWyD9OfpoZgb7e2rSsVkoFZPdHkplx4qQYk5QD13F++TJTpvaj3967H0J+FTq2snE5McEreopkA
eJHl87HmH1LLX/WgnhZZJLwYZUqHQJ52xcvea+SZ8OGn0Jk1DgqvUgUaAmc3lzMAnXG+w78A9OyT
wG/dk5t9VvINVMztlfA8glAmAigDlu2GL2DxLkXTEvX94ZhSvRze3gsE/PuAmRGVoAzpdvmBaBpT
wEKYPGtLOJstTUHOWYO6aEkKY1OP+BjSWSVGJL0uxsUbtLrGtw+6ltCS1UDvOK8h+KKMIME90fIE
zjhC6szrDYMuNIsapk0Wvc4H2nDnqqi7th8XLc0YPS/H0pdX2cWLqpDHK3I2zJ1erCvJ7fHcOEfZ
U9c7VI/Sf7bHiAfvnCGGSeVVMsAqdkarAOpMQhrabkMC6NDTDYTTtrYciHZXRtjhPHh3BtK5ho7J
1QIxeBWch2ALitv9BPGAIsaRixOuXF9scDq7yOo0R/sVLelvAQP8jAOaxPqirfqUZlnDDtY+hut3
0Q78IS7rEn6hCXuO+A0CvfoHObSFK6z52EIttj5XlczquUtxJRDrk2mGczsG+gQJ8qRXQP4aL9HO
+KE+4rk1ecgobIpdEu7NT8gEG3xjwhfrZTjIKvZKu9M8CACgx8h8dIFhdBJv0tk3da2qnZ6Xq5jN
Rd0VYxNGP/qpmoZleTjbHlVy3fcj6Pfbh5HXPGfrr8yl9/lqp+ddCV3A/sA47h8kjpPke0EnW8+P
aPO4A2/cXt/0NQsuBHP78ZRFoSovqA3TFdEfokQXo3NMG3rxDPilE4w5E2/T5cTubDWxrJzm1vrQ
wx9UCbAWjVMq/ygiaCpx+//c7Y1JSFgzxEi4OV9WysoqeCpz+PSt2ylkZB088n2U85B8Y/IjUmQz
w5NGhnHvobFHhDHADsIQyFX2X3uLFNDpA10l5mGWSbpbK7Utm3/RYeAsGc8DCNZs49nZqZp+Y/Ug
jdMOnK7o8hhB/OD3Dzwcr5a5q3gVYNKxHrYV+vPs5g+sRlzwKRf3P79OKvge44wAE0Hw4k3Xrbx1
poHjBQbfTCRJnM34yBLZWeP/xxnNLBpotnVEpFgzj02JqkzvQ9aW9NkJJmT+MqSJ1r9hAX1Lh3vm
E1EeKlFLRsEqrwmdsA/e5QNrUv6f7tUGDr179cx0xcxEeMkuAhfd6PMcdIukwbQ3OZYz5SJaO9F4
+4nx2RngvVJpYNUIFvDtrAXy127wJchHcg71gIo4kOtvXufKu/zJJZc7rIHWv5HY2jCgi0XKGIdS
7/HzX3c7qwJPI9qau4SZlhAojXA+uVh+TFvHcv4rZtaR7s3uPC0qxd9MSIWL4HMZIxZZg4ebJQbD
bGr28bU/exnVsuLsnAmVGQjb6iS+6OJRS1Ue/ZH6piRoriB9NI+ZuIa+LBVDCnwlHSDpIkho+uSL
ubjkU3gQpNbmaNVPfIFFVZCSp23G4D/FFPc4FaPPy09v0EgkZjFb6fawyl6GNxdztdWkXkRBgHvT
qtF3HboQ4lvElQ8XweEm+ngfoepX+4+E/3R0jPHlxEEZ9cIvOA9Wg9uQ9k4TrIofTfdwSb1w8sov
sj6FC4+nvjVgW+91OacsBLSbSRK9e/h/gxsKOePVZT6h1+o2RyauwYA8qQfyMt0MkdXgh6KdDOlB
uXYdDTbkHQNEbhq1n8cuLEKvUg9q+ImyBIUYmWWtOwx4HhrGGY9/mRVS3sfTAYM2YqiaSXv2r+Fs
DPhKbTN6yMcS+IFR2423wFRjH/qGa86rMxAOP5ajsFZPpkX7XKIUzHJ88ctUsz0QXF3TMk26QadM
D5CioZfTXkEu+Yp0XDTt0ZSA9v/Ku7wN2byfyPl1/m398jSQqo3gi9v0DU5B8wc9xWEO2LFCxooO
uDUObxQpn9zDNyA+GJvtj9Y+Ti5CPijxk1IwhiN4ouJbU81F3YsEjqncGBIVVkhWPiTxvKolkE23
LAZpPyu8imZljeXDqhEiLKuKpwhjuk2e9oB1Z7uF0Ik4Q51Q0HX4EtPWxzMx4UQ7MPPVgdkLGkg0
RK0X0Kd02tqIhFE6HXxshqgo3XqQXkptnjSbY0VfPZE56llchcWdL7zLUBDt1or34FNg3dQeb/pm
InPkn5vBgc0Ehoi72z633bQ9OBP2bxnc8vXk5q0Jl119aAAPp4NFc6Xhq4bcqqC7VG+ZoZvzDA/z
MGjWlGNIYc9x0DRoGqUZ8/WLpHVA8UsZNp0AB/H2vIhuT7tMKURsKZuh6gTklmbYwvAOkM3KBJci
7M9Jt+vaPoxCjE6YumFpTbslcbyUGXyjWwPzH8n6FuWPgBd1bpEGhkLSv8ajrG5cRGD4hWievjFa
IGTm87pm5C9glPnzgNMGhQvW20pdACYjL/xGpD/i+6D6Z/kbsOF+i44mCzWIzZvyDvqV8cCXg+yN
e4LCBM+6wl2m6Pjfz83WHS8Gc66yUp/+soPyvVapM39Xuo798hftgUvnpUUqeQr+XA87SQ+pSD+3
bd9cNn9DGylFaaxoG+iH73g0V8alV6YvUJiGZTgEB6lHQt4AW4LgQb7aMpfkIPiDqQIgc+WrzL76
4uZfZCziiw/LucuRWUmD5sBM4z0rBhGywam4EYdZedybeYpU+mX66HCGnECZKiGd3RZRB3fgpf4Z
+wjZxL8qqS4J/TprYFdGWaVRKyN9Sjh5YfHT4TWEcDh5XsK2+XGvVRWIK/WHe3rImILpkl+Xbcjo
DO6oMVKUl9YbIiukeXbGRVYlc7TU712JxBBAWRmYocobN6Tiq1q6Ff4tOyu+QJPajR06utzT50If
hPo0hOAWiEp1gsBCYplPa7OMgnC3EOMWDP4jNvAzO5cOHuxMsQBs80P3U4OcbQe5JUBApGM2HB5t
yCycLoc4uKlv4VNFG9HOCACpikuiIj+Uzi1/gIRbWkgfaeprIYTe7WfzmxIP1OGBvM4R1ofsLqBP
jABHzjcgbvVjnuWldgcvpwQwsT+yo6EHsq91+XoO1XDPqxfHV7gxYXVUThbpUgt2oEo+GKM+eEYL
BT9UC+k1Z13vF18ndnQc5wBjzOQ+/dR26EgvLN+KS3fL9c226GLDYYQkA404FzMrTdt9EbKCIwnt
3Gt1eXxw9FQDzeEozMNl7bO+EcvvwPaEAmBz5w65BfYGSn7Inh7Vw0slJAqm1FpsUy9o9kFxgcJh
i2Fn8gtp8s8chYBoq3uz66WvDR55y3jMU6EqEz7XCuXPnMVLhtEMlIdIXoXiGQJuLhwh10g/XaEV
guTYjtslJ59GgrFHshI//22OrAtwnC7L1dw03fI1vRTNsMpHt948D09durSl9follnyfmBZY0xQU
zHloKvMbpbtrZyTgzE4oE4HjkuGXSty+Cbf3a3X9RWgT8dBWVkh/5uXy1PC9QGTEuQAhtOmYAQPY
0ow8FDK9q0XEQkXTXBWNkn+I9J16EHxNgDBHUaTLrg5qbTzllMvwxyeV3hqZvWDRjW/ZWM6qxCbh
o/ge+Arbf6eBxAfrRKtsEEFsPTF1ubCH2JLgbCR1aDqmDhQtQ4kRvOXy9kbch7rsSpPVdwIIWP6A
v4uTOjzR5BBNUMS7OOqWrOJy6wm/LTdj4rDoBgoFzLGT0RquVUv8qsOZcEEF3uWuFfCMfNRZ65qc
v9+38CCuZUC8Ocf1IfpAlv0lUTV5pjUDzZ1AWerNbc14LrbkcQUTdJ18OVd4qO/dsRgSwQNDOjzt
01j7mUSCEZ8NyiwjUDiB37t/dN78l3fGpclK/KClPSEVV/EAdPyEof5tZ1D5yVczmO1t5VWevC39
SHCavrTVHwqzHJG16Ylf7kY35WTLYdYrk5VhxrNpwS+k7OnC83DO7TbaimE/LdL4yj5bXryH4QpS
28AOZdMWPKOHRPlsYlcXXoSkfkr8m69WoXF86inSxQrmYO7lZMh4s/I54xUTjiqOGRM2yuI5GaCx
x5PYXOBiLQygivOFDBXim1FBU+CpBkozq+jZLK01j55L7/8PUwfs/HCmIHLJiQgj2YMnj78HpJqd
WQ/5nO/uaDDH+YT9xSBZzrktRR7I1AiM9+v1as+uQJhFQJ/IX+M+usH28igFclLQFCb9RbzeTDNk
lQk2UktClkpXfZUFZJK1rTP05+jfNiksCIbik9Os0iEeMcYXaFK4v+rkZwKptRICIlemYdbaTWiX
C1iU88q77/6db3ONfX80+5khECYeS1uhR8Zm+oLFrCn5dwcDiSDtCYpEcr0o6FSQuMu7VCFsmXZF
kFT0AmcKS/tD7Gltr7hmRzUBG4ksSZMwosHKlekh1HdaElGbBe0o89WYXWfiy4CDQeI4yPRnEZv7
bfUvTV4xUOtQcq4ATI1M32UqjI5u6D+mCo0J0FNjJAEZiEaGLrSV01pKg60YVrG3L51M+Z4LgL1o
woYM7hnaIaYbYOTBeLphvlBa35TtSW/SANsRtPvw6uG+/XQgSCQF5VnigbD6baTBYr8WLFuiX506
YYqXMCs0t6JwXBgO5CBVpD6VE2rY30tVGC3KFwW16OKrhgu4akEbWJmGaVJldFiYk7LaQs/TPnBw
y3cB3e8ZlJqqzUObj8YNkchp9Zd/UKZzAO0QYra8F5yPQkbUKnPR1uwgYTMHOUiYsHvG5t7kCn79
h2mvuXEO3HO9T17+YKAKwUu6ZkI041oyhJUvSy2tpguHoQAZMmPv1Su383K25og7GcqpBHS92XHS
uZEnIE5eGjvO6DsE18Ds07iYHIEC7bElq0T+fQbymDqfXFHj2UJmKvTFCpvdgF8R4Ir1HDdwK3gw
efqKHu2zBATjFUwdLBtd3LOhwpp1g/N+vPFr+ABy2cqK8IcLPuZIb/pLfStJ9qBmrdYrg+HYd0ij
YcYEfssuUVRNLe92BG6bEKA2VJGOJAuGInnEHKM7E7FFRVEuFCn0+lddz+nP1GVnmuW++fwFpAjZ
9oEMGqZSsPKIyfTSxXY0hOSnXhN+I0ctWO5T4Dr1VlF8eFYvFSKGbDehOXaCNTdPaC2NiW9EFHbS
HXgNfGKKz2xlC7iHJaygRUtKrwDASUmNsfI++M/sGsnCGWHwzTLTDkHrwT2gZjXkJaMd9B30dt8q
VfuJ3WcT3OltmrQmq0QO1BZXU/A6VHZcs9UhvEaj4RVBdkx9W2OOTJ4OgaL5tlpki8vAElO0iqNT
N40Ut5snHpIkEoi2V5fMo4C1U+8Oq2DwfBNdHXQ7woCdptlzVLEy7AGFyBxaLq4Jtjg+mzaauxfD
YaGrGD5CVLptypC4Rr1vCBvorAzWUA52WecB/NNJj4f4atdUOFu4p+ienUwXiM0aQ2X6GcYev26A
0o1GzPNA/edDLEZ+T+/A/5LAJJr7LE+khdBFo65fFZfq3sA0g3MuI0n82W/WllEG6IQ317UFQwGJ
NfMO0bKEt1XIF0VKtySozEAJOuVW6eYGziM8dsQuVw7Hf8WEcDhm4/Lakf7Srgyhs3CQEeqzkapx
htuTbLOv4UFGLg0nrNzuqP1AsdZjbcKoKq72XDK+ta7CEufSS1NBiqSx9rhToDIDupAxctyjW8le
ygS7MGd4c9JtMDhru+2vKV2wVndJI9tC7TRznqw83Y0vXXYTJokVTTPxfraub/NGswjCA6alU0SI
uCdCoUZdHgxrrv+yQQbBdz234G4UZ0qaViZp/+pxNMtuMBQxEOgv+CHiSPguSiCg0MXB/RHDrooH
ufMSPvnFitxPYbZb4O4vIqQkyRzzJbNum0dZrSTYhcmsynx7Cu9ou+JxLuc7Wx82rJC6DK5CVTOH
HZYB2YYoTveDiVIcSBMYorxrlEB6H3rD0vS1mrRCcS0Bt3omORHRH5rosa4Kyfj9wQgMjGQHNttx
THzjQm5iwl1eAXDCnX3LHJqWhBxoESGZcLNx5PImRq51MBa7pSHUWOTpJugIT5toel0bVOtT58rl
YVpSEeFxb3YYGvuEjpxQqu/vtaGZk9bRVIqicUe6yoR7Yox52k2Gi1A8WJiSSAsUgYbh1gZHwgQW
do9qdSrtaZvIxAZctGWKcYsp4mBEkyO6EQ9oIge/JQxddr5PXHQTcsfmd2dPpVREkXxvK91UyRzV
1ohJqR5lTpIQIixpc1oICEHPdquAXsSLgT1pZdLOPvLwr7FF6ZFM5+Vfg7VONkKE+iTTXTINBu+p
vdWLkEGMZ8obw5aBK1Ce9c1rYCE9jcI1KZraJlpzzBm6VP5rY7aIoorrt/c2QDwtysud+blLfyyC
NZdVdTmwVI1aPwlcejL2nd4izdljD+p2l/P0nlLs2NgI7hqtTOU6kRfYJ35N1+22qNiOD6ckXpgQ
Gs9UoqbM18ioNkPbNLgNQCcCqaumPrbfr1JryaLjS16IDt5YeqGKb/iaRywV6/Yw+ncw2JxcL9+M
9FcbsbFdNPH42MhEZeotpAUQfGrYEyuQgxjTLRGCTiG2nfdO4hV4e3SSQ9LBDn7FbKpOzKj+tuh4
Q0TIgSnlj+zjmJ2TXovyspP8aD7ceef6h+oUD07xtqj3sMZSiDAA8ygyiofPKRcZ8quT8MsCnQzH
4eoSR/XLO1lg2gxx2mZKt+Z6V45qyH8Al/cLThFP7TGA3qBRnCnu2NlRi21skTSrclQsV1IjTU48
R8MNVgUguY91p/Uj1+bc4mR/MFh5pE0tApjmIsNofZiT3aAnutFcUfyqFLkQ7y8WGO5hDZuz+QEZ
U8eXE0uBAhVoaeUdL+TkLh7PC316eFsx5NcCL0GiDQT/Rmb196hV4hHCNlSLcFRdsxLLWAspOc0X
G85YbJUHuuUcma87ib0V29feLoYrKMHW/QUaBnkuQc+Aul7wBtYtq9t9oXY1OeB8EqCqacbzZqOM
f2eBxe90UH+CcyPiQdEZTDUfk/r9EdCx9uJyDR1ul8+966X6taNE3wOS7qQ9F07e5FVP0ctIcsjp
1J1vwHlLZ7SuAN5TN+8bj7qSfO4gXZm0Chje2TkHAvbP9uwnhb4GeK9vCl/n7G2WAECkKVeS9zvx
RldJO0NdhXjLILDNj59PSup0sLj119X0ZWNa0iC6Nbm1DqKp7AXPox0HXXK1WRdg6QPXyJTi4Q06
R79QHaD3GusDfpiFJ+I2yof+iyFJDsKgDfBqS0G+nzp5kslHyGe+h/xyq1Be6Wf9CGJ1yKyk0stl
dpQobVqDJvGdDPeobpGF7vl6EsBly4LeNvBUFcEGOvBRj6lsIt6i4RS3PVnQhaOtWiyaLFs8jCCN
K8MepBdWofJ9rnCsrTcfWKyVZ9QqeWj9DwGmAkPYnJxQIb5GQWxSz8C36L9tPG0klMm2cqLDgL0n
JFPJ7Co1tSw7f5HCFJYm34vfs1QL/jtLz03ZLL1WWePnxup/JcVC29MXBhpy8uvK92lGLuKwVZZ2
+an4/3upLVXDoY2zqaYembEr55WgfycSny+CRUYtUTqtKGOFWDU5/F5zU2p8MosIw/5XjpWyZ4hc
2g9UaqI1Dul8w7jrbn5hLqO2DuUdGA4KWi1phpJ/tLP78+xy568yIJooCAE3t+CLCK0JJZbEdE2q
dsW9/TR/g1M3xkOXPT0zou5v4h4D4MYxdT6yC4fmFPkj4H/unuT0PaZtfrQJs3RGGzTPjKJvNXQ6
d7Xu1GHRoP1xyuU4ph1b48Hv5lUGiol9G6phN9eu2DAOJ8jAUu3pax7r74BmNJ4D2c1/Uqxhg3K5
4wmCAffVgdnv6HH6hTCnaWQfzC5QxT4eDHcmpB02Dd29GIapG5HDPWkFmXTDSaqNBUSbxR4KvQN2
wllUoZD4gb9QQ3cemoxssmzrwOuiIY8lBYyT/09Ehk3dV2IWJCQF2HGy8kKYQFq+rbHSkLEPgO4x
3QGzVzoFGAuOI5vHW9HR2FXb2P55JlC4Fk0kPjL0VAhYWHR60oC1ZogO8MvmKzB98xEAT3Z+weOO
rXtZPwWEN5AVC4NR9CsbVeX4iNHm01hbFaVbED968pcGSzPMJjfVDUaJrUSgPI7KXFKN5WtNtHTu
QOPl+ddSiY1rh2fT7o2+nJaNflIrTNESqsZ+s0jhSYvmtRSaY/LQDr0kr9mnH5lkO72Q+JzCWUE8
9Tq1gNiJXQ56ydqyQlhP66TZ7fy3t2CZiqFR/QK39FJpzdSJfALZqq13IZfQtjHhcKRzoMIY4jAX
DmHiZXYL9SJJC2UcSShKG7zTUpP/AGQPfkvL3zgEnG4HGN563nkcRTKoC9Abcr474DBaqU0mZ0fn
V7Phfk+ZqnISuvoHC4ut/kxWZCkOxHR4Rz5c/0uHuiclLNJLdf/J9rZvp0ptCGE0EWVNh9Xti0Y5
mNWrT9C2nB+z0eMMtGqJYMbjkhitz3p8oHOlSQ3voaTIj1xzn39WmtZNwIVVJyrwwM5JjmICa+CT
K/IggI+CH9Wwr/MVyIC/ui8D/iK/gDgWkIxR77/S8Uamt/9vVh/dhWzAURZp3O4ZUF63toss6Asi
GylosP+eQ5/ikWxPoV3XLuxbOTQGFOMBETPmnC7/1Fs2Y5+hk2mZ8Gslm5YTSqHgn7jkkuF+9hxE
vzWEuCud96LD7jAerRvRL5dFHh/ZimVdjpmNJgnFNTCbIi05kCB1IRH+r+uMlme4a2Y7ViDEdT3t
3NCXmnVBpe2KbuLCE2ienmMqzPVt4uHE0DVlBPs2hpNklPZjVm0VLDfnp1pI68qXNMEoyZWNBUuQ
RuJk7JejB3H3YhfZBCMTDGMw0SQ7GcY5btlnM3Eq7Ee7C60wsifqdbL3GJC4QDGYNCm6WaLJAYSa
XPz1OwkdSTQUfpIFyFW3AaJTpYFd4D8v+guGiEJntfS3KTRcR2hkj1Get4cw1RSQawTEjPCjs7QV
PRRUQtuJCwpIEHr6DBtyXG/LP0ZhCJeOH9yNaHFz9yx74rMpjfQe0VwUzHWTILzpy5ZaKpUJaLFF
VvlHfNGhNunI7n6bDfo5wZt+Lauxj9fck2tqiCv1A9OtBhmj8WvyYQb/q92cOQnpXiCRds4QpXQe
5dbqeUilzZLT2DIdpis5vXCaMgzgrmvFK0qc3TMtSL8/7g6w19vz7w8ap8E6hKK9xV6C52iK9Urw
4d9HYYIuSBfOElhej/4sxmc4d2zd3VawDY38xfQkPLFQZfK2psufoeTu2LI8HCI209dNAAPdvyVG
TbGi0cpo5GbneJcQNqPiSSjCRRr9JCiPQ3Mu2xkFC0ub1jrcFA0xOSndYTMgtUlnL/x0XKZm3xwf
HH5FU+FoA/je62xdssvAKfTmuI7ToQdzCVIEuMq7K5dFw3r2hOl7VPsS1C4AcIn4/LutmtJGhjwU
a3mhrgUF9Emd/D70Fhtjr5CoIOiiDAK3YikExzXT5Tp4nSb31fU4pf6Zlu7XV/kR0nvP3ZffHlXN
fuf527sRN25FRGmmcqsfMTb1sdS451s6vMCfYvIt0V9ijwVWEFfvQAKQ4RO5kpwQpgREyw1py7yA
gXVa7PizTMfHRPBbLvkV5ZK12DPnH5uAmqSD9h5TBsf4TqwxGVf/XhUr30IAX6gTihVeOwM5uciA
hyiKAsVSAUBwcepFdOqdizYaYkJM3UB8Apj6H3tcLLYNZObf8NGh2hpzI5kRnxH/Yq6nXbip0NQX
JgwWpzb/vByaMSMM97Et/tygcskiXv0WzmscKr3XyfuqfuURas8jKVGGAeOar3s7xp+uujHvfQnS
hVp0rDY/zcAbwB5oiWIvVRhpAuPrah+ywSFRvrlsuGNDCgNXWuaaaH+pwaSButDUussTCU2j2fWQ
3AtzwGrffzQhgp6b4TI0dbxC+lfdwcpC9BG+NsNV2X68CpV/WU91gck4rM6uXsiJk/39bH1kK9bC
IT0wXDdJbck+Wb3fgDamZK62db4pugvhHQ8YE0LeeI01pK8oGEAlXL9Jha4JhgirqHrcW51HMmXe
rXw+TMH3yEKk6FDBcxO1CsXGfuuCEh8XJdbhbYr3Li0c0fMdU0X83pqC7wcXctLUrLoT4BWya4lg
ibdtsxQk0khTVwLPGR4VeOFi936eaRNAd65rgwW/aA76NNtvy4kM94/Ln+HkgA69kylpvC90Xoj2
HQJPUrTXD3RfH84MPR8a6nFL+VsdHiCXUIbo6HLXzh6t7pJtiD91pCOxPdKd+QHTpFXKX/g8cTy9
4nogCpd/u5gVSGl4B6KfrCnN1tszL+FA0GQe7+aRqvEQGvmyjnyHqirydruvWMZM3UuW/mziJthL
Ry9ToObl213QcX8StxQBUAs7N56U13U37VOhylwqsqzFsikMUQ2pq7zvWUT3ZO06TJ9LocKD12xI
L/GCWn+5ndWaXpYSArUbeq2WTO8ZgjiarRemoWoZnLX5VZfnikeKbCr8NUxWBNUaE7WOXw5RHNF8
yQJ8XsSMPEBQJ4Dpdjdfw7dMO1jhK+CHzHcHekK4DyknGnn0y06rXisyygqE6bdVDZBu4Oa7iTnk
O62LUCq2N1y0l9+yxg1gytqJHH+uICIsCxXDk/HZTN6JCMvTsGLjdzg2b1VuBgyHgZ+WBF6IiIz7
cuyCAuS+OeVEFGoe0VmtxUAp42XmtpV3LWe+uyzJP8/589GDDNsNaD63KWvnAGMmuFb3ZCVO2Oc6
q3OJu9lRXr4idorJxAJMTxjEKLLzogxMfUsZ5r4XGB0JWpYjT8bd0//f4wJY6d69UgiSbmbXEGxQ
JrH9CG6h76M07/0ddf+UZwqOw8Y2JyV6oG8Y2Qjqf7JswFabTXtnD60qn5M8YMnucmPucPE8Fl7o
K35g5UpFTqrfP2DuqgcnFPcz+hjdl03g832huIOSgTe7PGWQU+mfE6mfrmkxaZMXHNeUhRGWI8lk
tjc1ZJeKNUoJZAmkKR8MV4FggFkYoM/89asnyy/vOgJtK96gbQzKdrxQv9X+37qC0feHQ3neYhkx
NHMDdMIhhZ2dAp2D6AWEByAKPJzzn1amH2bGtX8B1YbGrJBAvCCJXWlsTxiLat6pzGbg6OJl/u4I
3xH41+1wNf1M+PtDYZzPryWtW5jIhJHM9TdTZzdKPC93GG6mlogmsTO6HpWnhs9WriMkvm2i2Glo
AFBXS5e3QhvlFQjpN1z6QnRqZaMCtThKeFKKv71W2EI90YmYF2YqK1JN7Q0hPG/UhtVkXZULlNy4
2O6AecE7F3A8RkqJYbjFU60JuytfauSNUWVsUzKzxCR/q3VLJ/7uc3VBrszvFI93EQzSuwclCwl1
TF/KDJTux1QWnKZ3Zibz8+RBF19viZq4E7bjJ9si/j2k6u/iTyU9cp/buDmBYZ9XydyW6beq800u
VDtZDEwL1ir1ss8k0237IBZpRGrrpWSdyGwDRCYP3dzliCAvYCfl5RpLAihWEfrIXDuNIHdQlfGv
5kdzht0FPoT6yPotlVzD4yajGdUmUa1H3ScC3Q2g6G9x9uYMk9Bo/paC99rRBkq4URZadKxJF0U+
/cUjRSQ2gYxkB632kwbShU5u/WC3P7QJBiWraJ/cKyesY69qpEb2N1fhagEaEqc9Wbf5aCnrfJXW
aIS55snYJSxkCJOAy/bcC2EKNu7LzoIF912hOjQ4og4ZD1CtYdmFJ9isQPmXjv+HDj1ZdBWRpyh/
yTjNIqFqYVZ/HifxqKmCVpRSdW0T4HzDKg2mumE8lGDSOK2qc3aZyxTxJ16S8D4i3umM9FYGA3aO
UAUp1gMQlvkXOSWf4fqtd9EzSCBe1AXFCMM+Tyc4K/zm/vuf3QObraMpgF5l/xOAgT2S9Sf3nAfD
BnIKNWS75ZDbn8ydgckBtNyNGaoHCS7ztieDYwLy+okoyejWdAhumfLkDmw5xRQuYsXRKoHu7rR/
OySvPs/eLVNgLgkmg0TgFuktiEr6p5ObqZq5OnT+u8wKh1egtf8mmb1sOgr6pwB6Cv1AVmCnfyOT
nLeD635YSnDdNfG/2VNOAufGjQtCPLfxVZwySef2ES3FGKhSzpcvZinSpr6hzeXP3zJDvK9kYnyB
j3Rj7OdeonLWOG++gCkNClbVM2G5N/QGZaGEx2zJDQNOM7M1/5T/inKoOxZpuUBsvs7Ac0nvQLjp
PE3KmTVJsEAwkJIt0C6xuI4b5WwFd/mBaNOjzwe2WYSrouKf5q3mbiypM4cOa4f7JFHHOzOifhsB
RjD9wanweaCW6Oq7CWjMTDNmA/TYe+3pI0v4tyO3k4gDjC4GKrFGsWYRCesW6BjHezatIBByZbp1
4FMhmcfHkXajurqyLkKz9JRmV3IFVpw1elWEcUqS/lcsUBx/C9PttCER1YwClErdnPUgANAM8LVd
wz+KBcyD5Mm0FhNPoBNm5aM6oyNOTY1GfbBZPOiHvbDEabni60B8nci1BSBC7LSkSTfi4b3U0U1A
GYKuRud2q7dbIbZ9EFpHDwI12NsKQb6QfDeVoy/0aq7D1fX4WfozlwqRJeQpyCleZhRyOIf4JUdZ
qeJNu75UlTlE7dQZZmUz8azM2698/U8AOEQ1O5w1fIxvEG092xTRIYxuK7BLf8e1XtU97HgH38f8
BJ38SDxgVxV+W3820nU1e3L7l8mmPK8BEcIwHU43uQ6DsS8Dvxu9534J6WGkc16dUlQGWbTxA6Z+
s9tYR9q94H89ofVXwl2tbvktxvD4IVF/oZpdvKh1OrE9hZxalHlPt65w8j1mKLzP6EH2lPoRAxEs
7AA4et/4cgbs5dwgPdZ4Sj+GVn+lXn83TotwLjxb6YFUf/dsVDALvJ/eOTYYei+8SytxQcRylmPQ
FgJfr4ETC3AehUJbqdv28L7JqgTzBOv5z+ptOo9Ai7TnWMJxX417l4zmIMgUq50Z1+IwiC9wOHJx
/TbiBuv348zf5G4/9+bdzcI55tx0z5VQiwV1Gs2fR8WhskKgFxEh9CP6j8woauZPXjyvMRGFqw1M
2TGy8vqkkBgEYPGNbrHXggusvLer3oc8o6e2clvVRybXtGaH2bkarLIi1Xz4FEtzutXR4ncTG9kv
cy8gZFZOA7kOp17tuCooNnvo4YBgQFIMo8fuxq7d+GVDax1csj1uGkg5bdre6hRpGJnzhQdm9nPs
Roevpvi1wnrr1yzE/wDoXw1jQl2CM1Hi3iqg6NIbV1sO7YcvldydYuXPLdrt7NQrdbbGyasHejR8
vGXtqtfR2IUsy6oVtI8juB9VuCiuwnKnWJRIv3WrkvxL3aXRiNjYmgOFCEnXJvSptoKEMKuvt+J0
kArQhGFncUUAfk/Dl1DgnQJQ1JmJRiH7GmWRFAkdbNCM1hiEk9lVs/2kGfukzaTioo1ZcDkuh/KH
xyb8+GxIyvFk3zfir4FBDrrNixn2ZfX67McafR5tQzzkAcw2AycX/jBRkFgd0TyXHWtDjdF8kLeZ
w9rzH5uEXynMWLIb0tgUYFJBy6zeNqUBthFdmskQcyxzX3+tI8se3Cj2WbHttupWpqj/Xu84+eIn
yIjaSFLrilnxEolF1JVwy3KgwT+TDW1/kAdQPlaVue2WbxE3+HQOWgVYXIhZVM4W4bOjiN2LwAEm
pJ5WBKF55J8TUrDa7fFm2QB2/S0LHnDOEhxnvyEWgNu8L9UAFvGoo2MhhQ0rlSVfIic9JtC/T6aa
tdgHY3NFpy2ZHCSu6kMmWCvIixxrZN/FrKD+AQUKPWSYscTGjMLVnYE56cUVALTgpwkB50ZxZb/4
boUxFfxH9mOdlcN9raoZmnzughe5FZkarEgUUS5zeOqIJ2FhfS0YSxwO/OdV6DzQ8rxhk9J88NSN
WVdTi65kyeC9nzmMjZwYYwKVcgsQIkv7M08qDuSr0bwzNu6C1wXSPTSkgfvT+FR+Ry6ySf2AL5cd
U60ITV20URtZj9v+NcoVW7OeYIlozAWaLvy2A01GeFYPOGnHViYPbaerhjtHW06bJfCLyEkUUq+k
Ya2VV20I5WoSm4Az900UwACLIZiXtrQZfn7oEoMv86dew6VWS8MUw7Lq7wgUYsixEI0vXIFR78td
AwGRnmn1H+B0MCVx7UdWgfgJ4IkV2rMHu4tFMyPmJs2YD9C3zKZWWFNuJLRllvZZRRFbcu/prd3l
2vszC1DsZNMGQeMEyFuzWeeD9DAEHnqB0pXdoqaL+tYS63oDmDGCl4zBtQ5yxLvarS0v4eL3po/q
fRwhYJfznk6lUuIVipS5NcXXhgWRyJ6ufvEjQmoP6HFxgUFw4cx6OwtrPlUM6arupiaK0HiBWimC
5b0b1PgTmwTYTQoitY7Dsb4VqSJMfC0MLvzLgptABTQ0EuEqdJpQiLH/2uwi9MtzVIxfxfFqOUiX
EFCU6SstUAVLjawPu2npJHiTez+aSOCONBpWv9ragdtAnkm69MdeKLXdZXlG5k3Ju2vDRQ2UamcG
AVlyEirnMoDgfGc2fuQk05WBiPWodMOEm1JIr+rGPNy8KnszzeWzLL7KoArpmSUeoRrq2Q4ocaEF
jRk7xLiZICCC3qCvd1Cm6HL4rn7Z7Cyry2eOSerXOw0VJ8pqnMzHEnsUdsrb9vTPAISzk6M662D0
Am8UIiUuiHoXfGW1/RFRVhWgSgB2HzZQRZKeuKxjAiojaa+YiLY2K1btnXr6WOzvaMdXguTIThqg
g5Is1nqxLb8Og3KTzMAgsnPfFEQcRzYVZjQyAFPXCLGzcLx31bxvshRZMvCo+yBAReD+MqPhczQk
JYYDOGWGYcv0wDmJUu0tfLp0nh6o4nPyHXp9TtNiiFqOAFMLtUTfs3bwGvEMNtxzBK2WAmOxbYSf
yRoCjpfmWWDfm/JMvd6H4aYRkog0KpJz8b9LfX5RI34yoacaUntnoNE9h0GVO3RmbTjfM1YT6oRG
r+w93u90vPD6fUou7fxUGlkpBIud4hMlhTc5YYt9+nTrMH7DJglQ7D3sfxAnmIL9hqyvs1ahlqwO
ZLdzrQcNxjPGz6bXdpMFPz4NevV3IuL80JONQqVl14ZLAgWEiYD1KXmq1H5irpzb/ZUKSRGaNJz+
A0tjX/dqhv6u9z4mEEyXWUQ63VIN7GC1vvEfUYXEi5bt11TnP0731peN6Z5d3BRiApo/vMDCCwfY
udmfjopiw0fm/zgf/gWaXgt6BEbtWGqmnvMSnkYlpJDFClUO1QuV/7jHSHTqSrDqvfhEQuuqhxsh
9w9IMIwNtxB0+Do0/DnK5rJzdSZsTehPe6AjBfFdxhu/7cu0wgyR96T0XcbXTMCMX1Vv0QX6V7Hq
vwzzJzdaaWYCk0WZXWKKoHWP2Zhw/+KjTMxbaZsXnj12ucmRI+PEHr8c1etUHxO/D0nXVtt2jvrL
0z5BGOy0HR3FRo5mPehRnzP3vWZyLGPBovecgcfyiaS8VEETT4bY5RkI2+GYdu/mbMD//7GTm706
L5Kk94GTbz0JgQtmvzAhGb5ZDZglVts8L/DYjV0v4ZGffafn8ytRwe7iFOTh4bzwYGUB+O1A5J3w
d5bzUSWMaONLpTdhrje/BVroFyZF/TSYAPVfAB4XTBF8TzPeZXPOkbq4yzeUhzPtVaVAXe8aVpc0
uIY2j2kHGpZ7gIgSpUeKQcBOAbCfOoC7fi7/g3jT06BnWr6ytrWR/u5clQlU7o9h6SHzNDV1NzvP
Mfbo0Q5gomkcER/aFgJh4FsFKaA/5fFuibRCuYn1czEJgwTMnfogmbJ/46ArhFBtfoR/Hp5DDwUn
7ltR0ZLixWCH+zOK2mmkYO5dyGhK9C3bMowx1WHkNHzf06gWKg++5XRjNDHD8ogeOilCpll+0VTP
4Wfyunz/ebJW51uEn13HEej3bCNJT9H0/f3LEP5Y22CqBbEk926Lm1pRs0BznUVNcWf8ImDDFrBy
f5Tp7rTP1K4sSCVYYm39RzrNZ28VuOfJqMold4XrEjmtBrLU1ZiQoxusIKRGpxf5sBEmQ/YP1GLP
pyK52xkvF5d49lLcvDBddyzbcrW4cjApGksqsnizCw63JmQrrFnQ9U49P69VtdEIhDl3WszExmbv
39vHayrjDGhS3ntCxvHPHTrU44E5xd9lTYStbVGZvPiiFayqJwF36vGDw4HH6b0hNPG9AgUcdu/7
TyotE1om1pZwqKc1m2KyggPEuWfbU00qR13raBytM6WgMmil0IUt0QHUa7En7DUj9SJZJIcDnlCE
HVH+Pz0NqHNFFtQaatV3vfOuXABvRwuAVOKvikkGLaKC4o7OA+rvNA64MeXDGO9Uvu/O811p+C2j
+0AzI1RuoBVD0hFiqzuri/dZeFRgjoDI0OTD1Oxrkay7can4sv714Uc20//7xFKp33+QSLBiTEpv
v3bnDPkllc7jbosCcD4qmoYKihYvBtuncRk3UIeiniGx3ic59yk/uOlEwJzR7kby0eI/Qzro0EZS
1Bwal/VVJis9SWEJwZg1R5wqUrDSl69J7FHiBajy5X/7JKfL0Y6rW30MdENdkm8i5b8pxWoq58+0
J0XoY9B2QIxBckrzXjnIEVoaQ741r1JDWTfXIzJN3EBSbEv5a/W++VDw17C8Y18sGaxNXFAezZli
pT8ZlIgkajtWcNgQoPd0m3Rjisa5PWmBNwfVvJ72JXFYYFD7uZTZR8qPe1nJ071/spspR/UhSK3F
SQAp4kWBfgQk5IWb2MJfYXzzw61Co7Vx5A/tavf1MHHBo0xAwhYmEVE/wW5r7jPc+IeEW8Or/pCX
h16QdsZLQy6H63zqREEh7zWQW7zq8+AXTj79rxZanunY/9oBxtuS3GOv/TtGbMT9h0NMhwNSYfw4
b4SPBKXGscIxC2QvF29vKFX3cQW4HKAF79DXP9rjiew7YHSO+QlDeklwNOG7Bz+2HXs7qVjvJ1Uc
JNibMwEFqobr9UOiFgnYIXl+CLYn6N4RrOzNvNUkFK/EPaTTUJE0mQ3zxfaxjLrojF5NiaCSt1cq
hwg2gDWMdzo52EE16ks+1c77xn3oPmFIm+SjNHCso4tcqW3o69lN1eOwPKsBxJMpB97+0g+SCG7Z
Nazsm5J3spr9avBWlxc5az+hSkQel66BmjO+jx+WFKEyt9I4mA6WpNSGXksN34EtXDnC/hhPAqVy
S2bv9pNDSQdiGL6y5S2bePnJSeq4M52eoLaDitToSDNyUcXfwER307ZjGjUoDB5vhCOrB8Umjnyu
Wlde/hyl7pHjM9O3GxBaRfZix4AOoCukIMZIhR+YGlelvCVETSh13VyWdUERd3y0FFaNOSOJLp3t
SDyLKN/FyfC1hX4BKv90Wh0Jg+RV2AROIvIUMZRTENyMNH8xqaouiIvk/Hkuor7ZejNU7y/tCr7c
kKEBQ0lJxZjw0R6cuCBcQ1anPZpvZbzH/Cj/CZpu9W03BlYOKYL/egz6FcTAk8e+OPQRa390Oy2A
BClBVaKjHXQfkQ5KzHmOcNMS7JDsjafrFvts5Q/pteeKm92LVomrA00pJCVKhd3bw4XIAnIv7moM
GEizwbZIkPdstPxaNl4Nqvfa6aEwRkIfIUh4x6YqMSVBSYnOyNCWzy+F5afJLNQHWmS9p4Xk7/sa
mtBhEfe8DZDWKMmK/E5DO/2b/A0+gagIY52nJ8rtwwKBCNK2SRiCcCMSAIaYL5LBHhQiV/W1OwPA
E4AD5LiAGD1fILxmQSTR5eiMLnIRIk42ZKIKhtbvmEl8jQ6GpfQIaDaMe7FJ83+wUreD8Ed00lzm
WyNd+8mPmD5ADWhtMtlhlmmifXGpDif6zJx1eTKSAV5mDVgWXOCYodSB7vl6d/Jlr/JI0/SqwIr8
euUpYnaR4R6EsJ17mCZvDqkgfExeIY7y/bk72A4a9G5QAkVeavOoiQWtjulBA6w3kCC29l4zwMp9
00oYFttwriR12zidjaB1RY9UxLeeQpyJG9T4bqzUmiKWABXvJKxHmsFGyC75gFC5DyPCr4gvyba4
VAM/kw+YxO7P27gRWlj6RS6ww0o9jp9tu7TBWeiomMZI2YR8ZY+w3WqAz/evRGigor1cD+ZjDyyU
2M36FAYfle+rr3lbSfG+43NcqrwzYO8Z8eq5mP6b0xuCKnyWSwQgL3Vo89Rynr0aENtGIWFjgTOg
bkJim7lz9Ch64tusJk5Oqc3WKf5YMnh5kORja6/m6vKBXd135JPe5pWGAehBQZl9PGnmynjMWgmB
uYuhNQQ1y6tbTmH68vqp55qUZ6zkl7VJ1/RsFTv+oAYC9ylw/Z/euDEeX9qCBOLKLTq05Xve+fxL
1uGMvljUTiTpk1+N975WHo7kCOuW0KpKeeZG7l9xY7l2KLIQP1u52u+d7nNwrC04lQ3lZTcpH9VK
wxRDOxirZok3xPXiTL+mnRfB04LWOzYZ3waYm5VBIPaMeQcbsMuKWF6ub4PGPc8Xf8CH+nuD4Q4h
o7bbu4HSTNrgrKD3VJZlQjE4x4kZQWh6pXvfulqLMGPwupS1bAVtdKcb2GUJwba99NU6xVusZdx8
PaIVtBxkiY5JbnIzRRTldpLeQx8enRjsYScu+zpS9SBprXtajAvh3PwD6uM7UezeNPPquh8UD+0l
tgkCN8wvvRF48TviFlt8BbNEn+114EOOqcttpg78peh9OfEB2bjJkbNUvNmWvhsnEe3EBCL2pQCe
hgkg0Ec2iVaLg5OCgzszcBX2oSE2NQrqZXAkXjfBJCYn3UAP8R8cGDD+sA2/DRoIROQ2V5Omah1D
Gx6+nxjDmInsn1QPywSjpjXbWohiK85P5M8ubsxEuRCzUw1CVxzcV3YlYoi4+ACJaREfbJ/fhSz+
l2CjRRezv6Syf4eXJ2xQE9n4vEFcpR4W2ArU9QSyS+cmq2CTn3FIAQgG14D4iHgDDZELdDGqGIKF
22t34VLaTqVubUoircKK97EcvkYVCWjnFT2zAdVeDP8ocWck4Jv6mHAiEizJihzhT8SJosj0C+QE
U337D/HUzWbX/jOhjNI3rMw6PIEngWfLVBtrKvEFE7FKBSXV92ihDd6nuJsRyIHmWREkfxOrpuvm
jIWWEfKnJ/5iZ6SoHQzGkBDotWAQMLereKLeItNps95y2TNKPxgtxvFqG/0aQBarTB/G3FuQIwJR
lgW0S+LQDv1NCUO5/khp+5OId1l8VLLP8JyQHd5K6blFUVVnm1iu/1wnOsdPFOtNnwjsQwuFeYoO
xmrSJemlrDaRUNUc8X5aWItZdcyo1n+z1yhR9YtGaHEw5+f1m8g7nSTHsvQQFW2Ya7+wqkj7aIDy
7mTMtnAzSlI8gdCEzJtUR8Mxm6MJfgCNOtpXCKH5dgOUQG/OzE82WUOEf2ksd/GvYSmEcBmZM16c
UDF2pBLLBDKLyEj1q7J8WM6UWYVVIxafvZ2CZtjtVXZHF+XVIn/MP453Xvw9/FcMRJvZ36thMyV6
jr2Ydyl+ng6AKr7/tjjCj+fW5kk+5UnSctcwDWabks1HQLiPQwUVpqSRLWg4KSZ+23aK0iGPgW+m
YFp9TzVbNETv2MCdaxRhXx6xfBlTyihwmtrL4MurN7oQRYJ444mOCFgcrcL/u13d3AXVXt2yMBHi
Qx3EKryZgt9VpuDr59b54W0FFaSahSY3CBI5h8Z5hso14/uvRo9ZBlrAYoCkEjNZ32p0sew0pb/O
eoWKX5B5seFelySSwfy5G5JBDLocFMHc8k7aAd7uZQuTvZ8zHUTZH5PXGEOeBiOrkSQU2bJFCawx
c0B9yaRc+e1VBn+JyzmioktOhgXNSJeTGt0Nn6GaoYygXHow3/lgVANvMK8T54cI5s/uBtexC4ZC
0xLHYHfTPl96uqV1Q+MdqhIy9e0Odh7W3KY4fttUpAHcmoiMlEYYuriGC3Sy8glvqxqMx5l9cYOS
7iOVEMMzv7YhqMKbyat/SCgj7ZszDe6x+4BB7evCCH/YSmr8yclgvKBs8eX4z5RZoCwvEOnDh0UU
mfjgeM0YSNs9BaispDxPwXOC49cXMbki1U2DM7dKVYp797uoil3Sxc2wW2GpwRwa9qIOLMff4g86
VItemY8aAETgLDlyzoEq2LpETJll9a2KWUyVaNnksplG1wRXC0+mP6iiLWDUJ7hd16jNmnZYcL52
P2FYOIgkACKkdEGcMnGzIM+n/pSklDpkbHiz8x9DecJsJJRTx5nA3bDCgaQ54zoPm9FgT5qPZYeu
qFGY5KSzDfrE744DdY2fvC2Q/CUX2baE1lQbYVXUPxqYbYkrFSRAy1UDn3M061gYrDO2fKr+airc
mvnqR/Gld/2fJFCgGVNEWn+9N9OpAI0+AX/QVsaRIhCTCrULFVhAsEDedJOuLHOueBpyScQneN0B
cQ+9mnmCI7ZC0mv6OOlc1eZWeuT7M+v/5V0Ib2c9Q9QwWILl02MTsJP0BY3pE6DzppVI0BQbZ+df
y/VZU5XSQob37lS4kPpWlpUup2AsG9+t7at7jjehUgSdOcisWiimKSdwktWvkWn+vEvfAKuoUlqL
MBrKvXC7tAJPTbWD0CaDaKdvvSELj/8WQ63xIEF3itm9p0U9pu71ZFBJO4FlbavNu6mPXyy2xFtb
Lrm3kOkMKFdt4ZmZu/JmHFRFuOlB9P5eTQ9T3c7AlYeDQUWprOf35LwSnuadSQExrqkZlhWPHrLm
s66c4qP03e+WwzQmgOBIQX/T/ZNWC6iLk6bXmnZuoUMjJj077laxza5FjBh03JMCdPCRR2Hr6TJa
NbExerixOHMszi3aKcOwbs7S7MztFnWa/XnzgskYMCupRw5FnaNobu5Ag0kqxAJMbdr3iQe/P9sV
DAzTmLbi73ZNpuC3kH2PI6VzF0i63FLaAKGwI53u3UOHFQQIsemFFnAwl6dOaTW8YQjcpF4CUcT9
xdi6eU8Sqg+N+YjxGVpZd0UaQ8zs9AqKq/3/j2ctz9LaVrBLQc+qzKvxxxzX7ohht+6PMLn4Hrpf
/Z5v0uqLD5OKTYz04T939R+x+s22I6cWzCq4vIdgiwoNOd2awy3NqulNa0hrhUAnZu5zW6WILOt8
Nvv79qRmpr35maSuW8TnG8hMlGO0u2zQapEtF6PJ91K6D58jtGGdiZ5zS+TIcI0z/nWdCIeJSXTY
7FotvC/0eKI5wyfPBbrmFP5ma06S0LxR92m9HDsHwkN/4XPZPL8g1V0yCukIkSZfBCckYR/ofDn6
99yawpJB+wIp/J40ODOf04FZzda88IsWpc2qMqQBun0iMcJfnsJ/s0+XC0gu5VfZEj59q2vA4//Y
7r4HfQ18G4ufX3NOYNzyxTt/J1E4fn88QYT8UvS0GX8t1S7oGW2RaSsc7VSOXvHVpnPaqqteOI1a
2/tH5KKp6/Gnr2p1wIGQ4Do2l8UK8KnsW3nlKv777sx31vPh3dDerz86Ovm3FFdJVTTZFMkuPVTH
WuzQiBianRS63Ds4cey8hRvUFfpj4j7sumrBilBCBCls0qbeKn2WbQ2w0QdLabU8xLwcF4w3tkB1
AR64r+hEBir4P32YOFu8YXrI3Gg6SKEMLKouum8Zlfa2QQ4giwNka6cciBsM/Cgo/VQKh9lXEauk
5v/M3fKO7pSxtqogkcbqeLUZTBo7HpZ9iWPWA6es0GtiLh/x8dsyTvCHGuHk/oPdrG0h3TzdSL2M
6iZNLXnmRqFRMefJeSWuAMoH3J6pm6GIe0jl6B45M/9yZqxy3HJfHmy0sAwC7JVwXYgXjrS69zXv
kmnxWHdbO9P7Yp4ed/jC/elHtLQ9oIfmWSmXb9F86BMa5KcmLCrBHoDPgokVSoDlxEwJm2pLKWwL
2RPqE9F47ItfLoKaNU/hHmYIx3KNdfbTgm06ruG2SK3btCntJqocx5GtWfySJnVpBV08AsEa9I2W
hO5MObGsTgBO4CNpMfNdmlIf7itpgE9JLk8vp0S4u/2VV5tRdvowHoStnG5ZzTDL20iKhia5phMq
rv4AH2DpFaSs7y1itM29WixlN9G+u7FwQ+BcXt3Awr30JZPxK5kUgJyVh73Put60qjU1mXZkMMip
kg77TpqC8pn5R2ToaBhAk8FaP/OjQHbG89ThnfJ3i2O6uvbX6DqBggkAKMyWVUBI8ZN+phIUjWe+
U7LPPhEJUUetCUCsYppfYimV9WS+kgxbYpWDwrK3x78bii1ksFb2vpGTteBsVUbF3EP3/YqOYJt7
H2XPt5TP+9vu1Z9pDvVUg1SHxTkRQIxvwlHJ69ZRb7WMqYoZFN9a+BW9XTvNTd5qVBMg36WPgSKt
m0gAWwLb5yqSV9O6FP4jYZLWyIkUWIv/8O3+8CNIM/LOjT1QD40Qbi9u7/E3mNxYXjyi3vxMHnpJ
SgK3Q2b1YDFCJccqk2BObNu3a+1QJXHRK5h0qhbzPpUK22mybZriip0ilTQLNhQXbhQWyd8Mlf/2
/d56l4tl5tHM8xtEbr4bBT0AnMCE4h62tJWJhWufZVip0VZwOeaKAdQyJdyg1SJZ55LmTslsBRaq
+TIdp0gr8dSQv4VR7QBj9f18pWmtb1/BQobODdN/4dJ2Rp42hTgtp6Bud1gquvsdsdUJUsuzJQh3
W2Cnc2ADAAwFyu9C/YhffUHTWyBDx5+WtwjgthCleseAXBAzJMiFmox0apLBL7REs7rkBlOXrcKg
pBj7tAFzf9S0vC+qWix99RWQkbXJZEF0VTtJ4c0SWUL7pfhN5HV4M6e3MOitsN2oNzrkcemKZX5e
l88mV83ahROwZHgEPmJpIAqQQ+lylAQ09ZGPxNyBskHRt1DqiXnV8tCGxIxqwdFNnfvtafwy7tQE
ftYnr5TebY9xrR3cVbdJw7AgxV5+dQZkVqod43DyJ37OVft5k/hlnUFgyjEQEpTpebNY2QOA6xQq
lPmPNq3I7eRdocNr2lEVkjegBEwRO0ILSM2XIvRKXkiYVLWwy567QPuQA2U5Ov21ZG6NgnW8bbZl
Lc1zdBg8iX6IxmtuWPhTetwtml6eKuLfxjXwqIjM+MWTJseff96R1KQ9JIPPMHIeb7SlN0rcb0jq
ankn2KV6ca/oI8M5KmUwovl0HD9eT8w4nEQlMyE55qxQtn1xTQeFTpwWmYC+UuGAoFPtczaxzi27
5qMNIBeo2tOSN8uCxNmSqDwImP2mNf7ZOh5xvYz8nHTnQ/2lcSQn973p05twIfdWq1LqppWh0pfY
0/rdFuq1aseG6oyOjJxthSqgUxeUCQsiUg/Zz+rxpHPLe87VZCKQ/+yW6QxQqpWWDR/vpEBw+RVY
C8OPPG1SCVpbWhsitcm6sRvWFdaKvUzlEafcgco1T1skei5jyaxq1BWVvYYMqiX40xTbLGUF4vu/
Hmet4d0izvK7KuVuH0pQ47EbLRA01dsEdwOQn+/QNa0CTz7vRXiJaHKsKCwd/MShEL5Scd7gHO1A
1SOHCZkPJH2ZDkJtAbcRkyex6rLB1ot1CRr6hLLLZxKuvQUIvjEeWVFvwOSIji9kJkXmHQ4WRDWZ
eQlth9pPGUFFCxtsykLwBA/lN2lMCu5IORYeEp/woAf4Cx0/pIhoSxaHeZmZGWbO63r0a8OVbw5N
y6UmibJ4K4tyMJqTZIQFr5aV0AbwoYj1I3G+snqFnM52PFJjaD8QU2/GmenH4L+zipWfuVNYjOdD
3toOP3CwoxFTUHbvcOz/tvboS61J8GZCDHcQoxSuu2swOn8uU1WHHDwliZbQI4Q1OskAIbV6NCvK
ZoTyd5AMQZiOCTOEjhHbNlfCKVvTn4pnxrcVDgq4ii3vdpuNdjW9Z3RjtucxezONsSO/WZpAbusG
1eYOPWQ8E2AMf7p2hrPgBjIOnnBkVWMfPABC8tbezKmOaicWcb5xAh+5/3HYh2Gy6YwDOulWdwGw
QAFHWcXVd+bR+BiVnInkhg8CO8Rz5tWp4doXRpMaSUFPt3yujWx04Qjrgv6541rBtfQ3+MxdeMzL
cVvOACV1sa5WAPhAvs0aeFc8szSffwMLOhY/IIYQxwpvcIzEB7RMww1e74DlvwciROgZ7uPoEv9W
BGB1uVwCpS2P7AvVRVEmkzDDRM+AvLlOMmatKGPHQNjLYH5+v6dEP1iTjHDQKfcBwzpccwT6W28l
hvtRDc1731zjfDK2vDTgVEcJLj8uaGcPMHsKZ4LhBkkcqEyKsl5r0L/rSwTBF+mgBLMjNeL7kWmM
YV+P9cZusvO7Luj3ySKHA8e1rsMARhwG8gGCAviqSIP3yQ8CY09uAcmUkj+4RcvsZjeW6tuvzXwG
BoSpMypiMGEAGaO3AKfvjkMGkUR/lhe7Zm+gACxPGTz0Hm56LEZ4mQtav4StE0pxH0RMVhTNF8cv
azgvylVsUO5uc0MhsshhUf9E00e3qesWZg3kgPUfEFeOvl+J05mceW0GktPKLmWektDOelyvftaR
BPO5fS6LTY8vBXO+a0wbWobFWwwXddzycIP/XB30elpliMVd2X3B88z4oVF84Un7goUf1T+NndRC
ETkNsyEsL/+0oD8mrp902kLRZAEsUCqyjthUlSU71D9ELhmpKFlZASUHt/hTbpWaFg9iKi30+EEK
cwFfQuO6cZj1BPQO109m+ApNc1G1krhP7pO68gaxjlUibSyhnR01ZEvAF2HpAQ+fTySqG4LPNmu9
mGRmj4PssCqXLaH5DmGocRkeoeWK3dAoMZREjLgfuWQGubR+Ef9u4gupBTZbqYAJXTEaZIxz7vJu
q06dl/jmG8p2cWCyJhLjBgzU7VM9KZrIUlSRk/CI2YM0rUzc2/hMXEHj+li2trw1VA7OOq3qEfw7
YsdxUz/YHF23sLqLhJaEaW5AYU/zM2K5utRrRdCn0RIxmB6LxfB2WoBEx22RZmoxGOsK5sHk4Hn/
ixSWwTmhS/X8AC8M4AbM+TrQnbaSqQa9q8cY03XGPJ0VYC9saDwHD60TzTNPlpI1OoGP1IOOdWkS
8CXTlTkbwM3FB/Ibt/gLnmJC/ZI56ScOCC2TU1720lPsAdgnliUeF63H6lPTD82f35GWOHjnEy4x
Hyao0OYP3lPkYh4HEHB9wV41tYiW8z0AM8ilspDpVRL7nCg5JbQZgHS58pTKPiIXG4h7B7jS+99t
zG61wOLWwwoTfphzy9FRa1RD+nk+qN8qfMiJmfTvs5c2QXqvSogp245VBzB0YPJPr5tH1GZqGh+6
sdqBdvkOji3qtkdn4bCRS8tlvhBvfrBDyZg8JDHki5+4q4xIMGCRtu+3pAItKyOVIlrVxM3t2u99
Frv/bLP+/TdoVRaNks5Ipq+Db40ydsZvK7zK6rHRuBA03BOhGy7vJhQRntlBPDbYQ5BDI7WbZOmi
IUFe4bNAoCBB8cnVhymX0M/s8CvIa7kr6oTqH7q7gAJtGDmG+PA95QsTQgWiOmNvJFqt/PQF+nnL
WQ5OsklH8mOSBpxvasZRBYgux567w7GtIKBm8Vja9D+85kVvck2gDvUVCRH+pGm4ctJRRO5KPdKk
irJSq7tKBwZTbO74gKTFqf+9B7G7BXygxSVJZ9zePFP/WhftsUUeRH8N0F212ELyxZ715B8YyZz4
D6cncP16aGGq8FxERrM2DngyxXMtewvXjkZS76dvrdlnjFEaeg6wADxNz98EOYSZP1Qz0iAybmoL
5fPpERUcO63q+3CB4RLJTsogEGr8B2+JCTK9Q2+UmdcknxzLYwdOp3/W5t7LJfP6KwboNztAKcoz
xezLo+B0D6BTewTZ2idqnR9L2PPilYRibJgki3KbwP1d4pDFPkXz50EDIqnQaLrGIHhcy1tla2/j
iHjvJ4Wp5ilgvKqvOzrYlEICuEQ7I1WvLWeaTEiDyY79qa6EFhgo+PeJqC+k+1puogm9jUb7vmTH
SgwkDwQFdGkJBewh7vGG/Aw6CLFrL4g/2+cxyXWgqS8kIcatX9whYROaO+0FDfLfGtKazIdK3Vku
I6bEvGGnFqUW+/gIlhc5WF7HoVbONuuE4S+efDkuCuu1feH5eZJZ+aTIiRXbVsNlF2fj0p4nLweM
Uc3t6UwHQ2/sZc2sIYTBRiIkI5De6Ii59aIcn2f1IfIGt79+/qNrEURDT5PYsKRkfpMJ6iL82Xhf
t3eyfbc6A3SPIoishhjfESc+km4UxT8OaCJZShvVFaZPkJmwDyUbTOuO4AJJ0895LwAVwOVdU0eJ
TpPtduTmYlFXOcxPlGh5Chnn+W0IN236NSe2RiDFnXjGKklTyaN+vLd5zuiP0BcCT8OtbfRoj+VJ
MQ2AkocijfmfcH9jJccvpKJfc5nwvl4Eq4gpVf0Eqr4W8VpiizmwiwaDCQYMVhCW5bxqTNag4rR1
gr8jkgPXANyxAuBfanXUZUGwlNF1tF98jbn6tEOmEkOqYKKIF7QGGKIVAprSZRR3PLtMheHku6nB
iy2Fq1PSnRzXSEuyhq5v6xs+LyxEw9tRKFd9Q+4h1NEr5K1qbiLm8KooaXjdLe803nyXUOIjB51n
O17PPD8vtdShqMowpjARtFqqeirn39WQuRDRAUxhBho9SQTxVLkaAcKWTJVkVgHGbmjJcpp3now1
5i3bJMRQFalECWbQKINJELKIL/YEPa4pMxVEAMdsZFI6ybQgcFMMmYMdWLw3oEY8gwm8YUGKeqKc
e0daW+26KzB9Ox1k2VfNqV3eA3fNnlk42ySYnrT9LRU8XoAZjdCu8FPBDVJEZwT91FgTPEgGsYBV
ES0Ds9MLtAiOa1ijI111QyTG49DzGo3ECJeJYVgcRURhI3eK+//PndDWXmY/fwuaf/gcBDRYMOiP
RJZrZH8mdX4jh3mURoFGYZrcEmIKPD5gGLmGfaNOl9BR5PnlKvl7b6vbIThLHuuwdh4ZEjnzZGQE
DZGq/qYdRqhI72OeW6W3etG9JeSpagPrk8js/DEeS/HXxRY6auLSe51IxBQfHWHOL3vx7GjS3rOx
lfx6rs7/HLbTIb0oHZ66AFnOpCp8Xvgih5jfc/6K2p/70qd72TmZyIM06bN7hmsgFncvc7smY8Ux
0bSzfhbB038as5/MFhz3bo4gkSkwXswq1C1rdYwJqiqhkxf5rpV87uvjeVnmcuv0Fabu2H44ju8z
Hcp/fJE5HIAEtzOqBDb69zgYNtyKrdMMpKRHimIVSYyMM7Y1SIq4d9yALMwJ7SckVWMz2nWrumoS
6gEiY07XTEXAA/myxSThyM6hdueUqAgdarLOueoS0/Z19HM9c6OeNhqiR8UtbR4YODgmhUtjhZIO
TG8g8GQehuApkXC0ypsIQIEBrzIRYBs40tEOtqouEsYoxM0DmsPw0WgV5fZYv/8vKi4Mz/BmaW7g
vnpG+I9DeQSBt6KUbfUnvrEvgEwJA2J+0l1PXHQE3sv8bjcChQyZMaImEfp/qR6hJvfN0aNqRlAN
LCCkiH3anRvD3ykw7UV9+JiQTG10NtpVe6c/r5DclOQY4y3alsG32jDW/ljFRsMI+8tA0VjC2tKd
1L+V6qimLjR7GfxDyX8QMhcg7fTNlx6c1VLAWLA1hbBMg1aa7SluFyT8JbSTLnbzLZe20pVQQfa1
lX301MhqF278ZrkPKN01bvm9puFduLx6tGTdLlIADGGghDJkbTGIseSmAbwxPZsMJFCngCCbSaBD
XeEqVYAppZgPn3TrW7QF9fkZ9Gw1gJl4NO8HKBV9LQq2IaEcDKI8LdoiScUh8e+Td0BdNyVkObxm
Sn2ZZlQANtarr3lOSfnGv2NGBievYH2xjpTJRPwVPSjE0gv6o21MI2Aluo/0X1BDh6c7rpQw1Vsh
Yjs49oE3IhkweFlYTITFZLx9troYlNaCreju9fedMEuh5ldLIZYxP9WoHfn635pTWPcJCfDYkYNx
zjHgcCTGLk9y2ILWS4sPcxH8JFTL/wIUQ0YPnilgKdg1Gfgxsd5NA4pfhgUGhFm5w9CYk4hxHNdr
rZbsf5k9klXr0jY+N/pZDJwK5BlompTshgM3S8cyRj4Y5RyEMhXQbdXRawgFdilEohUvExYjYmmm
TmnuZoPOZCRov7WJWzxzYMEVETRvVS2/lXLXBMVkPeWIQcRxyYAXqh1D/QA8gA3QqC6QE70LA1mt
TAhK2XAs33yDiWf93ZsenHfj1yuDdLWEferZuHth7Z260dIxLYpwuNI1bbWSBF0c7aRySmGARHBv
2WKe5gpitC82TtQ5ODARbNR9poQh8YQuqRd4AZ+U85GA8YiQrLcVq9Qa96CfmOCZKhVQ6Psp78sd
sGK7RLlieM/xoeBjukkzAmYhfQjueY0rLmwtAJFMxyMiPEWRqtJJRlTQl1qp8ott4IJXCm/8bXUn
3ZgFzey1etAp4yEtMLDV4/SgKCql/FZBoEicGPrE1Ytch3uydbKhhJCxDqoCrSvhKoRj1v3Nvci3
QGeqfG+dWbhMRE4uGI5uiNwizgz8ZpXN+/Ft/19NYxc6P7PGGeNHAEcXPDwtGQ5DkiFtKKuDVuv8
5KRtHH0XzEn7KWoLxVibNJCcLavnK39veV9BBbseQHHAOCmjdbJ+h+bXQ5xOSvg6HxyKjy6zExit
TCfo2f7byNND0Qr2HVheAzMWC6ytDieINnSD+4DNOgHEZlFQonyQI643LshKgfeXBjcLTN78QPd3
aKb/Z+w6p/6Ugp//gb+zn6hIe4H1cQMSH0WfwUv1bezgcZhPGHkpiO5QGNIWetV7Sb4k2RxUlaY7
nEzbwm24mSGlO1GxVfQIFBK2dFoSAYZnMYRVv7Eu0KhTpFuebgb5DDQR9eGRvghhGHkwH7opnvc6
aXW2EZEVAe3R7vMl8L8kxp0EYkFhl4/y8adYKT9HhuT9nw887uP9+ViVQ+ocAGRY7eIT7CUZ2YWt
3lP3403DjY1wLnNxDgN/eG9QjOBiDqbkfoni/wf7DlYAqPe2HWS0LPCe6HcSOavIo+ScplXFkMQW
LejWBO1CQKbLZHdVkr/QeOzPejK4Y1jK3qfbq441ta7h26jxkxzgCUjumM84cySX+MYs1G4KEhi1
0M6n/wd+/ntxv8rmov9CaGdJitRlw+457uNsPQ+x01eXD0Wj6h9yyHH0gLXUFgcPYAtZ5OVz6FgH
vLKLV5D2L3xmf78wozmzQT9DhKTV85DaaGWa7SJ7ZSct4csIrjVd4V7I+saz6No72+JOqlunUH4V
1ZAjJgDovfDzUbGFndj+GWM31W8LJIrVYKA8dsOJOlPz34T5AGgrknGqRdETedBsCxefP4fw59tL
NyLJjoxPySOy4iEiZtKIRUtBUpU0b4W0urVfhEPynUx06qt1zM8xIO1uAjZDT/pqq1++DYCKwCB8
B4vJlt0i79WETfE02EhTHt+Y+ck0CpxL4VBZJjc4HI1LiDTjn6Y3yWBxP3M/tCDMM7Oq+k6iew6r
ZWp5QuP0xwzTOYBI8Nf6TgaNaK3f34gXbVyCUYFZOo9HK4dHkYC8JHueGiq/yJAw5vWFtGpNw824
ExvZ1qSbHjo2jKxdgo5bOQv3DQLJu7unGhA6MIMvzp1VR8KFFL+hBS+02Wvbe3JHoCYB8koKb+Qo
HAYWkPkrIULzXtg6Ah8PhE5cN4qbgfXDM7+Chiq7Oe0IFiwNljd1iA5xdhPUlwWZYl8aSHxAePn9
1CKUG232AFwVjq25BHQRwPcGiDanumziMSKsj7Njyafrkpyqh2oMDgS5VFVPQtorKGzIsMAOzcwM
mcn51NarzCItW4w+2qL2ASND3oDXtwFMxqEPvMNHf6eFeZXk1CZezLkE4/eAnXV2DEhHDndbB0W3
8NO2DsZQjG+YrgEhLTH8BR99us8uASfCgt43HC8GDmqV5wKuv+qfMu3omZubL6bF9BUNeTT9VGiF
e+3wKIhAz5kKxfUXT3DaCmDieCK+RtzWco8wWCBZY8TZqSGRFEdk46+p4joL4towoecBzhwQJUA8
PaZiyniOCoVuSL7gRNsis8Taw3r8wEVXEIUGaGh7hzPMOd08iA0jk1dlWoC7VOpec8TGDlQ7CRHX
qIPejfW+ZsYnaGd1d6MEfH3ZwDtgmdtmODsBvKGFif9XmX+g5krNM/xZVaC+OT0EFRjsXx1RVkJN
d/ji6dEvFbhsuX1HbiMnOc76e/sZ+2sIYa4vtBxSW634kMb2tU7XSwAHnmDZlY9+thRBVOheCc5+
Kh0mifqW/p9qm0mIstQpDaAIEpGPoeO9bwmFvsLChDMTGNyZeTEJhhrxj+Qs+gGal8jxEQtdrUWu
8XOSlQUvCkhN9IXxcLolP66xWaStMJjwxXBHg/zZTuYPAvXDSiaLcbM8uUarZJjAbM7z0lCK+eEy
qnE7kw36c431Ym8pEw0uPYa3kuwXre2+crOSinq7c1qZqX8w7ae4BDtzEN5fEhBL4C6hkVhTEzrs
vZQzmIILDiWC28JgGjQnwMHRkiS9nqlNV7hBR8L5WJvL9OQJwRvG3AgKZiMYuDI4q/k6sfMfXxOg
JUEqMJlORVelRdZU/vgbE9ShNr57ALxCt6grYbJMvegEuzJ4dMWo+uAz25ZHvgoufHUv19jGaC+T
7xjSpJ7RqGLoKqeII/OUxDcXKm/7pDlYBf89kApEw7mlam5qZBWVbeaMpnjU1upOsB0tj/II3j9K
6l6gUS1RHYFlITferH7lUWMl2KXcOMiBxnHN+8bZ/yPkT7qz6aFwg2Otnb/UHSBkn4Vuag9PcR6D
ryKpDTvlFStRCz+gQ/6huF6548dfgIfCYbR3XO8UxAU5W/hEiSzSyUhEnjjCNALZpWVXGGny0n57
AsPWYAyAqcRcwWgAiJOQNzdKqt0G0/KJNUztmxe+Mk+rMgmq1E5+wqfVYt5xa4DzsoiZ/KYF8qRr
f8HSzW+V04Emt4keNrpgNdERfLNGC56Vdy3guFkLWeDAfRLZ8m3GY/36ZnHjtePqR4DxHC+vENsi
ZFQPh6kr/p77gEXf3dayRjhwamPCfIbSvP3IZD3+4FacWQNHuZBIXsxLkJTXoONmVqRCBrp1kC4K
TBLjlgiDscq7fIS8iU+Fu+9A9oadvbExWkiOPUa2/DjiOb2uej2aNN40x18kstM14nA+FjOJyuAb
9D0M0ouDKQx3Dsc4oPZfGaJWryhEn8hFelR50Dkg/++hRNdjYMIINAgV0Ye7VLWBpEPblVftMOWd
LVN7LLxw7SUEGfwjT/ub6fCJu5/Ix+I+S/p7gpNrpQNKVSO+Tqn3AEfbJYDEsL7dhPnL1MI2wWhF
XzYhAgrMmN4YpFnHQSeR/h1nEOZU1LKEMwjdm8lgxd8inaXTGUlptPAfup0mV+UlqWHiuS6IeQvp
M5AsPUQN/OtZnIuW3scl0lqBdEUO5CWbZNd8vvXkRNvJTD3xsEI5miosNTbhs/6XDuMNn2ZnpLkG
RgFSv8i/AIiuBp6/iuTl7igbOuua6Bmp+96olYPXbZYnNl1C+5NT1EAznI/N4oozEbvKPyUUJmB6
yCZNzQclqNBINbDQBSzLhACNqJiCDBp/3nKVMWXHVMUWo4QHOG4BPy4YJNuwczMo7Jjo9ucNsIdV
AJXoeNrbyl2XfAmvs5ivV0Jp8TSkIiUYYq2wOrGsxBZkZkj2pNp+UPhonkGO5j001qDqa3nZ02U6
RuPFisqWm5j02IupKkjJ8qdNr6px75Rgkv1CwNuccXhdhDwMC5QZQmaRBTJSknk8EizyxiS0FN4q
JopFL7wGo2NLrcHw15R/TS+pQ97apUnaz+mtwOG9TpZdnhBSOz/Z76qOmMllfrgxSlCUsUPTUe5H
K8RJe+o2cRDFmi1AYLeZjdMirC7+9GBt1cUEU4JoOKkWOULb5dlSQJxxgO5PPYGMPpY5KCr8SWHp
zyckl4Lc2dBl4J6SfbTc0qQeqSIyMqrs4iqENR3B9CSBYpQYexfT/kE1LRaIuhCx++28W0ojumXY
ewaJj9ZYjWfmLlG1l/myphR9fFEzaSuz5R58vtl1D98t8EfyAJgpQy6/aUHbH1U/RkpKFPGkrvNO
gwA9u8BF3Gk8ay0h+pM9MQ8ItuSPpE/RVA6+8njKnVTYDMOAAc0tvuJpkPUH29sU7Cy+W4DOzu7O
PQu/Zd/+M81IusKh3n2ANe0aaLQx8Xte37avQxyq7OkG6brcctdmWzYIYaFeGNpuOt2H3bU9oPeT
ADHBB+Lwt8FGDstIXRvc1EcZ7UsnCJoPexTJPJrru7gc/ZxX4VG2np9Bbhz5SUZfva22FFowwM79
wDYf7SrL36/Fiq9tv/ZtYA4ll8WnQHHRl/4vzO4CSMTm7Godjp3g0obegqet9H30Lu+Mo1Bfj2v4
gjcHQq0BEYxOBbyQDjlPtEB1c4wwARQESHjt4NgL6qV6JqFOnDQPPlpwE1P4yoFfm6SC4e3HHEXM
Aj+hEFVHAgBbk/qqcsE1a9zE4tvqU1nuSPkD9iE4+VdyWQlb3jIXr8FDOyUFSZ+IebE8MCgw4lgY
OTxc5OsFHjJEagnwtkhhzuSEc2k/AqQsEGsDj0dF47I67Lhbc9gnVafrq7vllAQaBrOR1ZnX33CS
yT505YSqu7zpvmm4qO/tUkUPgqGi64tlruJUqVtJjF3YNOPHZUrXiKmXtfmkC18KxJ6IWsro+I7e
H6txdHI05iFmTY4bB5DDvmoij5yI+slXvzdfAslA/aivMEa3HSRMfdWQDRbO98s0UCfLRJmR6RDg
uIlvtDLYsE1JDa97PQKiHJ03nAW2K40IdAoUQH7y5LXqvEjSlS/EJxeyy3fKSmcYmgFbZhO2HnFL
BSe/ZeCqGKLcxzRUYtibae2F/e6dvL9Ua4w2Z59BxwLB+OE4HGDbsUYiMXgv6VsPHRkXeoQwfAOx
bRGASUpvlosQ1ocHSKAkXY6P7CJSyeCB9EpX11kuyu5IIPkT4cT+I7kzUlkp6bEltY7tLilfYJMi
QwoBTAAG98Y3wa7UGNV5fTy4aaMpPe33O7v6GrFVNd8pMOsVeRxLmw7C4wf3VgwBwuiViaxjBplv
xvbtoMvOMY7exuoXyfgkBu+XcjP7D0eacKFFvBp/XLRBr3c24NZje07THtUvGeRJoBYdMBljkkte
PDvy2LVMtbo4088bCnr2b7SXCXsp7gxjwz8o3ppAWLx8mr0ck4VSlrLFGOHlLFVglKUFbw5yj1aN
nKSnEZEjooW6BixdRXmwx1SgmpOoCRk7f5v3mxo+1nfIy9LK7OqIVLm6kuq1x3yKgCCjtrNmWYnA
CoImElAmcxsbeHuWibcUD8nFJ+lXHiLtVjaU8ZJP/kJkzCIoMfQuL4RtNwrh/U6cAC4pOgEA0WGD
+0vwr6J+Rw/p2852uVzpu+11G3AWiFkkvHYObN9ocmR2+dw4jMB1nYAp/k9tVc7BNgSXLVq+Xy1v
8GQhMrTKFb3JumMauhhgL51ysn36AaE0k1yuwzzs/41y1dyeVgUqRjaQK3isSyzXwSBTcWTQi5ZT
pMytk6pV9kMxhrWsazbCs/AdFHYnZpvCTbRvIQGRUB+XYLuEbJB9EN+FQpoXmkocnLX/Lsyt+p6x
ASccKzIs3rqilDIVQH36Xn4IaeJWYRZ8gxgwU3saqnzqeAGHl6fWuqthNRSrSbPbjFRg7U8vyJ9k
sBepI7jjDNnVVTxa8PW81mwnXfwBSo5rHdc4Rgt5NVbjNe6jHDJGk3pcJqPg+QvhiH33ywDQ1vz/
ggnYzJI2ISxdQK7cbSlxBZfLn66U9gYjo3fLROHPxB+jpvWdg4vm/GbNh44IcbNGKtXGh1zwn6pl
ioHxe8bLyLNNrzQAUWcHivxrGVfmwlK4XQY2PFX22HsmueeMtreLKQyM9HdjILRL2G5C0T7UlH3b
gQaEFxfPNG22xsIDksJJRaxccV/Qp2GrBaD/brBawOn+7I57n9mvY2NA4wgBZMOzRUdu3DB5auei
3b8pK5DH/05qEwM7Vwo3AtY5aWHUb0hQp8hMrdarBWynQVZcJIcXpi5lAepWXYdjXoJrD9pBcrbX
qAfKuhMxQOnJ1ICHXm1r0smMb9rVlnEOTyT5wKgIsk7+eEL5IGIAMU9nASnO70cq00+4Emd6+zeW
7U9Ykycs4ZpT+kc63HMo8PMTmNTTisME2+eHD0LPCUrLVkmZVmHPi7jR4JzND515fVDvtQHeKx/5
iEOcGFmYwYIWaJC5nHlLA7i4EOPmWss7z71XbBZKB3UCYMru2OSF5mAMmoufUWN8PkBEOtGJVjNH
FuZVtev7EyA0VrLLlAU7dN35Khrm9FThQgBCn3YfF4q9FUZDljq2lVPU5AuLBGVxQ0r3XmGx+K/6
wbY8XrOTAJJR7q9Ev6dGiMv4s26kfRcUI2X8XheqM9JZLGhjAtSRgij0MwXyl4HsBrLYxdXWgqyB
+lIY1pHYjKggJzgw+TEI8qtTK8I/vLDzrDb+AjJ7FvCpkxfpxCjJNfY87DVbxi/dSnpXsBhRFnmC
D4+45iNv6anql9afzr20pqe3CJ6zHReuISoiCnXtZn1TUJeXuIuhtgQmwBM1GmFS/qwTxyw1Etn4
CXFD2e/gld3zrh9sHvwVEkOUpQB7jF7NQn2UVocsiriFwSzg3LGKpNNn/qiWSQUwtfNkPvCi4yzg
iBKnkd3tF8hGQxxZHWCkiJUGqXJ52ZqfxhvMVDxF8qwAygZYxUounJjqrN8NYswrEv01kfAtWXeV
N+mN8tHi1hZ9niUmFXVZdFRWH6d2XLH2SVPU569VyoPEFb1OZNUqEuFD4Wdgz5kwS1PEg9WoDBNI
/Xb5jqH3qNKp+h+F3QRCRlE9KO1YKXBeCIaMF3vGbCnkRKe7cWDCpemP5d78dxqZrnZ8RpOkzQzT
O2b2rb1g1FiEmdePxb1Zx3vKoB9XNgB5Ug3gGwgC1MjzpG2yBpf2BFTkhkwM6HWYFS6Mb+S1a7lf
Gr1TWswdAwn7JA+Kh26e5W2PCt0R+xXk6WJU1/t1py4x+DmWprkZAJPbFtTV4SLd82HcbOET+CiR
6/1i1txeAnISpZz2clJzWuAgZClYLUvaP1O3W+ZAde72tMgqEumZEsWfdIK2gL+qQSoOyItmwM0q
DFfdajoFe8a9D5ZlJM2JD/7LN0tJ9sFeM9AAVoFPHhtBpSubHyL2+HRf7SPYDd84LjmyFw8kuMYd
EC/NZb6P9FV8AGtvq+L4SrIoPLOYBfkGYBNyKwMw9cMfQHuExJYL4YZ5tkfofVCdRVuL/i3uGXAZ
SlWfJ/VmjxHL1aanqqeRHvoOX4wpV3Vy1eRlRozRezgWoSFix+aWtrYLPvEPrNFvgRfKyDgKEjMT
MbiM9PWXsK14kb/DIdq4/wYl/VUJ3Mb2GaGFU3+yZMZKdPmPTdUZPgyUwZ65aKQBkoEuDOgotFr9
JtdZ80ZeqStibeLO+G8PfFJKs/ffROsrQGcsYvfCuKlpdlVYfccLcwyoKD4zKYLL3DfytRoeQmT9
Yjxl+Se3Y9BCM481lG7Ka6lmIKlH/FlPKlxnPoxSCNYJIQQb70s2ZBpbWezQOt0e88slUCwTebsI
VdHo8PK1ODZNqe3RQ76ay0PILflkcL/J0H6N4zwG8+jUHpXVcA1CvXfmF1deafs4zrDXZLxeWN36
n/jbvxV/sRVcTEpZfo94/GJ0Tb6XGjQ2N5bxVQ0tUcexNfcD9f0zJztZVKRhD+4ON41/s4XSy2gY
Qb4/a9aA/To0cIa9UiNEEf7iQgY4bskxx0UhZA/pgqxujOGG00onCz83vNpTvYldYB29HQv8x1/F
Xe7STejeJfU51VLwQqv3JRzZ7qkiBqbwzLF9Smh+wxTT5aOTWGdJPsrDmROP10qNeFGfRuhi64lx
ysN4VvYtS2ma5iAs+yDpV8Rm5Xqkp2QcYWdyy66aq54LCOkoG33wW41Kif7dkTHUQtaSvN1JCZGG
2Vw2hLmcwGpbY02DAbFpB77xpm8Dh8WzXXQfSJA2NkjexdWtRoQPauJ2ZZjx3To8vBbb1JAe3J4U
vsY3lmylOP+aNsU5f94UUtUMOA1Gbi24UErEVeTyYFoMUDimefDY65Jc7o/nw+c8WSp9mvY/cbaF
KNJPqAtLsuyi1k46SzkuoZzU8V3RY49la6NcetMZzvHG46THnTEL9Xw15tgyYBbrIEqeXN7FsaL4
tITEsaHTOvwza4B7CC9g6DaCxSHhC18RpeAuibfJbhUJbIWsFe7vgGU/kosolnB5+uvgnn6A7gJX
u0oUxMKeOH0uKK0DHIU0L+Pm/gKSVZwdw/hlJEmrEQnkxRK8V7c/icYnx3lrfTfkFUoEQaLx/vjT
67n3ZJlOkIoQn23P3/TxcnyJlTyyPc2pl3hkXb66ldbcTncJFoHY71e6mQQ8uhD37v6mpJB99un7
uhXit7tAzMTUNgDqfmvK6lgI8EnXsyrtMVzdNnVINptOXJNVqNsKOcR3xl56YIv38hfBtJJslEES
AnSSWbU+kWbxwl6CFpBSCm24nV47/HnHeH75j8A5I1NQofrEIV7ecGfnyHqXkKy93G9dGkb1vCZq
4LODnJQkmdGGJKN3KYvGf/jmHbMb+auKWPTV5CkGPg94FMDc0SQdOMWo9Og1AZj9s7ookv1kwWMI
RbxAkuZYU/T9cx6XUIB5g3tytpkH/5EbnxytNgRobOMse0U48FnDdO0MAQ/XIGjKvnIjdnw84WM+
TrUWST/vpX0wfw35UNxCirPjiWsY1DG/9D+1b6meWdgqPJX8aL4xiwe6Op/m+QSHmUcGYwAafWVC
v1/Ff/G6d73bMhiMZQv4Vgq+bO3iCy2pjRq+IS1CVtG9YWTHQf+l3o60ODoeYPva0vYLZit3Xn3r
58wa5wstq5Vn6vs0f5W9GfTBeQU3sNQCPss4Vu2gvaOt77SevI7Acoz/OePfnO0NGQkQFilLo5Rz
RoOMpJPW3SZiogz0zmFmbb7ShHsaLnMnHFBaRNCHNLQ7qmL3Fs0lQkEVRXkcnplErqlmyylsQC9w
GzTM+QjjNvtQQEz3ZD/iTXv860A9xlNZzI82lqJTlsO5R+gTOF3GOacv62Mi/gnbVaEBcKJmL15t
+m6vVR+77jhKiB+AdfUCCVOCySzspocpDWTTzakymDQwukUsmO6NGhLVkNLSO5tQf9jZ2HETMrlt
NJvQDOMHFgJQSKrdWmn5tG3rM+DW4b2n2/WalcTqUwgbcoRdxbZu7xWVw23H1OjEy1CMZCVxUi0d
IkL+GBxCkw7saSELZMDH4eb9d0nXOIGx/+2hUmA9uRZJVz+Ad+R/N8JCu5uy2slVYyqEA75XeBex
jfSShCKP124vnsJpQj8mxF8ozonY8xfLWhMmS9XF5AyKNxQfrnT3ZYmwwyN4/KAACjgs0i+y7tbt
h7uqAKwh8TRpJHO3R6gXZueUGbPLgUXkkdX20+JrL9tcKYhNX1dy/EzoTGuVJ/gx0TPKLN37z9mK
RHRPq+ajAF9MbABoZaO7bEBC6/swluSHuVQfDu+rYBYzKMO20pJ6Ilb5HC85i7r2y+IUkolfM82/
krdYZcXa3QCvrMiZQuC23T1tf5P2YH60dH6xc/aMBDjPmRaHjntNJehmBEIpI5+XCwbSFaTaLkAR
eZhOk59QWLtQPzXD4KayxeLetuCfvAxlwcQs2yjie6Pyrr3YPjNr8KOcpR6xrIViZroOwfesSw2l
jwrgZy2REn2uj7aDgoQE7iB4A42gz0M7lrpvjsAuekfHuJ2tmt7rWS5Zti9dKLCBLMt1ulIqhkUQ
1D/lnUVMVM8zslZGW+APKn5qOX7BomTXsStYskDQcd/UYpid/QtIJYN0Nv0jZTBo743kjVG3CZA/
tkfjJpsTtX3yjR+POFCWHKuCsaCpQgjn2d1hOAGrz3sVXuAtMygbDP1vIgpydc/REjGATGA7ddsu
lNr1Qs2FrMKlpO6dmgA9JoOOUhP0tEN2bAJqc/AtxZi9pnkfOEgCtKCZa8O3EiLHX96yO7A84qtR
Cb8d65bez6BN7hEmfOIHf/lFll5SmES/0CHTVEYwHvuEC+xvPQdK0VjWTveZxzVrVJcDGsg2wrQs
BUZi9M2B7BK9sodtjJ4yuAC73CQlqWXmygOApbpAe+HKy8fDIYcajINr2gNiQrob+w0GeyI1hjjW
KLsdl15kFac8VqdwwU1QFqpCVgi827JX9hxNm47dZ6ZjFjXOPu86Fu3L/eW6/5yHjpVzSZua48B1
2JKVm2GI2P7490fwuh/rBSEesE4Li2gi90DDqF7pazJxNnvxNL6ZXF0Es5KDIVrfCc5629koKv7x
1LYbRnGNqTpTsdJqgt1sfLCjCJdCR3t9flg8O2KOcJFTqnuooaWS3Lm+/tq2Vul7e2TCyNtI1HzM
Pok0TlZtrFV2BP+PfMLJI+dOeSmHJsq/7QFe6i+ejJytOpPTItB38y+hjrsfJwAIhYz7prXQGhTj
UKVpa2zeVQ//50HCioPLY40+CuUhMg+oqCmfYzWjfbIskp+xGmoXUtLcqjSz/zc432PVyv2wtlU1
g+wGL1pUz5EOt8pOvmZdJRfv1DVpaF67v8WixcPnONYDSKMShGQzFxGUL3SNLO6JKkHhuDaRxXLX
9gY71WBEFs+h4GQR5kbUp9C5o1dOiT6LIwFk/HA4dpLoIqpkOsoWmdNfcAbJEyI57hq2yvciwdv/
wsMfY3oLkqEL8oT3AgN4TF3VD7lL8kXMyfG3xye4g3iX58tJtI/bQZzEBttES/2mVDOueIrwn8Vo
dvu+VjD+ih6WMidF0EEDSmsUOKorvaLAEuH7qrc+AdcJB06ccx2v5Sel+l6WuSYvR60zea+ZvO2s
8GibmhKhFUiutgu/eYOuoM+SV8mqKGr105aMCmqRzyLTBYBOrTcj2s3F52q7X9eOleoLrBaW2ho/
c25RUzISKDVZIAhtL3KvR5BPIS6JQb7ah018T0B3Z58pCIl6Qf/F2Z4nnjM7oeYf3ONEQFySRyja
jCQfT3Ec3oCns8qEGBblbVewAfqPzk+JntuHsfvKwzHdN7y01S09an/FDUW3NlC1zPBSbJXH+RRu
WPZu1snEmjffa7kBQ2WV7LAsRtGA5OXehgtY20ZgZhyDk3vEHIiy8XR2YcC+2g3k4T/ZfM/NneIO
29FLmDvL/wJYPqvp/3ME369P/+bpDtzRJ09nUhEbFhBg0M0ZPgxqtbEV9sYmmI7xaejRGZXE8ZPV
aZxb02kgy/jCjjBvmH5WsaYVUDILJIMja0iQIZMKUJqn/pU5n7oqKGXwDnvakcCY0e4tz1hMg2Tl
jc/oOGUZbFzs+HWFgH3z1TfEpMRCKgoybGxYkBEQfibe1LPo33AgsMegI7X7V8KXTvi1tltLeQhK
jnv0cOvPmhhO18uLbQ2DV2tlf19ELAQngR4HnIfas1RgCaQk57mE0WAxOjfCNh73vX2Tkka31C+i
03KD16Ig29C0EUFtkHzdQHyzH8SmwQbz6WLflFyKTiZA0rqsOIwlqRF5uS68lMtmMG3RxQH30mUC
/wEH6ViRXcr3/SgpKAX5cqnEKjwbu0C1juZrBgGud5GuMCVm9AH3UehKR6rDJZuWyhyYJgvkCxxT
uZrExSGbOlkZso0+ZSwqmW6S4D0K5yj1tiF2GPCC0lzRerda2OHGu0g5uiImymY3Z/iHxoBLayxp
93hlavwvbWpBkXw4iHyPOk0USALhM4TENo1UGg8GE7lJGQgQSRQfkYOgPXJMkN5yLWBq6ri0Q3rW
FnnQSG6B7WRmQcMlGqjuzI3dgsTrjnXmOe6UYM+AEZ9vN44CqWVwmHXMkoBstDez+fWyX6Ov72pT
dz0qQCpfZOzFGgg7ntfooffbGUmmKh1U6RVlr1hTD+Xb3JVMQQ6hLVddMZD61YwZHU+6UkTEsfzg
RbMYCjVJHFjunziGzPYFoG6auKK4O/OgMF19xeSod8gqtxGaoPb1v3X/Ocu+M9WDWdHBx17Iob4W
pNl1tnIrOEK3jWWhFrH0g8FAoVOYsS/7xk/xQBcAwIDRcTeh9xFuOJXU6UMiZMl4MISRlJNAgDlz
WAPypFR+Ng/tBIQqIBh31aTkRfBNqK7Aie1/cxrGxS4DaFVEfq7wwAkh3uI9j18eyX8K0YpmCzY9
E0pU+uPTrr3mwm3WDyyiEYra5g5Vm+c3Vi6eCLnPM4IdjbCijmi3G3LRv6nnVnqsol/TsOPyTNjQ
qMr2SykJJAjfkoVPVHi+3TZfrT2LiZBldU6LuN0TTbvIFbOjGHSDE5RLl2NciZxpdsI3q8CH1PGw
RChkPhn3tJJ9oEbIcQmc7UFYgUv7iknfMwTA7axCiGpBiXwD3JV+Ul4kScx0/dRcm6ynaGp1omDM
rjHzvALLFd9s9u+1a0P324aXABNK5OkGwSOtFmVwXK8CMVxbcCSDEmHp9SjkxVavDChStNYOQHZO
lIVdT654IUp5ICcpvCotFOxzcjXdxuuEQSEws95I0fV0nCtuL47JKE5vydlP/F2UTl2ps8c62o8+
wMWT7Xs/OetGb5eLvAWBFqR5GHd7FdojA6EcRUv7G7eX7LMkgolWcTfpu8uWKSpe5I+8MD2ZjDhq
dVbnyeVnJ9Z07PxwARCk/wrzxjIS0Pn30owsQvgfSZ+lirL6sA8TK/by+GaC2I+b8BKqx9sn9p90
dyKadUzhaMz9WmRp52QUOD57Jg6EB4POw+g47aXVrTwiQ2TOuTgiiVgAoYC/H8L3sOT+0qV9OD23
3nrKadhEV9EOnQMPDVVrcDFxGPUe6tiCmn12VO45kEpINBbJPvDMfVk7l+XcHyZvjCswruOb1ajI
g7xzrVZR66BoKliBTQb5SQKWgJSB3cKdJ6HWC+L26zbLXjK9knxUmPQxuWlB/s1eGw5JoQYnfUbq
HkyZSn3xOBtRBAkDTMBaN7x6c6s3g8AAMsE/F6bgwD5A3zjnnes1gVw59t1IYrjDp7Ptsw8DFDJt
Of2Vzv1+YChlJf4BgP1e288io1KmcWHoTcvMz6r5GICUblXF6806XU2GLviTb9Iv4OY1ZUuG0lQE
UtbQIFy5NZf6KwiSgv+cD4ThDHgwL+t39EiBens6HMliEXSHycon0opepPXXXIF/mRwLiYbvsh/6
EH52C87hg6NX5pngXxKvI35kb0kPqvrPZt5Gj0Hb3RzTKQA7jVf3oEsNozWkAKfFOaYYBcBCFyCT
/oyKsSPHmDSKfWaB0/FlUU5TMQqTPOeFopmIfWeUqtb2RW5NLrCK8OhFkPi8EdKwOuz2AnqoYwwN
LobIXj0IA5HRvTmEEOANquy8YJBdj6SNIhotBDp0phKWcLAPeBNn7fsVjgARYNsysOcIEOxK+2rr
RSlKpHOdKYYj5xv9ZXv1lIr+8l9TXXEx3L+m2wQvKC23FuIOjJ+eTlqPHF3T2LFNCjIo/uBeQPpJ
fUJ/HsZGXdyT1g6242ciB2spIROhFYQtJeuwB1gbA0XejrBSu9SyjNrBDHbMeMFO+IVjMWw5kf7r
kDKqXkup/u8OBCapkNukr7zeu1D/Q0ahuFq7fxPYxkBRfx3oF4F/c0v/kVLg+jpjsOQbr65b/wab
Aqy56gEe7AViIfkbN9rkjpiZH4Jx8UDTy1onr6JVmffIw/qgCg77uEW0VBoZPUSbG4Z9dfWegG/V
wi5qpnfeDtzQBmn+ipp305lp2Vs0J/DUXmQT6kvch9soqH5JCJ45NlPlvBL4mU4wXd7pWzeLy9qZ
GwIFjcX9bZXcysOgUP4C5grOqtchJr5jQsdYXFuX97llYYp6Ni/0O4Jy/863q6a9fsZQOeL+OAyL
US73PQXtql2/THjAfuJezD8HLY5clsqWmbLPOC+an0BIgSNSjTWx9RXPKs2KXYyai1/1na9cdvVv
xU0jrRuAI2b7RfiejmF/qB/YRgUl1b/qjKJdPUGBLBcxCw6aBzygRmFLGhLcC4BZb2AAGrBmkS7g
dQbkaJ//qyZ2AQmHtdNMIz7IJL0hObuO4fZ2s+NXNnD4U8JI4YJFGiF0N3uHJiAiYCSMcXaQQvYi
daDEiR5J59F9/TFtoOwjjTiU2E8aQhko4vng5gESK3/btN+ke92idD/6uKr/H8N8zdMx+EysDE6u
u+Fkqy1NTXJTehu7oIiO2NcabULa4Qmse5dlVnNeRUbDp20YXeS8IrXMmEUsI7e3PeQJ2WbIBGit
De/8pzqbyobdWBDmezrONJ/5qvR4YBLxr3aFhdELEsR4rpyR7TRcyRR3zwcBjnUCmkBNL/REftLW
08Ar380dm9byH9xOHc+Y3qm0Dx+a8XY6LdqCC0ONOGOjI9g/SxFEHXHbLy8WGyLrk8DF8B91OrjB
rM1tRVMJmn/h66QEv6y9F41IucOvh/HA/yLh1Ta1Bx06V7OUdSL9HmG5x6Qobfkv6RUBT+72UE/X
nGN/PovL0xAmEo5mGpDnEO+fkGskZOFaHPQ8NLqKeIVQ1Xh6s5cf2mKslz62pA/rI50GWPiAI1nB
KNvOcLgvgt8bQAplGGQGi+nWRf/OhstX0aPnD549OwW4+xpxpUW9opmGjoF0m+qjKxKTshFv0Y1c
66DB/HvTXMyHoJ5YgKbQoF1U+LJ8vW7ib0ZJJomtacuigFIQRi75RV88v1Ncy9IwGbFFVK7RMfYG
ynjZkm99dRdRLoNVK8n1oO8hYLCGIseMEizzjfbXooCC34ExqfXSfp4yiP1yiEhTG7vnMip+pLJn
o0d1dlrjk1EUBu9SFPSxoDSHJxP0C/brr4pHa56aSE6qQcH+H+PA7btx4O1067eH7I3CM90Fkwbv
kx1czToGQNwcc8SGgdUURigehTVoB81qDwgoeY/KMenH5L4TA6PqmbpbS/Zn98EPRw5CkZ+YVhpD
PTsASWmYQkOaDMoU7IZ/4v89MQKdfosrCbE9GY/vlLR915Ckt5hIfi08wKH1pVM7Hf6ZWAQLaAih
cKPB6oJLgslZW3flt1sLAEkKg2ibLfgXpNyoUoANwVPqCI4CVbjJKr7q2sFtlP0DlYphAviAvA1t
7nQ2MJ1lcWpLz9RvsDhRZP+8l27LKwvXARbFT75V8TBL0PPanjeyySaqJvFN4wWdHgF64s10OsuA
+01U9EzdPRzQys6Wa9ahy8IzQo0yEFDbAZ8R5xD/6bkfD3dn6IuiwZUTd4U4cYsvAsAT9du2gEGI
yygFwwBRedZG1n7h4Kfb4j3K9uwBJS+lPTJLj/aqHIfwarnUqUneM7BIQ/HSmBPg4BiR3p6pp3+t
o1DoOLi4wIP4+lc5LfvP1PrDlpNWm0/52X75ue/aOrbzr3NCRJ0l64+dj53BMotBs9TYKiZebLRA
f1G9SpWGwqOVMDRayEE+O51uyspiyr09J6saZt3ndocEkjqGRPMOgq5RkQrMmF3ky+59B4yQbIVF
sYefZrZe7G5mPdMUfqqhJQgtGHaW9/eBcrMVfzb+Y+Cfd7VBaDbbu9HOIBhMl51M9f43N//olMO5
kUOdsSPWLgofMFWzRcV1uiBmbdc1GjRyycMgXIL/NuEKbCMzTySS5ZBPdNZuSDUAx62KK/470USS
GxKu9fwIMTB3mTNGXWmISZW0PGrwxMgf/HjYlu5xrnqoUVishKPsxneRkiwStd3v45jj9MtNSsFD
fmRPXDtwbHEVPqcQh9zx0lUC23V6MNm8wpar+SbZ1plNTKUQhTgOosPGldEsUfqx7H7NShSPG1Di
yhw5agpY78O93VqmWVsGXNkF1tIumorCdUgiy35fPV7EKpBPoDFVEF/B1lkWjvkY2Jfuc3ipN1Oa
TpdSfoeL7KmLwc0sTUlZy3PvQIbktx6Tz6kHOSGw0m3TJc1qjM8b7OOluHx0llSlv3t7/ObQg0VF
ilFxJ9+fnyLBIqpHLLNc4f0ckNjB+iubb3GnpbwVT3SU8HgahX9IdfC4ldQW/ysDqNP0r8bz4dpJ
Mt1B4SnXdTN73ceRdYt8yJrMHDFI3+lOS6mjZh0ygCJP5V4zwl72O/W85QrWbp1OIkGNmxN3VB5u
1XIyPouKoHxA7IqiB93Axsil72xuqxgsICchwkXeSTt2qNSWtyagnyq0rMAk6iq/7NyO5e3cROoo
Osve1ApHr522goQl3kfYU6dZfXkOB/lW1XfHtwiIW7CL/2xCfAMm+LbddkdliwsnbfEvlGFN9nEO
taQ374cp/WTPQsaCBFPqFVHrb8xrlsxYQ18tD8oX29lpPmten7MyE0vmjYyV+ADyw/6VCGZrovaf
imbXYj7t/qTXHijaIk4AFjBd4+xmzfuhWyjeLhrtzytGZRredN1eGwQMkvDpOaFj0vOw99dkoHmr
QqW+wz66eRrEdDFHMbonoCpj/FD+KP82WVTHXjEWLazf3nZSGFsnPXslm7ySYQ76U6HzBhEOa5KM
g+KLQ7Ng+2zlaYww25/dSfIedzZ/L4MPVKBZ13oe7VtfXD9+WbcG++HCPB9giUaI4cMvg+fYJfEd
Ac6JRqzTNNlKZFs9oWrmZpiqvMPStUxUdtUtBPuSdIUXZLWtHsla46vw6G/VzMAmNge4+8G7kKwo
9k3NBMEfbLR6/5or3hFQYSH/5pzXyV481r3VT77zExk/bGCGQJnwWIddxMUvQ5oU9MtgqKulIP9E
tDrCbNuG4OqvgZ6Ki5rVLj6IXk0MQDtQkxRtLbQwrGuPoEqpSQAHPM8ka8IsXDHX/g8nzLWLWn/9
rNvh2a9eXoq/RQ0hU4EV0AMp9LZssIxt+bTAwbZLO00yMzsD17RTdcnTbO56IJEZSV7sVnM9IiEB
SDX1+4G8Ne81HRPCbv5khImWrmucOgyf057x4vcGf9SKhTpDDVh+/BwaeukWmSiWThf/EhRX2TUJ
Jy7ml/ZX8VkzDIC5KlWJuqW+pIH5iQVf3SXJuiNOHQtVTKj+5xxP9Zs9yzR0ZjAkCmvHdqcz0Gsd
xLkW+RINiE4FPJQIVknt9psvkyXRywKjjf4mGi3CiMk/mc4e/ZTNetLk1VwBekQXOVz1QHYwHozV
z6jzni9S2yGd53dOKXwPTcEFwMS1R7T5XiTZNiHymM6SQAYIX0+3Zv/AbtGt1PXrOSBOJKHpOVvI
f0WI8EiRrmIKvagsWdswvNbLG0UzgXPQGG7Wa+ezB6n1HMyND3Pl7ux+HL0sl5Zv2S8xu0gLueg3
iPnl3ZuH0+hmrO/jd+9RNrQSphuy4+oregKguE6a4M8r1j3X/mw9Gzuo/WAwnQJCWzydgEByeJOr
MOw90akmTsWhRdGqjGSeSRq/dhRTDUoIzn++5C7mqCD/BzLFGfUUvo5HHLeoyOPN03u/mFsjhbeM
crgvxo7FWIvDLnH90fMJPcSrfQR+IJOR20PnS2ExF2tW7My47tD5yxGxXuGVorJHN+D0t8KSSQXD
7mB3QqRE6fm1Kqvu+gZeIJzfeAXe/UdbVnuZwtinCWrNIXOilokgcjCsibvdGEq3bd1hVObWsmy9
tiiWnCIBMdDjByIrzQtOM9pHHy6SuqrZEVDNrrytZ0qbzvgIVVUNUMh4vGdxtejvUlvL49smxoRY
R6MMjOQCyTRLZVFgAl1PcBphXQuMlicPI/naiRmtfniMMA5Pp7yryTrHN9SCevpsPWi5REpSFUjl
A5XhtHfjMG8TZkwhYdXlwryh6tNp0Lc5Rs/iLFYVZlk+UayRkkeWwM7AfW+ggJl36pvB+OgIZrig
NDBEBGGNpI5xW/elVkO2dZropYKqS6Rug0btk/aL39E/FEHYbhRR1LjV1CbowvdaJIo5lxJniiuw
6JEFaWiS3B7dkSrJPEpfP0vtmLVNXxD8+qQdyBmWQtX/n5Aw7mGJ0ip5aQrhveoKXBUnYfVBgKuP
Qdv8/5/9jwtpptgUCA5BVr+b2+B/ZgPTb7YhvXzNQvt3hrddSMzSsLBN4CB5eUh2SdVXbfE6SE7g
RLKmuiRH3Ws07YXDEgrkaOtuDj5TYCPoyH3GRHevXI5vTYW8eU4S7XDcRpff57Wjo9UTBC8NWULp
VlK64sVs8hWvqESxi267qT1YXHBHctgAUut/INTBk1uEp0wco7k3MFjzJxsdaw9p7FMylggVebQs
wgUgWg7bZPQQtpI0Ksc+wXeyx5nPo/EwQK9KDCdMaxs13wT0FBANI5LL6QdrPm0KdRwGR7TOEyfB
AqUyXGO8/lWv7H+SO9dj3arMxDY8T5QbYwFxGDB62335EhH6cTqMd4Pk+EstSIse0hf9C3YbecJV
IeExdJ2QshhnSJNvFBgw94fyHtkCcLMx+EdWp84gdtiWzBYonpo7iU8vb90WtEwPDSXuhX3jZif7
RpOVZsPR0Sel91CpJXdrzZ/fxv/5Ov0XUxqhRGRxIqLNSMneEoFqzJqUhK7KueTti6jjpYp9Okvu
ckOFL1Iqa6bDBApdgVtYy93pylpclctvHKEaioHAtVoaz+YYV57libGVh+4tXUFh48E4xui/qDR5
3blE9zKL1Pfby0pTSoArGS1E9g1PxC8E+DBSMognzyfs5uru2kVsiETg22GlkRnRXW78g+8C3gNl
ZuTExCRy2pHeY4y4NE1MtDe9oB0pet+i/t1V0kT/OLAY4BGNIqXlVYgSJEmeLYJj4jH06zd+sy4v
ykduO/SbbvmINejcwfVCFHjJKyZ41BwpdX79UjVJZ8LQmEy6XdexnxrwnB2j1yYW27pOOmT4w1Jx
a3K9EGaftxC3z4ynKavrOCOi+M+88dv78qkRIpBGLc8XZqt40DE3eMnmyNCXO+teaSkykweJqSla
u3VL9t9th8J4BH4J6vlZdsKw9W5uV9pvT7jzfrSZV6dqtBeq72tu/IYYxiP+XxVRS/1h9/UYrlz7
ysQnMZq11cY4S/iM1m+geEEIpO/l/Bg5TxV4OfwWsbl0tYshxEYJ9hCazyyEJx30PdyZLh7J1cZB
RPT3D6V+oXZMr43YzkH8vc2mIdYaCo2XOx2ctFioRGcFG91SFpjUhbsZO9clhBKOJn2epKr7NWLn
dOkemOXAeAkQGilAN9UZ5OZ9cDjWBJrvlGKBFX9S/XQea9ymOxhsTuAUo4OKk43cG+OGhQJ/xWv5
USWWDdYTGH5OdBxYRz5Q8yepUmQXqfWfJPUBtzlEHecjNFGEdDSW0YmrcVqBMn/0tvABwLt91IkN
+Z/YayPNkpmLRjzWD/UQ6k2fkkLBt+4kSoWfuKHAERreGLznTD40u2qvBVNsyY5BHBJQfBRBq3iX
P888tV71nSUcGa2BgtBqAMqZHPXLsxPTqyQNdaBJ5XoBQ7Nn26BtARZMU4VXQz3jVY2aHs2WSZ6a
euHdbCx6nc1fZ/SM+LsybnH9nQkE8DIpOvh5EL9oDHQERaSZvoTqIDspvVwq47NQOqFGqa8Qg5oq
5QdSpDjxy2hZka3d+Mp85Ofbe/bwathHvE8zMJCS9YctzhgoN0SXZq2VCxcUixw8dRv5BbZd16gE
WdAJpXRaHLH0CSnaYq3PGOJp4azJmNq8oOAGzjiXwnAS0h3qJt5yypZfePfbjkX1vAtBuNanZXdx
u5FmGriZ2lgNGvHDlmHHwLREExHT5n926rcnWlE/TP5DdxFX72rg9J+tvZgEPRFqSt3HN4pwih2P
sr3uFLrclo3M9Mk4TdEptMSPYqUKqMAsyBakYWS3z0HIFNwVdb83cf/7fegnlhjB1Zhp0Kx9vfLi
8MIldOD6XpVDxx783LUrBUTgdedvqsm6z2C+CXI9SLqLwcBI438yGV8m1Cqb/5uCi6vpwLERzzsr
+LNCFwWTAoynN1DMEv6cTNLKK9ZiX/3MVNc1YT5knWOjWzZ+2CrXhPC1Zov16nHYupbrXmWqMDyO
Y+1XsDczkgatX1YkJuB6sRV0hOKMfXE03O6OYbl1dWU3RkSpuMJBlO4GYOqVA1o/ZdjsmD8Dy+h/
kvPsvqTSbpXjfoP+MUV11hw6ZAeMO+ebZ0KHwP2Q/Gq/9VI6RgNxCLGCJ1V0NHC6YwwkBklirDcv
roE3XqR16vjVf7hIOJKDMLrTzIT5wi9lGEySP1mPfHvy1xwTRhGJnndryiZAk3jiUq0pRzgv0i09
K2ngeLATpHT3s5noZLDrJBM0tecTnf/XOv29N3hkq5ByFdzewqinubSOvAlVFmqFSeavbXpHRieA
49PWPMIGbJgfRgujP2ibKunQ7Odtw+En4IRHhmGEnqnwhLnW/iSUxHJp6H8qcHDkmlOX2Q+n9jjg
CaXRKNtC+Y5vQpz6m3ohFaC8rwiYPwmHnigwcdsn6boEX+pxFfErLIjAIMCRFSdR3HbPtAbJ8u33
+joAvTjC2ie5D96jS0RePh/ACEVDciowtEJzNMp1PJb0LOfF76pdrEhBiqJPatrRFloCKnI/FHxf
icZYtqz3ze2RADk9uR2q0l5t7+qen+3FzHOfCxI2FoJA4iQV1Tv45rrsDgGFz2bA2ZsS8QquTjIj
ZTR7/kne7Xc9LpqOck9aGIeSdUFjCKW8inxe0vLBpvdMAapHfDozyQxZ8Jo9crQNHHFpm30a+Xz5
vYsIWaSrjqNE6ByO5liH90h1N2RvLwbKHM1Def1VMT7HOTWWB1pQBO03nsZ+fb3gRi0rBYdzYULu
AH2bNyKWSA/zpZtL5uUEOn+qkc3gCzO/pblQTwnb20ztxS+f9fUi9jw7BXCsUtKzFpbi/S+J++uZ
VYCord5c0U1kCThaci8Xp/a71Zefn60JspaGDO2bnejey3qxx62uq1hbaR0nb7TcWG3FTfZyFPg+
L9voxAcbm22KtFP4v42CSpjIk70mW0R2+p87bQBTlm2GSG+iM4cHEBPWBroJ2ZaslwoSlabf8bwN
x/y25rIq6TO3GMR/awpZahcmzMxkccgCSwK7NozO1sCoU2s1kFjgw0kr4zWVO12FG0DAqnppK4w2
4rRe+hNkHpaxAscVlaqAy/inyn5iIbKJUMCbasI8+AYOuRZTOIjhSKsCxoWPHsu4d4uuhnGPoAtH
boR3qqQkiBMTTWcqqjZD3KidJdk3jD5t2HmCfMhegU4fRESTnL5KrVzuhmHrqPTaqm0h/Vf/hTJN
/QwhsHa1f8fMd7135FJOsskB0V1+YV5sQOfJEE6OGK8jePKtBiU9LNGwH3jUDdmvtAzmaAVtu//x
x4Wdb9q/qEZbn3YrwyhYArDdxAHBhrk4yvGZTks+cEJFw4DGILNmQhIaUO+7ORx3VRK68mh13Ug2
STMHGrHAT0ijdkOzWRRZTInDeh+Rt3OiN9rYGa9+7If+R58eoonSdx20zYqs/S0wzbJMY7ZLWxbo
EeT+0kwgfMxIqNF4eSNpggL9qO95Ddxm8itLiVMtqqUo3DXYBEHLEV70kz3xp/RgdcJFBs84akxQ
fRIsAv3NI0gCYPJAxvJFCehBYp1UvZwWsmb7Qhv2HHxcH522LRaMvfsl1ZFWS2lKMqkhgr+ff01K
CuegEqZkx4pyLsf5KhqSwU9bwARSBQE0WDSbZThxVVFDEuUT18gaAsevQg6etarJbOZJ7bTmXxEl
n5n5gPkrg8gdxba0opZFNhXRtGBepMyhGEI9NOkWVYX37ay58kjO0MEdZyp6xatB1zpM9xPSkX6Q
mwq4fWd9kXHN2r7j29RKFF2B3WGB5YRAtPYsuhzgOuDVwbECgeybQDz9gzQXidJI33KQlKxW/H1y
vyumoLFemCX/AajdNDhqaAUSujwocJ/hlYKmEIzkgyeN3Kb3Z0pWW/GY99l9ZxEJZMFdtf0pXNsY
ywy31NcC64pX+Xc41nUwqqcb15liPq7TL/w5iEdY870UZNKq+oMjBHduKTHlAcGtwMtG5DzQ2qey
V+yeV0i7u677qK6wIaX8zhkOpdDDqPC/U++B53nxmtFpxHtmlrvv+Rwmavr5QmTv/yt9jVzwDDyD
mwc3707ExUKuPQpQ1kmgOxpuI5wGXTKSf9d9O9HI1DBGaFUTE5N2n1SE3RBzknD/9G/LC6A6HtPi
gPrvkubkvLrrPy9fIq54xDIo73GvbqTIvmb/ecZupbsGkXu+djMqL99C6Cp08+evoQchI3W9oAkY
Mq4xyIOHdvNDpkitF5yCdOeaemMz0SIguVaevAZvKAitd6dL4abqF4HdrTKk7loIixo0oRp3juWV
Ex82Nsa3+XlBG5we3Xb5FNfZLtOTrJnjD6pF4GJv4o1FdfXevy8s8AMYpIooZhT0DOWVqxBHO9z5
PZuQAnaD9Hx8xBrjjI4RnVORl/sQgbWbrtvFdj7S2DwxJCMj4PlaRvDlwzn60kK+DorekxABoP+F
hMLEOslgEW7mrGq2TLQaPfBp2qGZEnwqW2aMTwnbsl7rsLzeiV/hVnF1MlOTK2AiqUn+9lsLMzVx
dieCSNbx1ZMjcP3ZYcXHe8UnRRcCtZt1pxJfBw5vpKsZ7AJl6KSqp6PFFGVmZwHoSTSWx6lOt+/x
6PixhXH8XV9gtqLu7tpYMmHEhTuG/1cIJ1Yv+fS6GrX/3hqv/4uEACcwMpCgB8p+6eOOMU/UBDWu
t0GuwGDwRHK6RRek5l/kbLuJS0I9EX+JEAT99j4CeD4edgJcCf7fwpOqnRmDmEEJzf66JtmYEFgl
Lvucw2B9N6sqMBMx4Hndjs+LmzxMeChi31QWBxQRXG301RzPbe71tHM/0A6YKltzVNmFoEGlVfIn
O/TC2oaPYhxkd+t42K8s/U8nG5qEzp5t8sseSC/4sr6JUcyR2UoIDdeD5NhqyPtTlM9M2gn3yTVe
ZKoIil7uAhYdMsmWTiQaGb7hcjVM1ieDRUwLQwLq4nsnXfsbwqCAxtQxTueoFrHWxGjuCYhIxYV6
31e/47cTbsNbFXP8OtR3rNkOphlQ5QIZEZ2lmIZcXINrVlXAeJzYaAPQhRPOajj7OupblREl3GkT
g4LKEzBH0f7wzy+JfkQqc/aNWRoumCqCISKcC7pf846sKH1VB0SOACOAPmi44a5HlQ11vanGP0OU
z+FJIY13YE9md1fjQXw4hoZgh7hH7E0n/71R7tmYxW/85cw2AUDL7lsA7nq7tV9UR7dayEc5dcIf
DrX6K48o9a5QsJmv/DpGv4BiC32+SqGmY0VF8C0BQuETqlnStE4H7A/D7N8mk6s/YoRElPzyUb9M
+gO102kJUk5CRvRKhYmxXKi17zxMK+P0CJlzJtycDlZQgfjo9kfJn8Zr+vHuyS6Ww3VENzOcacZd
d+qGvgMxyX+Irh3fIlnoK3/lb3U6LfcphCxrrW0O7+glQfvECQ2VMeLap4lItYICu3oRzURQP3Ry
r/+c/p30OsZqHKdg9e7DrgigAzoufj1ZDPwTwOCyQBgYk25SnLIAzXzKbvH7B3JBvwD/c4eT3K8o
6LWaVvFCu45etaHgLDtGCMIUbknq0QYt71KTymNeR2en+CFz1k5rIU18+sRicMmqCm8dq055UFNm
hoPx4ZOZtFqu5YCEYAXVJQPhiH0YhVVVh+V+md1wo7tbs2+aJkpwWqu549LRLpZIuvrCB7TeNwpb
z5P3QsbPWGmgjgjnW/bCKm7L20swvvrrLR4XWFLhq7dKh/aajaZIzVb2smkVPkEbcCHRVmK4f/dU
S8YmWZoqlR0xwNkCGSBVRfpn3rdXvdXk50sLooJ3NcoOwAsbaOBOh0G2k8QJtSzfMXoYGe8Olo/6
ic2Y3AJ/g6iiXB8laE6wiGXVnrC5zeODND2Dgq8z1ROucNQbHeAYDDqNu8ItJQ9bkKvqTFqiIfOI
hd591Kir1ekwxFWeziKmNr6N5S7SC4J8dcblfm7vorVJtEvc0t78NmbOozN27wOOPOKFsi9rDRVo
dQ5n9na90OT3mxONnGiQZJhXFLg1FsDvAlljL1W74spwFmCUTul39JDAe2lIKRDbCyfl8crGxuP/
MKu4HT/Dobd6num74Bienp1tiWoTWpKYDXKFR+ckz9cfNHJi5qvdSlb1JjXAVuYk53VHS1yjncGS
qbQFrl3zg0BE3QypYIwQlMzb8cefmDCEll+3cKPUYNNhxH0PEEghm40unMW5h7kyBk4fu8xkbdLR
8APmOf77yyb0UhjIWPRAr19wxPa9UvydmigE7phqLeQxLPZfQvYa6M1B+lwTaTjT7YGXdu844A0R
wUEeV2VvkZoB+/bk7ydQE60PpjNfkLNlQ4WlwxVb8WM/AA9wm3Friqiifa6HEjcT8IQZ7CnEFq4f
2tEFKcP/MOR33McdsB4p3iATvvXvJIQB+zHsk0t7WdlEY8YDHZJYZa9oim/bXRZ99smNneOK9P9R
aQhesStT7yPkX7/7x1hVxa83w4OsVPNoYKGUsH4SKlWyDD9d3V8ISfYt57FfC6Mj/dAxAL3DJFEU
bRgLZygrjV2Ubpa9q41ZlcG+9912AugRd9HlGAdfX9QECEdOKmHw/Cur9RNhyIlUnK2RmXfnm5Ky
tma62AwHrtLUSDFyTNGs+lxxM1BCtLEMjOAK/BwrfkL/q0Cvrh8jASRR23p1Xs37GvKZV0ia3HRE
A3C+TocEvfERlIpm+z5NWGQYCi369ZSAgQ+RTEhryG7CR0UQKtGA2AxFv0TWJ85kiom4U8Jnvx/F
yPqzatAIDcyCVgwhvudjuLA2I4Iy6LkX1jDhla40FcqNWOVcTYn6/f1jIaBEG0wH9Cp/zeVJe08o
ro3p9yEGcyO5pOC3pxeb5Uo1ikG6B6DtIKVfUvQlWNQs2diIurPUUbcAAZ4v8fi1kDJAgkAjrXl3
gAuNRWNztiUdk3PM0HLQctz7cxnRQAz/qYfZdo9x4/BkRP5QJEHuJjCWrVWkCfUUZSZ5UVTeSqtK
dUUYzloiWNe/RZGmY/6jtyxRlTnsxSSFo6gAM13599fBsSOGI34OqEo7shKVSCI6HOQ/BHgZxDp7
8U7UXCe6c8ea8W4iOMBmNTc+z776ikwv+y0B8/9N5bXs8omZKkSV6fAz/D4Wgi4+waCuaew0esZZ
B7YUxeKzMYuUVbpD7qrUk2maYaeMxYMYevWXyn281EnMUSbgb1VANQUaFowtHU16rTJJs13IOdCL
AS1PEuWgtFexQhkKnLf6LDa9FmzmnT401Ff7z2eAF9N74YjsrWg1rtxH7JQO19csTJN85xgW3ulp
dUPf0dO1auM5dfL0xIL0Itq6TFbC4SoP/bsi/0tZXAm59nihr0dwxw6CJFDTyGOcGpPaeCdjhuFv
K9DHWnq1nkF093QJO0y1MyKnwTBPtic5v1OswLIS8Ez51Cl8345gFbFq3nQ78bvgp/5PuaJgOlhy
v7kwDahMewJTH7Q4jgoQkuI8oQ+7uS3lrMrfH9+afcChdNbLUaJ1khykE5/bRSsI/OQBE1tItzqD
9i6s6sg4+Capj94GcyAdb+/4wb2crw1Xi4315k75Bt2QixTfKEjMR8BYhrezRPwflaae9aYlSQgY
lP6p5rsQB04NmZ9Zs3AUKYWBjBBVbdSSkbvklpv3NrV4p9OyIPf5E9siZ2OquCytk0EcC0vT+iWr
02HqV2fYvoTKV9TPu4hruXTrmqlTYv6/s7CO6OoADr0p0lbwPYf62aKOXIIpyf2FfCIonxWmqg0H
Jrm83iBfAv7+4sO77ICOw4kfN+iewL8iT9HuTy2GSSTHDEREbmQoSsNhNu538xxVB37y5TxStvnD
XcvmfxGFpSoh33ll3U55c/myNB7aZ2W+/cbQ2Gw8p5AA8ZkktAB7XVP0SMUqwF7wm6kemoNc9cZ0
im1ckmFvkK1DmyzkYx/VBRjxawc81/+XyV9/l5CkXXO8IrI8ijb5i5YtncuxHz6p/VLJB6phZu0l
3HtunaJOAzdFJra3svBuHjaNsGrWGikHj5z6R/piir86ubFBtBiLjDYsQeQUoxbYJGoo8gjdgrl7
ASfpwQlxlWoWTgyiSqNgDscfOcYQ/DzSxWjOQkQpR+OeWIonQ0MzT/1Q7DJVb49Ai7YR9N2cplqe
a0agP7exxJ0B6Jp17C2iq7JhgXeGmDBLBFcuYzujp5NJegdgopzcrOkAXZV1lCp3QlWEDc5JydQQ
zgKQabJGp91zQlD1HJm9Ca3sPj3lzI+Fjd5xcXBYvy5yLjx4AnoftfzuUK7PuDg18YlMDzNjdzhr
B6TBQJPUwRBNdqJjqAevqAsqzwUkwlZR5BL1XGtuNv9cMFYb7UiNPekXzuO8FzrK23FKUtyblpFG
cmP6AlBioxypMSjc43IAnE9or8D4tGyk0ctVNMZAIbBeC5ZVUXHxchjYdDgvzozjj5k3N+Nk2hgX
+SxUTRTmYs1Ap5TKN2jXxGBpzWxu995/LMsYFzDAtmr/RchyiZv1mwTK8AwdzErGwdw5vBTCiRde
wtfmWBySbKHWN4Jknl43d8VTHrJZ7biGuObhPLA0oST+hpNmJ+telXXZP/cWAdhlQzyPP1BV9DSH
dIRhSic61D/wDXCBUoKj1BW3rCP8vzFPuS4j0zqeYQCbMRZ1sZL/YOkkZtMxYicpMq+OscJvIO16
juKUKce8HiFHSLWgjf+MX3Iqpuv//f+StuC5flbPq5EghuIyiflr212bdjz4MuLlwsaSmouvfYdQ
USahM1zeMjnZyVpkPO8oXObIzia/iAu1R4DfMZ6QsCJHpfUF4ojcbv42LdoIY878tOn3naWsfQjX
A33IAjCshPII4yiGOpaMPfUJWgPLibs3aBUOgVJoLm5ecFs9UoHqJEFnBbsaf3EE738oqbV+svKd
8slTNowDbre25KiTknI2C6TBRHdODqAjDcOn+5RbVWivDwgdxtfRxqZKmoU4kXsd7Icr/bLEFU3U
msX12BMh/ykkBO3Kd23Rdeu4Q9kXxHEEYc3ktb61d+gPxWeZpb9urKEVavHJ5U/MuBzd59Pn2sIL
iPK505avgo16QFHTDk7+aF3H2r8pSq0TYQel+SjtWrs5IV6F09o8tpotflyGzdKbT176m6v/ykad
PXIE73kHRxx8kEVxJ+02GCHbQprgKFCuyGGF3LWoFUcRA3biJkuzvY4eC1LB8S9ICTTgaCg9Bkxw
rToKtPEaekMcPvJAmqs2CdDQ89XQ8mGfw3ECwNp89Vz2t8i6W8HE/lqKhn7MA6Ft6AX3Q3KlP2p0
oBRjCPx2dswmLjk/0q5DPwIRy4vHfDnTAUh/0oh7Vjab0/NTsXEiMQtS7jlnvpkbQkuDmVQCBc8A
itU86aMXK4/3hYGuoMMpG/7Zm9BjL3okkUTn4qRWEoMlVZFYmQurcLHWoND+469ot6krHLdGZ+tD
1vA/rQ7B3kxjWr7hmPs5eJlfan8t/9dLPxbmdN75nVd0REVrDQ3j1JFLDC049KhrrQWDMy4MVXuN
lULcGVtx1i5E4t11IaK3AH6z/2STqqK2YIMVo2RKCBWmds0h0RgB5HcNd2mCWReeOqpcKmnu25ss
i7U38m/quZK2bWn/Ru00nFaXVXz4lN/xi1QfVY0iLzqiSrTEL8/uz8uIfdCI7tILr0omm+yP8yGx
FCkVIf/uUpI0axWGBsSU2d76iYHs5KAMfskxQbd5JebFJNBugIVO+JBPQmyFXbOrRVkCgTgWD+9c
nmpICNbb9o0akqUXNYTduu7PxADbl1fqnOjk1DVapxpmT62ULKtKd2yR+/nWbron/jw62kovlrA2
912K4yjAOIOuW/MvubXmpV/5MsqhBBVTHtLRVti7SWAeoMkIy4FfVJs8hphYAO5b2Zc6JN/MJjB2
D1JkNBcOw1bL6jjer2MejzFRxxDb08UQ0AB0p4ha4J9t509KUBpaqjXL5P47xdrDTOYgS7WW7Y/B
MCYOE3qEGlT9ZrcP+Py24fyGWC6YIzZbAzogMwsqKP39LvjHfTvtycKVYqQE06bXBu6xNwkMsRJT
QMvhFepqph2lqEVW18f1i4OOTwJknRbs0Axk0O5pA4Qmsw6J9DrSjedgxRTitt5RfjTk0PmzeG/U
GYFYOQ0KKyrWFuDG83EqHogPq4FAiW5n+ZB4HZ9T3/7HFHTrwglhbvr0qkJkvCKXijkL+lpql5L4
3hccE/+qMLp0QzqpW0KfJ4dWWdQfFUu2tSPJZgd3uMJJWDHUNBG9LiKpTxmgaEzk3wpFzLjzZnVa
/elxgfxgWEwwhyehGObR9ND4gcgRwB322qLI7UMRRpEvXNfo8w6EQUW+Y7+WQzOfElvMTNvuR139
3Lw7N9BWjfxz6Nx/cmhBDf5qaDnJlbqVeiIna7gWB8gbOLEKiVt77b1OC06gnRlFUKKUQqWpb8dy
d3Uq+cwYyIbfimp3Svxz5Y1gmLnjAWk/Ld592YQj3uDV/lbX6AT+oDzNGOuwHSRMnkVXj+NEDQC3
9BJDvjn+82SFIfcJZ2PrQyECoWXXIJqhHbHBoRQJp1LQRfwXW0TNJOugukhwX7YsEge2ICefTwt+
tzY8On3MGYQw/1IUp5i3oW7HUmQy2ZeK2BAfxrYFY63k9Hxl2uE8AtjgfxzswlZxG5u20YpTSQmm
tsHL0FoLxQ2IUnq1SHh2w0hU5ajGYAzgOpWssAFNaBKdlja9WRXjEUsKmAqJx8Go9o3I8sFN0tTg
J+yONnqeE4hq6lFJFT6Qxje63FwIMVYp4EnTvaD/AlCTG5yzBvDb6OyZ2Ia1e36MbSYYmYSEfXu9
NzITwTUK2uSm6Qa2hk9DyseJ7niLOB3SASKVQrc7EX/t5cwSlQGhyYuewULuVFVJl4jKKyIg6D28
aSkPz7YPX4i4XFiLzfG4XtqhNaPp7DQei0pfTX2EgCBQZge6QssUEmJlzySVFhN6ZZfc06J/1T3H
hCwZKSINyBDFCXQvFPe2F7Uddovi3dRmC0WNYv2AHx8AByT81Y1BURnyxR8i7Vgw2dlU8hRYGl8B
y007IXWQcDm+yARtYd4g6C4SlGl37k890XifNK6swiN75eCME081DrIUlteSsSOosIRpCBmhBucI
+v3NF3cOomtAVnbRi/ED3qMw6j3t/F5WYXLeQ5LU8vyGk3FaB7Irfty0pWGb3njYT7FuHKa851Af
amkAzFyxfaOVP/VFf85RoxwGQh/pBFA5pMRFNQDqBZW4Y+At06uKDYlFCFYkhRgfQtfox4RpjYo8
H43kheo4qZcUu6n8ui2XHzEP5taMCqIHcFQ4UMwpDMdx6JyFCTlNyAL1M+UOJ9OwFTdAs0WFtQl8
3X3y/uUMCC6Jak3unpm8WRvRsRcQBA3Kmxx6LwLmR6/GPoy6bFO4WDcfHD/bFXEpbla3Sfblgnpw
V0he5sclHTy5r8AQWvky6rN157yKMGkGmtIUsAFE0Dp9wD5bbQczMvXApK5XcDxKJClAIc2HgNSI
ExbvhjMyunSahZtxXThHJ69we9os522wVFmomb4bz669eGgPPwErMEHWWVSUj1Krk7Aud14QkIR8
86uGba+xxOW+P7K2ae/GiKqRyQOVQaTwvqU8PBeHq8BRrxmN3WYLpVr9b+BMXxvMU1ZG+ywJdcQY
SXGkT+jTZdNuDQnEcj0WI9WmpQ9C2EawV4EvnbwqAGxWJ6a2JYD88pTN7UyYvN82LR3tlEqo3e8q
c6rGaX6GyXDYhvas7ub/W+PXKnBfG3hZaCAGEo2ir4wEokIyyy5GJ4jZArpbbupQ8qUh6b39moGN
X2LHsZD4dK50T+lW3dLwO7uaLbOuKD+YJz0IU7PNhyVHE2ogZAap45cT+2bv/lPdd3/MXQhlf7T3
r1fxWfuUxHSaGB7zWOhM8rv7balm7AL1c4jabUm80uSdnT0RYl1OuEuf//ebAN1e8i4SyrF4xiCQ
m/miIuxRhVP+ezfRiHuK4nfyv1bZ1HMbrPzd/9DZEJglFK7uWPnoHCKJODT4CPUpqQV7zKsgdw7B
jOefvlQOr2osC8ZN04zs8py6/b1gkKGJQirBjCP/VNBeP/X39uryHScuFY5HoisA4HP074lV5hLC
ULkDsphhJGlqCUFg4QSUIgTye1leUZ6MgkxYyZ450akS9oDcqO6PheRWIMxRlxDQEJrZkuT+kKTj
U2fv5hiEgbx1C3d9z6DV5D6Q28lTNYu1avbP+5mkM2vvAJpBYEp1bWEbIKqdn+YzsdPXCQDN/jEv
8nVaG/UKeRxqLK0u6fJ0+Y6pbnECY7p4L5gIS/TZl2gHGz/zQcZDHBiPlQ5kVgeP0hMvLX7gIukK
rbBWrGJoMSy1TvCSKqLgua6KFOX1DDYpneubmQtgydqsc1oj0AR/kvBCa90332KTHvwC/XwIqGjO
euItVzOIJKgSLDAV4OMxZp4ctlntnEOFai4pxwILekIj+0qOa7hwbLqnyfUwUtfeoxwKNeCJSjYv
Z5zy9ojdiIcCZNB53cgJeb+AhC4/6Nb4DOFF1vT35d6fIKBBePAqdQg++aTPsN47g1bJewnPjZD7
FMoi9OGpaqHrRbTyL2DXprA3twTkbbz4ZEsfAxvhRsYWGsd2ldPtU6Sz6bmEKQtohHQeZUyia74r
54R6QbW7yZNEK/XpDnSyRWcttlgILqf+aQig8/qp8w1PbaQdnqXQhpfT7CAAGCt4guQhaaRt5BbX
/RBOgukbrQaBWkv2kTCK97gHyolmVDDjn5hJXlPGhygwoIlRzYxCb1UuFS1c8totgHdKgO9AOfbX
l48kpj61oJNloRbmLLUf+TZfr83IceEdhM7VxKQ6gtoh0/7MUjE6mI7gDgX+WVfUQlYKusSk969s
tOgCT9ypBwmr1TNIpucSdA65r2RvRVGunPx465vk09CsHEqmWVFKQHcW32ZYBsG7kRC8ng+4zqEd
rueRfUz00Q25K+107F+5vn03scpkjsEkqIy9DjwF+/cT34gpNd/f9NMKSG1HA4CuzdUEy75EacQz
crFHfKxXFqAFYBOSMFvMhhEIYWNcms5MvCYAXUHgkRQZnC7RrtXgI3Ao6T6Ife+dAWN1trlMWKSC
S3bZPlsCe4ZBF8HypUhPX5pB44D3mM7adJ09RTtrSeLMy/nyTtjTEncNMLJfBDLMWIfICAnkRGoD
kh+s/OU4DGpit+YrRH77Z21bQ3og3de2vgBtWtqLfOiJsmLy43GpSkBhF1RQUUCxaoc1fT51vNPh
ha5RACZeHmDC0slKgPR3coJ4Mu4E2zgjE5M2krDai3+zewdyQtK4uH01IJHYup5bTorrkHqGoFmz
a+PlAYLYiKmzjwkLhEcsgpZWZLkxz4bvKzBB4MS01wyiS6HmwQYrms4fpturKX4X+eWIPo90wOTI
eqzHFlUd1BMLc37mqXsibe5SyuLUsjwOJtN9Kfg4vZAJFihAfyw3rwDd+1i1kTfPQwbn9GU7PIST
Tb5ZvTCzsPiKL9WvAHPuCLMhbNljhLEuwBHVNKkL8HOBkdtACkx1c00OUQJTTxGZWT25gF2Nia9G
NrcjJIsomXBx4FRl+0cdzBdeReR2KZ+oe5yyy09v30PgymMING6hmIML1+BKUzEVcbSx1SkoiisQ
LKKQEwDhvBqLhH/Ic7i68Nz/FE1JKTxKnToZXfpblg7Yq7yQ4ABaFK8qZGqz+6F1zVHka1Q8E7cc
cJjnpFzjj9H5Yfz/zT6XypEsUmUxxdublrUZuR7gXjgOYBdq034vFj6yNEYO5Own74d1ySWN9D15
YlKw7mHmh1NXPvmPd1UPWznFUGt+yvBuA6Q/Dh0i77cyj2bLRGhYOkjd7BOXGE9de/Tl6FqpmD8M
J0IzB8PokNMn39ThBYxLEdmgkOo98aHBJWjgpnmqEzPcX5EpCw0FRsa16+LUV8913YRFnoGGGX4d
xvBh4xqaWND9uAArbdjV5hgx7VnioaKz+tzpZjrHgJJlk4fH/Kcd+ZJ8lG6XPxUwnV64bEVU04w+
kwbDGtha30Lc649L27MdLGUfprawn2h6EkTfQgaelfZPPbZ/dk/SEDtv8PLfP9E3JWfi/miuouQZ
4swGvcNGQwMQapDBzYrJA6Z58mjIKFq50D1jvKKhoiFJcymOilNM8ZnQ8lwXdIRS8HpxnpoM2vAs
MGVHK3sIef3l0xf/LmPm51VtaJFnYikkCMhuJzxG3QNY+alt6aRtASfnwTYmlLD2JyGp8u45BV5a
X793ZRBDrUmDCZQ7gW7Nqe834K6D98p8lc9jG4/Du6Yvv4o67yi61uQ1LNQex1hxpkT9PdWb2ScK
pPNVSEIghITpZZPJXQRy+UtMYz3Msexn6VovDr4XROOdvepJ4DWYAy/AbSJUn/grJs/ScxrzPu76
6+fzVYDosocoytSuRBXBIiMBLP7PP6hHJqy4k1XhSlWFggz1UcrdAantmrRxI4XDV2V1s6xunrCY
ng8eWMdnXWypCulItL/98jZOMbbdRz1O9asi8Sjs1RYSrGF7DExFjuReaoIql5nluruUbx94nHrZ
47uTVerOFec/TGK/BkyUE73wMj1DpoT5Tqo50buMsthcvijqqpDosHR6iZyadSoY+9DS0QApeDc8
n74GzoFUdCamkocQWs8ruIcwIfBTwpiAWsHUWijO7a7qnDer55iCYeAFSBjG8ErcSBn0I7UCeSBI
nSbh6vumfL9B2PUHkAYKSJoLCRy1FQ0qOC0oUvoa+DFdrLER1kAFwv4fK2UQkfWwmG4t5gAqAV9R
WX2PDIoicx1if9pn/Z+ZJJS/D2rc15NjzZkn2u4RPRnRnZUy64+vKQ5jO1BrZ9bRcb6rBwat1XT/
YL96aF7W5gEA+bvApwaW0nR6dvDIUwLXH/6+2ZdavTNyirqVx1GG6AazNzRWf5Hrh0f/4mZ0MPFh
riZnPysv/xGM4TJ03uAnhyVkL7YIaK7eSBMt/y0ZCj2auqLz1FtWo1co/h5i9iiI8854zWnD9MZl
KPX2X6z2i3LVCuX/tcFZnsWDq1O79laL2kyK81av52jpDej2VYNIdiQ+4M9vLq057ZH6gIiLE/4o
/6GYUqV+ZVNoFRzdAV/nAlKz0bva6Vwiw6s/jrq+0t++YTXCKcom+iCuIwqohqvdTZ31i0xyFkAU
9OpMrd2CH0sUhaeGHonddTejWD8lP11zJQAjO4n/OL49rw8XvWPgiCjW6m256NAj1MHYxRgCzBeL
bDGxxIap50QMqfHipxosM9SvyoNE7SKhqwFiUnpvYocakvAxx9y20WEqFi/i5d6ZpRmO6W/f5Dia
WH9aDZ/pR4ahAG1+D/xPgjJnUqq54TcwpsLRmbHxNjWLT9XsY1EXIUboQXZbMOFTPhzHkPEopzfT
pMVhulx1k7qtwZ+npf0OVkkLSHXPD4QqYok5rKkMVKiO3dbss6yQ1ZVujpsjzOJx70Q9UaBD2ure
qcDP8m3Ma7kwNG9Q9KPXvy7o97hxzEA7W/omyy9TOOaQAj2LtdzCxcmKrT0qsu2xcXuuMf0BasXO
rbDPlD8kUnAS1zGRUROJUBnyBdcpXhPnSICi6SN1dSWg0h4Y02uJrHq7WONg74K0ukGw0c30C/ac
ZHRNmYZgoRzWCLvuHF/T2h4W2XUMkCrB52gImobNCobTy8Lz5xKobTLd6x+DLTgNrxD+FIWxG4Iy
58LAhk5c0TmCsRgd4uPnEFukvyIucLSU10pupRJgenB4x1js1kEcOtFL6DOm821lolOLZkAN0dzp
ywSk30NBDYLkMpINObLsVrHy3wjKjKjjfRawYudoxhS8GOMSfV1PLRbULhuA1eDCAdasqghzg+7b
3JnvdyRI6GfBeFoMBsk98CfjDB4Y7xM99kf0jkhfdEL8nvLMIpdWW01D/PvOnhYZFJSzJDC5VFGK
8oigGeFJ/5dgS2uazCXCBJNbiuKklG63XOU0WzjGBoSUgIDIQwZYNAV/UWbv3i0FwjSz1uGStziY
c3CAkzFpRFffbwQov5bylgvfN8qnaRVKGXu/Pv+uQ1r4WqRbavZhXZPLyhsADkjhG01gSuxvharI
sSEtBfhxRJyMFgZuMlIG22s21HiyKtshLUjV66rwy7NCC10GWOQDHu1WdEIHlrb3c+ybywbn7NK9
bDGFB6KOgGmf43PwyzBnmBHfrCHHT0zBKT4n5bMeAUeUrZU6wzgAmLh/sfa7oYZDjISHUeKZ30Kb
B4D3tqHxhLt/t9cTB6VPDMGi70OJplTzH4P5mqsks8YMSH3CV6J2PDOtMt7UqLt8xtIWhDvZNmpX
8nQPxCh4gWcFkZWk0KXi76mibBcukkzUEJKLjgsXqsKSGzEh6o9YOUG7QmfmOcyoJdMoB2itxiIl
1V5kzd6Hur21ZqVcULiu0StgFqLQbgAENHwSwiryUjJFZQ8R06ygfCWO6lzPtek+i/780v+QWhvO
+IEVEeVDSm434gS6B+KFKo8HVj/NH8GRT2JdSJHJcdLKvp/vN3p7wyPFJ5/Ne/qRkt+uMs4fJUoF
/iv0W7saovvaCemy1utq4T3iCSHTqmQxcIUVJuoqN9Ii341xSacRMd76iy89qFXD9tIdxuEb8pEk
/TnYr15vbRJemnj8dKTWkkfyjvXVEqwSLvVwL+i1dRwdG+4gGl6tJHJCzd5tNc/oN6WQj3ncobg/
FTdazbFFbW7vveJAE52e+LgL0taHOuemV7/AIDr6rPbhNK2MBAOt7SWFUpsHs3LPJ+wNDxoJDkDl
JFtQb4jluIwN6t3iuyhr7ywRfvonKCe2wVuQkyd6SdLb91gJRgd3roTKZB6IirDbOUArxuYf0trB
YWBU9I7ZBRthSf6bTJbeKQ6HEt955MOBwP3EhT4VBVNm8K6SnK9HJS+EXTwAZzNDOAezKx7uFiRG
fvHIjRm7+a7BlG/k6pR9tBB8oVNoUf2GRG3R6KCPQxi6wbjRmFNsI0uZtbP1vohfILJOtJgy2lH5
aQRay+pl4mw5q1lSgw6Ccyv6FcSasG5Ny8qb9nSDOyn2DnTuNQy2ZgOoGSbjlkoxnBOXsBD6aPtc
ZqNVNdy3HXD/vMcg6hle0zf3n9777mOBKJLJcr6XIdgIjO6AmljL3yPTOcfjj5UoixJveHxWT0ux
3l+n40MOu2H8TvyRYKkQCcR07AD9+usmEEO2phRAvV/E659ZhaQwdTDF8sszmF7WKizUj0mncPcP
xqtIkPhxIpiS5HnvqXCy6t8NatBOTGkn6yAXH/YE4LgBXLWyCc5eyZohKPT9eIh8OniEE6TspkSi
qUM0rLfrky7L/0eytbRSuYBNsjUTft9gsTrs0vkXueVpWd35OxgYpO4lNpbcpDph5uqnL35Deayy
QJltXayntP9W36g4GZ7RC7kIbR0MTHOATx9iDOi4kC5s6TCiToDFGcjoeA6zxU7GUS6LA1PEzM5r
UyBMlQLiaREsifUlu/lYnwRW2sGmczzDkBWAjAHVlJ5MdOn93tNUa3kdV4NDXtBARg8L6LukaN8b
QsZsqvn+4ESJyzxep1fN4DoS0ui6tpMdroCYyoj+ASVQQSwiRnYqQEtbEpb3WD3i+m2Z6gPc7Co0
FciTQvJYycgYMoYH3SiIfymg2dFpv+xILGqDKch12fYLOGNwE1zQ81CWTwCvWUXa0RbBHfaERt2z
FEOCPB60f0I6O0UEhcxeKbfDpd2PugurK19hetQYdSCSVzIRFU3QH8IGa1Ql2iYY/lXxbIRN0v3f
FDwQRsXV4ODa9+Y9bXOFg/XygNFHu9fEn8NnBORy/DvyWET3sG/0nj04/bnStxAdhkvgF/Tuy+t3
YfalK8d/mhPcNS61FKfED2gUc1mcQEhPSwTNB4XOshpdscKgiRHUFRN2p5voeesBmzSvk1ApsqbE
lXkEBAUouAueBQB0+NlU6ZBpzBjJFz7XyBudzdTNaBbH6jUOY0xiDnr2eF1otjpdbmh74SMo4W5P
5DBp1SRZ5uQg6ItX4ATPmUstwLW0mqBZbZT4EhsyF6KMvr40PiPOeeROLigxXFK8wLT9FELsPB4k
xQBKS0XW7DAsepdmnG30Rjl3n/3pIDfM7Ci+ay0JXVj2dEMbrNkdrDHM5Q9mE51K67MMTSD56/+v
/bVC4541jNs7z9n50OKF7ElgCVdzU0Rqk0a+Zr6nprNt7a1Rt5RKuxfT5g7oJPLLLSBUyxKgepTC
GJMAiQe05rhANLwY7Ih8b2dvswlIJ+wFx20+N6dvZ+0Vojx4jX6wzStjUuZyqSvgdUz9GkLbr4FJ
Ke2XYeUz9SlO+m1OHdCW936+smGycz7r8nGKC1djhpTLBSDrw2QmI2oKl4FjVJwmgFuJaFKkPJaQ
paYlBWCtjxp37FsOyMpqWtXIvLAyFI/paNJ82eqzMjC12krL3InM23CcmG0OzVMHvm8jLJmR90KM
XaqKXIxnrRVfvsPCEKgNvsDhHlJen/mB56Z5DATw6sc56Dqi6/LimbmGsEs/LMsgFP+egmOdbGuT
p+VEZm5n0fMcw/2ttnhC0Eub7TJ2HpqmePGY3Nm9I14ugTuK24EBPSVlY48uTO5N6XzBz0uqh+3O
FUeq167MeJBZw9TTNmTlnPAniAcbptFMS34G2edW9NfWVpUQss2G43CTrEg0aPj9nlQfno2A24/p
r3oAo8JJwSB1FnQWVLvANHv4bKFWBacxklWUyNXK9aVRJhLe+7rs1n+bXsZhSqEMBr/NlVC9Za2Y
24MM5bFudF9rZCQJOMMQHnHQSReyS6Vmmi5SMLio0a+h/bAXR8ZlE5kI23++zEJg9GwCQe7UoOBV
MqBItDj+QkLcxbGYPkgANgXv8wPkN+sP6sFv+L85TDF6JogQzviVDuvozdiBdqqdnSkQr2pAOtoH
TO8OYu40KdAgOiHeJTI1EFTUMr+Pa/KOvzOxhgoelWkaLF43xtUT4scv96LtCPfSipEUcVxZwBd6
UoPmqhgDmHYRh/sEvpviWJnNjFCcElEVBH5ROcdyqCa/XxUkTqXfcejLcAay8K3MPkHnca6mxygG
MFYmyBQt4ZdAPFcMsvgaMM1uDPgYmkxroonqQpMLwf9emvyojFvSDQGH5S2QP4Lg/mS2Gb1RVumZ
KwTiUdG1l5LYgnb1eIMqvWhhLkI82L452rvL3uGma7YPtUQ9KsZrSNXq76rtWEajZ2t//Nm5SC96
9kpgDelBX2QS6Sqj/Ofx/FFZOlqhwo53xpAtWWI81UhLg4GKTpE2vNy4FrTZyziPlK/IQEunj8d8
n7J712RtU1ctzDaANNbMeyOpKsLUTljINlzkVQ/KYUQWUx7+tj6Rr5ZMKfmSWGvWfRHxOnzsuela
ZN0itG69Tj2HErhAuSNv6tvQ8jq/irCTw7PQUg+eDs4UwUuo8sK98NbDIHZyL5S2vYUvxrikHzXc
nCsCHoDgnW6CkDRERcUEftIasQtSVR8a//VGt235DlzIB0Un+7XxcL71+PaOhssCc6t+ZIZzgxRy
b4NHATn4lBio3AE0OL+r7t9g3rqezgBaoxGtD8t/eHNQV5m/NHLZlKGvhiuAi8WDOw4ZxBiVDlXz
ebkoB2xzRuzHUFSmIfptKDNNTKLB4DTi4aC+oZVyzfleImySnFAnHBkHxZOC4aFwVqFX/xK4HEQR
wpf7YBBzzhYhAc8bzZw3i0gnebcfElhirrBkf6mFxdJBWtbAIMzuMb9AhShthUhdYqoHYruLW3YE
l9lMtup1LHT91Ov5fD7m2IYN05dQ9g8FIvXRTasB1j3Zq8JUxflsVsr3WE+iNlrqtAV+qTSnLtF4
ItFW/djTb+gyGUK4Ti0E4Kn6/0aZftOon5bIS84y6A2+M61amA64e/6tWNrpyGewMoGxaxU2mGAU
5QEpAbU1pitPoEjPqPx1tkpqXmwzMTI99XK3HY2vVBSdDderM8u/DgH/LxokMvDNG4GiFPXc2lis
N/I10LLg7CteAfLTQ5JNyESXwt1ZbN1kaESH4Dngm6i61GC+L1dulzbCIY7WtfXPSTiB/slVjUNw
7ZgLt7u3oDqYnEKl+L3YvM8XQ+DeoiBkFamhgDpV6cAt2+TUK1EC8MrVGBJsUMc1DuTlGQqI21ji
iM2/2KnGYJzrgqPO9lxWObqb0BgcO6VvZGc78wfV1YFeOTe+bm2jYC4MXCV852GOfHgbNVPcyV68
9zJuYZ1Z/nDplB95X9V+3hlcMn7aSsIHAP5ZPO6xVnsI12HlPITt/T7caF/KNp2IIaNvU9r1BeT4
KOYaXO9axNUWscqEMz48ccX5yBQf4CbUrHyUXn6aRNbXGVnn6ZCQQTRP1rXu7jkspB+TO9MVttGC
JkOo11uu7IgeqOM+SiTfNk8ayYUUgSDe3ixuXWVQ8gu2vvT3wgfJSJphDbtGvTkADhpfblp8If3z
onikbL/FGNWcSfE5AryB75bJhRq4f8lw9a5ojuvc4gADUbkbQKxvCkbR5le3c0aj1Mlzobr87wqq
QZPA+RKn72Z7jJS6TJtvSTRRuKrr4ebYTuY1KQPXVdBw9h5Gn9GKlR1VRteggPzpSzOXuFytQllW
itqxiGqk40KspB4bJ8nOIP5nY/fvo8vslltdDW7RyvEJOpyMpKpLIEl92k5HApOLYpCx2InTOxwD
zCx3LWndvIA2MpXurbjVbJlhdnr55eJIJoeExzsJNQjSwhMRxeOTOGacIGtKlGJd1uqOYre92nAO
Cp+Olf1d6ebuc18TxEwRXEjosayyRbQ/GU/xTYL6ZxLc3IDOGzU+vWt8n+dLBPhcWpzFvr8Iaif7
ZqPjc5bcGLkL08uP/yTvnMbN2yJTUgmLgnZ7l71zhn6QFtYmmL2r2mFxuYKjjaJ309F4m4+ezVkk
cmqiF1mze3y4Cjya9SEtLIJXFIBGmjv49c7RhTFZkXlB6s/cXFL7xic0me3PlERqVjVCtJsaOS4Z
fDq41EqlkFlJeo9nUxsVYjWWCj2wyb5hJ5GK3udGUe0RP/X8PurnXN4PKCqF+xH0acVaBrVLyXUA
kAuFirZ9mOk7h6FJytFMuPOvMt3HuyVMpz6J/KyCRwXSN0LLyQrkIL3e6nEYLHm1YNKpNqn5R6Uq
8/gJcNoEka1oE0QS9BXVtepjXJueApTn/Y0Qo2WoOnXS4kjZMXj9WVk1BYIQTbZ2jX7XcIiUojKW
tJfKJc8zH+8B3Kl7bxYY57UjNFCpRSpPJml6WoAVzqEeWDq/a7oDDUWwLazoYW1sktj05teLh6iW
ocPuF9vuY+DEiX1agjsEX8Y36l/rhccz45Pw0nxlRGGQPxMWfcvrf6+JKDlqtIfwnK/7DZ0nKq/s
Ml3nHUEalrmjTxAYYJO+yRedfT94e81rHwryb24GsrcROap+um/HhhnXwyFhOqrkT2y6TrVGW9Xr
Aph3sLnIrZuvf9vqZQaHSlPwzivvB6eB+ovNeVrWWfKF+DgtbLDjrO2eRDxbOeyiYqTcp3zYwoWG
D8ixK/H6My2nsU3yHhdqN2k1AFsVowBtqcKZoaCKZKO6jkn+9dWF4a1ET+YlrsLdtXaZCslKbGga
uIyNfv5ujT4HjN6oC1yZ5RciwPcV/lzAq2A+gVydiM7BGjazI0bSL7jmIh3wNhg10II/lH2h1QIf
lcLQhdAImx6rAvGPUjRvGqJP1ICcxLb9tQ6uY21KJ79V4pgP8jHj4jzBrc+fdVzO5rzHlBDi70KC
BThqoy20CJGR1nvvB0CV2uJlR+oQjMlYnug0PyGZN77nYRLkc8e3xAQ8fx5dU5wjrdfqNs4VcKIz
qEv+iWRDFh2yi3Ho18oU91KgYI+QQ6ySPasvxRXDqo1qSVhTmJ1nMGGw7qFeguuUVUCgBbbGlLSa
4J76yCbZTORApphQmkPeFsuobDuZZt9WUm/eUhsi28wHY2Ci3+hi9N4BAEjhjwo2JKoEuRCtl9Bj
u1A14m376g+KImN0ok7U96NmdVT0wxCzMG9KlDvsMlpB51enXD9k3S2qWn7QwWhsJzdNznPF0Kk/
mMTL9RM/o7u+vx5VMOnyKM93EmGmXVIPGX3TIMvRkbIpiUwH8tVOqhE6KYdLYznAZvBncU1szl3W
E47yUWJpwuPF+KtPZW8vHOkqKWEQOhBDr00qAcbh69oQpbvNrko3BD4vAGPrqH9DE7bK5LX5K/8g
mmAg9shbJKbxZxOwLsErhQRaSh3tY1r7pJo4hRZ6aweIY/dfgcq1QKwbIsHd78iazltkxttuRJmQ
r0zmJEu3S1Y24grwf7tysAnwF/86GbHyWXZfRQGa2F55whK9xJN3NxLpvEuhla5HsMMHm+CPZj19
rBniyVbJRAfk24BsShCIGYYP+xveAuNMLvGo3Tly7hb64Tv4BbR90e8yAWgSJJ9lccqu6Vkr1vmU
JwdBAZpLGSFzJvoKEH2cbjGSICQ7qOBv3rvCFelE2CQOaxEJNzCuBEw59YM9aU8zZCih8AN3GcUi
fiaMe94In1hDdkz2CUuOnfjApA1Z5qn/ijwDBC5mDddnRUSvpm3ylhWWJG8sPp9q0gYkWNYPp20X
emZ9cc8E+nZSF0+xfI2mOzETnF6ejdisvOmeu3LaP2idxu+PXZFazBPkj68I4SUpFlrV2pnqumtb
clPkTsX1M3bbmzKka+LzKgAdceJU98CjHduw3Nksl0slFGIl194tI9s2Ug+Fk5/UQVxvpoE+ZVOU
IbyHTLQEZ0CqbAkxdTHUGQJwcF5gYA0wRVdVvar0HpxevTvUS6/rFaOJzh+Z8Ew8W+G9Ikqy7w1v
TuJKxT6fUUom/uqwYLBJsUS/sl0izmAt6+ARE30m6f7nRnXwhNzouPfPH/pzlPtA8fT9KqZEA2VF
ae/OsV1lPzCaRJ3zeqrH8cDR/e0mGn389f4it1Ws/EBXSVneBaRC6dNjk+O0g9vsnrBfbuR4Lx5Z
ueKH9zve5d28bqt71rWtDblA1K8/SONnoKwXPilmgug4r+52cztiqgQXVDB4BIerHkUmC6gZjhey
hBWf6K+YyIOFQ59e/ttsst8hiGIWxQ09HnnYdJcfxYxQdp9izXvRUWrB7+sLGN9Dkjb+CDnt/ASC
CEecpRaRL4NG39l0Y9ID6G3Z1D1KAerN4eAaQ6Efd8XUHQmWtMgZTOEmYSVYRsz2zKQYE59owp9/
o4YXc21pn1bG4BolcG0IeX3Y4R9xvMbC8+nPhcyUCjnVGZE6req6f8AsGaIfui21HqfzaON/2ZKe
a2sdZp0boJszqXb+hDWcFrF+NEVjCgANH4JPYI08pLz6aSHXEFVC0b4OTccYIRrWfdRSLEnwfKLa
Kyxn1dw4uRq8ZQ4QK55k628S+R0YtRt5RXRFd8HIBt66Tl20mg9N1WKex9Cg6aW7GxIOgImyA5YX
CCkT4v6E1s9ws5IxyrI26nTbkZNlMsgMLbSwqqM1L82ker+gnMDKuzWyn9FCOj2sWH5Thh9X5zXb
ns9MKanNftB2Q1SaoDv/epqnktnqsLV+dNDsDhXWFk0IqSKSX4T9jbDd3ELQl1JbrLaFv1m2LFiQ
MMMAz3IEHXotLb160ccifde04Vt+sQJ3Q1AXrX3yIwgoqV0rje3YvMDvlZSHntN/oaH4KVCG303R
L5TQAVdRih+2AnrZuSzFcInyUdaE9DgYUyPqimq+Y+an55KYlDY16/6aAGFF3mQb/BG3zFXeL5lG
gNiZ9JhL8Tf2vuuUGMlavMFq7P7o4tu0amOND22Cug2ecrLvdfPXagUTRw94XgcmtGQUcK4LBuFk
rCe1rwPbCnyaZYLnjbKRo0WwU6ExIjWXpc0K3K52wUrynWXhRaIKY2JTAMwI8sEGWywVE+5EAnQ6
krmt+h6lYhL9ZNZ91lvg/QF8Ka/bvGNy54Cz1HXM/mbJ6c9rcCw1Ess1QBkX9qqZ1wDOyh4e4wSg
wpJuQY7y3i/gh3RNapnuNHJvn75Nova1coL6DAh7MKd+5NRbcV6UiYv5W2x2tpiQlHBAi+TnDW+J
r9DuQoOgrj7CxpuNX7Go4ePK06+CQU9j4YpgTKi5efQRjl+QLtl9iYtFoAfoJWO0DzHnbLDw+ggj
0r14WpcAtYcvo9P+JHUUhHmO7zsj/Pm/3di0adozeHq8RNEc6sR3BP6QiIIG7GCcO1GjtSrfB3jH
tcL5dGi4pvYI13T+q7zVATbbjXUp5vyppeqvv2QzQLeKh9GMiY6lpWmzQgbG9h+KeRkLSFGhXgzO
Mp6OYWzR+cy0qPYn/pKUvqobhp89Bcjcu5XmzmYmXuAjJkQg95QG/9NqAj5GPPat1FYFeYwS2wM4
1zyVddCZVETCU82EqFVavNu5GlXCYID4WSrR7jd41yOvpPAHIWn312qsxRuYWK6SO6bo6/kPb45X
ZlrrO+h4B7IwlT3vJwEg0fSo8Q/nzBGraAKkEemSv+ulStOQrNkSz3gim9NjxmbVkH1J727EQaOP
DOpftlCzYjgX7Pw2sILevHZJpcDXbeR2zbfyN1Bg+pvTHCGJ4Ib1+z+ztul04geXk9zJ0iWiK9n9
ECAvoVvV0DwUsKFg0xPkRPoZa+/kpokJ0GEPOkFy5rwdzVicw47qb+Bsgu3teOAjTrEU6dq088g4
9IKLla+IElHTl/F/YJoVMKKlKg9qDkLxVaeruell1+HOi4XrdVptqotJWmJucAjFFMAI9luk96t0
hPsyOxMc4u4C1k01puWfi0yccRd9Jl1xM+5P8WXhJ6rI6Bo9m12wcFlFz/l6OBR95dvewnYQR1h7
DUnawxahDGv8My4NP4HRl4H1SMKG9YeL4DBvc2XZsk+jh9KGXb2UzzsEL9NJ42vkhGIM7UzP2abB
gJ4RwfMmHZphB6xpa43BQLxsEUNocXx5/RA1rp23nPSWjClcwd19duyyiY6Thk7coyEX9VZzgBTs
xbpS+7r/9u99QrKyn9197Ur00anVZ98THGLcJcTzLdwd8Q8850imG18pBKKdNUlqjFx/bZGIYkXR
YCdp4dg3OlBpq877+bfxrQnsoZLYYHjU0sCyXVurqqvdztjd9PdYa/gO6rCszx9Q4IVIhHWVR8Xs
Fa5Mo/zkH4j824V4peuhutbhw5zw1tK4BqQZQpneuVn6zX3UksCcSTzgaaQ/6LQgoqdfVFGAfrqw
HK9QFnQ/Xd4wVKJ75+N9e9jSh/mOH7/QBgDbChKzmT4NV1BR44P/HAy/CmREEEqqqju20oBYS/Ob
i0RPTgfj8OlB4RmRQdAOD8oOGEwcw1UUE9QtQI/tviwoaC0K7hsHI6IFlmcDFnGRm5eW+cSFaEm0
OjCtY6RHOzEnTn41X9oc2QiKnP/V6bUnpkHiJAc5dZGUmTnsjxWa9t+gad2W8NZGRWoRdu9rP9qZ
zZHpUaWc186HA9OiOIM2+KHpAI8kPDO/cdVKcINGeLRI2tfHQpJg59q5h4skGoeu65/lSTzTdSYY
EFgFxmnS5WBAQgt908wbyGbyc9wyP/dEnJUj7Sv6tPOt6bgRBCB0HYi3GA/yBURhMIsU64Meo2OU
Ygi7eLxDjmXj935JdvMaw+k2Je05uynqonCgCZU4zeMceCW+eTfWb+D5zJV5TBKgLv0/WobtAsjS
EOJUc9wN3IGc9IIjwM2KgUcolPu0T9j7ePEMQYJa7J+pBoUZCjf2S2e37HIwtY/SwRzKxbbLxEmK
uPOo54tHidC4zPJHAMvVwNaqh5UysCMHZbn7e+/4BgqscZ5uRmDV4BoW0m5yztzD8cqk/Pi+KpyB
nZEoSV2TMiz21Fp5VllwDpk2ATRwvCJOrwY+JtEzDWpCDvqpPfr3NyU4Ss5xtf3ZlB3PAl/22H4d
WWE4QHZR8WrO1iz1hm4Ksyp2jAGb8fAr5LOzlYoV6tyBEKffRNKSZG/Z7ieQjUioa3ZGv0WAjvKx
1HpN9QaX+asNfTVIHmTlmaUoHziMwpV0R7dm+XJbbJZC5T/Sq7w30E2wROhZpKb8lm+/rMPFsn6L
JScpy7RkbFxrQoj5yi1qFIGEB9Tr3KGef2NSBzREjObGk9Syay64TTqp7f3UkejpaUjH6YbuhA1R
+zns81AMeXEABzYkfksLOP4Oa2WLRD7nHfullm4hPKBOD9FjbsvlQflo1GYC2wgEeIssdE+bpiV+
QRyM2GZrZMDLBXgtyvdbXlsIUm98HUujUFb7zAJzMIDokFXUnI3vPLZhhl4rFXKDntWmHjA7StV5
9r4crIbE1xVGHlhNA55uUlQhZ3HL3HCNH1/HkM58vZ+75QiYw9vBIUvIqDWj8ptBl+1L6UK7COTS
Wnb+OZk8Uw7JOkquTaIEgFZrWNkend6K0mbbxWl1N1FQl+wn+k0v3cZ6bIJ6xZ3t1qqg3xbsObT+
BoPOj9sJH+coYsWYOjc6sc+9lNzZm72JR97wnkugCIfK1y2dBpud5mgxV5xWCl89UjRhrWBmLuqa
ub+OTLqCPpFJL+n0iG4Aq72Fo2cj5qEu/0kf9f9JrM+ubLde6FX/iw4ZGEgOapl0ArprvP2ih5Ch
x0oDQ3Ruzz3yU2fLmuqNo6kzvO1kGiQJdXlbt9dFwOa0oK/pYko5m3c/hFIgKBMFyICmsouLPU1Z
3KgbulqGbyVr1WKz/QhjGTQbZsvDrfaU264W+FmVhZO3zk0bUBa0xxz70cTTy4P2nZzox5qB2nFp
z5Usl3lwfW1AVyw3ewg9OydG2TAtqppyQKdZyEOxelDItn6VBBzTWretthbqoeEwdroWMx3D8QcZ
di4tN0W1XNeQHWC/tRHgzmYGpR4jvqREL3dPLM0qyWsj0qqx4nIFXqzpJp5BLRRyFkQ51HrJCT7V
hlNyZLMOqFrrzhAPhw/ELU/8np2TArOAZRy8KRfkJ/fSmF0GnAVAKi96M93XB4fRC5cKq4EhiNOV
oNDEAxe5zJuCqD7/IT7cEQriHUpGYN0M0LzmOyRVRr/+3FD9+qDVx/s5Ebw4GjiWYyeiKZwhcIUF
VhM7M0b+6ICGgmp6eP5qepIHmukiS9oe4+y6naybuinA+vcbO5efVysyarrIft/JV9vurFakMI5S
o/ahB/9SRjIFgHD/ur2Z1/eNOuEEWKxJj2rOmP5MzMBUpr11EjG/CQ6OqG3y9EM/xjTitMHDppKp
jNsM03B7hkQYLKeXOn3Vn+7wG+hwPmJX4xhmEsKpUjL1XDkS3JrXhPUQgJ7yq8dJ1JLj3h7pVkxe
ym416N3FJAaX5e/omeWQJpxjvyCe20gRRhzf0tF02GoIK6MA9tp47v1RuDwqWX4EWjCCOVxP4aJ9
5DKgkoP5YvKdBgxXo/erONrogAaaHHTGk5mBPkpHG9Uvi7CApFhPT9Rd42B4U9thVdSM7t2WJWWu
DD9Rt7haZBJSqOZEU+2KsdTiU1SexYqmeo82LlLX3J3SD5xqW/29hPKXlRSzMMgbB3eX5tMmxEFu
1Z6zFlAPs9Mb1TNTfxfcIoxQH8M7bDUHygZ7OraxEgaI3BjoH/RRoOUJ+UhxolUpylSeUChMieec
u1Yua2XnenVWhJ9NVUN+6bY1IFnGcIHONAV3eCjdeoT4Rx4gjiKNxhFeGDih+HQ+2Eo2+lB3HsBo
VgmwkCuqFh6DwNoGxPdYKkOGkqNVuXHr0eogUAakp7KOUimBZ7b185DqQOiOZb2Xrnl1rCzVvOw7
ePl6zCLUKkPL7GD4ncmgCHm+LMj+qpS1CO03S3LffPIsQW/OPWg8EHKl33uC0DnBMBVR511tERFY
iA+ugCW15hN8RjoBU5hz4aKZeiE26Y0KuYaD7d+/1cMelSz8Mr4nVKEaenQKetKbaqsbUnqcYILl
HrGiBrt8oCfktMMoRiJKL0B8Xcteag0BGnCpkaZ9SxDRjl1KWJnhdvqwEqQ7gRpxQX5yKRmy2YSM
c1pONYeFF+ZYBl0hjATsJFTRIFwtf2L8uX8j1M6VLSjTGWjGpwKhALZIJJfiCJzfcTK+7Zu7BbAj
8AbIFw+R6EILMmoaA/KPsHi4mXHjoCGysijjnQI2M5mqQ3GBJx1JHUdbGId8JO+UX4/2gyz62PDv
iiRc1KCmkQc+0AkTd6kd2944bjuQVkQuqRGBPPRdGcjk0W2r3kSd5vBea6XWpLnHp9gWWhdFK2Xb
6FEfoSv8VG0/ASdvLsvLLBq0MTi38cUEa1Wk+bSR8p+2J1AvUzLqov5ScLNTcYg6L3EKI2e6KRqw
5jio8EzCQ/fVQvpq1InNfsFjoQ8gDsTrkA4QoD+zQBhSoV3+Msq+aU0HEEbaAjH/3RHeIW3SAKSK
jdba8EzMNyfH+V+vfN29/PbRJ6x5Yhe4b566q+Ec/zDqItkkL36is31CZ5l/P3yQmm6vXGHLDPm2
L2abDg2Nbt+jdlZa+clpC4tQAFZYHWJrye+9N+hP1B6rA62cn2lCMA5zbElTAMLAHwtL57wRsMdH
7FvGB87lR2yeYKP4NbrYRpXmy2JfEqMfpiQmtM2H5x47Rbs/tcudV6y8XNAYlbyWV/VoJcjzVnq9
Qz73D8Kiyll/cYG5Ic7Oi66E8W5FDvg2ckUdqLu90piXVcm3Tm0Y3zAWFZVEequqOkoLV+RvYepb
Uu9PsSdAjPaAQnSD3OBwNqeabkDUYfGJvX2c/2Nln9SRl9mp/D7lVe+gHqVTdn2SlUR0GpbPQpt9
SHwtxRrzyMdMe9Y4XeqxA4F02VPAn1YF+x0ebkzXIboToNxOoUQ1F2Tw1OVCuPNLOktiWPzWhmav
Mc671RAvgiDyN3BbmQr0d60tcQuU39QgVbFsQ6ZdipgOGyqCYA3x5cRMruqMSR/PST7+WNKD4HN5
bdETLCbt/P6EdGF8Ner9co4IFoaEpzLO8QQJwb24e6IBIv+Fsz/pqvczwrL3TZ1efVFBAGRdI2Wq
yB0Vkqk53TosfGx6y5YENgJ0441MOhnJaIHRPH2flcx3f4EZnaawqEp6fyal2Cw1Xuc2DyFIQQ2K
u4GEljzncae0w1F4c3/Mfrz4JV+QSuIcymwJ5DyCS6UCI9iR6txx1PzHIHyo/8RTh3ZJ1QI8U5+c
qdWmdkkYUJja35SrTNnpmSGNG6+o4R0hk6e9/jvWpG9JiOJd5vCZs+xYWIZpHGb8NxI/hRejX8T/
sP7J4lOB3FBaSRZVWfcQoEr4k6rJCglwFb8og7gynEGHERCGNm4BXV2PknZXQ3ADIlr8HLzmY04l
bRJe5Fm6y1HQoaBeBnu/U+35t+HpslLXZSOlN1U4IUEOQeQPVHY7CuCGH7qZmbvMm6acKwEatsEj
LOOSEu8oc6D6umTRf49qCKFF/99Oa+AXVVrHsmH2om2umqnoUwWxXPVCfUBLa+zkh3YbPfOuKJ0o
8E7QSyy9hK9x9+SNKeCzOpgCG4FbuSYtjrmexgBlnaC/K1EqCW6S7dE9qHDTT1IuHdIT1FojeWkU
/qcAS3lY4Fy8XNoCF4lq/8otc1CIacRX0ZmcK10XTBi1wYIp00t69D0Al/qr+00Lm66QMaQ6t7jS
2UvVSBCieIonfH7UaCgUOr9IZcwC2xwlyDixEid3cUGRwS5a9lfJowjG9eCxzXLx/BxuDHWSNGF1
l3f+yPeD3RQHgcYtexVI6rifiZjuzdLx/oMwQDdPCzAKWWZ1kkpp3jUrAOZW/vkhxi684blsS7jS
/0uwWEMEs63cI4AmWtsKDHprR1uFnMIKeP2tnQX9+Hz+1+F2+aj2VMgL06RlckqjgbjlTeL+viZh
fu9Ew/xoWE16zDGy8yYH1QcHoh31cFGldxlzW387SNP9IkjgijDaQWyny+AKiCRk0mTgSHehr8vq
Jk42QhENVl1FpBE5x4T2KB8euj5Lj5NM9WFVRSY/Lrer8xT2tRrbKoV2/1bbUfkzUPz6FVSF7XHy
S5G+QLnSP/gn4WUi5xPVIpboIPfb6wfiB6irk3dMbs78SvpFwTd7KNvqDMnEqRoCOZroHT1veovR
rR8OJS+gHmX9V4wGcjGArOoK03IfBGJX55QKOZBQ3OPPpjxvAAjV7iU7iWcGyL+lI6uwk8WQ4/uz
YUAmwZq0O3/09Yd/EP7MpVFtjCoAz2DsaQ1G+r1mv6vDmiWX9BPPW/K+1myIAhmHWWq4QEdVEZHD
Bs5KzcEMXqB+uavQggLjkw6HafzTmNYGek6hXjSrI6U0GKjOV4GgVPaMB2nRAY+U852/c5hQG5k3
9W6qs8EZXKomqjFbVn7FNNspPyXXGCc8pUavHcarwAyVd07Y/Xuyi2U+oZLI86LlXXUluIUOkbbR
wTDC7Vcre9ezNRM0mX6xsVUI/oojuptUse2/ULIzeG1ABbfGa5IxGNH4CG+NPr+Ec1ur0bSkDjy4
o82vuaHYX6xcSWYbro4gWlt+V82PNWVIQUrYNSsS6AjsQYUkko0Unb5I8fVz0qq+dH/ewimipFSA
0/UdR+H3PfO0Ayb+vyH5HZmlaHSIzoI3zlgqhhQWvsX0Zvy8RKsH5bcnNkjEn1LuqC7QXABi6AKv
7IZFAT+Ii6Gf7uwBjI7chsPQ2r9cCOje//pAZf3hf4NH4cWS4GsHyUlRjLT24AoxjfLrNNoaHfY0
5aapDJcSU2AIYFyeLQjojyCwvcdgsV8F1xacgMwF0/A8rdiuBrP18uFpnC4IZwV0prSSpG6IogZ8
64N/MJlwQD7MQdGAcE+8bYmtnuRygW86+dmOYyWEih+ftdFPFImiNPUQYPwr5NukvjorKPP2QTyM
pPOZLKC58fJRYwAwwOvhcDfCp7KVvVNxwU4xVWX1uSTVkZTzCVtCk3ZawTAxyXE810zz9tcZOkrQ
5PN8K+ANJ8SG81ESXrJ9dLHaQhcJwaFKU5MffFYswERA/hwk4FMlHi3XlJLN+I/8GTCdmvJYmOFZ
hBpnZyeLAH93TXteClsvsAtED5wubrp+TtZW0cnQaGaNwqkTvkEycdU/CoEzw76Kf6MtJkUfLHxS
Yr6mgUs+Jty3V+8IGOm0hp7ZIycSHyxEQqwmZXFIccLpp9/smED2569H/kvWoGhZDoWkd+7x4FYX
NivykFBlNuGRAHn6LEr8RVSsWZE1uUVTyUgZpoJkqf5dT5cQZIe8bB2R0GIJkt25IhUVGPx4mRyw
UAnF0tYhKIsq4ilxqyMXide4BJgpGlOeGkj0YaGTO4N00057AJ4YmIuIfXK4eWvjvvLd3L/VzWOT
OnkfbL6hEybzRMp1lT9BkzfiA6M4TGNwtLrgUfFpSPd6WnV8fqOoTxAnTu2mCD+fShtcS1Kvs7Xp
sBE/PS/xiv+beij6Zm3rC1gGpJJHyCIjC7/vKF3Nihvqr2wG6VxZHbKFNO4XuH+dam8/TXuoGAib
Ttp+62FXzN3MgbFCa5PufS8NHqPsFAzErsMK5VKh10Rss1fNfNuTTdxsEJ56KQiq8miUrgM8SKId
uZCMVkDONuta/fnP2EKan1HTWbskRP+5x4VaaBIcf0aZYQt5PtfTS413wp9LwkddPKupJP5udZRf
Qld1PKsc9Ci1oRA5ckluTid0ji3d5UNljRCeWyOE2rnk6f4NLk8P9HhOs9GiCAjgbDh7tUYqYcyH
zvtjIh4wNIJZytot0pHLZgUjV/oydN+OBSHcNhwLNTW9rxfXHrUDuYG4hbLaWA1W2A5KGxUN52L1
aX1Rca9yjEsE8eKvilEcAhVnYuVQ596PuyRswFtCn87h01b3Raf+xjp2oiCXu6Kmu9NU0qflX93t
teiXXFhZtu1iOU8TGL/p+bQe230OF1nVk2EsUNDZFD9qW8ELpkjzw3zTKLYTUrkAZT6x5xd/cpG9
Cyh2GAo2LMwZgo8TYa9yn9Rp7DGkBnjIif4BwGsVosjxvaszsimUch6avQt4TlSA5nyXmVf77xcH
E41xCv01PpR+e3+u+kI+Zvz/QpLwesh2NNROyasSXU8RvEYRhNflZCUIQaHcUIA5xPcjZAP/Id51
Ipgb+Ifju+5NrqZwB+QOZ4oWmkFkMnBUO7bB3FwUJvHJXNm1ZXVCEBm4Xt2r+QOTQSLxEGDafsQs
SNItQf2giJ6LECIBgD8zd8MO0qx5JD9JvkWl2LYr9te0rqqoPdA6S1jnhisNNCn0uzDeBgavQeqj
vX9+IiBiZt3JIiSXeXuk+BKa+iKBiL/h7G4R7TLJf8TxEMGjb9McXsyt5eSRzpDesxfiShYK4k4+
p44/bkk5M7DNpQ/nt6XCMsEy5vz+d/NWoS3Ln7P2uiS1t/3NKqqo4AkDxQB+caqH2Pt97P9T1TXS
m6HnqzKzZANYTiRAMpK4TXKMS0E/pzvCOmBF3iad9BT4gP/u5luhamJkanogv+4ZVDjhQ53ku446
QMBOOOETj1cb1D9aZJ90jI5emVL0D9cokk+un4qsVEcBqH0vPUxNOil6FKTpI80JbeU8mLac4Jhe
3xLEPzRKRk0PQ4Ica82QKtNBuSt0OreqjCtCJ7vxCI5flsarGyQowW1ZSUBKGsUpZAyk3MyMLnWI
eWDzlfpJHjNcxYz6Gxg6ych9GHiZqfClSVZVtq0JDyE1qwmeXfZqbuLLSeFdplTBAtX1Q1TJOgx/
2zo7DmEfsb71L+XkIW1AksOJXnJ05pwARpSSagGBm1yPcmilkm5DksC0Nm1xON60koNx390XoTl3
QjD/Sgj+8mmAGB+Il3CUvsUv2x643Rm42491wuJ3sIXMrLY7SvMLKRF+y0amiF6UHNIo8Gsp1MEH
PBHLXGX9d9XT0timt0UwBsHUpPX5PP5L7ACZEREaqMYNfgrFneI0L+gO/8AXrlMhpGTUqZOHs2zZ
8rhB3NAFnl2PSJjU6Mj/0FXtwJ/hyIvVz1QBTKriMQSZcD3HWyM4lFkEBzHHoD8IL5I4K9wRNcww
K16Lx/8ACpfuh6AtoHqsi3Dm8g2hTmEhLoG/iHKePKm2OCIphfyQjfrq80Z59Fv5XxqPOAtrJy3n
CbsXy5Usc1cct56Iky+GN8Au6sXgN5cOtQa/G27zL40m/9FDI98blkOyAiM0vQwMGe/PDlD9EQiF
NMPnJpp+Jb/zDN7D+y1tCwMxG5eCmhiLdFrLOE00wDvO4Oi9MAHLS4f693f4deq/EwHznBre1SJe
CyGI6OEm+RLi9YxyQCZb6Q2Uabn/UgZEFUnreihHd4eewzfkQz/2Ps7m4JaEr795l3/PMCfG8E1x
4/4FUpHVcmPRRUX3two+9YtDdjLTkS1ISO+hWLttU2/qub9rk7XxPss/T1vr07VC7ijED6Pq7jhp
lpqJtXwKMCpe9XDwW9Q7AzoCya7XG0oOAiS4pag7MrZdqGEw0ztSp/TMR75OthrAvJRoidr+9l3s
L7kRnHUyBkTbYFakxdHEoEww2xvYitb7MgCeVUL+o/g5KwyHSPVgV+0a0MA9OVE0h1nYrzXpFBd2
2Ly5f59ljHWj9S1J0NV7smsOqe55Q/1dIP1e13FhZbNOm4yUL4U9NKqn6qQ6huxio0lEhWztVzvU
0HYGlnOC6YPbz3QUsVnQE9d4e9p0OYM3k/ucXAryCEkeAw/g6q/EepatQxijs6doaqAA8C2szJq3
PKDLXc0Wr+rZWG4sR/OBzswP7VqXpSDRbzrr0ZT6pshzvBNWhsu6yfFXWLdKTPdccGfbgXvfhcOO
7bu893yiuQjONaYkeAnhp25flLNHMAHlDnJFOLu3G6/25Gfaet45fOO8ywnaD8M9FIm4xWbRSxw+
LyVjjHxoGSbpVzqc19LiKKkk9tGBIeZ9V1eS2zsyolg3trp281zyhL7EdY6EfnQrgPWuuOfLH7Nd
hiSpDjzaX0JHtmuXig9HOrEBUR3uascxxAUfgNCJBB/UzKim9G/dnuzO2P2q8VCb/tm2eyZOntxw
F7tVaWb2Zh3tXEdrhjQxQChn+2DmMAJMHcKB1Tt0qA97vps73i+9E2MpFqE+G63+7rssS6DU93MJ
lfhuSFhOCANOIRijkebUXKf5r2ILcl41jigY+Ogejj3YdTptqNioypGcMIbF9yvcqT5D9qjR2QYX
9n62H/e305/Ya6DuX9toPgdYfAXp4ILyH+GZtUzcMo/dmBMOMv6mlt6QrZ9I8HOnX7HZtqkcrSk0
ZbghdgqYYZj0Ei2fZZ/w/INl9UlhOqbUaypBOSSK/nqWI6lQEXjEbLr8mwtXgjphCMZmzRNCRmgJ
eRlEt4e5WD3BUEVMa26tclxCRtc04r04bsPdEiHJpK0k5/wQT13bN9zl1GxVkBTc/Ti+DYA1O4dC
oMX2/3kP4D08WmqIgZsMlc3cEoDZ/8OPYNx66CSuGmYRgfalbcqAedeqcedol5R5UG0S8nYKFqUf
sW8QIosLlM/n2aF0G35UEmma2CeXG5Osr80o7x5L1bDUg/A37H2yb+Fg0HZeUEVhGh016YqCc5SF
yGk7ei79/7gNg/T8b7B47oXExSgZlUoZZ8aHMilZOHhmi5nYy+9PDhh55S7cRcsW9d9Jvfgf+zSk
I2HCqhhKPdWHzbAd9XgPeX8vlT92QyJgS4NsG79A1J4XnzD0X5hg/ar8lIFPoD6muXSr7PKPA7sS
KEj2rjWy6iEW5S25DeUNLt1VcCIHnT4mR60bcpn3aLpgDsWOnIPtenrnij9j+0a9aRipGWuQ7ipl
gb1cB/qgqrEldcxGw8YQ06fYuloQ8x9dkHi9PQoaUY3HQTwbUA8DAtBCAfSBFKeGGO+rvC3nKpDi
EhbNIgkIT6LY8mMhVFDl9NyvLmKtPm1/erT74HQjDal4OJryoPBH3BeSxSwquOAGS9fmX/dSRPHV
EOWYeWDYb8do8VIppsD8iBrvZhgoql9W6zM5cbbOgaV1IsTTHHFSdetjkGmeRR6HGVbGGGbddHuS
4wemPXky9JipZtsFqLqlL3O69XnBqliVRPB90xzcMMhB2CYXJpn+Q9dzuyFUu4u/EPk1E/gx1Afi
GU1kd5bJt4eewm2xCQWtnfVuYQMP1kWAx60sGFR7NMGb8j5RwOddxEUjSprpwTH5pRM2QFGf0EM8
gGEiHGShAWrWCUv5fvKvb0BqwNRo+b0+yPHD5rD/Dn+WDIWUDVntY+XnBHTwK684L3ZOVjMoii68
Qnat7cBkr8/Xpl86LTwCSTaHn1qnZMCzc6pfOJeR46v+gOpj+i9r+ScAJ5rTo4oHall2uw45l58i
c4FMhiNA6ssdq8ja8AtQMMSOlHxxQ9XsdlsFzTfuW9Ns9M8fLkUhcQUY20PWNkYMuNoebCCEQuIL
ifaL7OIs1d0a1HXCrYWtLYkqvpr5e8ZBCk3sMdu5dOsOFe1ExrXscYW935/7Ri1AhNNA0ZL0kR2w
M0fcXUaQv4vI2ft4io651gs3DZPxQcls7JaJkRmsXFKq4ZsbKsSJXWN1teWxCvRapN2I6EnxNLfj
/t38K1ayGR/jJELx3EEWF+oKIT6JumOmNcZe8GeOqAJam2WouoGUVn5/7UW1hQMItGg2qoggUYpS
miwtH/1XGB2Oi+JrS5reKnRzgEbn4x+FB6/v74tTIMgTO0iG+qOM9x5wAwqTFt5v+uLbQvV6la5W
CRf4CUvE9XDVGdHLYT9fBYzTlnKUpTP88H/zYhZ8gDRVO769kegl18l0B6fStN+hgEsu+5xum2P9
LTD6i8VHokhya2e6LGJA5BlhLbi1IfSeaISV+EYCjCqbDG3uNe9rAUCpIh60WWR7zyGW8LGvXKWQ
97iyS0IWkm4Xl6aitraxk182Xx2hbvgm6ZV5Ky6RHfXQyvFR3ZiQT6pqe9II/nw1/O0paYl5MjaQ
nVpF9HXlJse2egS3MGqgG6QLHo6zfwssQ4TGsoyzzXiK+Grjpc0kIHv5J+h/zUxG8DPbPWwO6iwF
ahM9hK8SQL3axLPnr5/veOIyAaUoRENX1B/WrIly5mc6oJ/Q7o424+7C55IUtEY31zp9hPGfNw2Q
B3CTHGJ6BYJukAW8Qe75ESc//DSxUoXw0/qGj4DDHXUPE2rZFyB5ZDJf3XN4oyxVSeW33AJ78xLH
B4ZURK90VK/RETV7kWtrigdIIu5V/uAZVuKBzSeaIL1Ad0ui7+AV5R97VxJoKwWsrWsSDuOQQ1l+
/v9DLLeyNkoAP5K0xHQV++BO4Hm/MtaYgSaqhOZ+MFveGSNTG3Rg9eSkcDjYypSbjBykn9nLlwcN
375a1/hKj/HBPOiyZdonqloLoi/043ik+JnJQjgzQE8WBjx2HkThd/R8xV0n1QAXq4ee0ttXrHdV
P9s3f6rDUT2FtzqNB6KdK+oFxNCirxc/TFu9wAW0awlqm0WwxEPWQQv3sLIABxGeBHm7lZClhh5a
tOEAoDrGt4SWHpRDxjLA6eiPz1k1Ulbz0qlywwSJSFWv4jnJHGF54feXDhGnFY9gYbp6IyM6pD0x
sp63EFImJ643m75VFAySANKHTwr7rNqHYdxx4SXz0ykp/rVuz0QQc+u4fi1HumiMzXsT1y2wCTs2
6z5P2OxUW8Z2paZtCcoTxMvb1od3El5ZQSDj29nBxtD+WcHVKrQWwf/mthnymyA+3qy+rjausWV9
ksn/75Lj1o+f3GUhQX+NUtsYdSdjmN/91qF+2ConMOea1UIvWadXrKK4vNp4+xGfKsTjmAnpApnv
cFqo3sNWmSZmuxCUMYnP8mN9TL9k/F+7Nfmc+8L/NTfJqaOiZM730VxGsA/c8feBVXH7Wg8KTMst
cz2ornEtnGgRYzPtPEEmXqoTsCtJU782oXnHkOmH8+mFKMtF/EJAQfwQMJs4p/ULrlKVn8gcoMol
UnMhQwJDNkXJ0GSWMqAIR34BFZKXbBnG3Bl/2eHXqhAxQrvBt0AQLRQQTeX5lZ/X2caKo6rjuwtE
DUy63spmA/VIizZdbXPjJ+ogY7UQXt0cnT4LREn+9KFi8oOclFjSrYhgcqB4nKMpAFZlXa1G9WG+
k7mNh9v5kZaqA1d+u7OVkM9j8NNmlbOjtXzOurOa4crV/uRe5jWBkulXvbUjQJH9gRRYZn7Co6kF
/G4bvzCbN7n0F7keW1Fthgm64epxeMBadNcQkZgoCOw5WNgJCZEgNn265ZxUI+JPyH6gyBFvs77a
8Ni0ZKr8SbopUyPeuamnbZPKjDzZkJh8TT26pBmT/y/35ngqLbees+y0oOkT8oVPSZG9xLefGw1X
WhrSc8B7UqBWfy4Betds1Jaf3jCAW5ywRGOT4bWL0UukbqDdKkDbZzCBiBEX3eu1Do8oBfSfTgAJ
oIN/KhVO7N2L7IPFjgOqF+ZeseAg1UnW/2EyGXLx9gVlDaR2oO9uD+sWcwYln89JsGR900uLnXfU
mo/6F86lj1CzvvUCrZjcMi9n8FO2UPoqXQtOyEiVI48jYRHJfTBfBgnrYBUBWyuO0JtGlKu5sqwg
evzuqmIjZD530ELzcfZf9IN7WV1UB2Pevb0B3KeOcFQWdeK9WERg96umQ7HENK5BOQLuN9NlMBhk
gKbAWq4IS9qgX/CChiSmsq8Fhi/nvuHDHZf0z3d6vDxWJG1jC1Nl3sRp+CEK+p7BheHIIxzInUYe
2WWeykMlA8X7WT4kshYmy/jhsBaWwVx7uA/WrvuoeibqSLA483+y9BgEJFexHsvCANomTgOCOyRn
3YOkQvP3+/tANXH74co6D45bXap9IG8GFQ3Q6y4p+m4U9Lk2kpv3vcbrT14dFR9NE+LleN3wUdmd
B4b4ni4hUGaoQ8D4ZYB9z3HvDEcDbM/Afvd5Zm9VgfKlVg2i3KtZCJiUrK2ifJCc6a1MknEFal75
gyJSn8Rk0y21hnIOOqFeKEEgmbRMisK5NcGdrnxCfbctwvhWyX4P7ooXYz3I8yQOcKpr5lYURT4T
hBf9Y5gBKFM596Bm8qwWi2/WYEX5rT83IyJOgZJK3FzyH/5Z0SrbtQbjxFHVz8NHmlqwo1USQ+ys
37EoqIP3jzqHR4hIiIcyGxzbDQC1QD6g7t9F5QFQtPmBHwAOSjhpRyV8LV1pNMfsnImdl3FXcY/m
0dzTvrNikO5WkTxCInSDfYfo4EmmrZaZ40N8b/v96e18atXe3Mljf0TAGOKsBH+P7IxGQ5CD0Vqa
8Gu34wHZGqYreajFevCfXA0MgQoGA1ZigIuFHavTTV9qb4HFxmLoRns3k+tc5NITsaUVUq4gfyNz
4tHH9mWf8HojXuwUWwFgLMMw5+umt+LJpw4crFQzy7wfEDukr4q7k9rDoKQnEXzANzkSfxClZ/1O
umo40YZ+UdLBIT28y4/XEMblf0/oQ3qgmnPc70rx1be5aYlkLZygW+HjpORwiY6BOz9shYqoSIsX
0UM0ie0Fw+E5qGaRcIAHRYnF7bue91HKx3+k+Mty/ea2S/FOnPvMin43KQo9VjL2gwWKvg+TveX+
zi1/+SKXfv9cDvGlD2Zy+VQsE4NoHNYmGlmm+ck0HXaZJlWrZdcVuEv98kstiBYVnZAfmOspcqkV
28SFH4hYqNGjdRmqNzdlS+lPPxAUdx6e1LDPikMM74vUPfWYsrhBOV2RPs6PUfXmUH/ojGeTqHWn
b8uQQL26OnhW+Rq+yeQ2wYt30WKKY9qxFpY+NQMVZ0+6mFcgLQrBGNTXym1HfpXZ9BzLrSWbRDxI
KCwbUGf8X38Y9oV8N2wRZ6rhAAbPcdcKNLmLSeT6MRV+L3KyIvIyCukNgC6xq15jidEtjjtT4WXG
TEmiwU8TBzyjjR16DgIB7zNOtdaXygzj7ZT6BeevwXEB/8weCGS7eZ8+soxL75tXxqljlt4NSzrO
O2kDQ41cTMlshjv7VtGn9BIrSW8CUMk74ZIxRwy5kHN6jPmxSGkbJMhtoykUR5J70qOG+8edsZYZ
8qaVp5roMJni9r3eb691mkoNGOZ5hH9543yqYGIAhPr6clPjCGih81dhPuWV5r923QFidsfzHqZ6
HTpq6ujvEjlACL+0BhBSQ8b3FMXWBHAiMk4XmOCOh5Cko56VFFo2tiXmSVhEKExOE6UZEjIg82MU
Uok1+qua1kWomyvlYmkVuBAayMNln7H5IMxMgqa+0NfzeD5qrNOsdS3Rw13AX6vd5JmTXY61Ldfb
0S96Nsu1zmyrK/UPOJhlVUIpibjtkhj9ca/yc0DInM+gj0T6N/audguWPBazef1Oj+i+OcT0XAF8
SApKnjGyUfH4YB8LarZalZmygXZda6j5ROYiFhkrPmpzsg9aV4O69jwfDOaWiNE9nFeSmmNR1ff6
utA8mD6z0Jrm4An36MUhzTbHJ0ToVDg0TQ1rQ/IO5SohdSC8+zYNhggoSpopcflOUi0bO9/mhUvK
XrtX/irvX9GYdbXSiKFIpvVeL5tybex3P0WAqIL2GD3/LO+dkXRk7MyG4yh6VQeeizskt3jaFdq0
wJWL8ICRBs71Q2rXcQb8zNutLGniIEDWcqZg+CRDavvPRGf6MRaQ+mWgRBXGI61c+CRfOm5VsJqQ
OVYkbZZ5NSetyrD6X10ReOvaP7rrCAiQRyqmNuWG0XoMRWU0W8hzBxUA+3gVAeWFgM7Di1T463UL
T+ekeoUcIPJLiUFKJ4ribNKsGi5Cj3D0Y1LdAQ3feGB+R57gpxxJ0kWJ8YiKqwEUuI71mGbwChP/
slrIxi0ZPk0hWRhDiSGe9FP4j78N9ResIIieEKwCCzO+cdygu92C26T3aJRntmbJM997SZbUD9HY
MW/0NM3qIsBcDtZa+LYxnFUvJDZkZdnEgt9RNU4ePm79ehoPv3ZiEep4Yb34bdaD7MxjCZCkZfHw
auAhevmzHfGGz0YBmeWVMsMat4ajtHNCz6UhyjsBs9xcU8gTOsIOfAT6xan9xUu5I5NoI1fSO9wI
YT6tSWjDYlbSM/nGMu2iGWjZZRhTA9JvVWRqW2ybOxwwrnbkJQo3+PeE7RJuIbGJhitwaUd7xAl3
hAb88HApyW7WZWg0ifvNE5YBiTEYVP0fRqo34cXaJHWD6RvWPF2OW7j8P5MCf3qDowWdeL3NP00/
xwThSpz/ad5rSlroA3jviTNXqO+MesUPNZ70CpeGUcVDBcR+Jm6S357tzeSFuU5AgCOD+jGZGxzv
g1YxcdYbXtHw7pF0PlB+BWsb6nxulElC9q5utSTMzabLxE+oBMAwAiMW6ncSLUPEHAuxKb83nvC7
MuT4+MkpulGV4SzAGYRwuqaAlcA5RcrfOuiECi/kUhKdHG37/p4kUXYjSTO6yifVRemBjJ06sJjo
E43g0/KzuVp/PKi4xRxrb41K5ojDe67eh11pukq6cVsud3RbE66j9ng+Fl5djK1isysdRxxRxpR3
huHVgdjlDjpe7BMTDOd2vlxSb0HTF2q6zwm7Zwcko5fgxsyo0Hp3DGmf0Oq/hSxI7mF/mxrDX6w+
v4iJfBOOaN+I5DT7dygKDy2jeC59yXL46NF5DvWJNYyKBjEXL7ldLs565Vj5kgcKxSHVfMrWH6Eq
MRfhL0mv1XxIL2EUN/1IDSpcSDt6BQbs9ruttJ40C2jxlRFawtcDE/dZjea6i79PEKviptJZxAJz
Q8MXjaUG8FHvHx4k2mEWBfozsJpRm6ZV+F/uierdsFQY4e+a8DRo8nh+bJcXXGkvC1wUalW7yGTd
aqncpq3PfKT2C7weRWjXsvokKHO16Vf+lr1r256JfJ3Pik9TCgwzCmGR9BUEdV9aY0174ddmoHTi
3yZYVCdUo38TGrC/g+c7E1gd4ZpMI4vlnGZdhE/tdrlg5UGuY6MCnO9EhyUj30QLDWwf7aoIWHl2
HCd3VmAwe6hjXFnmrJgGK+jYA6mqLLXO9KYr3G2G15Z/gntU9smv3nCBrSwSfahm9x2nCdPkFpzl
RIaBv1E3Zqyg+kTF3UJZa/DNDLBSdoMxBFPdsC26JdDbDD0srb+kuwzjQ4zjvXEnDfoqsXKJfygi
LQmOK4u7DMq9NGXwjpTYxiujwmu2Zbn9go/fX+DRumFOp2sTxQpTvF2+jr4oFxBOGL8z7ULQPyP3
o6Zz9utBgCt3lAF08aeDBrLrrvh8tlulgrRxqQQZypI97xmLwb5VEEJ9Ca2VstRz25aIPcmYpLYE
Iv7hvSS7MKz6+IS5AyWkl7EFZr3qWQs1VIkZug+Plfmme0U2NGP9es84V6IQWzuMmWlrx6XKgwGQ
5YFLirF03MevC8viu5+9swMpQelpgFxHFslxW1kzyfthhWKhVBjHSzaJozIcsElUxENU5ZQRzoJc
s4WibZVOkdqg3hFjBa1ojAGu+0IGjf6lm7AAPkxLMKSK8Znth3J6sKrKEfX+iOrwYhYu/rx7zEWa
Y+zyEjKdYJpkVKBl6GD41YlyM6q5BCXEcrQs5O4huKODeU0EZCBzZjxJq0pZNkWLCG4QbnUpQdTA
jhuaebfimzpxgYjrO2+IkBcWCv3tX1jk5YzwRGPz0fTbnG4ux2dno3TvWWRhMcfzxkg8M0ea/gwY
+jABIdMg9zj6lTIDB/rmqTO8vZo7OXbUWKqpm4FRbWyAtT4huuFuAgnUxHI93D6LT4L6lBBdnnBv
MTu5EYt6P/wt1LwWQX9IjrDlZwSsSBl19nY2TsCXkMOiPeFaHMSkfsj2Y6BN2v5Bp7NxA1nJ5hZb
Z9po4FmzIdmoF7wCwav/OjZZ6BtbyceJHjuqT1r1f9LCpmCigmMYnv6CD87GGkufbZZ75T/UDwbs
aktMksjp//N7S/Hc0pxKsPKZCwH48xIAO4LdKdJ3YXrhxKLzlieDyREEizQbN5p5VM/5QNkNGpbu
eZfsfpo5j9UJb1AxrEXG9f/eGpV5oOYktcklUUhVq1g4V02GA7oejyNPfpUAOUt5SJNZYLw94B33
xF3aRr3FxpKNW7xbLnF/qcVe/pbD3Pdlakb599nqYZfVlZhrI/64yH2Knan/QYu6EifxafGT50sP
91bxtf9+KErn6pp4AkiOyM0woT9SXi1K5lyEvd6Qs+3iWxoyWMeLiwHCY+IkzUD/FfoX91ouwuOC
tPdnrdE5K7jGJqMuih2oDfqqgQbD1VMo5Q0r+fUttR2Cqp+s8jZj/9EXa3WWaO/merN34kUEVfcT
pVzaK2ygvh7JzUaWUr+udqczgEChPskiIhaJQkTPzyZuBBX8x1vn7vA8IR2b8Wt3t2ICZ1Yq7q7c
HgxJggs/VdwfJrt4RDNOfOkoaWjXK8+y2qE+4109avZ2sg+2piSlf25CxmYj4Ae+mYc5CFXAwieG
pOdM1mBvo4LoX2sp1r0fhHAsclaRCiEMOEaHhe+Y3D6qeqotYR3/S7wT0do7c0qVsfGfS9zYXg83
3bRLOgNqSz2RIbCK9q62VOlUOCgx7cI7o+ksng6k3eZ3/rQI07Gw2LFb6xSGyGkdg1S97HxWN8sO
mMwf6r912vjvH257mi88Y8+w4r4gQzKlgqahlTFiXhofor94fJ05UEBjrApEI4pTx9QV/Ra90aiF
th+xz44oJ9la9ICT6H9tw9PlGCvLMUqhVCZl46gOokINY4nWJWfht4VbsjecsDjDwmWlNpwZ52pX
6oORgbQBDRfjzEt29ypAdvD8VkPSF+oOvj/0HtpMMiumHT+ewC66yZs7sc2XHI9hHYqkwBas5ViU
qHgk+zfe4TgKnASQhEm2griO53R7JIdpBKspsKfC4ONV7PQzd4woCVl3h4omtBkZQ5s/ZHJKGewc
Jdqdf82UWmyzJ4/0tjABSxSXKJKVb1h/qy9+4Tx9/G2wMhMIRUd910ydm/Eh6ZZl/gS8NY6E4dEz
XoZ4DsRO3zutC7A7yfVRubrY3nn+4Dl9YI8p8KXzSun72AVYQ0ah478lRZ/LtPrpKP4HWCxIr455
fg/RTAxg31UVbcKIDJDS+iS/fdb//fcAV6kQaiuj/CTmh6T7OBMqjnZUDIEqMFW0exgW8Riru5lh
t9m94e2QKWvq4mkbwE9mxJDb3x0wi0WjrkWoH0pZsO73/onVokI7h10Kuv+QgzB6hSEVWnO0Hgvy
ctjD5uYJ6gQYShMySDRXh8PpMUtBKOVKPa+zSjhsj8r4mQkyyx+PXPrg37s80MDjw+kbOM4BBP5M
/ICK6bmyRvijsaseNn4ah/4n3DwPQFov2bIBkr+ehmGS39rSGRIrAZv7vsSDTy8T36HKN9fR9rQN
JCGctIlZC0k7a9UCn+qANwK2getQSxv/RSXWOt77dz2FxAfmCSB2ZqMTvj4opddudjC2jS/21P8V
LDGnGm+gKU9Kz3jiszIaNYkfl8/4ShjrSvlkzp2kM9zJUTZyhoAtzOUev3KiHbca5S872o4ANnlD
VUiuvyLLuBTNytONIS0JoRfIqtV7KTEqniox8rvKjwzrXOlwf6gmWHelwO/aOR3iQkwdKlb3WGFp
P3I9hr/e8D0PQSWomXyFed2oenTc1dCBkJLrypEA5ymxfgUo7SVPtWSVj+qdfcXJrD2F9aN7rItm
qmATGiscgoXObRgEikjatsDxnplbDLNYlpFev3gPXAhE3Ejaji4I0zRRcD34N0USZV1JRmFMhPrh
bOXMCPf6rPUmeh2NAWpyIDwkcK2iJTYQ+rmr1qU7MJd7ORAzU18fNp2oNR8MvJT+Ca6nQDPVBrz8
vNtJfDbt4QdOd+1mVdlYnGyjD4hlp666lXhov5ErCZaRmp4W5gRYAGln6i16qcRfMjvKvNgJFxOW
wrx3XYkdbQgX5X9v0q/vF6onfqC71LYXypuZaZZ6XAJSRltytcg9uWxVu/ATbBGUyIkQhRPnWtmc
i5w6gU24yhuAQBKvPbYu5wCkzldMGobsb2eoST0oN3cHUFZ3kMG7IL7QpjaJaDWhgFzl1bkjS71+
Rrm9dKDSfHfo+6fbkiHP7sfJvmeIrBzK5mRpCWUVPw3ytLUWhESPBL6lFpaG9Q6JqOA5nNYT0a++
9VZGvC9++O5aCk0aPOYtHLLy+vrHJiPJ1cdYI05hPlXzRROKF2E+IyXHGOvp1TDQs/x63u5/GtUK
TCirIVwy0S4+nUgf9Ryljo0Xdc8sPg3otn5S5gjI4/oHLrSmhJLqEL/M6GCbRygu3DxuBFZ+a/Dm
ShI8CR6Q5nruRFELtsjEaKRBQ2dDjzYs+NoRBSQBmvxhwWK2w4iZyXpOa/u40fxoFmKQc1aHrAiJ
vER/b3vxG7cbZ+3c6SsXm4kIxhSII6EL1bFk4+9cbggw3CL1qj1/e96Zqfna6N1C/PtBAN4ZOaHF
NsN2e98fL3+9eYDn8jPnB3dOxWncxKo3Oqb/VSjqHBciGY8uUGQdDuqOdseQWsUpYtxwUo/Kfl+c
Q41bbOYhXhv4OlInRkix1zQy8OzZsad9ystgWQkJN1R84G9Xf3bhLDZkjW/z9igApis1Gdw77bvi
Rqw9757+zDuTz+NBdhnQTmFxsUosFCsQzCI1cVzFPSgHnzpXG7aAQrDJlymE9fpvgHOARw11z2Gz
GPNfFNbw7ZaTsCIeq996aWDWYK1vc9oTJLK5SZqzw+HkqR0ooPY0U7tQgwYuM3PXcSVmFaQyVdey
B9GXcgUKJMIZhzjIH4oOPUTJk0r8qg3tc76rLWsjjhUiZEutiFDZlogCB98r9rdljMgfDsjMRpRg
6kqx0NO+z2llQviindCBKlmKr5vrUHvxTowXmqpMLGlUcHJEUCrivE7gbYrqZsQOcViEu43ThxCL
TVb71erTKI63h1JlXSfVhZ4eapH74+1o9p+VTqjckOJhUGAx9NnIzihlv8nFS/jjsmzYIhPCXPmh
G+ts8pU9xkyTb4AxqPyejYC5eFhDu6WLPVDcpoj3Ax7jrHSLUKOHH17/eFQUTZGgx9pw8pJMxWv9
iW4Y+jSkmN3Tf5TL9xFT9UMGHLbUOsIlFBQ5KKTszBCAJNQ5xqwiasGSSprKTkJT11vRwUmB3jED
+L33T2M20FNprOjcy+38Aso3U/BKdfNegoOkbK3m4BJzm3IkJN5anJP4Fh8JrRWf6bIkO+Arqtzm
5hKZJBnGuv1PkXahPupPMdo6u7wWFeivPzaeg/xJJBfyooeh2n0Uezei9edNOkWaowAwuViOlQZp
bPNT8zB4f3n2hdx0EEsBqaPaxqLyh9tzgL0o1WtOwbMh9x5XQW0OOMB7fuVXPc4jALEq/7PCDkFW
zSxdSfv+VDp05wM8pabOF4GY/2IxoYw8fCUKEkOqGJ81aFSiCpvvCT1APCYKOKKuaF03ke5teJFz
FbxFxLscr8ULwcPXY2iQT00a78hy5knqs6WNUPpFHiDGMa/u1NlLpq4aKuHEFPFn2oi6KxUnNpTW
ZF9T2efVph5s31mmRXpRMTs7QavfLja6DdgWitkLtJMciSLg3Z+HVSnOv6n3+KStLrhvHivIoIvx
9hAnRUkOTy/U4ekAyHQVQ2eXpzz8fzXYXzMkmc0fi8ToN7vovn83kj2yBOTMiW4rnuaKzES6LPYn
7cFUB+6Out/exrnA2Uk/sIr/31H+ne/ujH0II9FCOx626hWRKuOTPPVQ22nf6WEPZpkdy5rkuSkT
cKvx3asGwdAO+YI96Xk/sa2YZ5rGezxnf4cvCqjbww1usTaOVazAY4QLLa3bOZF5j7ptJXSt79jq
luwx5UhBCCUHMT2UWzgwVXCuw/sMygXFQkzPXelP4pwOK5AAp+dlAKkDaQEmhacZgdI9ms87G/52
fZyP7gjmjxOxJcSxEUx3gHSmQTYzWp33Ch5e612LXImXyUALY+ypLJ/CR6e63o8CaREZrXQsnL6C
MfxJYpTylZLWNKalDNMuB9z/MAZK7wExfFVIp19QHPzdYRH/t8wXAm+ZkL54YfsN3OwTLjqSEj+a
8G56dWTioxson/Y372JHDILrxoMZOVlyDz58Kw4gj0lMEjljubD3m5430kbyhjz5QjnygXDdFZZs
mE+ULgNtGhCj5tWeNmX+Vbn94SJQpsxPVMTRzm/b0Lx8vjMgv4cCDh9Du+GqAXsQi87SGpxB/gjq
Gp/duhq6/hkJyxbOLeJXGYqn3lJYE5pdJeRF4LG+rEtPmtGVdAQ09M55abiCVkATzuseBfEHtnp0
CNY0tE9duMrXkkPJGlBGZ6Edd0k9DIGpEj6CdQVWS2iPPhWVGBx5MSKQ4i0rv/eeUAnjI/sSKO1o
adwA2tS0DlRRbgfXEhnbVMOwiMm77K88HaTRwAQfj+dS7Q31O5FKzLmQdDYbDXoEhsZE/mQr/ngd
utnPEFQjEe/BcwjRvV4/1zgS9sVhDt82ChG/80bNvUqggbTNxA9Ql9pg+TMyLpiYnllHKzjDT2qb
5tcaKwoQ1fD3pb8r/T/4YWXlmRUaO8g/PQLFqJsDtrUX6BQXfLhCVesdngmq+xTjZFKnRxRDdiI8
csWjuM6d4sOInYnJHt9P+u0M9IBXaCYYpbBpmOtgMBXexrtBWzuKNjbzdqOZ1xtfe5PzqWaJybWv
RYGxVSK4uF35yVC94avI3oolz1/s+lT+4a42/f/qn8Tt1lipA3mGfKUYKKaGrLT2xdp/RmGe0k7L
FDZIHHX2hLMK75EYjB6hSeq0zawiddBTdk3iFLQydP4E9nAvS03LtLGsUimIyJbW6oHpvTKCSYEG
UI2xESTB7qIQ15DJFDX1EHbEhr8F9trgaWeRSE897fEKRO5BsQ6jTmzD0paTKXX9XJ+GBFfE4h7F
RkNGueir8sq+kz+VATNDqc0UIqu+mqaV0slajKMNWGgFhTS8YFeW29InQ3pe/nSOpBPzVvHp22CH
3Hk41scdnex1by+Y9dD7FjoCfWqcIj8qfg261kuFjPfcOidjhz+qLDanEX3IyU1wtmrdPdNhOC75
3hJe+OOCORmVcKD94aSH4FEKOsD+Rn2etmSvPWj39SKkGnUi8paf19YZ2dK78rnC5QDAtK76BFqe
zsh50+5rYjmPIrhel00NimPSUK2BbsYkH+JBwsq3/Y7TSLr2yiVQpepB6HP3I8W8iLHeUdYOQ1PL
HjMu8k9tEzasyVLBoiCEbATxmPQbmH9m6gA55DRUGscxei/qorTHU75rsbJkAQ8arhK4ufZQoKAu
MZzaZHcNb5unSCKysSxRDAtaNKqR95OgnE1PMWvcptwQjUc9qJmLKtCa1nAPdqV6BVm5S+NneNAa
Y7RfhFNEc4kFvF6mTRuergzHr0ZtST2vvH0xXei6mTD6jdG/X6rKcPh5T8uvteJwMZIKw9x12tKA
GqWJVnYWfQFIcX5ajbGM+HK2eoDFi3TPWRxIznTqr6chDTbEWeP81zHFaBjyGjN7e4uX64w3MWx+
Hy6ddLgaZHWhzWvVLvJHupMnTf5ni5oooHzTlkvQv743k7NhItbsrd57QO6aC/QcVq0Cdm6ICWdg
B1EreX5FDRZrUS7r04Sp4eHA7nLZ5Sq2oVdNnsr0Pwdu3VFWAYLX+qx3IOjtBxPn+cWmgLKlpzY0
cuJ/XFDC13sebsvRg2zKl7rLhoEWGk5vrg7HVGhpNbJBIxb/ZYn0pzMFj6MmcbE6oYUorEgwwOQR
4vlqiAiuHwD6hkVpeBkstH09uKdMBrA1qM5HtU8EByjswOtFOr8Ot0pX45JlZ8WHzSys71Rcp/c7
P+3EOKywMlYLEmMwy405//O/X2m/pJZWgwlujPG63UF7jckSfdhtlxTJqipjBDZLFhftNI4gFJP9
RUelJIbY5liTWn1bFV3nVF4o00BJDl/J0eehJckDyem9UnjWVTmh2wULnUu69WvPzOLZTuBYxDJ3
/CAKOUocvOiTxI0SL8tnk1rFaM10HccW2Awf6hpt4emViFoud+idf9PGoxiSbJwo6682eM3w0YFw
ISVE78f/uH5fcjuSpwRL0ysE0LbH101gZeLMhTwSkINZ4D5JeBrz3nxaO6HNf1mRO+1tkXE1QHTa
QSR0UIypVYEmhhNlK4CBjqrP8SgPl7OM6JSyJa2QU70yrIQWT+IihW3A9fg66hcPLQGyhxA9Ngzu
a/mO2bgw4Tvc8xRN3oHaUo9v8PKKun3l73FCt3X1wAe2cCZFmE2R1I5ZnEzCyMUEOJFRI1UEoK5J
fiJgviDsgzJz0uT5etG0Cq87wy0jPcIwLj2SeIsQddbEziUXEAJxLLUFZj8uFXtbeETWXk67dznM
i/FWJMOTdVZsda1UaWfcl0KrfNaCC/AlUGwI+5OFh8PL3qvMQof1qTaBpOzURWP7zDqbcIkmqk5o
6Dxyv7WFLr+vaINW8gjEP59pkB2R8RdZKT+3XgBTkQHdCH7dcEKst6tA//GVpVr7nCGkj/C0401R
F68amJVBFNO26N69NR7Ah4fOXLTsfU17r9kN0Jam+y8vGRTE56/Q4IB6tSFjoL2JQ6Ij2Sm9DRXh
qOkVOOQmpAmOP24Ayo7/0bPhoRcpngLwlrzIyK/IpOZAq2syJbv79Mlb6udNZiJ231nHaJ+S/HFE
YbC6VHe4BDcNGCNzVsc/NQQxP2xaSe9cERM+7hbx7DwWCtYuvbBANARuiuT55kjlV+vMG0jZ0+o+
fzryiS+foSXOZYBo5jZEu9c+X+HuDAj9CBmieyMXCZAre3MwB004ZvMNBWeY7PscQeWjpC5q4NIh
aPGEZIvXmcFsa4euKrVXI2QMgZT3uODyrxGhRXgyuBZ1nkeWEJ50VFEk3KovRjOFEJWR7oLEqwQj
+sSxbretk62BD6zKxYRWdHc+vyl7hl9+ZWVz1ZbM7I2D4sD/S2l3pMbEkN1aYow4Bvb7U/mOj7Pq
x/lh77oHIOma3RcpE2os3iBCnGN1/A3WrOpuccxLFKDXy9b81hv2SIyByC/Qgy9csKAkompNQoeT
ElDovkKyvEUw1b3BhXgKM8A/SqQAL8Q1EUESS3di8gK/Ws7ORAnKW3ULZ6eDjebU+ayfDhDt3Wbe
6uiefUui7mIJ2lPVBiblfvxq+xXEIzgpQ+lHekazane/HSpcL/qkE2CS9EMTgcVmsVsASEzATX6Y
gunOjSMsIFYnYc72hcnp4Zb2KHcSV06okNithjgwNUh3a1r1c616hJn44aZxVvUtLXdw749Z/Q8P
CuRk3aPkEeNyrZBDutd4oeZxCozJhczq9imelqML6D7uW8euqrRVHXGZtHnIqvlnURxBV/C3qcYB
oQAx2EqqTUXfsedlvZPi2IMpuckgD4tZg3bxWzbzFuJIeG3dYqnlmiAZWC9MZRj1Uu/Al0fjNUPV
4sDlzUXyWzrDfnvYUdzVCYvMOvrjCCwmDjP+/DNSGu72D8oGXbzYXp23OdSL6I4LHDuEDmb9Mdzf
qGPq/b7VmOhawaEdnjADdmnNgUn5LgvxAe/GQlZw3kVkMrHv59XTT1QwM5+S4Kn72PM5ROgALOgc
bZ2I0LKkAZoM8eWXfR43wnXtikDRzm2GDEj+agrwKlHJJTMfyfM8BdNA0IJgarN9319NsXYadM+4
LBnjIQ3uF2gLk8tZz/zupvc+aaSqiN2KuA3lJLF+pvXWWEbeKaarNLuX/ddqwXFrpvOud7wvz428
zH5N7Fju3wPed7j1LXG3rbq+gmgyZLMO1bD0pnfbWEixWiR3e+F9bOk0S8y98V9MTPDgRaProDcN
rONPPGHwMmXAxQ3Y1eAedb+hbBASIJ0w47VA3nl3Hd9OR9ND9NqXBccefHe449/aXwL2jLzhbDxQ
nBqonLWafOV228JqeNdCN99rgSFDA5whn9UG2ar6W+1CfieMNcY/PBCaGHYC1vuTFSuyEg6EJPn1
ozifYrbR5bW1USOy0wqvcqUsTYcZxlZpY1TFmifQTTv8VSc77ZX1KzybU3EL2LllWqguFis65g3g
ae0ojfpCYNjrNHgU7Iv3491wC/YDEtR31p+ofaFdmAf7CV8ai88M2XOSanQ950q7VevqOrD94Lh/
qlUEf9Pt32nGJ5Qt7IWb1GPWY6h39vTpg9vArIEcJiR8fBCBHK8RunNzrrd9NU+HG3a5iWLx/PNL
81lz8HoYh+RWd7FcpcPDe3QAaT4ngJ2Mr6aGbqu0BW1FxukHGEeoReSVPP0SSykVMR+YRNUHyYCU
j0o5Ac/Lt/Hj+9KxPNL+5n22K2pRkfGyZ/Q0d0DdRhClAvKXD7V/mItkmV1wtbmPP1wpCT1Lp8uS
DioGl1G8ppO76FJ2d7UnnZGuWF5EVSoEXtny7zae3auXDThAZPZQnBLhmG+qtB2qkdIxXw/3xr1x
U2ECfhf34HdZAGaK/drB34rpOnudzbnrNZx+V8PBlIplcA4PZOdyG+HaF6irNpEFdb3uGlccTJ0+
nw1EV/kt3keIW6fOXTOloK1kJdPd9bm0N36uJtBPirgOGOnMjbP2ugdt7iQdHNR4geCtnjfhh9IW
GrrHgnUQ5/JyJlK+zVuWPLpsNX2XHYDfugLvIm+iIWd3XTZTKaKKQFOBsVQlMdn4wZfcUrqJeIsi
oV0Cpsm8r0kwH6y8O/ldXGbQQDKSlV86dkQSyc30QD4TJgZCC9yTRbwaAHazCMFhofk7kAFYYHEK
kWDT9jX8/R0b/aB7ZydK1/H+KPikdxVsTnKQcZq/lO2cKh4e9x9jTrx04l2hyPM2lUXM/mYtv8Pq
Z95ow9/1s4wBWPt4f7k0cddNIf3pXxwMhRSeTWXFyWU808XKekR62mFrHgSbtWwS56VI5k0cD3O9
Gt3cjDvOl2n9kUOZyApEvINhtBzrt+nw20VXHcGjvEd1e/boYo0zSA77EV2y7m5CPYxpvXCX1fN5
TPzI598juv95vU0JI1BtdRvEGmsPZsGZWAuQXfKuYdT1gJSFdeiiPnCQdfRyklpRpa0cYH/vd8Lk
n4y9enZDmDJC7Q4F+kJAhcqkF0DS6kFOWy+bbyphjd6ZprjmQJk3tDM7bYPEVSmMIPK/GcSckX8F
KvxWRkqXfroCwGoDgka0lklraPhC5lKTXu6lXqs55sdGSYa3oV+N/jDWAXRRRBLZaOC4jquAOXVG
/kY1hGq2MNn84EQdvX/nvWEmI5++hqjXb45x93v7pj9deECVV4NtP4QPhvE4b9XO6elxuGpMC7v+
imKh05mu10I+Rguq/Jb7Z0chSqTxKH+O2JROHYbpnY3h/U0VmyO4Ih0mv8qGjz+q72iDvtUZ5DqP
I7oNLXCnssm0nTif1kLKPL9rJDWHVErGWn7jYFL6lovzcgE/6QV0oUIKfr7OLyBTwBQ5E286+JPg
KtKFzVd0cTcu8m5j//StUDmGhxd5nLxTk48twUfT//V0QUauziCxU8Bni9qlX+YtfaaAMMQq6FIv
I0EHcwsgBCn0Qvf3R3/6gaS0w0cYQ8HeS0RJpreWsQJQrJS+n7WIC58fdqYHewqtZWVTdwrLjBhe
ru9gG/86gRqYTMA8xHZ7GHM8IvII67C8MyAJ8nieUalZDBN1IWvKuEwgEjfFgfqTZq4rCtNjMRKF
6f5uo9Fdxt419z1X2ccvLBzAFlffhm4uPokVggIuANxJRVAmssn9WlUxqh0AEJcPtyklhqPBa677
IqQd+yBkU3rmadd02nccxRqGbVcavIiBDy+qnyD1DawGGGVNlokyUsVRpGzdMkw0PNZ/tcpj0X+m
ZbDs1fkgw+mmqoz0m0fOR3AvcrzTJw9mo6KHR3n3iP0DFUxB+Wha9pl9JOpVEp6+B9FMgA5XhMUA
utq6+Z5+Up+hKymXJrVLzTfuNkO9xluVMFeazlr42kVPx2OfE2k/If2uhHkb53DGYsUGM8IdFid0
fo9E47wLX8KP7PvtSYkFfLn9D6vi7dcP4PfvrtoXpAWaiwxGXNA/XbPPY1LY1pfA7YUgbVUUPqzD
AkDpzwGN9LaOAIf/WDIhp+LwTwgB98XAZ7jvb4ykxz409NDgH8xm00z5m4ZBJHcANZCBlT9mVHVW
s7q6tJUfigqWhCBVmWBxF/Rnckjj7Uxeh+G9a7JAtXg/yMhSJw/yuqPwjLiKY3etDihWEOtyDOgu
N3WrYDDgS4b3ahb9DeIzggVbrv4UdSvS3uNbMFAkhNO5TGkw0Ol7lBsysf7bMajynBoINYUPgPvy
G1txsdGD8nx0+98l+aiLMAGATbzx2Njxc9sF6K6OYFjApg/K1uIClQagtuItLARoJpxMbcBGFoEy
O1j5Bnz64rjTAG34tScFyXOB8h4vCSVFsT4zNrn3mKxWpalquEELmnSVfpW4Rjs9HOdzifYa6jWY
LJOiHP2vqLADmBjkdJdn2/sSV6eOhKCZQN/eBdezwM777/dSArHu9TeUSPRWc9RZepTmq//v3NC/
s6gBx6FXGqEMbnwQ21gn5svGdYzF2k/bStYnu14Shfum+o4VDSGN5TMI17qvovFUOCjvrzIoZXiP
abH/sbXbA1k94nloXs4cgqisqxd3wSipL1/i3MklRZtsr7wtqKY7olc7hyOap5yp/YpwRkRnpTre
taRPrW4eI7AGCQy/nkheWTKgWBcBu8+VLjIadRCUIPUBmOBluL34Sz55pXDyIW6Sa0y3u9ZyugNC
Jlt6F5tUXmLxvNW/QelxhQN7liALkI27dr2sQ0ZOO6aGlbCPbeJZdKz/qx3P/1OHg4ZKJ6ivoW3d
bf0PIiOFXVLo8oA6g7fSXGORGVj2DszwZa0g9Nd+FYk2eKF2ukc4exaX27KgXjCxk0axYsmsOAe7
xJ+yjfPLMSv9UjW+Dd7gJqGA1TJWVu5n2Bb35kaE74mQlhkAXLdqiwpD9z9nJVeP4udbNFYZWaDQ
LkNZCSk5Tmr1wZwL7Qb6leRX0cOm6Z4/T5W9/hY4c3nZzeycnujXVwbP5anVa31p96b/PQoGwpkg
otGNAIU0JBFptUzBjptu3ixRVugBJVjUTh2qb4snhEfe4YbR6Yxp4VnI+ocyZMSMo78l4xXWa9Hg
LCluZQk0Qen9yjjP2r4MvAl+JZmJxOLf/hZxCf/M1JUsWBc+qAer5hA8ainxYveLgvbkriEKspXO
3kABbqVz2oVk9x5Mjv7DIkS+NiW4eO62oE4LAzpjqC+xxyVqJMYVHHYB99cqQNnVqcP1R+wY/LEC
bDPfd+EHjgv3gvHMbOQfAyyQGJz1G64cIcLKL3ynFdx1wuxUPVoSlSziuT5/9ONeESKyJZUv+hRJ
qSO5eo3Q7s3xw10+DFPb7yOw4+s3fDbv2ZpWW+R0CiTtoAXyCgzPv6sZY7cUbV5VFy3g78chrfmv
+/Qf1OWW5UVMRxbvVLj9KuhCNkyWbweVaEpUs79jrp1hCIECMkTA32Tdo2IK3XSSgZnDhbsl1Q3d
lPdKBuRQ2+IchuxANctieS9V0iA3OElp12DSu25n2lvKjwGyPlP48sj/+jed9J6z80reT5XI04WT
6f7+fVm80v9+ISA6UOVxQgxP/CGPZ4kvoXpR3RjlujK5E/6KDNnNEOjBLbZDEJPZqDCW90eL1V8S
A9GubvGeEsbBDK+JzI5p4d5TF6hk+5h+DJW+4c+CiMIzU+e5Va98p0QPuBXFhCliI0B7qvrymBV6
j4okSeXnPwZHGkmJs/bjzQZHsD5QmV4XwgJwo78y0WcKnXTNPOBfSc1Bo9de6WLwYNxjwWNXpzRH
kQdzjVR6ax5ku4c1JJu++wR3stsAoa+ok8OA2Zcz+siGK0mv4zlYeRnpWNYREhvAeoblGNxFi0tw
2BSCS6ugG/k24wiEme8khu5j0kDLAspAF38+MxjB8FmVs0hYKRWWkLqI+Dxp/KiDMvcnaeqXcTnq
Sx6r8pc1vHnDcSIoroAdtHaxwkiBatVQMDhcVCBzacIuA1+fr0q3lYgZGZTIRPY1dGh0wcYHSXv1
AbGjF0xv7WDhyZUPRNhPYhYF+bJXlQ1byCOeaTE2tYAJL/XOzben5GrQDw4lMYU45HWoVJTc3Zze
mzt9EGVx1tySPMonITDrHS8QxNv9YaT+Xpw3MBd3j5PyUMnopYNj7c4n76wdoJd05JdnyiZW8QtG
r2hsLc3zJgQTVF++bMQUyxPvq9Y6BcBqI/zKMMPLeq7Y0ha3yNiOtEd2NcH5XqZihtyIrYd3yHhf
35RmpRP9PyMAeKyN8mnYM4cU5EbyBAXEwPoJMKl7SRfIXowkBicIYPZMDmSD6Mm9K/ihN12adAts
ma+A1HdntNhkd4lxu2tF9uAfJCRtdQ1ICT0xR2ZjcXogJTi0IQtbYwrxTBxBZf5+lcdvdY682ceZ
SQApMYjz6EabRGJmmIowJsznfwsoAbk76N+aT/tsDKdvIXoriHjiC8+JdQoRV0lydvmxbXQlnzJy
yzjj2w5XMEr/Xwo3fh6Q5lTy+7kL2QU5NyrJmcn5wUNwG3FJ/9RTwUuPxTlJ+L5JzAhoUjJsqY4n
Xnm+Rz5WKHzTGvw0xtAQqA7LcGspKkWFWyFmas+cveARVu9qLtmIPsAzzPCovLwVDOuLGhezI0Eq
+/APQ7TQo5sdT5Znni4+zLI4XC9ivP+gl7tRNU0UNwPOeV8+XcM2uvpbX94mnQI+ZV93a7Kkcz90
hETuEVeS5O4fX2dVnBGireuQJx5BYfaMC3KgmOCG7bkN9kwRg1emmHZRRtqOyNI16xz9lhKK8ILZ
7z4x1ZLNIP302Uos2zTSHqiFYY1bhlNCttD+JQcD6QZPgNKS23xBC0IF5rgvMxKOc3zDj7PvpAKE
GuC9DGzx4TUWauG0N9Ngq17vtPP9EkoHV1n4L7f4NEiuMmbQo/FmWe4wvp8jMUQ5OTZbQSCK5DtS
BRgxFJ0dVH4B0VCuChQ6jtiJCpvlyHXgpmrPNEteBpqt/SsJz0JBQeyJBDckikWskJ58FATrzItE
ShsR59OHfBg54FLY9iKOlbtyJ0YTSgClimgCTh+8Ggo4I7T0m8G1WS3aEmHirzc0OxZiD16SUWkm
onzAWnGTKiGKhFnHuHy/4eaQWk8Ox5YOFCG0EGYtQ5aJKqUbS2ynMLbmDco1fwce+rVKltIitR14
dFLs1XyuwAhui+4hDgUiUL3NzaQYCfvRkoJbD4s4KnLJdMmOuPVr0ypwdq+bNnyVElDjxZ/iKtBf
rwPtpQZhPd+BZ07w7XCYlI2R1KrAp4RIa0pB21nlzMoRMTM+Mn8PzhrG/g9U77R4BYoTMTMttGMO
FyDtrd5uVpcBHoRrhfwsawbdSIHhTQkl7oNGVe5in8DDRJJHr1gDIKIaW8/EGV49AwIbKfYHEtWL
9H1DvhGFdqIRoQmFFRxwdTgyZuhSaccdw4E3L2Z1iRVUSDL+Wd8NM1/Xlqx+m0sEnu5hkWXAFifl
tYG1WHQHB3sMRWdCxmyBFAJcV4CM9o++XRAkhNk8v4V7mVp91bQPCTZoUqqswcBpBFdJCBLRCxyj
36iNL+FTgnSwRuG9ingMsdr3//ZyQGsbGpeZkm9efHqsABWa0Ep5Ufy+f9XId+mm1SeIUn2HhcTW
z3bvBUYZr2/bFVHw8Gs+w5VdTOteELsRFyrb+5VTyrZDkvA0WikM3R3G6dX1FNHqgZ4UM0/4tKzr
jFFMwGxcrSvmt7Nl0cOXAGvoJXNmwXe+4jQVB+gkwT7l+xWr5cLZo8qoDJInReI504kguvTss4Rg
t1PWtTCZ7f0niN8GoKWK6GppxHv0Pk2HbSQv5dulIWRolQI2NlE01rCxpaYaLYJn7zz6OrtSxvIB
yaQGBvP+sOm3zVYsG3Q6P3sjuDlJgMJ4K3Vuc02yD/goAAkCDGX7++2EsWiYQspqwIkduACAzWrH
/99wGdiHbKURyVSCzrSBr3q7bDw8EwcSQrHQ6HLsn7HrxAscB/j2xo2J0ZDHgr2PgAES+61Nh3P8
262siYVLNgRN/T+tDkAhQKHgziOorzEU0AF2r2Z/9ozqXqSv0MQJ5vqemBuQRomY5QW3kzR/QzET
n3cixx4JZ3wUQWZHYPBsk2Lvz5AmEpMRXinjRamugJ7W80lVG8xoTZGB+dWklhMkFd2aqk3nTMVm
59YTliUSH9fjthMtNc1MCx/cITn5g8uRX5M6NGlRDAjgdwNBszh4V5IqMeYMYVCr7FT960pBIgMZ
c2IumiWQ2CdvIEsB0KwSM4ShdQjqwhzJ4Ygf6mGycokoBZALXqYU6IGHmOAlAee6IF/YBT5QzOSE
DOrPMHGblGzyupemQXB7FkQNIOIzZrY2Q8q0DK+3DQ4kWvWrMx6Ssq9ubnnT3afBcXlByxWozkZj
ILaax/HzA1r6cnAp/N9vh+tAld4g/zP6OtU+WJS2BdxsBJruEprvcm5yrIhZXfjg8w9o1Qph52gw
HFEHLI8dQPPJ2OFjR1t6UBblZ6Gy5jJ2fgxgUIiITxg9BbuIOEWLyjl0Oh/t+QTGvDz76Byom8Xr
gj5+f7dDCSdIGclco3gWotmzsLto4kgYDTchl6QdlgtoPs13PNZaulg5sgr97uarvURfph4FFs0B
uwhdx7vTx4E9aF+XsvAvayQ7cNOYrs3NESGJ+Qnk2j+F+cMT+U3zGLtvWmQu5l1BgOPXg2vBXQA/
nx85fxHBMLbrk/OgT9320O6oMAgSf1SnSLdFSYt8AwGq8/1aN4L897l7s9W8WMpWSaWl0IrtLeMn
eLZWNldhOJDE6+yusITWQmg20QMaGDE0PdZoFf8dpF5R9A+Bk+JLgrsM5VbDkBowFzALvJR90nFp
rYPirWW/RQSLMwW3zH7JayzA54EAqOP2eDik5DonX6VtzRuAay4VawHd9Z4IU0rli+HWUPTTeR/g
/5nQBzoqXcced6uqGY0Osb1RuSWK4HW1w+P5ZkPZsuO7mmJ9ww8ylUqOu6DxzFlCNmY0gY43TJL6
QZF5gvE558hQ6509fVTePxV3T8Kuv1RPtWHKRfi8Gv3rdgjgPuQcBvUoI5PxvK0k/EIIVLjFlyzT
E5cYvLUY5aKuJheU34LzFU2uLkPkdz9urZvG1dL0nnAtlDKLZA3f4PBm57HwQkaQEHGw6Z6H0sbe
nDYuFDaM3i5pQuU0Kip/xU8IODhCiwwzG+6qdwvy65u0OlOoh7t5jaiBs1ElmLf+fCI4VB38gS6l
whsHqXH39DS+uD/EE91AhVusd1pHTRvI6HQUyzFQ1IRFhPlMMaQtmJilhbL2LBbopAZualFwFIAe
BMq4oWR1WOTn8EfhL/vOP/EHgD8xGuM6+o4OceUk9crO6CrCD7bEm/HD4UzA4tnpmXEhvaK2qZrx
ZxYO5JPS4VwVFo5LWEFnnhvbTysNZZ0/sjV5cXv5d9tgjmUJOSuLQtMVssKwekQ83dGVSEBVO7WF
H0qfUu8T1PMl5vUTBfKefuqmc2ZJTwmhXIm1QZOrdJEHMcShC1nveoQA3SOrN7qpwF9kPk5XsXOo
G+rOGeIgqz1kIQlsAA9j+bZ7HywEvTbyMQ6/SKpj1Rm6tK5U3Chkv6TzOABwKvb2ua3wIFopPVB4
gh79d2hTQCdK3KjLLgF6KCmnjaU8wfGtTyRgpDj8J/+STkcuHB0EiqLpsT0ny59OBHf9w7YzrPYA
9lCVxsX6Z7j3wNbiHt65JrcQL4mWcqnp9GoM83ue7OKNbFfSXxACAClW4oea7BDyQnTaFDGGV5P/
pvbr+XNODRL1SHXjYEfjAHIS5n9KtKNFR5hEN8Pna8NGsXtQweuIHz45hB3EWJzlgLbUIXN/nKGB
nT1UlmmtE4LliVBqBwm1+6VjAqYdTok7RuOm8FbFtKaUJRCAsDZsbryM5eBra1rUUzhnLyhLyRbx
fTJaTXvMaYj4LHy19jdW0d2YFzoW1ctYTobs8fY3NMKIsJvRr3UaFVFHBdmiaKSBF5NrIt/Y5U2r
Yem11GqfoUx6pFNc5hMjTp9GuBoXceecw6JI1hWX64E3tzdExkrl/gZbxZA07np3JMqXUfeDMl2D
yDv/i2k2041AWTmSMIKOc6jdyq6mxZAmtsB+JzQCV8kWmS61ZRw8bkLrUkUfNv795Z1/1f9mpK5s
PsNBmK0viO7LnIBeVntJTz1sZHD0YlliTmLraOyUM8BUneexfupiGgCNuJOLDj9kenJ0BM0RDewW
efqmtnqM6/RQIhl2s5LQrnO9gb/xaP2xp7RXk+PFCmxkrfCX/Q5tv6AntPyOnLVviyU1iwk7bSi6
Xx+fgAEEar20IbkZB8V8o5hdVXZD/emypaAXDoBK97HgxHFNVH1RD4Vx5o3gtM60JpiswL1erwLA
aCqjfl0TJIJ8jVidjnKGqblqkn//+xOvltRQnPuHRWksRnl7ChkqK79lkKrCPJQNzVS5APL1GufL
komWduO9n7AMHq1m26RyrDFXpv1YewNTnZC3zE9F1pZnBAVqYvCBOLDU1LCT+YPs+iXd+O/PQd1u
dTZV3krXvMCwatpCjEBlY9HQ8frgtH7kZkG2uWWjQISDT3vvfwQyDmapvY9MVtyY/eE0guRylnJK
hIVfsN5VbtatNjrTjHU7AsS9t1sQ24tWjCAgvKfIyK1aG++rWgLtNVeaneI+RMdMyvQ19MbVTJ5n
ltZ8Xiyn/c+Xem0jsKxa5WhNofQ6Im7ezlE/xHP9oBtADcAvpaYebPie/XW2fY9iS44HyIJzZerf
UOoKn+a5czTBpEuIeCVvaJEACUr/WPZHZ1bUqaKb0Gq8p+FGR5dtCLAjOFX3w7P4V4MtkKwDJfi5
GEZ6afMlUj7wAzjhrWrSb1RU2GEmOKG0//kZTCOkuTbXJQAQiTu2KGCiMcGvRI/biu5+PkKvqIHh
Y+4xFT2lupS/NLNcw7RKkLVUQIqa26k2RjU+U3hihhZHjO3Pcoq4Cagy7rNehZ69mZjo3ZHJDxxO
MXsC/wE6gOLhy+AoTylG8hvvgJr2pWAw671C+XO/ceEQvKr2JOOM7ycqKzfwJVev6/xTOpgEwIZw
oJIFD2CYkN2KsLPGCN83p8mvF5othRJ+jHTSOsjYahKU+2llQF9vE70RYxS91kx2Yr1toI1+BKa0
eKM3JD8AEjvS5GXpV0/vb2OqfEyUnL2w025pq8dPF9oFMtA19YdSitu6f+gz0ArlppodZ8dhMRQG
CdCK/U3Z0dIj/R61FIVW0RXf/OzCIOFdr9PlKJHzcGERS3vMwVmXXx2T0qbG3xK7GoDi6w8p+Rjg
w/8JAlSJDFNcOI7QnVS01apn0Pny4QfeQH6Zj5nnnNPEeC3w9ZmAQ0cisVtkcmlSvQ1oh40U8+Wv
iPztmwk+xi8Xg4KsK7Cu1sPw2nb64pBxVTv5O2nwk9wYaeaWJbtB+zpvJTpf5FoukP2WIdGaFzJS
kq0VAtX79K5KTo58NhUtc7/v/pd48ka/fjNKuAK11u5lSm7Y1HsIiLjU/+m9jfrpQdfLujw39qY0
GPd3J+oj2fcz1pgi/AHS5d1ez9qVoCOm3ODCZr27Q4bUjfXtFVx4PEt9jlYZ9SAMmHN+83gagHJH
A8n2RtK/dFB0lBw5Ez1fEKtiASXmTjlsXHGa+/1O3HgYmJcBfyhkx66TZvbIvy2wbtY5OTSHbfoq
HIXXw7KKbfgmxJigsUiWxoJJZ57DoVZ6g0Qhv+TvdsErpMTrPEb/CIiudEfuMFMqvqcRnktYpSRz
asw2Jh1I9XQ1kASoE4yFcbiNdiaCAv7pwUNK4WQ8YKE8O56M1QhmkeR8AlQfLVHmFpJZNO3Ork6V
D/ujkc3QwDy6TchRg7MG3PWbCUeGWlszqI3lc4/rGEROuukI+ODN5/cFgHLT/1HBCWXtMyd918y8
bXEK1ugwUlCi0XnrepgvrxBFFbaqPxZ/t3UcyjBieyB1ZG/JsYDzI5oRQ7BE7p+KxrWTSStmN9Ss
5p3VboWA/3hOWLZMa2hTRxoDRkQ16e5FFKgo31hlx19YG3UaI6+qT2dZ3GdyzqhAoXPaXWxrYtmf
QpoIiBjuNrRGAK+0AF0aSeJjEgjvKeAleih1hqt6tUkhk/X69neA3mq2GZW8Bfgo0fzqImbkGC+F
0NlTl3bnFFkUB63mVlb5w0GGUL9JlDnwK8sL+zQ6wboPFHCOCjDJYOpxsbO5GLOE2yHl/+OCbI77
qcuHw6XO4/9fK+6VnHcRbQuzP2Lb8QgR0aeDK4jtypfsnC+8ODR8IaflKbkeGFAlEaHYvTZx77bq
uGCzp02fX91zBY6u3VA2PmF4SehR7XaStjCrSReAlJtPDWgwI3H8r52hB1PhymPTvK/OV2iYefnV
VahT4tVSeP9mBK1oTqVWhHcN/bPSOdxSyYFqsLJ+W/L8jceOV/Bxw9FwSAZHQ8/Q+eJJY1Uv4Fwb
1wPMTwAQMHf5Jt4qXnLNwxqyix4teFA6IKWm5re+mVirEDNr8U/MzI4NNPLLs3+IXbLrd7SjFRo9
I1C2+pH5v0vlcHEl6FCDPWWyFbWzQzqN5Nidco4rMN/fPUQ8UcItXcIdt6IpAuOWPSg2XmapVKaG
1wtcT+Sd7v6GZZx8XD9rgTOg5+zbQdpDw8E2PqA0A1xKed9HJhH8J2VO+X/NpV+wxLr6Z3jVu3Ac
zJZqcBovU7MJ3MXSqvBdAG35JlGzWVyKf3UIepMrW4dya5xggtpv0RRAGYtCj/U2PjFQv2oDHqoy
VMrs/KFfWsLh/h43n8OFgdFXPRpfHr/FHWcw8b6+ejiIIiXZ2hND2cIAyqKchshVdGFBoBa3XTXj
SPkoCUHxVrWeXUTPjujGiPyqxknrjhomONdAZXNYB0rfN5UhnIfGiFo7I1QJTv1NA8IgIYUWO4WK
lY9aRIbpt2FcN6RQN1rmrlFB/GGBaKz6v+KuJ+H7ksAxqDCv33zACAbUgY7hwbphABep7hr57cBU
Wxo76g1XeUb7DS1u+zbJD1CH8311vOKe3B8lGCzJnMGTuDJxX7L5bkqzzg2MooDQo5imDcbYw0OO
9vrRjDg45VD3MWy/nPiQMEZ7MExIlrUDYM48aPpMA915VfxNYZKWtCLHTXs8N1+WrP83KWrzqwrm
9lb2psBxUmddp8KJvcZProD/EMdUTpexJ7rjNNmlcR01PH7i5674i+8p2pgzJHuqryuQbKx3kSfR
PpoeGB0CWucHjzXEe9ZnxIf6ZJnitJxh4Z0rC1Rq9LmWJlggQp9bBMvt35mGe6/QKqTXdxLO9J3U
0GGWsYTYHFas1WTmI8OalnHG/PvYmCht6Tzm5PeOhLMJhfHnG8kJaM3eOxlNSbW1zctu+gDcRyhk
xnydkrvX+J1jE2PdUkkPuFcty/YZumb1fZ2J3NL/S/UnIw0tYE4waDN+lqtLrwBHFj3AVknXV1zs
3vwr03/q9pK11bLGeTV9pA6yBoBbk2J5OKJuLKJO9WHmOhr6gQacAtEB6NN8GIROP30G0IiAc9bG
fzZ4XPVdBfAEsvBArPbGmbhI+f8lz/01cqbiX3QTXkXMr40ZRNjnhNqAnS+NnigmOrUrt6CoDTyH
N/VEzsCYGzOkZVNfgk4c4Sh77ZY7ajuD9u5SgzfrfLt5LGm9bmbXKoxqC9RbO8NpESTrFwjeIKQy
2D4zzz8atOY+47nhF76fubuNpZRmGhCckB43VaYmIUVzDOXJn+GBowYcHjH+fKNWsZLMSoNJqidW
7c+K08GPHxmHi/3EJzLjgTfxcZSLQDzVu4Bsp0+828zJp0M9cPDyzy5LnUkONIVQIAdRW41A+G4s
T04E+inDd3lIpNfdnoinFOHN4XmeitltPPqCKbD4JTwYoQ3zEgko+Of+Sv4tWo6S3N+subsVW35g
f87BIZW52amar68tERMZikurrxtzul41HbrzbWZRM0lwLHTIlaFP70K38xYNJgnZDK4Mi91+E4Vp
5JmWTb6jwFPmNkhPZE79RIIlYvL5Up1Pzx21U7il+RlrYz7+3Et7Zh8jHiaTRBPc0fz7LOvVoCTG
egaUTbzVwfSytRsK5GM75ag8q1nlONSKnUHUlmXOY23MWO7Zv0js5f2sdj7+abkPDT28CaQXxk6v
L+Dtxn6K6Rq5592aJNyZPmdf1vsNgSkiCIlPSJwpo/4T6f8kiTlFYeg0ymzMMYFnhXVqQYbAk79V
HdZ3Gwb7R5FkcpFuVtTvvQx2Mor7xVUB4YhbGt4KqOhLJ3dqR8hw0yEJ+izqSD2oTGpK1KSs1lPZ
cCBWSbLQuD+srf25iFQZOxEZ/Q2FdJ+2EViAmXnkq0cfTNTUch9X0bAlu9bVnfsMNUJnkpM+oKEO
qTRBVO5VBX/7AZmlRXrIvk22TXqSH5CPLzobarbWhRpX5LAhm4w3u9h4sDdiNSr0/5b3oSc++H8n
mwJ2ZxFqsaK0o7ZAZi8UHKRc7sq7rH6QksHNDNjez4bjJyv9vDXxkXUtvAr2qZY5RKpoiz0DRDb7
A4IboGQGqmE97NJea4sFCmUTL/MNirBYZjwWRid7lLQsSO2VxU50GOUj9G9VA8PfRPa5K4RCR+uD
CTXnEdJV58lWk2ro2kWy2KxFyzShhG9Lq4eZx8fXH58wGi31vyYNUbxuTyC9SAmkfNGjhtTe0Ck5
1i5Td5tn8OQd2nN7T/o4vTqW+Nhxkh2L+cxqKzu23juQWpcs/T9eAwtumKdZ/P/xyeqv+5YPXSOI
DawTjgxyhsxdsMA1OE/ogWc7YxU01tA0HKU7n1XIOBiqRRR+x7kqHN5YAxzi4xwMHRUocgZhcXLA
0jINn1bPFDksL44vZgnZWyfxpSq8XT2MZRe6+M18dHmKNHno97y0n5a5ePfIuFMg/eHiWBEr8NmO
hycO90CCPzv7dKmH8m/iJzkaXJ1U6hotEjOL7Ud6HuIdbNquD51nb/LCYA2Py92mCT3imUB+BQ3Y
NI6YmSSm293GyHqVHHYCo5hDW3Grca1iznIy1PkU+6DwZgQVJby1cMLrRic1OnPalQNqHa9kfdzu
ZiEMGfmzh4nn7shDk1BtrPlYZepAaXAFzAJ1GN9Czs7g0rs/iQQNWc1FmsWGYDvFaoGPV+ppA97K
BEeYUQg3WBYUWds2I0EWmOkmO8mrKl+VJoxjSaPSAE9k2QpKYYzB1Ssn+3GrVqgBvcbXzUhri0Pd
XrKQuQ4mPIcjlJE6MU2x+jNp63idJklNNEBYP1EUClnZ3vKOcgJVbIHVWcoWVVc3KvyoMGVu6zYI
AUJmXg1bijxFLGzgXd7OWwnUrbTeyTgpgW11MkYj+4v8D4IjnmW5s6nEb9yCGnwyz7PGKoWhlfmN
J3MVNyaFRqge2A/2U07Hfp6KcG0BXRWrBTJfGk4A5IUJNpIt+vM5o6fw7z4qa4YWYA28Wts2ckA1
SHJSxkqJr5vWPyVoAxUgSwsUukiOkBxIdC8J6TShYDH3RcsbSwEpDJSTkr/XUc+53LccNn37pYGh
rLxnZdMFuuqyMXWPFVqYe2xdn0bJ6VfwraICTQKy9gwHvN+Y0i7pMa1cBEab5DOmZmkdztY4NFbf
L0A+95Est9pFiWg0KvchgIcq2XFE69AHDfGs98pVI1tf3AUrRDhriJfnoHEYxCIEP4tGx5i+vPEA
Twr3WFGAocoMtoKewsxqXdwBz/3jP+wCByZT4ouL0Ld7uwFOp9Nb085h/cTFpJ8fQm56JxrmqWPb
6r2NgHQ7iLfVf+It8vXy9qqpUizu5fceDnepjbJqnFBvfQBROKcStJyI8HZBfAZzrZh/gI73jt2c
VT3hdyfGaPc9JgY9m2ik68KTer4ovCetbVCork3HJ/pmOjxJJGYgvgSThRFsVQ/ZR7usJcvjJgZ2
HyleBId4+ZP2nKcoKrT8Kjo9sa8l8qxz527O29/5e5RmogKOGbP5kqKwV4i0Bfv4Q7tkkV5NN3aH
RX20EsfwBXShIVhj3qibz3R6bfQYPZ+YLKTVHcE6t8TEyv0QC/gz5QxBOR9a9B73huaroozh0/Kq
+EZWBKKP6V8B1LJY4F6iEuWamP/s6hE6h395W7JZtPAu5wbLPrgT+/bZqAn93DJdL9qtML2t1avO
OmUG8qdfNel9t+Np85tdJpatbhmyEcFiL3o61Qn9frXB3e6a4yrRglOdW+iAJa6/4MG/vNxv0Ydo
vbegtsSbkuuZhXxZRHdIHRmbmH3UFafftb8ifZLVODeVR2DtoLni/RXccvt1kwyUUstUhHARO7Uz
UIngv1y/M4IVmcQxhbn6sTB/HhkUDl6COSJQoFmla89Vei9Ub5JmeaWcIdCDGGI7oUWn6d3Eqio2
4Ie05aJO9EGXTD5GGucMD4LMx2dMF5qCIWTaM3p8z0R+2xrA3/93vh9GQfoqJV3JwPtvaa6+3XUm
GFRDpOIzfWUzBt1Vn8tgtgDrKafQqrMX/Ufkl7KpLuqlZdnfCl9Gh/6ePaRVC+iUAXl2IHlUHsiw
a9PT3s48yNdIzuLKMrA+dl9a/XY0jnb8F/MdfcAoaYwUwm7FTddG0HuyXbikJfyfuyOe/Uuap707
luRxZHK/c5Uwaxm9T8f3znX4ZPJDJcVX5KI1p4IvpeNBBbRoSikgZlNSc51+xyKSCUYpyfhmaRlX
67VyIWQhYJDnZDAto8YR7s9YUUYHXjc3ur5vA/PVynnGK13oqH6GSDpc+OVpnjyNCS67FuKa3Ylm
k3qy/JADmLAc0zbNcuvjMF1eFOAK9l4zFdIQTXnZdxnVWQyRvfU1dhlYkH3T18f323+r2f87fpjK
1l1vvXvWsxhPRiryxD3rS5n867ZbJHF/pk6WoQmXt78nO8rWXwMdHi5Fiu3mpAGJtHpLRdjrahhL
qfSobTZzKw2DDeAVxJjnw9WaB+1KynWNeKEP4Z5TSx4IpVZEl3MRpeFWpjGAXw0t/AqchSroVay/
vGtiYEA4hlAv2quwerafpfcJU+mBka3tV1ncBxGeYd67QqQBMvv/j+RxFGWm0CGoaRpsEgctL1e+
XKrmNu8XQ1yWBT1wO1ne/0m+JMlXIcFuP3mNkyG6/e0r1wrRHUgZsHNMChsykxRvE6aOss+A2MdB
kbiPY2oJvPb191/CB/28PSIMSy4MR9olTlNyh3vPWRC5I0QIE6O+0vCEysqNlp2Rb5IY5UW4Oopi
yhii9x6kfcLm0TLvouOx51lp6rb0EO5FXLtsJH92QMwygtHdXzQ2P9q6zoaII8HXCv7lL4mubcHt
mKhDlF1YUn6dRXPyBBa+AjhNgSnW4wqDIu1KqZbpVcfWjcF/iPq+B/XyLr5mjrwMR7mGzyEbMAMf
IDr8u4Mw8HkJT2ZZOcr3EEG0/ljpLk6t2xgOMV6QdB0qdTpW2IL4vY1TVLJJrO0rsB+kgF8ekZwu
t+S1XcOuCBO2f5JhOhGX2XnL8Dqi9nmVUqpQLTvxpzq/DcwIdkvJiEYcoevbBobQQWrDnZlYc5l/
k6ioI1gWmEf5EnqXxyMEFHi52HCIaHlOW6Q7uxcJEWfP3LXGWbjVz/ep31OPNGyRklnlDOZkgkOZ
zHp53tsq0tAtPumf7E/hG68db2fUK6y0U80K7FTVqbYb3bz8IKKQ5mBk5BNPHecSoVERZHwZYTSt
AXfJRdgGTUAVciV3YWzci4LjMIVNnaSF8E4BQdNE1OF3I3LGgfGytDVXkl+LOj1uLbgDCe8DChAc
hp/4Ny8utZ1exXj5re+jXcp/pOLiTutLpu+VgGSpxqJZSb8cMOMSe45WMciOeoxEBmZqs3iSYtKJ
lRIrU2pAACOrWYlqdD7HogaSpffqyBmKu06tlKTbO+5ibfrWiS9xiECmEyv/htqoo9GABWhW4uZo
XTNyFWSvSsOrFGRL+asC73LIKGhYVYGP7/NWHpRlzFxZopfxQRwlRQonoCbJywgBjeQjJLEHt2jZ
kz+G8eW57/k9rzNcNdgwm/VIXgM03Q76Kn+R8DOo7PKbJw+608W1W8aGh7d4hdzSaoUsoiJriGGw
vMEcYc+eL0izSL4BWm429XjBDcQA3xjkGUO2jBG0slhTGgz6HUC2bF20zZe6EJYwvJkEQXs+eHet
SITT//c9aPRUHN0HR/6kFl2iaBwLW+Rs2R8fTzstOFE4Y6i7MZQSfHQqJqsdM8tArH8Lk5QZ9gx8
at8udT35QQsNPO3AeMPU9X3F6YdUVgEvfYLp0VS+he24hNB5WcSbH/Zgx6xPz6wFV0d3uus9E7kG
xE7cmxwUv5iTXpo0IIWqUlhUnuCkIc3czn993CZkmFvQkhpRieyoKnt6Hu5HviM0ea97qo+p7WwO
NRWEmi4JUN0QmGkBOti0Kzb9vKEEnpW9+mco2NV6ZuP0GXHI0WA7Ublx5pB76rcAkSDimuQTl2zY
2ilvZH0I8Jdby+qyHJzOc3YGHZNp0PtEiobyoMc4cOJ0H5Y+M9SmKfjNYj5JeFO5sVsxSL2NLSmF
m2kgoemINCPZ8oLFpZKWgSl3WJ+BHQbZ1buly99VFo/EYtCwYIWFViHXkUncldBnRs2oKtVQPjHX
l4Yfwa8EWGR4M1szneGLAH/Dmha1RlZ9g5SY1XKGV8EtqFk1zNXpdJJEWPBkyFdU9WM4hU4ygUGT
AFhJANKck9PQJWpM2+O+Wua0ImmNXIpauNuDwYS2MRKPdfPP5hyIYvFTMpAEfpvrG68mATs3p5SP
DJCzJQAr8g6L4JVHIzZKesfsinF8lyf0OElInc0KAOSL71QrFNvVBgo5GsXtU4NVgcAC77VGVI+v
AQbOLlVNgrtP79icSa3BKbgan9AoBg/QzmVKLADGuv+vVk9b6EkX8QfDxgCtIV3YfL3OWxR3hQ93
iFLqwTuDYrTy7K2FeAvDT6ZWZ/rNQ3kNcmdmU1ctbRiZzHPxZmvKNmzzzF0UzXtLjUG00cA0HGH1
umYtbBT2T84UPErDGFAHl1J1jBRqBe6aYNV/JBmYp1TmmbEgS/TDx7Kf7gJ6Oqceg5X3GQmCkztZ
/5UK4ax3SfpmGfCv8WXc30PH5vTv+6XsRsoKf41nvN50afAX88gc9z4PUCr5OcvEiv+OatHqtJF0
t1v2ulWs8L5Sq8DZ5STepWf1O5JVmRyjjL75TSnzid0tBf4+zc4GY4fl3w2nB0B+qNGJGJEq283R
Ah7LMElBavN5xXlHCbZ9vEcy8+4V+A3xFu1NKAujYVcvnnSCd+rELktPzWiJ8VqpuhoHyDVskRb2
ftmafxHVH4ExTGixy2oAghDZp8hi88TaVY0H9vBIZemfyvtOm6NNN5rS1vJwSZfT5OUer7c297st
d9NrmFcEMWts2uLMIZ9QsDscwbEp3KEvItcwHe0BLek9v05nAHA+g/88UZ0qygffeZYi7UUK42Rc
dEMzf/kDwTAiLmJ9LXwr/x9fD/Y9RD8zlCwBbi6Bm9uzplgyaU3gtk6oTYFrL/Jpzbv7475kYznh
LfG3+66ORGtiZovXUYaqRa58USQ7vI8/GdiyNkkHA5IHqYclClxxVl8lxOHrbzKGETDfrf/AiHn2
QaN64x8tP393XZX/FHC6VNXR5tuFcKDMdP4rNXN6n+gyq/K6Z+l4P9/r3J1SENKytwAwWKsDZ2jZ
VZAN0QQh3lupMt0hdYYwoBLSez2anzN5RlASwzCgCu5VBCf1XxvuL14/WVncx/DrWVyj6cUTgb51
Fb7vdiq+eEyx/CVNAY82yXlf+Qb595zI1crsoH5XSVe1g1k1hQxgTLQGMho7kARkK1CswI/IJwfZ
fGGx1i11dJDKW7bBgCkKAP+H5aqEe5MnwkVpnJMyCamNJFu4dxs64B9MmlZNGzPb1ZxhZ5hljVJq
XXTbt226vJYz+Vmtkg4VsFi1EN0EWlJKphCR6GhHMO/gN8XDYnf0M11XNsfoBsc3sHlLjwt0QZ3i
xPa9IPfLjLWfMpsIYPY+YQ7VZfyFUqFIqdBADAK9PUg6XCGEHUv14sr6xeIdMY/tCpAELwaoUBZI
UWEqt3JtkxqrZP4QDnboauLZxscuukrmUnDZkv/w4YBo6VNej8mrgTvczA7hagfWcm/lgGkITUA2
3LDbo/bCTU6CNiJDXDvhfIiJe2BcvFilvG/oE611LK29/livZ9m3G9sZv/MnCeI4+jDzbSWTUd8+
iH/Tn0TR3R+VSDieztouMTEptxKFgkzYGrFd1j6FSyA/0HsbCrmWydl2gVaR6MK8J0+HGQXqaoyL
FRE69XX+YeCrrBT3/zYZrRmVAgff/SFMFAvoK+AkSlDuSog2K/vmuoVSVlMuEiGc63SbsShFx898
Y8NAbM8mamu0Pi9LNJEKSX5T+mudxxyWi6ZQwi8Oaeun3JZNUB3PD/w2N4hDVW2wJeP5zdqtymjT
DUncNQTVWaIq8xUVJtIELOdbaLAr/VjXDAcdBBnAZ232zgqo+jQMOSnCaSQZno/WxgJiEWktQCPE
pEaqXxhYz3IzKBcD3JgaVv3AoURM47ip1BkfW5Vn6xZefQv3q32jaMDTMIFMPACIa/nUzc2FmTT5
N+WTojNcD3JtPuoG/6eAIn2dPp+alE64qAUz7jkTiN6KVPuUukD0uTU8BILEpEsCGI00uyy9V0t4
NHDuuSPuxsGG3Yn7ykCbZdXnGPklundFlSpZU1kWBktX7E4fN8ILtUHsYM4GkHUZFtWsv2PPraYh
WVovIEL8KoTAyDGbGzczkCSRWj4yRjZ1ZKD0saKRM9Mjru4uxXPv6CkXPHJ5ndJ1GTID1u3iryOc
mx5fxkUubQTPM5oeUFcXdurP98SFDHrgmn1Hx6gJueAQMw4e/RWMq9Syv8Vq/3A4U8Wqr5KhKXzP
Tvw8LZ4K4oAyeZnOk1bWQ/6ReYrfekUAjU9jfAohaGNxYJ6VybZD6iBj+ZiTrv43K/LL/T2l3ffv
W0oasGV6DoF5PHaGid8n1Mv6uxMxZvG5YckwBZ7esLmvBJPnb0bplcMSmBclqW1tx7ERJbFKF+ct
FgRKOdfb9b2wPFha7U5rXuCt4JNLTubgolq9yLd6H+phfl4zD+F8jkMVzhZ7WLAqhx1PANR2nUTZ
9tLgBKIRmrb2rjxSn3eZ1mqUCXmuAO/ArbU+fDnTKCcDm/yQzWMdTeRnheD38gQ7APmD6Q34GlNZ
p67dp8LNI7aCM8qjoqPCZIed2cy1gAopHlAIRRdk1mdcnIu/K3yhM+mUTqQBbRgJrum6KHldXCVd
AZgeSz6WIxg60OFm1BxYe1FLJVPZM1YdOAlmUoBCGebZ/EO1nqiCnESco7GOFSGyplYei7EvKahT
I8womAxsl+IH94Mi4Betq8u7wgqkylXR+M0sJ+PP7RPRC04gdPJyEsGHVC+cPlQ6JhJ54vkfKClI
KHLsM0Pdhau7ZyEUB6aeunvuGPnoDHVeXi0laUzILOL7VM0df9oL/BW+NWU+1wuwL6YL54ZTns7o
pUaQOR3t5W2We0UAWl5qqFyFZDBYSg6ts5uxR3BI2+YvSgzP2EBkEV4Fa3jyRORjvcoToxy71dBk
StlNHqOFy2rnM8o+EYTyW+nP7Tpdfbl0PeZ7PFtcFakPv9wgfjhgTUxye/88cclEpP8JwfuPFaRx
RW8dz06dH1y/RzVLLrB1JKZDVjpohV2ZmVL+YDDJOiqDh2CQjZQDlu/mJJUTzbQInqhE3T3xPfDk
eKSwy4Gmsb2cZ268rVLlB/a9dYSIiQzw6P/cMPh7FXdmNBIpc5yjob0xLokMXT2hnTDp0RSl6ycb
1y3K9OPahHGXRomUX3j9I3gHEPJkP3wxroJCAyzGRoL3uITRwxndTgNd4v/3bx1IjgbmWN7Zsj/X
t1BbZWS+NdN149JpIwOEmKULjjV36xRS8Q97vJMaSgXa/OvE+QBcQsnjzLzU58uR2PvaDQhgdRng
9kx46JRGNGEzgg8GA37tYanvkLD4T2t+nhUrvCWIo5XZ2wwc6/m12ryCgm2JbsYOBYfykoyFLTS6
bcuqnP1ArTVRQZ0xkBYndctl8+yHTVg/Bbc87yxto2oeU3r5Mq1Mr+LnNjKvv2rwf1MCo3fN8a9u
RcR9k9X/tLSWSucndeKrR6HKpZvne3RRUp/ac6KWt7lkUI23cfAu62LUOYFJFIXCTlaW9FRifQ+u
LXB/04RvOpVxbc8/dqgqlKutIaVnmFMZEnvvf6A+1AhFMxFIGdTgV9ji/mDm5moOCCrz+WGnuXKV
YSs0VUIsDIZXyjnuA330/rTIzJRU2u/vu+lMYP+vNPlMsJoW/bTqE3NJsv53D9CzB4L2MskyDwuh
ZXRFdrELHhlwQVLsytK9pCGS3ZLSRaZb2ipYj7957IIOEqJx1KWq5FbBZqd36HsbEc4D6nu6f6y3
F+sgeqbzy6ha/RYBseM7e/LJe9EPTMEt1pes0Wc1hqXpdEKiyeMdTAYwtjGkQ5shWJUiC7sg7j4D
clZasSVzyeJdT/siAngezl6VpsABigM567id8y5vUfMHIntMQiRdAMdSZnokp7FkoX9IIcwnoNxy
2HeOIwAvuXHRkIYnVI1dyeSQCvNg/ldGWret3JU5MOKnP9RvJQb9flExrA6drgQ2DZr7Zeyi+Mjq
IluCN+WRWbE07buokw3zhRMVyxn+kzu2XWIgCvx1KKWumQ1Qvo3pzAxxow8HzthIu9YGBLvIpjZf
BQJfbXecRmSyNXuSZPkCvqrOV/h1d83d46d4+/y4iDKuy99bKJPefjtYFIffWJqCobrhwinibY2P
RmpOkKWhpVQrQthSrtfRN841r+FEXDWJB4XHumIspSyfoqfqI3kgDEdAKIH9jcn41DZVO1+lUK65
QMmoLzfE7+1kUR4urjaAPS1N+FHi3AE6qE4b1OROlaPs1DpD2JWQTVBSgcqkJ1lucbjjLUmZEV/T
gKSE863aVgInbe/WcH9WC6bdz6YMbW2h9sNFdYALav1hVKWJVdsC8rI79pYp/2B9cyTR2clQjRGy
k7NFwE+ON/uR7kiJ4hpwcx4gGZ2hQYF4tIv4nEz0Ac/HPSeOPe6F3hV8uNQUuE9jQflFyFXB2Gkb
Irc42q2wlINW0JR8M2QC1+RXhSA/JMbTjMUHQjEfyoTYWwC2WGnTOnBbtjZP/Qj/4MnxzLtkYvd3
4lwVmsdoi+Y2BtmiCIeEzZypINYdPIR4ITGHsd11WRxHXngGOkC4AO6HduSOO2QCmL0KxZFvIzX0
UIHgw2Xsuq6nPFJ0wR5d3cRI7KvPMmSoZAezMQ+idh3gYBkTD2STEBnYK0pAhGad3DQfVI7LeIwW
50Svnau3mCO4wmPweIbKCxRWCDb38ew0mRyAUMtWKKQ9PH/7b8n6JuIYA6aTQK0ff0HLlqEywu1q
eV39FqWcve9tfl88sYDalhVivVgnMVA3ep+f/dIjKM4ryLFZn48S/kbCyUiDaqAe6bUiPSyQoDPV
+zcv7Tx0F6Al3ANtM5BiCuAiqRVVt74f2nUS5kS1AhqRfIkLaWg+iBxTn6pOVsjtH3bz+ZB5LGVX
fNa+rxrKxfsbcupSX5ZANYR1EXWnqyIjyvlwoEI7j1/tbXoQxXb+jHBZGvGRz18vfIpzNW5TXHz5
GtEBgU+sisX8E6dRoIjzDdcxJ+o0H8assLPzZ0cNzuw+jv09mr5dyPfeTPH3jyvVgMGpxDc5PtkK
LzXAPNxTO7T9jh7ALpd/akTlMYiB8peg8Jyw+wJXodPE2TT6GZQRmIC/US/hoCsKze0dUcqI1NyB
vTO0o9nEKeG/2HOIpGBAtvKgHck1EyVAvz0xHwBc2ER1KvqPEFDVAssLHBefNx6ihz9PXFb1RmvH
v+AjYV1j9M4XNurMe3Fm8gSCGOUd7RR8RVoLthY01jK8bNnZ6Ds5OkXCJPX3/IoLKsZ6D4sv1Cfx
7RqpLbJDRV7hm65QwVIUH6vas+PeeCO9s1B7E9DsmL4f59tVUxcHM0d+AOwANk6EoPyiGciePVjU
w/oKqtJjmw6fTVnYXI9UAMEPpmXC/aoVmkLn2lnIyXfjaoJtJ3bAp9Vn7tAC78tNMzR4BEcEvkPF
aEkGRo1hFOQ3rVfY1z2PT3glaZXLdklcEgoj8M56DRP8BI6yV0YvpTGEI4N8a2mlBUBIbFumciOF
aftgS4bi89adxOVyqhYjOzC349P8cj3lsIjsK2qewHit27mNF6LVaeEdpVhELOAW1STZfOcIA5Lv
C3ib7ieNsms4jJxm4IM41vTRbCW9C5Tn8HqF+eO1QWkWLXFmy5blxP4yYYd+Xc6Q5tSixJhyLS5T
VxywbfeG85Z8LWV6MzvEMlDILdeqWPvj8NLnc+ItRaFEiTo2VGnosCqo8qWiXpTOxcuzR3lfKKFU
XE7543lI6SbbG5I5LQltrcLbCmT/p6eo779caNJtldBT0XFPEKkAL1w9M1a2/0zMqnRc+kNxnP6g
VN31mCPtIhL/otDU3uVHhYSc8VWULQNMEqMwc/ggCUbqUaNiqATcMuWaWGSk4csMGa1I/jnyQhhI
7OqvgxUW23wQzGcwFltE4INwhBw5q93jyYyzS8fKiqHBwKR2mFZUPy9iGVKsQwEyTXedFDzHKssN
FmYri9pq2dcCAGAAuJ3vynxsfHuCtC0/64MTkPn2IPqmntJu4GynAEpDCLnpcfcP1QhTuGGSZmQi
OG/DaAXgag42HybflhFG+A3x50ofsu3acAFKLm38/JQPA1Lx0IkaO6WSbFgzlz0TcXxieU1sAU9x
GDUTRt87nUrDYoXVOLjjkZ4kFSonJbJJkLDlHerVjETntt/4IvDRlNdDjE2+/MYlU4Fudsm2ObLn
7Has51fCFT2SfZq/3xyIdLCb+8ofwEOWp45FRSbWQ9WzcY9WD5dnPU6OMzcLOJ8wq/E1nNLGTamw
P7QVCoRuomAOqlE7/Erf5J+M5LRk0oRHR8AUI4cAfoMDDWneWNbU0gXXqn4JJ/rDpPay5x8sZHX+
TKSYw/4pfU76HgwthUk4l+hE2WwSP3viVJ50V7F8vWCcc8TU3eOSfX/Ydn4lTDShQu5k3LDJ+fYk
UovvZzJYiB7sq1k6ozGCgLQW51zSNiNaP7/7nV0jur9lDERNWpyHxlzZ3VH/yLgyRZNkSXFglXqS
t12BgQDFH9aWx+gKuiNK7fMq14rEADIPOvOfhn38z0zPtUKo1Pp/sarGzZj73ua5rFoOGd6/kTab
DjjSYHhgtYiN4JSF7zij9lF7UqLxG6TsRIi9kigLlGciMz0AF+En9V2C9rUvFcK0pE5ahRzHefqp
bCHfnE4qCkpUK1OFHbiHG94yW+yBx76o+FWMD8qMz2ReQqQDQR/RN6uhPhmbGKA/GVz7zFYZeABn
G7BmBY2LTCfQ8VhojZDuxwKm8kAkrHOP8fKiXdQhQEIDG5lrbQevBE+GdbEkLOW5dWpAnUJpyOCe
tQb8EJXP6J7nPChYAn91gTwOl1JyC/TusSCpVHwezEV5vbjzcUSpmQGTXkrPXNQwGXXVBUmkhvxt
G6sB0KFWQMcs9+eeULuIekPFox7plLtQ/02q4AVbpT9ltHmMItp+D3NjDPFtrV2Vl8NVQ+BT2TGC
3xkMYp6QPzn/Pb4aepDWzN7LSiueVPM0/edb6WgjxoBq3OLpqH/6ynNFrdV92X+s+pFgqZM0NUoV
U0CigZWha6rrM2ML/twotQQd3hR5733pZg5NAeZYlO89GSvJZk3T9jB6z7o9VLJ2zbDV95uU3Kez
UCVgiTWX6U0Ul61WlZdD6aPUQBfuZcph4FYWfMmjJGbqP/tJfRDAfWXgJ1od02q1MHStzBZxE8o+
ieMeOV5YHcOwmhN6o4+lNzOF++ecinnDdJK9cmhi6QlzET7pLCB6evVtwTzojQL2ipni6U+IjYWj
wzs/0B9FOFLuk2hmoAZ5mWFRFkI/bIDXRMIjcq9L3Vnf/VYizuO+mlcHaw/56+7TKIZS+3OrjvWP
rFyryVnQrResBGEJq7vdzfbZpi1kUdz/FH3XaiQ9pQb97QW+cpPO4aMcQ5R7SJXkx8yJxDR3UoZG
EE2QSHt63ck1JOcX7gRs8836cz5dZrTltiLUP3BiKwEAzh0KitAQFemmCQD9IxFhjGCYSe8+qTPK
4aMSD0KLxqfAZ5pPcGX6e0oZeaKirsUpMKGx1j1/BT2Q5OEyBVRG5uaRVQfaUU+uU8M7quCVbbAz
TcLqBhcv+iMZ9f0AZ3ydO1GKwLFeyWib/0F8m4+6A+9st6qTb04ojCQI6SFSOSkYl19OG5m05Es1
MdaeOfNuBKYPaL4jshD35fcT8tjojhd+QsPm+RuC4CO5SNshqUsgXyGU4qD9ha5o3QfPcyoSLNPh
UhG5S9xiQrfeaRae0nS1I8eirtu0BddhGwxXNJREP3duXG5groNTYZ7EFbVRA7LnUj4ruifszZcN
D4e0vZo/j+VqZEULZhcbV5oJ8XLR5ftjXhnrhHsnvTbqqAvvztVQPmpH3BsFP1zWXbCZNzU6fo6u
I+fTa0359VnV6yQB7PISX5/RGWEDzczhmoPIq78diJRFcKlfOOqgHkZ45/BH6ZSFi/LLOWO5eyFZ
1H2hOAzoNdSxY3B2UPM8ruPiBRYQGrOAjafEoJXOOUMDhqH0SJsHAyO2zRUt/n4c1JDsR5XVNWaa
FLTp9SmsKqwFS/A0fAYcmfl9OzVRtpSUQ5iiSKHZpcgVlMGiyFquYaGeLrb6jRp1Klq5iqe+hBj4
Mv2psrIP+m8INA35B/FW8+MiqLlGjcSijik2ixVAPt3TBkwdxVhgWGcjuxGly8fI4EWtg1dEPkkC
3P199Fn/WiKpjTLDqybznzCWIz2udhhxvFPiXJlm/rrDcr5M4MQJOYSS/1FCf/tjD3sjc4zsKPZa
sGb8pNh36Oq1On4gpYhckLSsNvULK7YHndz/moY9TIF5uhYzrOTgM+xdVlmMgc8ndq427cvBrbOi
ClQ5zsdyRAjI7h7lLizCTu1IALbgCzLa/hv3WB2bsKWx5oO0T6oaVKiiHzNhRC9/AEtRh0cih9aV
MHNr8y/3Cmtpo4JPsZWs3UxfY7p4HvaDHnA503gwLEgTHesWwNpiBn5ceEI3rWt2XvBtPAYRApoB
2t936UmCjwvNiREvu3I8g1q3tPcsTY2CdWenL1KqSqiaJxGamOLl7xZo/G6YDlD40FgbMId+j4nz
dPClxhHSMTXbcp5WLH5kSTxYzhDCtdJVz2wLWpq9FdyMLL+x1g+ObqiEKwFD3cFLR2Nz7A2mAhgh
RTVei701hmQBbvjiKBL2Vkffa+xAIO9MUtdpmkdXmn8Q+v/tFxgTDueqWVza5IJ8vzyxQkLgqwNs
gct76cf3Yf4SoMd00w+BLOlnbmB6nSbJkI62uA3izdtfFA0PuTjubcYUTiT7pXhmsEcc09E0+NQ0
8xj1ueGc2LuiD9sKu0RiiiUnKRYRmNvXDviM+HYFmBNg98da8SHN2JClStB9erhFDYuA7gCTjBGI
e5fE2peQuUdyhRHFafOFe2DBSnE4boCCtbdgLcpxcYFUOJfpQeyi/KlCX4XpdJLgK9egeWIDDd/V
vQnZHbrbSDnC3hf/ERxxAGSQHw+TBU7FPotq5Xo4rKDMBdyIaL5wZB8WI69zbXAhc9uLjakij0K+
nRJOezSXiuoYBLTJEDeixhrk5WYh/kjjDZAi9YF15LdHZOWaNfe9hL1q3Qd/PMpk5MAlDqgCJ/r/
RIWe7jS5V9Rpfg4mFdUHUzx6t8pttmt5AQNHIFjzICsJVI38F02D4UuaZW7Ntaq+Yza4FdDYfvu0
1rTClrQfYq+cx5i3KcKJTyve2RvaKX7qqfTS/haD57hvmidl440oT4qHnxL8vcBLeNQ/vJ56J7lE
5sAVBYZAWPqOXj+N/Adqff6YzrFwq0k3oT26h0ZakFLuBLdxcJdN9e2K15aYSHAl9AptKoDQbLl2
BmanUSn8AhJuuk4S8eK7V2+QgN9uVD+XaQ3n5cKCoVm3l6fvtQCIunkRKiDNxHRTabMcdMB2dA8n
gWLJQXNLc3uecxm+YB6A8LkQtQEeI+ryUsMd7S0OUZBISkUguHZuiQnTMiRN7AsWJxH2YjThmSvI
gctko4Ey+8LmPM/wfhnkFRT59gloPpb4RZQ05KGP6MQ1eHw1/43YWP0OLgEATp5SpYM0ceHsZVR7
6IDgs3wB66R2ICJEXeDE/EGn+/D2cEHiV9dZYxScwKnG0G8OdVS1HVAoY5sTp437U4HoeDuj84u5
UWOl6ieyauZHBLxbF35tydimFPu2VcS1G3tcBTOFgItqsVB3R+KYzEI7nbpqsCWQHUC0lIy3U0TK
1OQ3gr0u0MRboqe34jKCunoIne+HejW6HIdJoj1WSVJdPg51mMXApg4e0l8gqyCg1BIBMI9xiPEB
hXazBIdtHQf1HIfSKfI1pcaNDYVIMIgTQq/HNNKtkPewbwk5KOwGw41tfvLbWjPGv8OrALHPcoVQ
QMjVjo56G6xS+IMa0FprDAjUsEqFM7C/dG6ZMjj7nLfNUsAqGhVMR0hfciog1fpgS0kRzBhRMSfm
i24AAs3raJZEsqtvU1rFgSY0ek5ORxj35lw4FbIjS3vzHf87GqBtHoSS0/MasR6WvlRil2hcyDOv
3zR45EEe5trVM1fzHLUmO+GV+zjrHVxNYqjxV7u9d4csmR4Hgg5dM26fGBHBJGRRiRJoGXcK6GTs
uWqYxq3woLixpUFc8KVKkZgjkq8ROSl+29MswncoYxIs04V0psI+jXK09Q5/yV150ZsSC6yxDLn5
aEzBX3ZWvLsrPy9Hti6WfsN0vKpZPYYU/PxkeRVq+t9a3BO/sAej9jp8OFcx3WB3GbfPQZ/5fs+S
GeZtvmCiXvn5/Hhl+5PAgk+Dk5re1vuKSj/dwbXS8uk8ZBRO+Wm4w3P6ZGm6hNEOeLVwfx6nnyED
j6EOvC/BNYyafI+pb4HZoWa8RZAt0nBKo4H1kn4R8h+L3LABrMtYyt88x1+jziwIPL15O/WQO1eZ
godIKoeF8CxUqODz5YaN/jXaT1u0/SrMQ0DlO3I+7UZSzkcNvYAru+MuAA66ZbN08cl8TmsThqP8
MGBHsi1R/qvgZlzWdc/FT+0tCsAdvTc8uYzm9ASbqgwb1H9i16d3x9yyEHV3WMHbIP1UyukmEKMY
ej8en8EchDLPGp6XB8yPA/UwlRZQ4qUK0IOYax650EVR9R0U87dM3So0Jyh6ccuESCQyldqpZ5UA
St4OoOcMcHI9BLFCIo4+2ukidqPHvaxZrCRWajC4sINt3hvnrLQDTvkJtARcuduoXKEqlGsEqIlR
KqMDM9KyYXUWQYF4KJSeIkvBspXLk+HXhQjCkFtebrP6aL3RrZv4uNAe4UqZSXiKYrV6UMQ2QWYH
ySAJbEsPIInBLvbHDLlEw89KDj0eEnUXnVlekI2GafzWbL6D257iaNKZpLeq6RRVY4T1jw4PzrbL
5krQGZxmw8Ag4KkdgfvNWJhC186TarZSw2V95qDzk6XeqEo6fmCFI1rxHDSSkNf9hWUJM9lEtgAj
LXh/mB62k32bhMv1OmcKoHe3I6YkaP23GI1DYBdHmmYyQwLXpAsq9LV3K0lpu7goI3/D/jKFG0kl
MzRmJ3yVg3XVqQagfVknOBRrq7Y17vQtfV5kD7zowNaz57R8yqO7HpOulKl6kEQgOuMqBXCTSd4m
12oaSiGWfhA5UwwdYaL/ulerjQzvOEYUHNdGdm/YH9qEsABPsIsLU8A1JKx1yVLxOgaSt1AAgzHY
g7aS+YB3QhuwHf1YLtaUjJwdHwGyWDU3TaS4yjlq6jEoRY57fkExGcq779Ym5CopxF+KXtcWhUv3
DVysv4n8vumXzzWPGM2woQWRArKqnC02v0pxJq+jRuZ7JhuXxNEljTBu4UKc/LSQMxQzG2Yoo6qU
vxQxuyISUIdpLnrrblFhA6+b06Bt+8DSkV/CaIHg0lyq3NBqDm1rVI7xEk34FZOuw0zHM+Nria6J
tyZ6PGFwYW/gSGr53Yunbfd0C3AdNoo7m9euqcRoHasSzKkeYX+12l/fomgWPw3g/38LFYOfUEmv
eBYVkV6dJTaK1n+5ZHLEvxlvXnx5SRs1GnIa1bxL3kKR5V9WidFBJ7JA0CwSTgjxckMOTRViIqf6
125UthcYqtifFX5FKLz7c+tqVI/r+BluBNppFbKOhl+f08NxdCdaFtq1xecSaDJTsf+D/M9T5E2u
vjOE0JEJLxIYNkUIk7AR2iutokYJgJEeSH03gGH4erYovCsjbL7jdMnMRpkrXgqr7iCyhOFQHYvU
hxLlwsddyYfmmxGocFhb0EBoIjrc6K3cAl0Vk3wKhu4cZMyUmCXU4ei6u77kGgl3aCc6FkT9/adD
+JmJWka7Votg31Q5ZP2YV2sTLsqwEWG69spT/7wi9OYKoMh40zE65OSYRRUdHf3O+TmwRmcgt0eJ
SXACM8r1v1R+6bh6sEXLs5zNbpIwGRdfXxE8j/OSx1KH88txtZgAV5Q/NfR9ZAnv7S1KcosLoYXw
iMDVAS3tkHWQtHwS13kdk6x8a5AFUdenLgGV0FDW9lShXF+i/0uShve+VP4BZtYnCvWVZXHKwRyH
CeUCKpXKHn9x4dtPYADQF9IwImwgkcxPRWUZetnZ6RvI15RufnmAvkDzsjVeqg4QJ7TMy+V/GfSY
scm8ttpV81k5dDGxMHuYP+TKgnB6pfj/kN5oo1Jggj+6NbKj6jCS1cWVNXwIoFdu0KnUa9BMgeUP
OR4iLFeqiEtDS0eLrSBcOFxri8b+RYdqik8csEZfezHtWSj2C3H4xrnZIm85NlhnU8TkdKq2D3uz
eJ2OaUQAf2wfTxbRWAdDDZxcxQQ2ISCkYfADmpHNbcCB+WPkTCrvp13zPsV4wn6O2ryK96xMggOL
x7FA0qxIvRxuTcBumjZtUohCR/zMN/rT8cjAmgECFd1O6RRvz9J5c55UW+z8hetVDoM1BnzChUwX
cj3kgyiZKpaCQprS4TIWMQ+DpdPyUdL0lJ1lv/y/y+xu7LyTfwoPjLcVT+yp8m/L3PvMqvv5XbpO
4n+5vQF8+whMT2437ejS0hY913MPNfREHQqBWi5rARIHnEbp2k77qh4HPybFq//YVHNUkk+QeHFn
VmiVh2M2Y6fL6U7nmTOelnvEN4VCLC5EzHpP2KRyPBZ3asEK4tTP2jApyDaFjhRGfbsjBM0Onh6l
mZl+hC+a2XMbK7LzyFj2GX32e8MTydsY1l7Snbg4pVRYLNI4QPqkdgxy6uDDOS248R+pvPU/5AeA
MvhAY6qzWmKXwSIPrSJmCGTjHgIUn2A6NXOuQNfUyf0FFXbGpTIJ1il6t3NymWONK5sxGrKoay/g
SWjMeF+gg14XdzEdbU6DqN7OZx+q240pv4nSXs8rRnOj6nS3/go49SagUS9wb/9NZDDbRmQVP5lJ
kYagOlVXG+S4H9DXba35A0xN12eC/soUqRiq9BgyIfLLG7rtwDK4we6/GDmgyon6aoZRfpieHNu7
o5aFSti0fuFgFVMbo/crtgQemBVCw/a/1ZE6qbcE1ZWal9RnyLo7hPGWc6mqp4oUn+4XK9sQw/lR
kgZFzO27a5n5QuPu9PvvHhQmN+vlXddMTW5WuExYOgYPzsMrwvxKWDYqOIeod2/+e6bDKBdhwp1h
ZlCvnbJ7g5/dfmqjIwaeiH/7Zcy0OZygrju1tPVMszE0/+Uef4DVUOFlnN6jDEvSB3uFN4tquF/l
Ysgcv39nPzeC8zxMY0STPfKnIThqgn09ZhL1a9kfDDA5U6xMd/11onx/60lXZaWXOTsTQ0hCTzfK
4mF8MbPv8RcMRMrpW1aSD2JfOIFQlkE85ndDm65i1L6LiBUnwXclrepabpjIHLSNoAK7eXm9adgH
3F5MNOKvBkGnA95cvI2rzqeSFQTE0zWgaT5hiB1uoogn/RpOnEbvPe7mMcM0MVw3Wnb2aJ6Uje8S
KEwkND1OOq375dLEsQkwoN5TWCI3vZu8nCqVNUqYSy4CdM3Gti+lrVBxl9wEEKC0fuEideTTxiRn
uO4w4xRmCVEsPAtmI5KEW2lWe+ZgQhWx46xAl/Z+A8r6anmOa/V99XhhyRjec4QbL1s/SRNzacBP
o2G0F4qi8eu4zXsvDTQbA4nhoZrVVcYhSKCVvVqN0+H3Qx+eCol8sbaXfQihBHlLFOIQzEmoL4II
mNQLch8pwtz8V4hg1iFcpn2pXhnmWuoWnzw5tbSEvQv9gQ//ljEdfWw4WIl2WR9Lsfc7Cv+z6268
OmyouILK18IIzgGh/KR61cng7mwb6bx9nkRS4/fupYKhlcsF6DoDwKDWYm2FZIFoRSsQRZgbjCKJ
X/LNz+3heB8KC3qQ4/c0X7CCoLtV12FLocugdESi3kddI12GvxG3oCklsMIHsASVgpkspwGGOg6Z
yobpF1qfrq9vWRcvzGncViu2nbidqJssHZ+WfE6vQ6P041PTqfaGRdG+g/5wwbNFMdm4cCXwpvW0
0/RXAX1rtY3nsJ7Xcp+JpZis3FpJVjksjMjykMGtRKrryYW332S2vbqalMwx9/KUOafJxwjrOD0T
v5LG/CT0gjvzeagxSOWv3UnAQFlD4hEd22xKRRWQW+XK0BsXgG6PPUGyo8irAdTGT3pwyIjs107b
sTd3teKf6+fhiFiB//0xgR7cUo11vPajjUBz3CA0l7+eMTKXxFDa5Sa+76ak3pqEpsjjoA2HvrW7
FXauy8EQUChgBmRAefFSpOft3fnjkOE9vvMLBWxOpIZ1uGbKRg5jfQMWq6J2G4Ycs8BGPSVsMG8P
FUa+5PerpuIo+wUgMz9m14tdNfb61ehOZRSSmoyRdgjmxi3TTmmSDhNN4iFLYu1UXUJwFZFmw3co
b8kk34TPyvoQIrMQYYigbjEB5ZCKxQWLDqyF3e5OHsWVu/fMq595QaD5VEa7g2LOjEj3U6Do4Ljg
q+Wl4RtG2UY7TTqUkDI/5Ji2tKUpovielYjXxG/Fr5L0lje/x50QdnIW9c4lmVU6TaeG33qFSm/X
YfSh14gx2HibTBXlUBCeTZoJyVl8fhzq808AuuKMlVaYvTLSRe/I9eCcbxCUCkF3nPIVvk+/M6dK
l3VzZrlKVwdjKSPi4hg22XBbxOTLRuqqJzCMt3v4qlSzS6K8DKo+GCex+FINqFrs96hDHZSKvzmb
z0LrZqKMl5NB3AaP9o+0IjCiPD/UDmxQxevV2SmJj7aY5W3UHNUQlGlWp+hWxTV8aiFyumjzH1Bc
7WuIk6Bdx7fTzl45hnBe5t4422UFLOlMoCb50/mloBgbT9EHShW3CKe9SL7yTEfeY+iTa1NrQlru
jvqiblnEVfYS9n9svqQZDEl++Ajkifa01yDLRKrPKWSQ21Od22Au8VxSvOl+xSOQ9bZSKOwPWXLm
5+xyPnjZMYu9aJNUukialLg9TqD/8P39MIQ6BTLpTChVl5rWrBVqR2SigxCaFS4UhCFiqYhXKXlr
XfKkZkG51KdRPluYY1el4NlzAj0UMkhz7/x07XLC5qckVTDh0nxDBjhE29ncHgrGToGpxH1F+0jH
yMa+ckvArk/5NV1Godgheg1pn/rD8g/payzd0H+6qSpBCflgWmxZfiNeAEMoZzlUiOVtfI7M4k76
/ErZdlMA85d+dCuH23GOoWPd51QdFbpvTwR15cCGqxt524u/Vqjk7HFp4K/J3KO3+Qv3B3XEhsz2
eucltEm+mrr6OqgluXSqAfHNzbvm41fwWdMjtwbTnr77Ll671AFRb2QA1NenFXR6cAno9c2qXo7/
A+YPGzQW+bDehHcDwkXlXjKzqKHx67yENHREbKuYEFFalj7qrV+QS3RRQp0GQTU0wXTvYC27Ph6G
HH3JiG/z5acqzI4UUd7lR6IlPLr/qC0cW21+McjXMypcZP+f+Wsqk78Adpk3xtdLpx6dxzOQj6w6
y8rOsFVvDfmFtPfTc7dT6tySovpuqvuHBc5o4XVvYMR7qlHuu8BKRGclisIknoEqCxpXCJzGXZ6z
GtCsIiBu5ajHUQ70yOs9oWO1TdGQ/QvinkJiZ4wgh1KpAnbtrDVJ4KFbhMy/WZrgZWjNTyMOMvKS
UN23Ku2iYnaHE9EkrAjQlsVi5jINjB1z8KbqR5m3bjcRegMDtzhGwKmJ2AqoJIt8h5506K+n3npp
tkO5lTIp9nuSRg+YV+EiPkwPv3/+trVe33r9MCY1Kaeaxm+rnRydQkVCIdJ9rhsEVezanR5zM+R8
LfbbvWxLQLwzqswqtN11V9SrbcdaW7hTnvKRi4Yj4T7xTL5i7Vx2r4yurF7NeX6l6W3nRjxZcrh8
lXpG7u/Kb3+79I1Z4Phr5jVM5wHdopP20Z3oKqQmXT+/UiLai1f59LIZTLD9OZOXju9NpoH5DsrA
fJ5ha6/BvRQZQI25aJ8kLpFxPKxAsrVjHp/2aKBrh66iXV0BlcYHvqZBb8Xr7s+l7JyjO+M6vuU6
S9X6eyTCSRjFrw62dd+BOP0LBzfEYS4BtcVs5Yh6I1U0TCI0X3AbqZ1bg2DBM8uHq2Rq5VY+PZY4
ppz+LWPC06zOvgIMOeorDr9T4qAQcjGcesxMNNdCwhoZXVhW1cHxvfNnKlmefn4wkx0ud5IMjSli
G/kyqEwakakfmswLB7KwpqnwbjVTUUfQFUMzeoiEFph7UKbDpGCFq/DlzTgqfqkBYArXgxpA0X7L
0jqNAZE2f0tWkKlBSmNLWRIbrNXIeWI1k0gpHy8OudZnGIkxiz5NqcOZ4g0IFY1Bf6a6GYwIajIt
oBxX8wGnx7lzpffcar6NApUBTVuucH3InOvXy9oezx5wES2AubGbLjIC0K9gLlDe+d7e00ROA7ZY
PzlLShulJ7KNV4CsOKCxxo6yKOqzF27bMYgLDFspNGeSiQm2peQyyNS6tTt5r1i9H0D3XQv2OFof
Jvv1HdoTERt3MRbwfA2wrRAENUH97j9CDxg9lyh2TVcyvvVwnLN/e31yNBnhqLU2BvbFTrXpybhn
MrG85ngxgVBXWgOzySx1lvmz1LCAUm/e1gFiB3d5iOepnbF7xFtlw3DWUP09Ff0bFPq3eOnxYNcm
ItWiY+C8vn2QiVxyyBCeQSi/BkMqz8LxKYDMPbxLT52/q6tFG8dsAeBXx/zcrfdxzYJOCKLqj6Lx
xBKvAW6oki8IaiIVae8+aPCI9nO0wO/7PPTsSLam7xAEKxXt61rH26IOebVpoz3UtZ72jhAXFG8b
ztXvJqYLmGV1xEbwVUjgwKWQfx5hKgqmUyjFeLMvMk4LqiFwF5FtVjXAkrjwjH6+Rc9HopLE/GXn
qFxKqUIqLLtjszQIH1dI9CvH8CQ8TjLyLSOGYlF0/JsuW4uSXHclQHN6lAZ0HuXAl6wHtgopSb2E
aFNTrdrvSQagPhSrxK8y2waxvcXJ1pQdHoHy0kww+PMTKU5/KBtoaNE8eF1zpbTuwuF8am2g9Y6P
GWzPL1bPTdSHS4NS9Ggvqxic9b7Jvlfogr0DIBsxGlzraxzxUiVMWTf+vuZat3oaQ2nNRR9S5J7F
fXzWhR/wjJXaNt8sR+s9IzppfbL6JYnOwQTxWCW6u0S4CuOu7lTFzSfUWoQchypXxiH/7Y2AiDsZ
Sz52DURnQ0RQdrdpTIVV+JWYpJVz/+GKBSs9lQwZ3ya5iZipKv7llrmjdqY4QrWx1DxluJ8ZJ1po
kj92LIOVMSr3MT6Dk3HW0EcaTp4ZnSnDOGiKUcVfLfw6iNZSSIMqcYYf8+V6ohMGTk6TuOlgFm0+
ieIgJP10fKhoIYq77z+DJ+S3NrduVEnfK1JWhlNmjEUnQ3BQo8P1eMBu9IIOMFfqEk4NBa3kUTgf
UNhjoOhyl5kuwYZ0f0V+Iw6WmEq+06buv0M3uKS2wZrr5SuC+1Fg5tQWoTnOuzl50FTkwP2RvAOX
3fz8taDTuTQ4euPKmEyF1zK+L3WwklA9/ALAV5OvVrySc84cdJC4vRMNegbHECPIwg6H9lFpGj+t
7blnkDRHhnj4oDjFw3zj83xpnmgDu1R6rx9gIJ4gWdJGHKItwQncoj5X/QerBXQvTPR10FKumPUQ
Hg0tdvZVuhPSFNvrFDaroMQ5dB++H9AFFQNgXUiWjXzM3OHlsypPU23kdtVUeR8b5QR5lEas+p8F
IuTmJY0A7QJic0XjAj0/Htlao9Y1m1wC4WovLiTfu3tgRcvQfnpNGqFvCRhhnmIi4gNJioGoCQNx
GkXympC5h6gYMJ89exb08+M6hgPqQOBXPid8D9Aj3a4+/QBa9sIVbqHevm8QF053jMYFuecaus8P
AUJ8YT1b7vLm9Y1GXPKfNLtZzkDeuJpm0+MZMdCWV2gZQEEJQhMEETKDF2Ar8uQeN50c+Vy0SS+J
z3g5xYK9f7MROn21fzf49zbmesMyAoN2fsUujgFVwMqcq0+uNgsdTLqOEYOlLx9UzBPdjoJUEPAk
pYlWTpUqxGsDgMDfI/b2YlRqeXxCo3mipNSPDGvrOrOsHPC+cNv9P0Xworpifdjb0c42k6q2XnAO
KGwaQ6FvUAhSV+cgDYl9g0L6D8avXYHqf4f1PlPPFlo+98zClSpG5YmSFGyFC+jmc/GQDngaxEzC
5DscJJn0mXhfLE9SKFsbFDxrjCeIwzcbhmRyBi5KxOh2ITNriGyT9ADOumTtHuhirx9KZPWM7pPp
bcsVdbYw7WG9QKUMTAGphpP6JQuNjwpgxkGMJX5bPYycmkohuQ5rKYaanWjrOTgeOmQvjxwqmiRb
aVVQcV+arZOa1trABwJ2OKRcN6DJdW5t+CSr47Pptj/cuNHiSj+FejcEdy8shqtRTMj91KhtAbjI
EuO3Fe5apOjSWbMX8g44o6FdAW7CE+0Lv4mnGiBOzxnDXwyJFdlcftX3kzug4xyj8cfYDk9z+qXQ
w9TyBWwjZVBXWF8wms9L37R/0vJcrPq4ivlJHA3VLDb0siHlDUfmKP4ulXuF2gfHLSFdwa11p8Gc
/eNChWupvHR9CX6NaV+m+wiSu4dbN5IwnSAAKKNf1VRVWt88cY8jf6jZQqwI3MGSPCzoqalQsQBO
OBjYC9yM9UfXh+kbRIoUFwISaZpRfLfsjtF8JbtP2Sofvwtpi4cRzz4oe83NkgClXKAEGgx2w7+n
2rssur/1JtbmZ7j4ZpQfyvjJ/wmVheAtikc0Qgj21sgih6+GYIx0HrcHf8D+pBMSYTRQLoBD4iVm
eM+FyFXRWJkqY1R5YZQqWNxL9yGdmJPcnvn/dUl7LdOCo9PpMcE93oHoCuisNqps9cVueiVoawEy
pyw9JH9tkL4d3LOkQEWFYSOU11lWZaM2BtRZdjoREclvBV756NaDkmY0O29CtMHG4aOiqULGXHG6
HjU8AaHEGBZ2oE4+fZ9YX5h+15L0jrXueXsLwzKI8+YLpm/Om0CkStN8mbvsEvLpoQTr2tx1pbjJ
y9a2/RmB21F8A1UWLNNDJpuaITJUNUMYc3Y8RLkISdDVriCgrByR/OC1m+LRGPCDwndvPMwMVQKz
fGsLqkG6fzu3HYBvp6+/9hdX69TOMl4/Xle6/oKhu8MfAbCInj3CXbwdzGWFkqwvlXEB4VQsF0PY
Jj9foRcrQC6/YlcX87pO+AOy3jpfckO3IgvwMEM7V6+fg69qQd1aAa6evQRs3ZQd+KO78Vt6jD0p
7QPL8kch3Ulof1q23Di7LCSU0dc6Y4qKK72/4Gi2+I+dpfMV+qNXtYenXtw1XoPO/s3j+nlPO20u
5FxEpMwqWHqiXb9xq0TMXU4SkR8IQRm3g3FonsKmsEx2YNmGPwaIAY1NDSqcMJKxTD3OzkJSARyx
InuYWOxKOInpjyQr2txMKev+dJxx1ti9xfx9KsfzwSpxbVndOzgZzPcZDJ+g32mXuZMva0/MqC/1
tKaJW19Y9ol8tqQEWVntGwwb0yyrmp9TX2HRTbgdZ/nzzNRqNGMWdnUucKI0oZzHlblbrg461myN
faubXJWn6kOuVi9vThanNLj/AStcIZuc13hWK3ZC9WsM3kltFatW37EsUHWSzIseWMqnq+9mP1au
jj/n3f5FEsUDdFg8KZBWFgv6yz+fuPeKLeEZ53zkE249d8NUpkBxiZCvHuDDLGrcmbaGNXdV7SAg
bx7YwoM4U+5EKFvzuR51mDh32QeNRn40bmCXgbgFoiVLH/KzQI5oxnU2qX069mjvSoa0djJdHV8p
LMEiuKO+OnuaXgMki1g102v1UJCrlhIUDT1uSEExxZqvLFn/mr2KNg0GE7FY9ebCnpCxPEkzvBUr
IFPhXmuZ5UDgqS+B9NhxsBqng+c7U5vm6OMLiwajZFL1s+rhSyo83GcvGgSzDmD6eALr0nIjQn6x
Gk7AUxGTyHhl+zZ5OLd/d3M6BqAXXRZocM2HzAGw178I5fFea9GnPv+kl5Q2CgT797GXygKBp+E3
uzo59W2eYcn0VkKGvXaMMffFTHXuuAU44doH47+41q5M/YLSy2W7WhLOc7L5SU6Zi+JGAZnkWd++
KOoFOVB6O+h3EETLIx5tSERLa+o2pNfBypaxPzFPDFOtfORF+M6V5mpZuriaunxEXnhoghM6aZWV
+Dd+sxe/HDyZPqj/4vC48mo5layLDNXPFNrMLlddHFmRceG610d74YWO3sNldMjJa79AXiSLcczy
fwy2tfWs86sSjr+NSs1AI663Pf0C9b+TR2VDl1I/Jz3Qxo9sTVZ74QcUVCJn9mBGx+i2DyLXQrhf
sSstYH4ah9Cz6GI6cCKEVQHCGe6jcWkZqVhdeqs3TJz4KhuxAU53M0zR1URpiCcunWog960UCeK/
0no2NVoQdy/fnwC/4h5vGPoJOZ1e0KGUHmqLRA8X9SH5szQe0BpwGcm4B+DZTAuwkQwAE7R/4eFr
MhXZA0fhmD9BOPCDCZn7cKuMM5Z7BkCqZBCqZJLVrpAjklgcOqkrIEMHodx63CsfIjbQcZ/7vV7U
jEInvQsEP/14UU/l6Cb2KodDJHoudOt2c2az38gNfVqR9Qrb34AAWCnsQm+ajCoWvh+mWY/acl99
otc5yvSf4eFrmgoFyt+M/2nl3PWmDDRw0hYiOxRUoxvJU6aiOMB5k6mwqXmYjipRbQ+9vEk9jHAZ
q4ndqsSU3LbEzUeWKfHWOW6ooiBwnlMAtQAR1hjuMRaGXM8OpCJ42iuvUjWBFNmAMsS2L0GLD8wH
vgkbJDpLTkxNb4G27cFTZZ+hg3pWNBSpgGMeKfc0ibA/8iLbxCpwIsnN04QE7LGadVAb4vFkAHl8
3IZjAI6XKnYCtZWeYXGRNQAtgT+PcqOhdVlNJ9y5aO8iyAr2J4Q55WyhxexmI2RPCuQ2jqzdIovu
zXxhRXH1bL9esR1qajBa6SAHPoeSjEvMEqEGMLv/AzNdgLogD6mHFkPTybJ9KWMBloHqOB/9H6mx
Z9sNRo6fQYI+h/1lINFxBiv9Btx6079x85cyu+ZAWMTO7VdFBKqDmGHR/KOZz2KfTnokHtJOZ2MU
f1iaVWepfVAEKSI+3z+hzJ91NorEmOTZwX+cOAJRVvLGQxSVYoEFt2BJT53sjsESjmIiebkttn8W
rMgOFgIEu2Uf1dP9DHz9O6I0HcCmYwj4IaQ/wj8yGoG3tEsEXLoi/yHrHfqfhNJ49MmXFx3KnPdV
RrVoPNKTF0Hu2DCZsDluZQZAomtVU9yQXUV3T5dWlXxXL23f2dxdN8yO7jamoNy3vbjZ3DtbXqhH
YnFZ8fQJqs7q5PporP7rJ6Dcrxrb97iC9RzJ83aShYknQZykixS12m0KfFvwy7ulQ7pg5VxwscRK
Te/2DwzeXyrN5095d4Xlipi98hFlR2XVDArMaXXtT9IGVw4yJvTzRM65B8IKhq65u/a7ShUs13DX
o7qmQU3G+Ycr8O+utkkaevnkR7Funcm3FmmLljzGIT0HHlA3Q9hVjYmy1wxoVDMxpfHtS/tIgB0o
+xwZkWKf54lw0K1o0JBpeBEFFx1UH57u6DYoUJgFj44muVBx3SxxGQYqg06dg0gtjXSwY/jQ0boL
IAmUyHWi83j8lQmr5IVK4vd1tAqD+cGKpMp0NMfu5MukVg1Xx1uxGZXgV6XO6M3q1J9KrMKgsgTl
NOhO7sa2LzUMbktFDeeeu82jaQp2Oq2Zq9gCxXGOh+DjdfmW14NKBp8jVKapE9xdGaIhkGnnwAv5
WE0K9a1n9eTVl0azxPQVH2qctGlt0PejkMc5WPO562+N7p2D96oh+iWgI/KGr+iYHqiuJ17V/bhp
/CJYD7tQ4+69+KfeSOczTO/JH4olq4LcmgNPGT7syinRlIZpN5i3tdkKdOXOmEUW/V047wlwslek
O9CJQFe9uuudk54YceenczftLnp+ks2peJugCldcGe+imF4BiJ8/wrTEMLdVrN6GMuVXsbw9N0+v
tsSfGLxOWWseH/jRKfU5J9fSXz0vlggadI+Hn57tq+0fO4/mHOzNKZtJOI520eU6YFXvL7/kKTmj
Mp5mQ7DhAzvbIfYG1/QMcKeq3yH5KR2Yh4sPEXXhboIkpl3dWjlk9t1duYYatorfDYDtd6RNcDG4
Lpr9W262Kwmm3gvascHGKvJj3k1evoXHmli2t4chjwXyUjbjmRDoRzI7zPj8thHn4e7UnJjeasC9
tezLU+N2wgpUz3fHr5dJB9/QgR3TW9u1EtdA0/9p+NH4zKq3uMQ2gmjovF6mFvUJPw4ZPfdR5wrp
DExcqEIWbuDQsAVPkAnudOdiXjSKtalbi92/a8y+a1L/luYtYO2bMtZQfFFQ0oPaJOhLeLJg4TQT
gwrb3ki8jHMWTMDl5iSdkTGx2crW4jpEDoogJuzFy/yh9SrImXMqD2W5TTBB39uTRrUh8P3cGmLp
8d9g9EexxChLFjJ7pB22NKIQzTNNnypWSWeJA4Jud6T3ceZsMdN6XA1tOzUZx2oYUD0OF+oqzG9V
DOSAm/tAA2RI086ghhkcI7K7E3GJ3F6EjPTxgz1r6GCfJW4Po+7Awx+xYQnru62hIg3rwbyFvW/Z
649Od2N81b8YpJ/c5jZ6g+nN+S0iidiU0/5pmk2yR2vx3Rc/j0q2yDdRt35ycJsUbkwjaZnxfogk
yxjktGvZI1QU4dDiQooGeyYRX5AfBBLIUVnFr4BWcphuItHaPtxeg6HtfFezHGIO/eL8ODeRxY8j
vXo4druNqZjUa9Gypd34Ea4ibEZ3Z+BsHe1oBtJ+GwiYLb31ONwLs3et6MwS/ppYj7mViiy2nXl7
9xn3J52jB8B2THMCgiqofl1zK42Q8X1eazOgm/Qnz5TsUS1JXMn/ADT9xIi4ADIo1eFF/3hS/KTE
1fMZYo+F6HYjd9cpIEoiGtL71r7SwjT2SBbKcdqXMv2qycC398uTNPFmCaE9uHrR7eMXKU1Fp7Ls
r1sp65i6LeopLpAHFMvfeB87jIb/s5m1OsEtqGc9bxq/GyYMNzBlLOgAUqoVXhdBQdj0B4H4SyVM
pjv37a6vhJccvvjz39MJ7Y+x4vPNFq8Kdqw2eHz8oCg9WlRMWUmUGGFwvVbzmDot8HiJ2rp21+NQ
pN0+mwTahRgs5rg0fCKvPLO977X/LiVnAoSoy7yQZa0GGPV6uMZEC4m7c9OcbV4l9QuMGMLZBiwN
+bRj7msjkCZWX/v14hGLokRsCvEVDF/IAn3YGJe7mMeXhW14F2PFNykPDikykvs0RrcYvx3sw6QW
o0SqAqplgKpT8evZdbpIo0AmK0RFDDSxDHrudDPLsom81gptrm9C/jr/NkXKovcrcnthGDp8i+gE
f1g9THAYXapcEZ3WWJW3s3RZhKHgu9kyslDUWULhUTUecaS9frRXAagqDMCsat145yrnkCK9xzKS
4gzx5jfSuYxjSbXdtG9aXDj0ZWhR65I/M19Gr6QAHcha/zKDHCPQtk69aWrrCvi/DBujw/fFErz7
vEaRaeHmcdUCJVQG7oSuU9GwmYlO/0sMHV6OJ5zZtnjFJUDV01GtM7wTcnuohEiiz5N2m81hlBNw
OeGfYB+k8GKBoVQ5JKp0p6NFrmN8LlQZgtW3Xx8Yb3DhZHJnpq/rssb5UgDTqwO5rmM9F8052XLK
GDLbdJ2v0RBuPxQWeK5WFsOxnYyUrDh4hJ2Ybgm5RlDDqaqNoMxs6x+tgd7OLwKB0EbFK6v5MplQ
K37zOVdcFfAv7+yMO+vBebkRsZGMeqeKZFq6WQULm3afx+4erXWbTUKCJjELun4Rcf8X0GovA8CI
3LXqnkHfr9nd5RayEND7GBZL3QH+qZklqqP03zEIDCgISTvum2VHUFF9igE+qG9X3OMd8YSGwSur
jUjBfWy5Nh+3E1Nvt0/7JVQ8LAm4lHWetJvbetC7uKTgMKYFiivAYmrJNRzpP+c4cuvC+hevEfUE
IcWQ5VZjf5I17DJQwNCXtH+DQmr12CqH5zugt/rTNtFsi3jJpQyDmAEAsrbnBU4+DmUg57/38bMW
HAnsMccE+dtmT6Y3bRGOvoUzLXVyDgZR8ykdA4UTV5DCxAMAOkpnjZZhTFKSwbGEV2Sq19YySb1F
7iqmvWLoloM+M44C6SlvreuWWxHMVl5jF36ejISuzvNHmIk3kEaePT1EnOdwJD91h/rzHU7PHM6v
z8WAClRI26cnUxOHrrnRZQ7L1K8towzCTo/BP/QWk3DUE4M7aXo7j5zp3NAuooUmqO35uxo4LbHb
06vUeqE4z8H1hfWry5++YJAkyS5C5IVNf7L2XFI4Xfx/geglMH+pqZAKtr8Zt7rDx6PmlUFmka3v
fKugAH2JWT+KUMKnRHpY9uAnwWYvUPKU/9huncmTtkyzyfzcpvK3opUUbylH5MPvCNzdiWhFo9gI
7qgBI1Xl8cMpriFuht8sz0xzqLJC0zrWUT+JewWM4V97sxRid4K59rWT00MzdGEx0M1utgpy7u60
X/aa2mJ3yn9jdTeJxSM/dq0KONaEXdauqsLavzk6PAbbFshMIZs/Yu5OHkycmjPBxjcsV1LqBwjq
tQfVzTJSG23M11WGK/jvm/HHazFMohJkrmYwiJ0950sWxnlZR7hZ0pE5u859c6HUdJndFlJMuUQB
5buacMVwsAz8pCAEZ7PQlSQg8yXMCfefckO1D1M8nZUOEP9H0ScxWjE201dB9fSP8dxtCVp/emLB
mzEfHBQPXv8kuAc1dTOBzRxl4VKvUCOHxrxCFKnUpJkSDNM1XHwp1sCcElV+CSQzrx05uBjt47v7
0sBlEk4XknsGy8Kvjnr7RtSzax9qKG9AWBmDyDGbmwPRB/mTzUFVa3r+2vePFc47zT8fXCQaDEYh
blPTLnykPr3ozTEWXRGvf/61Wt7/Y2wIIgqqJH3urBgsp8xmGIwLmCSo3gjCkY/58e3Fkch8pqtr
WDHxsXj1j2Ze1sBsid3JcfH78zXU8l9QraPCrMlr/jucs2bp176fNiGTyUrBbgLuaizfeUm6b43u
lmEEPOj5yXBZwU21Lp4WkXrsNbjTUIcHrG5ia60739ZYKBni2oq8ulWCVQODXUvKowuA/LJxhfv3
Ul6bIPDcdEvf6kZW/7Y9bTXNIVSw8e56uW52mEQij+2h/v/UWr66nEkCBg+YNMCzcGhz2LJsx16O
xWTgy+Hxuu5JhVxEcBqex3G1PwIdLScBA50AhEDoGrNw9xHDcO7d7bVFLws7vZ4gFsVif22k7obY
dtFprhPTpzdQs3BCIdq8xecy+jliUtGQuEdfKsugAAvPUailokhj75zF6geNV09sJS3wdznR+Y5t
7di0VcAMtdgu5M94G95WfmO/CxmgRFuruqiMHBrSURLHtdG/8+RyLv//rSst95bckt3OnzkIiUgP
x9kqfLj5evsuvpnpZRw86rFOt93LgrO28zCMfhDEjmXGOUZEzDUGDxckV7T2eNODQKDUF/3U6s0R
OlmnqI4WSw2qouBJocuPtILmgoF5i+6ASwsAlvysR95/gmameZeFHzwjm3pRVQbAiSUOllH22ecQ
l3xqNf8iXc+8/SHG9AiV7SrjFgOrwsOJA+1f3vtchQtl+lHJtnyKFyZZoL88lGpVDCgP7WWQvzcA
4kpxEOXSQWn2uJznmFa4yH2/SA90msj95LQAtujmb08Q2l9OHviGQ7Br3Tft6arfdoEUwz+D+ULz
ztMefhJ22BCwVBN8EXiEZ5F/I3xK/NnXo19RRtXJzosfYYZVaixIMYQUnmBi8BFCGr/T9Gggr3S8
i7otXJiXItuklAgKYmhHsnMCNZyiHP7PciUbi2jpLf/sKrpnXE5IQslXovnEJW+pbjW14ZJxxbFo
dYFNTIb2i6snbd1KT28RRTubzqoc/nZhbycs++0dqfAJpp2I0K2EYS3xVqxbD056jrpMoAD2Yp2l
XIfbpaWgbivXuVox4OJWjuMFdBlKMdg1sl114Mgi4yojvUhP2Brazp9g6WD0RjTnX4oL2dDp74Py
y+H6+beh7RUfklkjtt0MBzftQkI4waHHfq9AZhYvTzv2JBB3prdxtVC5Asy2HRWaGVhOCDfCl82i
k57ytefi44n7i876o8tbr9l9vwkRwsZOSm9bonnDNKcSaahgrs5fSLdKAc0/B7oYica97r2jXQBt
wff0SVXvFJ3lmH31JAXm17+keQeVMhcahVq/l+0rDZ+Z7YMik2oULpuLzELP1ygtrAgAv4nbRC+l
tfAPvxUHoAr6bzoz8hf3duURpr0O9+jm1JIbdCM95BbzOYIciVzWY6WqJ+NBvecO1cnStDJ0F3Vd
uvQOfe9RXaDlXeJBsS+xmw2KrJK1smvGFA4nfT4yuZkm+gXOlhlvfrJ+XeyXBlxtR4T9cMpHKUdE
BSMMjhVbOo5sezstDI1lM/j4/gD3zSaPOVAbXp/0nctU70oV33u2eZVFK1/HqnPtJ3vBCdRGJHHO
oPrJHqumALm4HWYWJzetSFVsf/L7mi/9xFLLkVb0eBIvw1yqEyNummp36o7r6o52LhRq39atyZNA
nIoG0+LHDQVuqRr3Nn+NoBs0YeF0pHbJBpKo6B5RwDKRQ+mvDrL5UCreth+ECsFYjujNHtK634Gs
ENk0J5uYmAHWwmSoThxTO0PRgABEFj6NmT/UElM7l73GXWnERbLkMHzJRM/KVdK+ZuFrNoGcIiTl
Nc1VhwLfFTWVyI/yNZ2uVU49+CJd5338nQxPqZywDcm+PhZNE/iH2kyhM0vdBEEKqXL2bZiWEatE
EWClOL6Ls2jW6IRV2ODdfyqNC2+cE/fCyn25ZppVCpE4gy0Q0AewtG6SZbYtSTkkdYmM2eaQbIeG
LaxR7PeNEkJ6dtAqJdxakSNULR7ppvbAsUpRMkq2A478V39fELRPLPDbntIakU7fH6t6DAJUn1tC
ElAfXxl0m0wRKkTRI3GmJld1xr0N8t9cd8KXIZiDeeJzyVhkxPMfi00VJj+vaPN/8D/aZNqddWnC
KaOO1v42nugP+lY6gGiQFeg3QWfeNAnfjDck2wZAL2Wu8Cj5fVCyvrzxYNw1fqzk4xCSo64C3lAF
hpndLAfsm9tkoieO2Io49itw2KOWVhVEJRBqnWHpVBfdBap0IAZur0HhuWGtvr4Buyhmyk/+t4QB
uVLtnaVvqCi3YBvkCElPGDHFXnU36HRijhsFTxqeAnwtbxC2DfT5Wfz4SxzIMUhjPxPLyAyBF+UT
6dVyWJ3XK+DXgEeTrX6mLU5ZxEtonXJrYym2VQrB3JeNLJa/K6tJ1M7Ao1Gfe05lqJOXHW0Ek3BQ
bfWLur4rr52bZYXsffbRPsE+ecjZJ7p5Sonq7pbowSJpqR95xGN/v1K8ZzC+HlTK6+/Etzm/1yvo
W0v0XgRgE2ZPKc5DBHW53YAdassXzLhoWM3qNAXYoIRTJqXxMbDKdRJHbbfClgzISZTK63y/oF2B
KfiqkufT8QBsgN3jQyHPZzH62ymSAXBbAUzwepqE/02H4+z2jRtx2tPXG9xY0GOcqIUZfoJBQi5A
KX5HXYvr+vkHGfKq1Fl+LYxARmWD1ezmSuW/LM95jCt3QFr1YizYdVocIgSUZt/aAmthGVRz51XV
oHiG5BSgXBhyM6wqlVg2lflDX2ALQBZrcefMKv2o5p09HFFjIsjvFxhB0570qdjqZhPiAj9Z7WTt
/lnOLTlKLgdkGOk3wRzkb7Lb5sdodjiI/X2dqDNaE63qjAJuWCCyIIZ5tI4hYOBV7J1IQmu5btcl
An6Ilnomi20b0FbCVqQl0g0+2Z2uPl4IgkYHAFA31/9dror4LcQGJ3HVl1NeVU4uxGfoOu7WQosZ
4/34ThtyKm1psRUYCCNjc7hxZDcLip4CtcgHPtM+fMGibz2LKkGCQpix2RkCtknGiiDrptepmfI+
c3w+AjCTYMn2nkrdh2s1XkOyYqlaiSCCHlQVknG/39IZYfPRmFXGlm5fy8odzxCGXiV+yFkASaay
flrUIFkQLRh0wuUjI6BDJC+qH5efzrc25iY9BvF3wpmBjo3baT2/zVJohygiReFwmmslT85NM9oQ
dR6BwhlmqhZPqYLV7iTtVgMrgFvn6nki4cKVJWuWpALDf0FsGr/bI2z0qrOzTuCJ5Zk27tCR/Sur
2HHOsZLHFsEcY0pnLuxZyLufebPawQ/y9hz+B+Scs2cTxWy8PFwBzx4sKZlVa7ev+0byeycxoFJi
OTqdjJ5kO/bOkIMQS8qKtL8E6HuTK8QaUAyMdVYi9vIfaUte8UNojvqpN+RrhY34FPohgxOdQ7fg
AFZKo6veHC4nN/5FoTtYuNAlUjC+/y5ksHzaIuRRbLEVI81uw14zdnyYs74TBpmNVJkNwj5BmqdZ
mcKiKclBWx8KGkTGGi62NSjSSdn2u7vTj6jbBEfgOYvjZvcc/xtNlrPtLJSLUFPYvhfHn3vIjxsx
ZUaI4pV6FLrUplcSnpEyzOxanpX6M8A+ltsMJydpA5HIvyn1BAG8LvoA7DPtDhNXDB3lyMOnKoj2
C7c9hh0iBr3fHyBFi0aKL6ZgY+BmopWBp0wufVCmFXGzWKgbAAu2k7m5bDlDtysSU8521VbiKWC3
CTxsNUgC60RC+OfjbPsr1UMkNeD7EtBxdSf8h4a60qGc2OXBkjH9xmfDoVO1OzR5RLYh1w8vG59Q
U31F02gf283SNEIJ3HnFShfqYqp6H8B1VwpeZYww9uRSIEbObXbG+aH09lKnyhtsD1Po4us8s6uK
2uIHuSOrdOFYzVp+LQ87vCXim2Gz95B0r7yT2lfih40lhwc/xdbcmekICVfQPymlKH9JokZdwuR+
y8DQq309/f/ttVqDuurDGAIyPHwCnnGJD0ZhvyIrnAHoTJ5WaL/to8rZ+SjPbNfPo7XA7GjLcY5o
cuGwPcsRboap3YS4oy2ilKGyNWtH0RPuY4te7k4lYT9RCaBhMtDAhVjX8llGk1QvP7BFQie/DxNG
Q5DQiJVR5UniEMSN48F0qrlt/lqg6BES7KS6yaAWavitQxCUNOVO3eO7jQoRXeKLHuBbxjQodqJN
wL+Szr0a6MGNQmbn50mxp7IT7IXwpXwQmOj62GQi/ZO6Mfk2ZqiaOptql/Pa8fYwIlm9Yw3C2MIN
2Tef6WzfrqqP4UuDp+qXuiueEBKMAq9dvKz0sGRSVE4PE46PKqvWObdRM2msMFaVQlcUGvqtGYWI
IBVQg9g19K6Iqxb06oj6MNVhVxPFg1NiW6DA9pjHxg4mC9yZtGKUxZ9xpqlrEoTVnolpOD/AwpU1
Ho3SuSyVxkgb+wtntlBuEsoeTGLPfs6xMcPYaW28X26wRfiqLtR6hnwHeqhBtXfclGOhBTn/8dqd
uRFcyYyT+QyKUoxrHBUYMfbamOLLSDteVZ/yGIUb+K84h8M8hD/4kJyPsTVIQXTH01YzOR4O2rPM
uBNJwPDb5dWhxs9ebwzEXXTKoTWxPiYLMxvQJ7+JdqN1NuOvPUUmB5bxVz/d8fnt3JUTf6nZTxwP
kyLG7XWmHTsV3kW6Q0SJc6KNlnD1RC3A35SnoMatZqVW1K5+FDOEZeoK+NWxlYWs9lgCg/gEf8h2
9euXErG7L6d9NipDsXaqeJwXb1oInCBbQrJfa03qWWgKO46AiSK7t007xyWvtpNzHoSEWmRgxXsj
V44jzKroXlmD9eemYvExbEwDxHZAW5MaYWHnLtbyQNBZgvmhxY/mhXJY5kwXRezkDwmwQsmqJs0N
lIF0hwg1H/MN6LY9oDbVcP366t2xFQ/kqprtrNwfzLeXJ52gSpHOASk8Wryi7hTzM4RGUVU626VI
ShRC57OSr0nS+PUoWIhHQXk/AzBaJa1/ibIv5b0ER7L3+AOlzRGGHoSdeEhbRYYnwQmFa2elwQAB
SOoLo05JuYxZ3hGpIWzAwvUTN80GNiEqeH+5I5API3M3AxN/OlmIswXSKcBK9UtTZBqGAtCwzBAd
BGCbS2kvNDKAhtJqMZo57xZK/bLbhxR5pEeZ+Ykf8hGyfbMZiSGwjEihdU8xJyiEQSgoFT4ve4yK
pQ/Lwo6eMis6dmU8UlX1jR8riLfJ4241QMPngrcuxCc+BNOjjQzRt0UdhJzRPQ7a0HT+lYPIXE6z
q9e8gZPaEadgsMmZufGMFzN1uGo9ZQi9ffHMIvcayaT6pHBlI5sEVrnKII7BcAm+ggodw8Pogn71
OhvXuovhrYoJ95KmpP5T0+AAoo17PkG84Ljm5pBfbSpRjXv81CRQmn13zuJDlh5XGZAhpQubhFof
cxROUJfL3FCM1H5GB3kGrgnEDXkzkPKb3V0ahcu2jKoqYJWPleKjYERTqzvpLEHW+zq/c0lzVKNP
CPLCjKW/fjOHPImm8lP2bHWjIpO3r1NVSsL6KUljL90qYwjN/EX6TyJYhpFX1gEhx90d7XU84t5f
MRkLUjvbX4sr2XTYgFNkk3fMoLMRaDxn8e4TENWJ1quWi2bS8q5pfRNSl8k9Y/1ai8XMWfqX9g+L
MouiMt7DrHD8WUTt0LG8bbvSq5lrG4jVVWGHaCIw5fYk2Np6emytc5078hmzJ0vSEO+DdDGN+PDa
zkvp+LroAAn7i8bpRMnWKzdtYQ85HPOiwshmeoHfm0JCspvNG/H1lui7KbRnCVNlhDrnFqjPNCpq
82qP+yMLJFYDZhk94sm4Q4kq3Dz0o7GevoDMNfj7Nrjx1l13CMftcAk2/8wLVid68GACzNF+KMns
yAsSXXtf9gnhIIWk1KeMzgxX0WgVTQ0xjC7YuehWIgJRKm5iTIJNiXtkatT6TKRM7vmANkblDzI9
vBRJFVsXZ+W5qpBt/CW7uNnRK0IZs7wUaSpNH7+a0IdIV86CXPne/7ur2cmmoeOO1AJQYF6Lfj2a
XGv06LfeoeyCdrwuGnN/kGUs3KokieSwcdy9sBMFJORNW7X3yd8CGKwSo4MFarO80BV2slL0wVIz
c3hbkuJ6O6g0wdQCTQCbnSO7gCRWHuRyw5103ao6Ko20jyzVTLK24mnEMJxK47z1nxY8iYbvZHl0
9PmwmaLhHYcLa9kaCeB1yCQZ2N5K3hjhxOIqNwD4QXBwCsDD6z3hOf+KOFKQn9eIvY6a6K/fLIq0
bbPwa9B9G3nX+azduk/baGm+kHSVxYZIjgXH/T5/2Wt6ByM9gqnOiAR8NtSsolsaSJHF6qBeX3mI
db5FkMcay41UyQFwBThYm/oplFoj9XJaD64l5uyzQlSLAJmpAO6X2Z+vpdCjes/3PlZV5s2R+guE
iAi+Y5ID3lQh3uBAj8ejQF2gTB9qnjmUvuv6rKcLaFr9NPRTrosmMSUaKNiYLkebn3AlKlkZuYiD
3K2uAYsRS0zYyfX4mPj1Mmi6eDtSAInPiJzCArmyn75DZmm+2t3c99ZeU7IWimBoolVQ6BrFEqVj
H9LGlJbR1JcKP+I1sSrWJ6wwnhIjK50CvxFtFYVi30q6+EkqPpFt0zQsLD72PMpHcyqR1NVxZIdM
D2iFS3YJRlTKuwEw1K3Bnmymh4SpL9oMwhcisl/qD+WVp3BZbRq1oaCeFPDgsDlOdfSwiPS6i07H
vb9OA0toJBuUrQVtaLdXjSYX4YJQJhgBL8xytr6lg3KrnFLM/WFIuWAaOUSDoVvBeliGfjn2189w
xw06Mn06E8FttxFTNxpPUejFGM2A1tYaHrjZoOjuaTvEuYPAvXkysM+4rY8jziv0UNDfXTMcf95Z
Hex2JaFykBeJBuTQ8v44DbqJpo4Blktk5igzY4lB2n3YivMOhDsorAJ8UYGqi2NNseBQHSHJv0H3
vI6JXycYY+8ZdGqlJ3DGstqKdvK9C7aXE9gVPUCXVOI8a8QAYKakAH6WOVlxSa+2nSB2CFh02ybh
/LcKLrKS1AyJraijOGhTKOLdBIpMNAjxm4xsaXGmuxmzZZn4bs22spGj9SCaMjf8F/xTpYF/tm7l
nc2eAMUT0pTTr64Tbodt69KETebet8baUxyN1apWR73oTxDdx225LtN3nueD+N4K0fQbMkQ8Ac+G
0d0mdkt/yZu6+rHk2g8FJzpJ/4ZIwM4vvoE4hABfYtAy9WPHN+RA/BzksMiUCXgF29xeNYzHQQgI
oEZfdzV9sTjd8zE2GPORB782u7ydbIAF/Ya6oXAbkQhOqnybU1NnY632Jna5nLG/NF+eevHWwJXn
Qz8uEL9n1Z4Q4bfBvAqCSUqTQKW99s5r+BScEh2zHRMTnX8lE9aBTNsswZ8Hck23Uwc928mXuWq9
OiP5oD1Q38eutSAeP2l9ep7ZyX0dYjCBe6YtTCY6+MjJkgNPnCB3cne5ZtQcg55utZAnFDYl3B8b
kaGBIvsreCD/dtDeZmNCeZeTVeQ2nYj/YGvDz07+5nLz+ZJvEY9QRkX9QqVxVLhW5gqf1lXkvjIr
ZgVHnwQuLJdWS6HkN5P3SNMjiExAJdg9bSewZBSXW0w//Oy6QBSR1dKQJtqVLGOGfyCK4YveLz7q
pyh457BSQa9Lgn6kVVxwL9kmA2xJ7KJ/NQgsRrnlJy3YAhQDzWEcDkcd3Vvkh64q2rP3iTp2XkIL
uNndLjvUHnPZu1jK2Ub4dQJkY22rrRMaMO0DstoPFepAHME7OtKDxLmqVDjkcKVQxZO1PTUlvr/6
EXf/LXBOyMLTRa0is3IEkX6C5ji3DZ1I4nl9hZknfCeaTLyjL5FiesEPqLIN4L2+WU79oLU3QgDc
6PZ1OYNpAekOaZqELfFTnEw3kbFj8wwBAoF0VZpKSUufFx+YnGuFrYU/vA4hs3f88B8U09dqiGbs
LmGWgKSAQlB8zeDAjAjEtDlNvX7N7v9EeOPJm5bHliH9yIxr/PmcmG0QyKotBHanCd9vXeXK2HH7
FQttM+jmkJ5BFQPSFEJg3y/0Thx80B3aus9Fl2yxvLvJJf1k4Q7fVqG9Q90pJe52doWM3qQ+RiC1
nu/WMeM/xH9rEL/SKtmYTSOzq8r+DHuiMj2qWR3gICTcdevS6F1wE4tAVaDQ3VdgW2vEQita9fEk
SuPfD92y4GGl0tjIpLUPthwIwwSfTuXwCCjye8U4XaxkzFsL71sNJzvsWKkOoWtoTLaSadGW79Xt
cYUGPmBK1EFnNtdxWk6dP9cdw72AOV2ALWCOtoOrnbDKjn9Z6hX/9uNEXBDPAoEFP6WvPzcjzcgB
WukLDhrxOmRLcl7okg7VzeNyZhi3mOx409j60qEVgzOnYNILzqIy/buLdd7KHaZNmDw8RHe9utph
3FEKd7ai1XrinvGFzs/erijpFYgFU4+sDNXeo8YppLcuHEiKNM9Pc4P7cgJqNicAI/Qbq1rd3pec
TTIZC/NWf/xlr6EZjkl3ghm0cmF82dNya5zJuL0ngQeQjXaVwxTdNCzDoaoCSnxThyQgjKuCofBb
zBFORH6NdlnlETD4r+XhewwH+PSRBrlDwCmPUa53DJp1JlJOqDax2a7JvXBlPjX7DGvA0gC8jqCn
06KijNn1cYKYO9UwkSQ6+aGz3rJs+FTUV0o6kkQa0S/INRv9XAJT2qoLt//MaFwlPg2Q3OGRWBdx
eqN3wJoT4iFx7z7Bb/C6IF4XZHqSPmKp0d3DjE87Ov635Jb9DQlM8YwjL7f5vG7euQZr9LjA7klx
lL0nWl6dO1shpBqMJ25XJpVfhrLbx6hVVLrRv0alSPm1vDWhn4W9KCWtrIjcxjoZKZe98h18um7P
SH80NG7ro4ZE1+ybUltCkgUbtnOxmtuFHzl8susoVfH47Nd3ZMaVDBcQxm1744Q1WIKVJ6Dji9bS
4J9PIvFMPtci1+MJdKuEsYOsx3orb1TB1aTlzLsTTu/K7bmIpaiXdqkedBlcps85/VOGtHF+qAUg
540gXj9N0zDg4xcJraLi6zBr1oBCGkq1fQyJ5XFt2F8GO2SViC3uh1oISrasvwYZIGQeD9khSbEu
HlMmoHWzdhAlJ8OUcpuQEr8Xn+cPTQ5zKmJsrvJ+emUK+9sk2ddtnj0n/83XoD7f0DTHVbuyCDiP
0UsmwTAy8YjoU2P6grcnX1osdl0jkCS7m1b6WXw4XTkeHPDlczw3F4HiONaBDRVHkLI3SWs15JC8
4gIo5gTgcJ+Y6TKt2uOGKEpvRemzObgnE3ukvak10hc3AhgaDwbQ/F0vxBlQVIBdpp8XPZKbTPbl
GwVA0DuQL4Wti+R59TxUKnfzi3t4ffaHXPIHLq7OimF80n5T2zZletZEg+2GNxhFiTTk/vXTSMfe
pufZjMkcK9J0PVzBTsweD5Yx4NK7TJmAgOFoTgQBslQXedSAWYkKdsU+ClO6+CXBHcxqsGTc9oy+
F7Upr33zJmzMgpgbr04JuJjCywCuf50FtlZA9YIzqY2Jk+JE/IePnbaykD1YfKSS4xfXJ9dlAOiB
isbRdBz97LIoOlXaLSGEsxIjVuE8yUTZUR2oK5XkioX0r52sJQdKJdQHq6z8fVEmLaKSd7k18icG
DRoXLOt3mqIMT5zNxDLIleXAz5UtTL++Z8gMy7aGS/OiG3wqYDNm7B5tfD5WFUh+/3Hn8uEhMTFW
+Z7daXmqzCiIPBQ+nyRvv+RhndJ5YxWYyTBFGuMOazhn+VQWUf2G0t1Eoh9F7p+ytAjXkX+PKLL7
C1ZP2tOHi5xWy8XCeGfAZtye8U+HCgrPDTIHRtUQKfF2Jmq9Fng9UMBaGqhONbTRLUPdqtYGVoQI
0aNlGTaf4zK9ib7Px9kwj6L4NkMf5YBEl2yqVOWQJZzWHMdHVrxnMmH1iJYCecnQJz7fBIcqCPRh
+Um7ZEBJnV3kpJ0hHgtamoSrka5XHLyrsGQbYfnVeW6GTl4GEwCsU93HMi/ARt7g3VKzx8d2v+Dk
50B4LlG2Qp/35iTMiSwuySTKz2gXM/wSqEyiPgGToigTqycU0Zyi8FTFPnPchJrNzdyIsD9bvv0J
iovbY98sEF6PM/WRO7N3Jwm/wI2ZR5CuSIN1IAd1PpLHrRxX4j0Fq7VJO2EewrrpVIWXl/SwkGtl
aTxWz+7SlqETPUTcvKBjJVhWEyTkLQTfC6BDZGKVBs93lamc8sHWTdeeI9MoXA+ls3ue8z47zsAj
RRSnVvmOtlJiwomxE3unpy7CdinEbAcm8uJo/VVrp2F+kc2zlI1VB5Fj2Ae8eKjkgLHEVZKlF0B7
9k3K6m7dZT1YcWZH5WjBTT9DNhn6FR4I+RJODWrWsr+LQrqDXXu7lBIZU7UiolVQrk6wa245yee0
q+Nl2J/2ceW7v4kz4AyjpWu3qrgM0f016jyozqF6X0RHUGo+vjgrFT4rJzCb+6BAiyk7laV1h8WD
TAofOaxbSI6eeS9nIvelrH6Rm+eFGVxO+mMuxSuU0yQcWUPRsm2R7Vcj8t6MvfFjhzvRwsLNN34p
R6mxHAhAhN0uTD/5rJoploRoA3Vi4uw0jZwFLiJ/+OvSZc9geLO6Rn06oYaVyZ+BUUm0qrgLzg8N
WMU/tfxMCo4QzE2SAy2Ot++va4gD9QrjMqhDpZrDQZ0A3XjWsudll/Txsqj/HOnq69z7uNu8ZJEc
GAxYnyA4+U58ltWqud35NWXvNDeHqrb7Tvp8r01jkTCRFCpdcCyhk7TBwzD80swGKKhNUSsZIHrw
X/rSCr9/uDMIm++BQxx17jod6E0c1lHVawBXTudJwHIrj+nnw+1dAOMEiCfOKfzTqa6N3cV571fQ
fR5aEA6NM/ofEEeyP2DCiTCCRxW67o2fMFM1gF3gzM4CPjoMzhH/i06MTOy0+UObkaeWYGHJ7Cn3
RK4XoBTaj0/iQq64d0GWsHNOd54iGYWdqg17hQVIzWVU9CZKYuVzpNTBd+T0sxHV0WtsxUkKaDJ1
DWqu53TmNBHDHIs5wAsWq06QRzPbCIsCQ1opgwsf0qxFI6bfaoTlOP89dyyA++a5Em2LfXjryobd
UIylSOSpTJshAoy4j4zXom0y+8nBQGxArDsstZgts/4mV9w+w1jqTqb7n0FwdAJ95BRNjzfoEcc+
TZzigERbZKNnserOfS8chjtGDt7OP3Ysse/KLc2BmkjvXHc144YP+ItBlWCbipbweL8D8h/uSTZG
OxXAT/EPJsltC7vWnJpowumxstBxYUd+dep4UAq/T3byw4qOOcHnGh1ezAZOrGnJMcy7OTvmG7Jm
Fun+0MEEsP6UXNMcObH/CZyuB9DpY2HcTMdd0NluUQtwLeK53HTz/JUwLpGr2s0usBkASOAuUFp5
jRH7FK+oJHEE72NMrJuNlj2dGO7jVhDEcVZSfyBbD+jzDr7tz4RQO74bcst1SLnJQFFYTt7JPhlo
dmoL/JcQ2Pr3Z9qaW62Bk8UGe8Z/DLY4+fkJPElSm9IqRjYpoeZMzeDmob6eeavCe05FCb2Et0hr
BQ3fwXdfx3ysvxnulsvln91BJn5UpdRQYrvH7VfKstw6fZ7WlQAjt7lquInHtmtHU1W7hNvggtz/
DANuATce1xg5rMRBFzxvTsYPYo4VEvOdxqutPXX9MQc6n+jQyLcIhspZO7C8nMkJfI8KS9ImVjjF
5o6abAXZcimvqOmwRZsPxydenMMvUPTLxquD6qhhxKpomiV1RUPSGnYUHZntFZglV2oxnnIuuFHb
gX3oro3oaAdZ1I8CRtKeqvHDOgEYzxks+GmosNxlcw1lpkjvNZNSINKvvdoVBRnf0iPQgadU22To
FHEoXR25Nc7NFvuR7zzYyvHikQf85hDMYo8eOfL07++6iqFHLC/qmRsdMPLGYaNG43xig3tzO6x6
iydFUBZgahmL67h+j79YedXkscGDAc6WW4Gn+vfyhlqBpGn6K4eD2WD5U3fJZHySDpk7GrUMMeKA
QkAQ27KO7E4OoJpxm1SjUQkVGUGXQc/R15gPMQGAS/+MfTTM5rKGBIlVGOasLfXQ1+WHYEHV/O9S
IfuyC/VHbZIoJhBYYpe9RYXIpjd+AOlsa26hVI58SGffwmMjUkQL/wCY14F1JRrIlexfgadhcaxV
idA1fz+AuvVOhMX9ueKsR27PixSInmDSc/00ryQW5RH8IKNyxzjnD36bcI5IsRFkx1O1ynHjsLS6
+pzJFFnb3/R4H1l4OynJK7yPLsnt5Z138E+U2dS/C0/0d0NQSr/MxhggRvkKtSIbCIhULb1Ffa+P
lBP1sLX1VDDsgmliZLGMqmPEyDbG6KO7FEHzfAmbwJ8nO9/Fuio9TmU05OPLbabbOxlzU9x5U6lW
hjoEOAuuYQchN9FKfHajTR9BCZya1aLCVhqT24hOsW4RwT6h8yRBkXgATYUX8bLBTn9QPZP1bcUh
INsZ7elud44nDSl/c5hzKhuNzMcpgFn2yHJWycwiJRVGgIXNlyUMye1YPP6MEDPwYXWxVYI4pmcR
91l8Ff4nFulq5ZiimmAOQFAgxe1xPLiPChXaWHIec3Xxqzz2JVYy1iG1JNuAbSOIt9SKY8hAnf2P
DUEI9Q7K43F1X3orvngORgFTuq1nbvr0nECieNaCHQj0qx0nuvZ5ie0T+eg8lWpegXQfnkOkMecK
ZJ8lwaf0nEiIv9yBryF4k4U9CnWNp/9q3akZ1/2Hr9Cemt3mRtR/6XYvlJPJ6zSzARdL/N0xaYng
mIGU/Arzaz+tCnHsioYP+1EnF6AQNT43PDlvjizo96cwy6sb0g05ztPmSLjWwEPNzPAhHCz6oEG9
MzwXq3+QTW6afWhCgI+USzX7d5rxUxGHWdGROolQxZPFZSj9oKY5vUc86JqeGj1F3tj1OA9zg1YE
gn1PjocNWgLUR+0/MbKqaC/bjkCKGcevtt7N1jb4Fvt4IS/ANXqu5hscAnWf2w1tf7/g1TuY3y/o
qcCyCpz9QAZ0iYDb6yLR41yAi2lcNPiGkMZDXGOBrjLQmMErpPCX3KI7x85QA72WH6Ha5mDVRwOI
x/zDeD83QItlg28SpnKLeEHpVoVjrmYmoaa5uppmBdGYtivh8PHJtnMP7Zz0rb42sgfX5dwolmTp
nWcgdJOZwt23/yDkL1/ag/uTgNTPhs+aMCgzrWxzURuMC9hPW+lDv3LBToDNeKcjKE6//QKJumd7
48lzDqfFI1x/PvjVpx/WdnF0kFFbZ6VJOEBiwsfddutpT6nz867bLNPo1tjCXFUGadewMluvj8Iw
iGC0MQL1uXkAqcelJAW1DD88a6WvTi5wp3o+ZiqLej5mKc7CiiiLzsm9WgyF7T2jJZfJXXVl3KFY
gYyptYAw57Y+jv/2jkhbn0BPVoUaMbCxsuROmSqlYvrxDIryR7zidS+L5m5SuomwbZ2Jx1sis2BZ
c7d2T222biHYwkXzpaeXnmswkRfMOVu+8MBIl9P3bOeLs1ZMBir7UoBmbml4/0PzWruJpdLQBlg1
7suIyx3imICaDw+7bzmVsh0UHgP61BC+464mbsqKVIyjRE/dVaRgybEgYUf8e8xs0j8QtqkWwV77
GVDDXMSyRnA0EVemiPCTcE9ywhmGR6Ci6itBydJL7YHC1FB0MVG1VsXdM3Fo0uYKcj5fRN1qTNk2
qAafOrR7204HVMSfxkNpM5qJLSHS32Rxs7UAQaUVD4YsIoqZ9kGIYe9uUeu5iK1Yaw7l0qpxOp0l
S8+JZhAwXueaahuiPdpRS3Yz2+EpOnVpbUAswvGVR489t/j+lXcGb8zea4bplvKYSirIzpS9RnND
Vjq4llv9W0D/eephh7cOZvYzWi2C6hHoj+FQxKTOX7qMEGvVAv+EbLO08512tV9H8/Gji4Zj3RA0
DHdFRfLF/OnNjb/MYNBorTzLFv2VDbIKznaAxfIu4TMf77JbcjZbwiNKW2ObP3XklLSDI3q0Cx38
N+COA0KMP4IFV7MrznIOph6lCY3Y9qiFOW1nEwfgWKRKeb4z+8Zs6LKvESGPrXrILXs1za/wS44S
1jZVJahyL0J8gZ+dxLFIeN1pl2oAmSHiGwYpDBkmy9g+i3GUD+GIylV6u/NIIhxwgNMly0NNhoUV
wWIpF5Vm0V17yJPpwdci9OuKrX300dsxSUyKYKU9FAGEtYc1/+fraRcCje5fbdMGUrJ7ZZ9YdfXy
MxOcWe/9UoOaYWoMje+crM2FhGySk8jPYbE/FR2TpfS/oDCdBKEyUrsNII/6L7S1qHEfXL5k3lbN
WHPF4wa4B1YCOVg6bM5o09LE2YfZUfW47YJmnKyLMzt9BOPg3JjBRl3/rX+HYMmntcNudrmGoJki
B4yKjPey3b4MsvMPM6D0QTQSZ9NAcJl3NTXvumavwS5y7KkniXWL+HQBTUtQXypgIn7yE6obScv5
RlcqPo8I60Z0xIO8m/LjGX8o5GEEKNvZtyW4U8OLDlahYC7iOy1xztHvDOyFnC7T++vwaoswUOjI
HQed9nc+5s3zdjICgGMATLY4WyRjvPc/7P0P038sYwiLvQP5ZGcXtrFXb8n2doQB4HA8081LUhf9
IiQzCSZfP+vK8Sz0mFB1ZYazg8oD0AgKnHg16HxCCGqRqTkfUhBh5SJ/tFGJ+XEjxdfF7CSA698l
kM9u7Z2zCzv1H9+SNcWl2Eu3Dq5nkKdQzk+m2zfvT/jZbt+FepPM4QtUYcxRJru90OEA2NCn4Qce
8b2OoTMA0quOVMlNhhFPXysCx1U0yJT5XNaKCH4+ojMbOsVLqM7wYwvZNqpjRXfVe/rxvdaMG/3s
C+sF/MT3a0s4lgIzfWtQDH+6ZCzSvXL32vIzwuw8d2jfGRSrNhx9epzfiwpJBFaqTaCt6sLhvK3g
yCk82L3rap/OyNsHu/6cKOKpVaiB2K3cCKF3QBfFxAjdvsaH5Q0U7H6BUw+DpW+GCwc040kRuVZT
nIDRBi/bPYn2p/SFvVQI+FtiY/6ZGS1OqVJWuOpneLy8M935E2kwmL4VMgVnl2bS6PGbgBu35HJK
jr6EI2Bo9uWJpoxhJ3fOP2k6deCHz/XiJidzGS6yJOVp3vXM/Bo4OHQVjyXTuDPcQiBmSdAikL6E
Z2uZVJX2xLXIF6WntZ6HY3NsrKSj+SKpiZzw0yNfjP3NIJk7/O+qhUaqrrMFfEY93KdRQRIAL5wb
5bzvkaPh7JW7G/U/oEmjntg2GzW/8izgviqYyCwqLOOjEetEqx1qpJIS32/mpJpoLE6yQt0k/fM6
6+CPN28wCxqy3ns9hn0EV9aUeeY16QecZGwrF9XEbJ6Bf1x1aXDk6KGPW6lHWiplsoM4wU1Eh8DD
62oqy1fvqcfkuHcwmNm16zhSi+atVua+GZmI1cgH1dptsPG+RF1yln2JSLE0aG8eaR8iBFyRWXNO
1E2DoEEXqIlQzwjkRZwmVGNHTzEzMfeOlReXY7UeVVJmHu2DqjP4t7uTg/ACuB7yi6wWQ71FoQKI
deLzmPjYjZRtKk1uKS3A5x0QeAgTlGWX0Y0ncHoqgtIDqqnX7x9g0HZy4rlwRAn7yMvT5Ws90pZe
F5VrOqmoGEGpfEl5G1sttOU/zdF7SYT9XVBRKrXs0ZeDgCCbOfQKk7yapl6SBFcLlFKjNUZ5CwKq
y7nfPkdVWt+f7RYaMsKxjB7QKsGvRXGClYb1J/7g9ms/imj+YjFO4RRMbOYvtM+wsH2H3NqWIW9x
lTA+pww7wRzd4MSNCrp76NSJm+vhKAWjI5vCNZFx+ssQLIseap3f+pCpAAGa0mM50gbYBkf30/i3
+mqz9V5F/FPSUNi4k5B0PFcsO2JEOuBG3PkzfL8eZuWlSA/Pif0lIScJeMRT3uZ6zFm505DSr77o
YDBUoIUbCyNrNv2lKroYwnJQqSG2/js4R/3zP11hI7HboQ2pimo+QNgYQSHGfnwuuJ3cHgNwTSkd
ULZk6Gu7NQb/fzf1iS1LFc0hD8fCTgfq30mRe053cRdTCxVLM/pt6oLjmZ8rCnmUWymSSizfqfrP
5r7DYyKMTxQN4i4SrGsjj9Q8UjXrALESZ8O3UzjR5qUK3t23jVW0U7tRxV++5LBb0ogA8F2yCPov
4A4xYyUEp0/MFNhUpYsN5aA3McLqZP6lUR5lJHHQ4Nj4cDwcSkR/hw18YmFDEaWXlfDT5wLSQkiy
qDwuAquc8JRJwlJcbt9A/ZMFi2FGrrTaodwSqeFGK/qKUMvF9XEXezjbFC5cUP7ZAFOkSb1l1yOP
B9bB/oarR3BCHFkbq3yVicCLdI+gA/nWkj8V7QlhbB37Tdhuqp+iR4V8mT2vIm8b1Dbp7Wm2UFN7
WV1mgTavsltTm7tSB7J2CzWyyMIjZOUa8eZuTLGEkQbMR34pb6m6k4KTPbqRwLE+ccjRokfWSsYG
i4OBnK2FV7XrGDRZnDlR4Apo9qMdeYHPj74RlvEE1nd/Pr+gaV3UV4Q3tYWBBnLGYpfVsh2kSRBk
QlYBTmCB4lW0euOfF7tOHnv5OF/zgX1FB90ynd95ONvSzV6d6sPzQQnRtHZ/wLaqpyoYSuoOnFRI
HW27kwUMoSM4lNJYCRKqk0Gkc169Q5siFNaROTkgszYJZlKa0opfOasT9s35s7Oh+BxB8UbPZRpg
cEVbEk7zZ+B010BG8AJ26jS4NB0kw1hFcd+Sas8fW6k5IWIGvdKRqzsT+adFM5zslgFgGQHo8ml1
OYzK+Sh4nYm9/sdE4MAq1iqdpcDkW73XXIYRKuxBfKUYx+7V393WgvlkSqHKqHBpv7tM+z6P15Xt
fxJQbRCPLsoUSbVe4F8Bf0rVD2RBUDM6eRglMLzxkxc04U3REOs9JCh4rFDZp5doZc2U1DJgOgUk
Xks0mIzaAkqyFNQX06Hy5ZlqmIP+xbTDgnVWEH7hVDuzkVEByCflm+4CVGPl6KWh35XobwYCGtD5
ZmzbQ/jUT+wWipaJK2u5VKchtidVxUc6QQ6F9ynYS6u+hn9TmJ5BTZndkb9qJ/l++W5KjSH3rxBU
L7ACJSJrOCOxM7IG4piWY4mPq3nagIF5JEwsDXrUp+4mz8fi6UKagqfXHkVJkd7MfVl1GWJtoWhL
Zsgmm0HUusnweFJzsax1Dm3Ah+k6QsQ7joAyUf/T062W9BRI7CyWmXI2DkuZI4LWOEruupfCXsKH
jJ4ZjlA+fPouYhF6lL+Evp7jkc0mNA3ZjZAy+uzTFPGjeMtfozv+O2E7AYrno7Z0rR8xu0FU1rl4
vwp0hdbIZlRc3obyXAyEGvUpyCAOt7RIlEhyBQVMht8K9Bvt6tsnJKek4xfa30Tmxtwyqw14kgDv
kgckQpRvoN8dNrl9Bk3JvPBHYmOUTSZg3AR4UfoNMyvun0sx2AzCAVz9GjgWiQn2cLziYwkgHQCh
rwnpkpvJ11QGz5yqmIxFoN+L+PX+7Ynfi8TrnGN0bR5dJ64uapMHXaN2y84DUen6VjI/+jjkFR68
mUJflObPOwNUcABSXeEThrB9njFURVj4mCV+MIHAhR/1BUw8rGGQ/m/t4GCJIqXqwmBcJWZD3UwO
OAgGqva5z/KQQ/feHrGuEvT2g8TN6siqsv1+niw5leabJ1IDki3ofcLrw3jzGAzGPTh12voU2ji2
WXzqP59q00t4LLqX3Q4XMOniTkI8VtdMC7N9IC2i+MaHTgHL0Sn1CL7sORJmXx2IneREr6ffNeqc
nwu4VfEYFwJPlLCAhQMdkALLz6Sn+AYIySKjdHclhJIqzo88fT5YsuWMMkeITXVYkwsAzOn5GtvF
sJs/aXZoqM5zC5lfaTqpzE3CxQndbFjO5ufvFuhQL7mtq2JQhvKdoGZSa8+S+GsgdUrGQ2n94oH1
AhIpJRursFJHM4NAoSTx+uk3m7aZrYRy6DObYV/30tjwglDvsfAFutcB3m0T44NA9oayhl00gllN
be5GaZFo8/vQNsEMm9I9+R0YkXhKL8veu5kgnniZF7TodbcCMGrE0uJHdtMaUNloBB6YXpZDwLGP
sAn6cTXmgFVbJJBGGFfQtcvJEYqBDdWgIRd3sIzntBf4cjxGU3u5MrfFQ2OyBinOQd4LgFX3pDa8
pIS95Hg5CX/yfjg7PGLltplhv7tc+oSOjWcHQIt7HnJVrq7eZTdDAuLX6DAc2nlJt666vUebj+m9
AgBaOYvflsb6UHiyCmjnQWtmHwZ4pa5i7Gp9vOjdU4JFe5PES5ylfH/UvoEEG4Jhy5cKVrUV1t9A
UrUFsL5d7j91cQ+nBtL6+7/xh/vGwr4qykNLYrsJcTyBg4NGwEH8MtmA9BHPq1Xi04xpKP5UVHW+
gr9RGLpwypWuCUkTmmt2FvseMY3RYCGvK+KHbIfs43818T/iI7uQqMywYgOmbk4cgmdr19dX5xeR
ZBx5w5Ip51rcQFI6N+8sWynAzB51wvgkK7599hEjvJg1RL1zbH3daX8jwD3qP/CtlCl3U9LmrlX4
uoFknYGWVNYB4yPxThhGwVCGiofzsuict5wlw4xYXk3EU1/DH9q7DwbLjWgVC8OHSSagJux/3u74
coeY2dEGZ990523J2Hvt/SZN/7BsK/aSSB2zF9ZQpdxz8Biu1JpEOLY0dYPkmcw4itrN1PCU/w2p
fVRcjLdrbzST0s+ahRhUqe6FKJtHuIpX5ZCVxyYFXemRK5B1QgE//BGtHpie0/+vlmZ6pZYZg+DS
RxSaoqbW6oDNxREjYZibLC1QRvLGaxKMJiudHqIldLH/4khFODODRnCJTBze/HcJNULPuwXrO3r/
qRYEtiUk6CHZtcGI9hcfEOvxrDpBUPkjNqc5f/Fh+WMItRZ0c5LoRjNoZv12edUUTcpdwRIK0KZp
2Hmf8QwF+Ioxp2yodEoaJ0TFE8DTnfv5mcWQ7NdklyLSz6jBQMNLdlDzxwtOorf/jVc1NEjEeohb
flKrRO4u27kcJeyVNkh/rIKndvsVpvSG7D47ju8LKBNw/zK9h/43q0+5UeErOJpi11N7orCH3TDA
6sNkGM/y7JPxxYTaBrTWlQ1qu+gyGayWQetQizShKnOYXKzfUDPKjNMrA2CgLFRYavGUUz3jbl+7
XSW1mOKlgXn7gugv32pb8TE+F28RxTvHUvI5uMD7kfd/fFcTwnlXYXn/tMvD9qL4mj/KF4bLDq5Q
q9v2IgucbS5u22HdBjnVx8eIebLosc7yafA455Ua+5OwnKM1SO8TEdgp+h4xMKcNp9Ka7sPSxmZQ
bWYxs0aszIT58KOgNOcQborzzghpL8s1w38GupO2SpoJEo1kjaS2HhtxabXAFWZne8XFjzOmRgFN
HymwH9cDaz+VoIX+6FwjXqLuNFsHL4gOgjCh+23b6gooK4VWjTApvUHFEknhjRQv/ve8ZLwrmsBZ
1lHgRj/ngfaleiGrxxBe0YUZxctILLkIY68jp+4gbfNc7q2/HHM56iAvRfB/DUuauLrrrPa/7hq3
dGvHNcaG+zUDa1EKzrJTe+f7S45wziSd+UYSyhVdkqYLvPrKy/tciHoEHD5myugXpG2FY5A3p6WY
deNuod74hSWUQvwqmRYDIeQ1LCtlPdjCGBxmiEI2ChJte1Ge19F7pcmh8fecMv/LL2kdOqlsaSH5
nSJo84mXr6gOEkFNgbjtvc6ezkt6McdwpNzRuDi+eF/QxYngDDiEksgkiu1FdyoJXfXR2yDUN+un
dYJMApMjHMkDyCARl4iYj7hpDsaqGFnKy/Bo8nyhKT8kmWiOI+7sVC1zdgzaU15eJHO0A34/UuPo
txhXLNiapnoDJMm8VyDNayEh7F1Bff1hUltFqqr1TocvJY9weKmQmjKYE3r3s2xNWjIMqC9MxOg2
30iXuUK6vq8KnCrDCl5DZY83Kl7GFV3xq0pEeU9+RoPD22RCRw/P7bLk27Rrr6H7+QqdWR1Yy4Sp
QEvlPr7o/Y7f+c0MEcWUnP5WsVWTqBAaR3ciiN1q97tpBtZIPEZs8qnztN5Il12HS1/1fs2veORw
qQguQc6qBK6HWvwus5Uib+ppcksvm8vWxC0ECA4/B5xwrPtndmv+ihvINSM603JhY7f9BFNK3dnJ
UvJTvAJV4IxmfAf/hzOz3pvUAQ2tNsKE28v2LIpIMu0IruYrSZEiqgjuOwSJh4qB4D6IYz9imjkE
lGgYOb5aWqF+USw8dQEYDytaa6rYJbpoBKuv/nyKFEUq14eECjtpLTwOXMmSPY0hHiIXIqGmoiF6
3Ry1s3A+nIIpYGsnx98GkBXevGli2rLepcg1f2+7GT9r7X4yPyDRk88JHommAQZZUr0zeIUa3ZQ2
twIeTGyTZIZ4I43n0vffoNHfwdr6+J9C05b1YwQjGFoJESUkjbjNmqku2vr0pR4ccCWBRF8gsXTQ
c9LcSvB/kfl0sYj42Of8zeYJphyH5rGvYb058IwjHOOYcY81Mpd7QrVE9Ba7i0WYA9vipAQsd44v
r90OSLQWNEzCt8ldLAFr/Laa7tdb+gjg/khe/3Ub7fz/FjQt1riW6XadN9awlhBptBlQmMMkV1bw
gpj/IqJYVo76CxJm757A6m7ssXjMzgwgwvD8Vr178OIpvFVZdd9fly4LKXt+teva2BUkByJ/puNr
fTW+/tXo18jnKPDC5TMPygBECUDzHLtxXIG+sDH+HRg7oWAXawtc1VjtCBoHjwhLt9Rfqz6aYCAj
5R8yeh68BvpFrOleipu2k+EI3s3kPkN7EoJzNHPjMTuhqSUn/kUMKnQZssLv6Qc9quIfOh9UFxkG
w0i1GxalEqajjLKjegmQS1Ij3lhGvKcVKivBjLhLVoPLaK9GX7kYk5HBFDtWA3Ps9X6fKyiPEcbQ
utW3gHAhyQDgQoqQoA85F3NjNULuRvQUimPq45T2AD/K0TdNdFinsZPUSxUQetmb79i29584mgpi
ELKds0HcuWF8jJh7BrLujkt0wozw5AYKi8f58hlud15ytYFlI40pCsr6DteGvVxn5tpnTjs84H2w
jyhjc0R7fMcLEc0ECjn3khN+EHpGO0YXQGPASVudNgtP6gAJOr6kNSBEqFU5F9WwsIEFBnhehXzt
sPQjX3MH8sSCGsjHXXmuEBQCSOffccqvDmIrygjueHCukgiEqdw4wweQmurRxNm64U3wi8Jb6hZr
FgQJ3IyjDa4DenRwUzQ+V90+tqRhaDsHu3UCC7a/4jHmXjsq56CT5i+sgiX7ewi9CRc7yrLsenU/
1ftUP1eAggzxDgRKFSR+0dcUdRRaU9FVnBs6wmpK9HJRNZieAjxk7KfW7kkVf8uZohdkLDhe0TNL
wfbK5IJa+YjdExukLO+neRfxEy/NIphdX6DkHynIZuJKKep0jEXlEHoSSjo6SJY559CxuQMmG9tV
6T/kk4BNt9TcOCM2d3ganmTvifG7tAjpoEnZrtFBQdfnYTa1QxDM9Kb61uYswfn/o2rZHnjeXOMT
3bF4+iyfytnjqxY896Ez1DQ9R20Z35air8VyscnukznYciXV+W/Tpt+T4eybaZIpfM+Sp86TK3di
utpadsiJLVvE/OUZIkKjDoOVriZy9NqbAbD4g8N2wnVPHaK6KJ0hmCWY4Aa5INmQu5aHpCIah0EA
jLgpqTSacWwBHSM7WIxgrScV8JovbYgrUlBSaITNq2GuAszk/gAtIZLe1Rs97Tc9bxwB++NcefIs
EogHkOa5wWOz6l5+RzFzWEi6wKyE3p8Uol8S5Mk/0QDFIrw/z6nH3c5whUhncB5+Ns5Nm7jhSHd9
v5URsiYH8+JpwVODSGNvvGoiQHvPeytWx0lsqUwJ1mb0Lve1AzFod+nGhhoUogHdYZjkenuIiTkO
hSM3wFiPrWcAU/LWxJMS8ILqu0uoQWhtgZxJ59V0rlwJL/0/GUKTzZf7TCOESNwdJFMijpNm2aE0
y42Np5HRBT4skoA2yQt7AaXSYJ7DBNkL74/Mz+ciu929k1ZdkBBfURAJ6KYh5EgtuC8y6F2jvHwU
0Bzb++T6RDc2r33l1GeQJXOE1/JvCMuDX2n+My1fhZH7kecY6Ouvq5U6ZNMftbGvaidnAXM3nnQ+
cx+gpcmFYWBCjIOyBsH2ilmFm2xwC/mi2C6ZswnJ8LF48rKBc195c3tzPEXWgvVvTosXIkeJ7Ovb
IMl6PuHLzjHdYlpm0DPVQAgJh51yD0L/4jgGu1UNd2Rw8+nd+U7yKjYNIC3GupyHrxlc3R416TFY
uxOS3IPQcUNQoAjT+fbGE7VhcQABM49MyfEwJqeb91NaIu8lTYMvVgeaxVDVW+HnzPwFhQQDsLRw
A9xfkHR6U8jssd4nr0X0qSTAeMlrqNNM+t0vIQRqDiz6f9xW46u/fIyg1sNH5avxeZlOgUSOKdKh
YJMXX/+Gp20tuRi+uW8T+21BVXWmQ3IITvc1v/uqM+FIsBpGb7MNsS6P/+PlFMb73XIuHN53ijS3
BTtda3N5/B6d4P8IC0fN3NBLKiC34kTV9c3DuEPlAwP8gBheDGT/k9mvx6yoetrfv1YJTX/uXKsl
Imj9mqXxNOx6ATvOU458bNlNenfTIGQHEkV7O9rSLHKtXoLHuVk/2I7eVOw+s2vNUfy5ye8jpspB
P2BSzTQ/VbeBx6bnx0K0qkYCyMIWri3E4IdmDk5C3ISj2pZ585qinvXB5J7vu4fCyRakI8df6fix
N5de8FoPv/gL1n4r7TjbH8dsDrBvD19LE/x5xRIjTsIjV2ehP9DFVPCQ6L6vSuN5MxBsl4X58ay4
iCQp5gZMm31qcKandGJJBcz9AZ2ElwpgH4t5zkRU5GnnJPbCzW6EvNV2neIEpxuAlpYjMcPAFQAd
XgLXiGegV9VRwf0G3LS4KnvWgvMLXjlzeQAGlQu19grh9fsQG4diICcEzZ9ILfutiUALjA+4iuHT
JVTz6L8jm4/Nvm9kPVBR30GR/z5ER6wNRMKcinb0Au5suwzFouqhgtzOCWHtAmGtOLtQwlkNIdeI
ivjtbmzRvWLg+zknYYn+E7HKGYjRbvAlOlA3keicWj8RPh5p8JZQY5KUvGJ0LI/mkp8KaxvC/muO
P7Bce7JPRkTUjEjq6bn2OJmLCdWzwBrx6UKK6xQV/CbZcMl0EZt1aKSQarSnQd4/dsy0LkyvIriA
yX6aMNYDebOB0Kr4h82sixb+L6aUzVIpLUJmXITUVoWm4eyAwW0BHb5b/rfZdCB6+l/kmGM6gO0V
L4r1nnVWdVi82DqcZfUyQOhXd1wX9eCCjH9aOi+AQR5ubxIHCbQ0+FjFX27zzyfOVfg5FUAofRJV
3H0DNnNi+z052xqwJmpK4UnfS4PfYUuGCue5L4YiV3Dc8EaDHseD8DJOHqy60g0jNtiTd1mT0MPS
9K4fmDghpM0vb0H+hwMakFIXRWCyoPKHGbTSZr0WTPKLtNP0NJt3oKRZGPgwjy7Gj9wjPlOjp/z2
sQliDtbCUosHAOzlNfvxZzezkF0NiE7Fbu28sz0mrifYsHQqNttg79i7OuyrHlKPhyRNlT4iKuzC
vNKXbIH0d83sgbpxV5fNWeAq6Y7X/2AtbbjYVE7Xp90XdMCswkuOolf4JhWmtys4AZLxMghbuwJo
s+EFvnmpRvr/GbRGlyzjVinbiifeGPR9NPc+/V1WgQPa8D9LrqW/lLv41C2YuoEhDoSdIPGl9Gpl
oAnDVM0LUcUY4tVpWW0D++d1QTmrjyIbEoYUznte7vQ/F7xn1JXSUxbkap/7Y0zLnOlNXZiYcTXn
XrH4lpBLCeoBb4mH0sd6j0dnmFpU24uhz7lTuKiotGWirLIFv02Ye9LPd8oCRgD6OQgaA2d4216E
3RrwtVhInzjn1UuEsOFrXC3KBOQIHZ2NHqp0T3Bul+PMOxUi4YFtQBU+novJsXnx+1T7IiEowwY6
y8Q9Wz52eIy7lba6JVBaWnOvxCTaScvslRlAIvErv2OCfdNF8KltFTIU5z4LQO7yte7DBHpJCY+N
8LOok06cRgMGHHRTEH3jftlb+XJwdh+U8mIwBxpxe69Bw+95kl9XESCb2maxQMUgUwKPuKEYJZYp
Lpi2QBp6YKUO0YN2Ik/EXeiKJ6i4PVXmmCKzen1ceWGBRi4uKzfQCAFd2frYhLx1NscmRCu5OuKG
D0CgWnMBHDjeD+7N0oE+PU9znkMB2EbJrxYcYVOgcaO8qu2LZ2w/sP8/f0Xd5Cj5fiOOHE6r1bvo
BLCT/kBL2Dc+Xu11NG/vbdPxqGhRxHIsuHngjGzfFICf5p9yHTAr+8NRpvT4OoccGD81luNjjYma
jMnIAlK+Uhh6sf+kb16tmLm+eiCE5XzOpNr5nl23ENPLiNtYC2a1Q70HdqPZHgJjB940WegpBKBV
qiprDExBGc0uY80pVevk+5xWVmtrsB+WnvoljioAZGngJxzPcasyQlTZLCnCrHLoGQdMM/Ka1a2i
SdxsNU6UgnH8XoDTPDnUvr/fdVluIVoslSiBh1taeGqx6nfvnoRzb9Vhp9qk35U/AcMfaMkfW1w8
7f/pN4Hzg9vPPqGcYTIZ558qwm2GxPHdt8jc4BHAons8rMwBLVGTNAfM+4RcJ5laD8/5WLQM3K5x
jA6bOi+QrILPBUjjk+lVw4XPMa5UOZWANN1SyTwNkuUFKnVpVPG5GWVleb+3Rbbfz5R2MIF9hiid
N73Z9SdOVY8eIKV4jlMQMfkJVi+3zq5GdnjwKgZ/8zeY1Th34BA1upgbd5X1Zn4yBYTQncBzVNBJ
Y5/gO+yr8dSwmrV1f504XlfRjPepsSrSE+Nk2IJ+Va4HacMcz9mg4QhenEPqus8iC4ZfE2mpICHH
2SVEhus0AAXDT5EZ8FYk60+UjS7HRVHsl4d5fi5ZuPOuTbtxnsK43yQubKyaGyqB9muJN88FJTsH
lklt7sR6umAsaV0Fzz2s/dNxqZqumawLU/z3i0gvz8S5vOYQhnMhAljk0yRyH6jqlcQcojiOhQUp
d+y0HXguvJ7hFaqY7o8kHrWFfFSRpQVlF00C72IIfs+f0pYMS8axPL2+OQHDsKDc6U0qHkGzCcWv
S0fF4K9ArlI90y8OCXV4I3p92rhlGDDK7kFTv7im9ByDcM1ScgaaGOj00bSJKUrJe8f9Kt7500x5
oqfv9F/eSlnFn3q1REkq5Burf+lHxrnjU+P6JWdYL6rUsyk9BMpMgpjjssikfOxum7sv4TRkILvZ
aso1Q9H5nG6zM5vEJYMCz3glMh0Kg7jndbJJxeQ2FIbCUlPbLex0fx/Crnr9zIywLTLd/n9E0F1p
HcFr8gaZlam/dp+6qd7p98iFV9Bmkf34MeAG3jWMpN3Xxn7fk8if726EPP0rj871kqyi42N1Wkwk
nm8d8e0ybJWfQSgw0L4o5Qe14saV42FGusT6AhHsxiTFk5equm8ziM4g0ZD4ZnwEwxyQBqmZ5KMU
lAruiPItiiUhU/X0e7sfTFZoHBFa7yrmNMBhoU5G++5fc7jNjmRMTq3XfPz17tpsFGc13ri+YuWH
izryQVAXaOQjAmllzWwUA9Ac4LOrtq7hpD3dtaw7ZYEsND1x1+vNsYhtxlsqypeXdkRSTiiLY23+
XLKyhhoM6+7Z6+eaYsVldLjJmuIq3bqreiwEGGobgYtzTA8zsKD8H/EWgXwqJi4m9yb26iHlS2qx
kIdp3RyntqvzVMkPsyliYU6VVh1zRrimt9uczdQ94IvjAnevcJm0VxI8IJE9P9X+LeKp/ggHjba6
MtaC8rai/doljpaKWGjhSddwYgtrW9LxCa/FjibllPFk2PFQUkS1yYIA0vqE0338jIAGF8Dc7XnO
xdTIy0dZMgTbMhTJc9pwth/rzzpEqkIptgA5PNqI0WXnv/AGiRDNqd/O44mnDyjs0NfOBqsxHlQd
PtrLC5pFULYUd6zbc4j7KjBDBs/UGRsd1WhtjEMLJV0NsZxfnCFcmVyeAwIu5NQ/QABbjXGZGn2W
dUPne13A5iuyA0kTYZfWE1L/9Um+lMmpjPT3r2Ay32mx2201ITVaPJ0mfjQ4HZZ/kOpoa8Zb8WjT
s+vaj9rBFZ5SidjhJEsoDTtCKB7uimWtq9HVTvp+dSFg9UlHt0Fs35aGy4ZhO95zNYobTrE9O/Ek
bRAIanyt8jznv8XQ3RTRg6+qXQz5WfBJW00ADokmGq3F0PKFPCAzUgLPZCE6uZt8V4ozPwu/JyKv
FLM57yY0HSsGENwFMAgcUP5OX4p+RU90SAlYMXa3qk6H45ZNzC6ZYe5hKdHCL22fiQLnZ3VF6vv0
ic9jOHhAL5i7D1d154X9RtR2nKxt3Dhtt5QmR+w61nmBFUimJqYLUYsi3bOEnJxJBBSdPr4XhDvf
RKehIoG44V60c/LvRteZT1x5i3YLh+RIS+e8facHZemuAJDkX2dPvxKwaERR8EDvY8x7Q5OPv57h
88U6/d1ln8iRAlOY51SY+PACQVjjEX4pA1LxcbR7v/uphkt6GwtOMT2bDaqiAwLigtmbRl5Nw1mM
FIJzHYq3Mo8AXUvOa4oHxvBE7Fs6dM7ogjxsaZ6A+I9GQk6thE8Jlcau1fxp7GsSp1yvQoKWLvF/
MxAB/0ZwyV9/sLTsEA9sdcSkG5BhjkTwsUESG6KYwYGCOqxQC+QtaH/WnEZJ0747eIQBjjLbc5qu
HioB9xr2VsEo4M7VPgEwBEJJKjLMRJfREyDoSUwsThks5zlTeS058Y6zEUEawojQcQ115Noa0jSO
W6KJoCEs4pqB1WHcF8Hrifr2/heugfJxLzr8UOz4zxw9v0PphMY25pdoFDsEylFneLggbJ08jTuq
jm1epbZQO+4S4bHiKhqgtuO1JbnV0JOqiN+uUHAcKNx1x5pZei4vj6dzL4zncWwE7Qzj2m+dclP/
ZH+n5/536zFwqdHA/qLtpjrwRF+WkJQ2AcoM2MyXZCUD0lvT+HwQ7wwgJ4FN//mm28kjMTJ1o5yL
q9QiZfBfb9BH9qX1BjLV/xTJUNyS47TQYNVsLusXQl5H/sgaIWi09yEIRflJl8/ljJOBdxhZ17Dy
Ui8lOYzU+biMrR/8VNB/QF9MC1TayZwV5hlh8LIRFukZOw6gIobFovHx6nEHE8E5yl6xPvaY2R8i
TGPx/fO70Fp74gFc9WIblcO1kQMDP6qz1HJyXbA+9qBF4mJ0hTvl28/HXOeSCsm8Q9Lnq5/EGKdG
8NaU853vbzBh2VEBDiQiiu9FNRbO65KBbYRISPybrd9X6N+pK3noJrYFMSnhRJflq19wof43wKSr
/7EzEqpsNubnjnJYHhTADb938sF44jpQ/kyfQLGmf7LcDMl+75sYj8K5uSnXRLOhCvoolxTVknf+
TvuGAPlJXz0LH4wZ43lUD0m3gdJuN9WgOBNL8ObzTXCw0dYE/SiMQbELZq9P/rRPAynbR1y+Uf2/
V+OCK29Z07TVDuh0pPRsegSrQ1XR6ENK4U8CZW5F1FdpQRtLobEd1nljRd9MdxGn2fZBYVOOf8jC
jwOnN2RSF7RLGitP9E/gJxc8AUBYvEtGVy+kVkuPAIBnwQhnpSJKpACV2fBVuTvhY3kj2r5Iz9s5
K+m/lmAUkWDsqTfGXKA+QH4MkZXWg9M5fDWdRsJjpxaEqG0NC6AspV+BH6xk+9mT9GYrLU3znldZ
ySU1jdphgC0SkTB7KT/8U8Dsar91WpjWFwOMxvmsA6LXeQXRmCS06Uq1qCRJ7EBFdqtzoV0qtIO9
WzIIGflUtWSn3vEs58KIWCJ970L95XIhLwJO0q2F7gY4qQQx08cuy3BZ+cc0E3062lqgoATHxefT
NsPvUA7F9DOcGNeRQ8irflkIMg20fxKmAI4QYXUFpOOtfCG1Qx0HG/yaL2znH4c1HcV2LKh9BQsJ
SbduaPH2/PsCMKDNCy3tJkrq5KLDDdKU0Z3/nIayjLd5N0EpHahKAZg+PfNYFwMt70EPhwv4nFAZ
SQTtCC9LoDUJ5BSwRq3G109pujlmZC7LGGrCPaV9Uk/hqFpj62MBJ+mFjn6AxkjGiB80V8QCkWwv
lcVAzGQZ90DspJY/TyXBogFSSG7/qDcwMwmSdh8lgqW10XtWw6kPe3t7BK1e5+K56sUbGVGH/vcG
Lj0wMLUC/skJ9bX28pnhKtD+JKFRcmnRlyPbXIiLXRkdx5eiduDW/zkLgEZ2N9CYyl+YnQHuELOd
eV4TMrU3AECE48aLD574Ts5iwKi5ydm+RZMFfw05kNhCvNZzfJ5wbH1CCuvxIApzUdlR0yEyHz37
JBSoScDTBNiEGIi5w393jLRUNyq9HD+ZzyOgP0FXVOSr/smSIpGWq7aStda6SAe5ZIo4Sxd6YAim
Pun1sBxfgEMOYMDL9Gieas5lrQoiPe01M0XAH0uxtJm7HJEwligB+QjNROBxdZkdpwOC2c3EXg8Q
URxGgeio2b6tUuYfF3jKTt7zf5uE3bxnXVzDxd4MCsRdv5acqN1kcey/FntrR2ZvPTMdHU1vBXAt
Avec9xJ6yGc0XUn5RO+Vn9ZPOF6QkqYppC0E9PT+BSmS6khGVo3XmLA2gONy14A2mcVqSL38YA8u
rDGrbBwPDBONO73jg752j0UEtG0ioqUHnDv/O9bWnf4xYrOPKy7BkpmgxeKmyVHaRQmTVtcXQ8LM
XZq/8p8TwGxh2Md4HGg8LorvFP9GM8ONfX7ClLVQNXtI7+4LTL5h5mwTKkc9Ng6CjORY8Cfn3NiX
Vdiuofx9+LHPwMASjAm6LsUpMPoszRa13y+SRZyKnMd0+zdBu/9E/B8v2GeGMLOunO7z/9x3zuQh
rwq3j/NZofFm8QLbp+O/9mft8GQGLJyRvGq3agtv5c0futTr3MDYrvWLxa99up6KDJsrx8qxjT06
u/VJU7AQBlAqp+4UvQ1UPWfMUVUlXxrgJNtQ2VmVTrGnpoVB2lx+QGtdXwRKOOwPcaQnEJGSeXFY
XtbtIQdks+1M2DCCyy3wyPzY8eQzwvgRvKYS5mePA+71x2zVBZVkt/Fa1wcW4eFidaJk2u9D6Gjh
PjGhhyiPVwv5dqmaTtl4H9SOTEH84Giz6+fKlvgGB9g8xikid/Z/Qkl9kzzce8V9g0RlqGWYJA+y
oynQIGSH0qnMlnkUbsQXH9N1D4EPyB2iubiykYbp9GZBBdW894fo57N3WNwkXOh9GbkKAGiUhdnp
v7ttR35vrp/5SV3e61A0ubZy3gcHKO6yC2Pmxpo9Xxo5VnkTFEVPaCvjmxEw+s5CyY/ugitr63LW
+YBGkdbaJVdLs67fRlH/aiwax/ifm3gr/37KqFgQim8V+nrGBFs4xeRujS0dy4gw86etIJbca9ap
FZQx9POuh8NUEYeibou8dHja/GDYI7Uy2dmebZM4/TYLsbLbhUhH2tbR2Rcgpjbp5jK0/Cyb1Wht
uSYWULGc1TsIz/X10eO27jevHZbiU7TbMgOKI5C/mXtGCKHb4j3fRfaeHhl9PYBNlaKcTkpPD4Eq
Abo3R2RGjoSOOmXt4dxa6UrvRetz+vZgvmfIZylqrYEQYHob1hJtmNsPOKqZ4WfKdn3rb1PfPIMC
jL89QXsEl0lKdfh8zuDqybxUNQQ43kOdnUm3QMMrI1eT3MPRaloVk9ut+F8w1D9U0S+f7VeCoHj4
TUXzkHmeV3OR38OKApGRE63WrPLt28oJyelZbeUgw+nqaZ7Ul+mqqBU1QuxuMakP4dXa8nVceXre
Gm0ZbXgU9UA7nzjWCmXYGE88r8TsZcnLTSCVL+Ocmbh6PRaynqsluPQfeM+iWysKFrwVuxDQaF6Y
JkT5boxtREeUSlyADyZhVWbLAF/mYO6Id39DHZG/cNSKSm01yzjvN8H6EIu1+qnri4pdQiLXwvA+
WUspLZhp4/zx5lckdilnUoVf/aYNPEbEsPbrJedlofbDuiZBMyjw2wKy8N5b+Hu+FaMuA4MRIgnI
PoWKxiF0aU0a0GezB4pjSDKpXaOXNjfn3ZmqIhdKnPZR/NuE2ZnaWytzFdfcZr+ZUZdmCPk51Yr+
cMSGRx5qtED3kmk0qH0eDEGb0FEQ3138142WB7KMQOiZWSuH6bQLe/+x1NBrjWqJ9iutIDWUk2vR
uz1rFCqpgNToOjL7lqTn6+i21Ncp76JAm6GYY8lbkmY/Fm+2/WupZ3m6/Sj8qYNuQ7zQUFxfkOTL
d2S9uYYl+y+28H+Dpbd2XQEzjpEymaPga+kMRZuIS7Jmr9fJ9rzoVQFG6WYF/ZkOhTzPiCm1z6ls
n5zIiv0shewhW5SqiYve+Vxr7f02qELdjuLorlG1cChVdvfFTsexd/NJ8VIttmpM1gIiCYBSN8Ng
/l3VmtTmE6cTOhYSPFtiR7pcE7vhjrXy9XyAqhQpULpb6Oqhwv/LXIVHsviYEc+3x0wXlc4MZ3HA
Tj1c0DyIYvadRTDtVoE4wP9r67smxL7w6WGvDhpZOBxQBnHarA1XsE58j+qhOVlpDu8Q+dBE5riD
STbWjRDofss00UOrSdVEcHxxzcKqAnwyfRhjf/D/tKD59TjJjTfjBsKJ1PnCh4F2vNUFeCmUQAgJ
sBprs14PsBarBEIF8JCkyDgz694yHXffpOUJyLw2wcJjhnskBZxIJ08heUGOjUOkx7UbBhJUPU9X
8orypLkQ88noA+1mUWEtkK5J+gYVCbVb6+nXMCeP+Mjn1mV98RJh8QXdmhpxGcYMD2JUWQZr7tm4
PsadWFaEJlytiG3zERvOdJoDNbXXCjViHcQRilq/OmkaBgGZHOeY1s1Ze0Y6kH48mh81I6bpAZQV
J14IhShUjhHrVcejlJ67IJ0gMS3h8NTdd21QIUCUnqk1cVCKr9NI7IKn5GybAb5QpS8RPQEoebsb
a4lZd72nDbEdxDJkqofHxFVoWzIsyNJkS/mp1a2i6qL4g/3/0gmmzHJMQma+l7Vfu1Bj6vT+R1HX
5lt6xqB/HdSXOJ+ZI6Mx0FT/e0XEugFiGRfjTWQaaRtksf782pS0TC8T5jkBCm+EY3O9KLWaWZzS
7joJqXFJdxnSIX5Jx1/5SiPuCRP87AAuSrQECuiAI3CE+GekexwmQdxbEDcg+LzgyFC9b7cyuH3S
rqecHsiMtEdgm2EE384+L+IDxXO3Fu2hfVadS65RMEYB/i3q+cHPOGNz9J02yC5Zy5xO6MIs8Z1C
CAv3VGPJXR6wtVMHmfipJ+RbW+HZcGO8xBvU0TTHcVz9vpCZbpMa5MSbFoaoejNF3PIhrphAUhci
6ek0h4kjxosWRNT5RAZmbewd+L6hEw0BUkXFyvw6sNcm3zFJU1TmyBOL2ov6h6CMkf0Am3Zdk10u
8FNlh9S17kqjB8uweU1XGzXYaCjl+k11d1pllaXrq/su9a3KR4efLRam5xXyvHIHhXHwtoAKdEnX
8w5goj/NQ7Ufo6qtvAG+x4RjBBpk61hKwBFQSFfTzy3D5TO+Wfi/B9xDQUDlLEJUbwOPySAlpiav
QlcgTtDQr6R8Bh1zJC4cGImYjIefFKM1RBbwNF2igCbouezGuvJLFmpEZDqM2p2uXjLtXCsrMiwA
gy1tcyuwJlVluZSj0PPF5ChpHmUdAFqFA0akTXwTrKf3gqXslekXNksWYu0SCkSnRdL+F3VvvG3N
C8JK6PGOZE9OzX0vdq/aqyWoBjS6Yoel5bKLCO6p9oUSVBWp+qq3IZfFb7CDXKIS7+wiBvTSQ7Y8
+5fCAGNhUWL8ngUf6cbLJf2f12c9Lv4OCGAhjtuh39+khyr19Kaz3+tkQxhm29KqSMdNJzG9qV3K
aW8hueWGJ5HA61awId0JnmW2j0Lvkgh3FQuVA00NGBfLcM2huLlML7A0645LuL37jN7QZ3XT1XIu
sLh3fZYYBz/8h8NqaaFinCntnngJvGcClEkotItBCogsKYohKyMP8Jsira7UITxWjLyNB7fylxHL
XTCC/FsEDMXIxEmDUGVQEJtBquEmAe85lePDkzo4HnGfvo+Dc3k17y/aLFcTJaoWv3Kaqf/91P6B
zX/0Oz99GQIrrvs2qmvJ+gYxOXJ/AdfkwqgLVFSsWeg5VLFYvegjspQctpxgspAUHqVv5tuMpj6h
PmGbvFCfWAcI9mJvGm2RRcIz/oltdh82T2vpJP26vgVQktlE/Vg76d94jpy/NuLvdkH0gDEtnmHz
be0RUcX5XOc4BuSAzaf3eqtGPvX/jxAB0+XtJAe+Gm8ov9qfIYdV/u38nyN03Yb11OT3O6Tpd4cK
A/0+9qFUEaFqooEB/FrBHDOOo6pSwttavxo5G90SV/qcgxylCFgcWaKrsjUA1r6AVZ6lv2L9SBES
hbplncjvajt4KebLWe/jcicTdslxmmbItDM+Sbyunf5AkiNDaxtiUFRZr9v+M5dqv1rZJzr8it3j
LLawhI/GJ8UMRUCGy7T3e3dBmThZfZVCNO364ur/Iv4dZoVhkCRypRIMolrV7OSi/TAukuIu4/SO
S+H12mhybsXiNFEa1UD16UlMwFnn5giMzE3p3tmOGJOC2MuYFmaiZ1xo1QSpoSc5+rSEgcn2gNKD
+KAg7p7NJ2Ge5p/2y21/mEYDQmrjveYzXLR5rb89Dl/wpLGabD99yclyuDEWpSa/kdC2BNisX8u2
OwURg8i4KLz3aSI+mC0i1Tde1eqIpIiHCxBiMV60WLYNWQYEAyjg5tixVxPYDtAjCAoHH9+K5yHu
xx014enkgvkQKeX0kybNHHSSjMJGrXBB40iAHX/fVXIHRb5DLmDrdFXdA91aRig4OFF8Iy+a5D0i
Jwq7RlIAcJuwr6PW62NJAqUcPKxfgMv4uXEB6fP0jsIjvCSSTVXOlbgVlC6KnHLIsQtgsnq2i3ww
5pL80qIQAy+C8riuno26NWztN+ZjFNRh1H1Mvr6Eb3+DLlWi1TDVxB3hziBuEKVPZK7RzRNxbkjt
GQCq4g7f/P9hznucKsE2iEYN0F4evIqmSQE7uWnjo6okJTs9MNacvAReKfc8AIXORhY31erKo2FJ
FRLTvcHgzrf7RgrZRsj05mBzmelYbr+D+yKdOIx//e1FQpHNZct85THG6h3PHO9o+yPS29VLpNPa
IUQiF17mnLRGzx+zEj7yuxp5iwMpc1/JqSedr99Ay7NfRgeruiIlr3unJ4qh9evbMsevsDAAT1sC
ByVqp1VpYDX1s2MmzlAp6rscaw+BNz3BJMuSyRYjL4zdtfvJpOPuIDIojysdXB+Cle0vxcCMlpfT
y/BztVKZ+1gHBPZ4fBIE+RVGtoSCaYpRTxaRxg5Eq8M0RHm6Ijb3bSu/wYOb+SvIwjvG32vRkJdg
Z45oZdJfSN06BDMPmvJP5rgzwXWQ29i0niPm+fy3Xm4gYDrOe5iHAFmpdjj2ojrbNd239oLdzDPd
LFdEOMmcs+EIYzc0gj1HeaJmDkMY8cXuxD7eeCgd0cMcHR71Q+T1dXkY7Y1H/lUP6Lu2ZPWnXayD
4srvyb6MLTUg0gTU+F9VNSGNkYoriM0OboJg9eKaFQFVXmKTf8/r4HYB3IFcsaaiuZ5RZfeJFrq6
NFiobIwVN6hWzDxYc0yivnvlkyHC+sNsLzKHQsFXaHt4odSCmVQ/cdYT8TTxkmGywN8tWHqtb9q9
IjOY6yWNoyHP2pNHpsxI5SGlqSU3jUcv9As4pfrYxW/z9aaYYu2tqvfAt7+EHy5w4pqBRGXX7rxs
ApTZ42pHXZ0GcL9Qf0JfKmR7cVKgC8kSkO7kHmm3rFgH+RDl31RoI3bjs4MWXni89KPVBXz7yS3V
Bi8uVrNavn2MpNOvQjVmrCgFBfbt5wA2ywHshJUebmDcwvQdLOmNr+cGD6UK32Sc6UFeLbll/74m
q5xSm2U/Dim3pqZObWNDuFS+05V6ab+snzeModQY7GaPKNy4qAy6+YLQ+S3/3aRHvCAP9m9Wfhst
cuUAqFNaHNCmEZW4gzSGwkTNDbB1MHIonPPTMmON54rkYn9qMOMej4GaGGb4lbsADrCHpe1AaDiL
e/THjDTTnBBYpJClhdEfiHunEkLghYdOo40plLg9unm+qLSFKzruHe/f082vRgkKqnkHZqdrXq99
7eFFW1go3HFlvwsd8pvBUy6gzGsQ0LYpSzsOkPxT26eDknWr2uMSLjraZvrZ0B/vhjiy7oFqx2hC
AW2jOkLGH11OESmDx0JTBCR16J4zulHpTyInVc1e3UmjaEJJ+3pudP9+i0CBlNrIA0T7aW7Dxmyd
FJazm9Pk9rvjSf6D4TGlbqGnSNhtjWYa7SICWA46oPqa/bk6rtIEYGk4D8Nt93JZMk3fL7dYdju6
PJGZvGJ96P3zAhnMgqZjlJeHg0huj2A5SyHLhxuMSuQzWU2j5n4Ixv8/UdIZDTDzoWjhtrsyLSBV
SC4wBNXLD2FTNgjJINWopIpOJnQnHDpbwSEN2zPlaNwrjoiUd4OeDKSthGrPGg651/kR8zUIJPGV
6VInGyNVw1y0j3t2Rbsc2IHlJcN94EIATekhRmEDpESjn6lPm/lbzKVUOEmnFjNlSItEAwgfbA2v
JhNSKNOZszJ13qIABlZTxrfbMFkTbavRnMuTVv4bZnwlBNUsIIRwR/ZE3k2TtVJRhncPc/FPNCu0
4HuLfXBlYusbsJlsmTpbfJL30pd5YHGOJwfNgg+XlMHQBcg7LlyNlRF3fl1lSGKNNlrcykXrhgsa
dsaTgFwbtuynJoLh0xuOujhzp5NcDlnKS8+ipeRSw8KOmJyIGo1Qcbdk+aAoh6XPiP/NMDb0k4ux
l1PbJyTAtm0TuT1+N6x/Lr4tZrPzitKH0B/iLhWORGJ8Li5DSqb0AfKemqnqfbWjbozqIstJ09wd
lZdIJfaaLFPz42JDrg+53bqQ0mhQmjfogTS9tAiioqjPRs24kssUKAcb0iezSSZ3CSTDNhi+k/ht
bgtsQMZY25tI9gm1/MIoJC6u4oQvZsMc/kAMQ4Vq3a7nff0XiRzORl6uwQqeN6iZSPptQdiD6G8Q
dcrIZfIRvsmCIgpCsvAIjKBqCq4k7SDAAqlqRfBksulKrCnHYVamzQoom3l2o5rd+h1O4mdzRB1V
4nW9F7Fa74FOwkOYVURL9J25iU2F2jL6veJsXwhHsc+wBmgsoD+NwiE7gJLs298Erq9YTM9YMjSu
O0tkqW1Rq7UQpX7eMELh8Lma4wyTZR5N6fgKknKA06+NRXcN9/LvEwh2I0l45+sPlkENo53amrnI
FOFtUlZvJRU490wnfuoAi9GDdEwCO8H7MLRIKRT91jpIzzUY16X7hj+lC9a5oKeULuHuiQeLq1tY
iteAi0lg56gdJbAq4of/mGPdoQdrZGmZ3CATuS/UZb3XJ3MqLuy5ilEP3edEz6FZzUYB6+Y0j4FN
HxjZiImj6Uj3V7TsH3NqhXJnu4mukQUwLyGyBITSYCYsp9yUzQxZkh9u+AYoIPpFQ9CWN7cGMdC/
zW0EaySh3W4OnTOrK8KxKK5IACdHB0BW/86jEPrOH5o4W5pRWCz/WFUeGVNzHh74wEvv3vHJB8yf
09pZPc2Fs+NIbgPuTgB2QXTPuxDbVRLlUu2a0tNV5TwOfQMfpVU1A1fD9jFsiROPpUl5TFdVey80
TlZ0PZAml/2EHgjna7PvMqRbx+zBvuRqa4gQn/yZWHpYZG9Rvjh7eul0XgOAUotj1/m5f4eKpSyO
6y/NX615YqrSNrWt3ZltC1A9RasGZMA2RYJ7iGdAvixATPJw/y/2QQXMgJM0muE0jWi/Uen3m4YE
MOWX5AmrDygLeC93CcoDw8Awb8d1N/fA+rLAH9nw1MK61HIS8o2DQtsV95NLr9n/JXbH+2Oq0Znq
U1Fuv62aIPbxP8TiP3SY1RhfH33zwdEaIn0ig2pmetOhXDVBfajtZkzSKvBH3sqkrx0lWjnFimnI
+gS6TMpESEu6RYBUOKyiJ5Z/oEwju56Q1CmeM5NOFU7R8QphfwxEIJGxv9jlaycbG1um757HuR7O
XCyaiWbRKUu9P0Uf6gI61YsuSrjNcnkEif/6djks+fpNsFWeced/JhqvtEMfMlwyIrKOZNoNaabK
jiFQ8b3eFpjtibzbiUBPguwu2XlQMzNY0/3bzwFiyb/Yz0Ynl+OLY0RMyRcSzjh8HzBJcCqiKeNw
LIdPJUU3kyaHdXFS2eS9cO6YbOjm1FScAq5aLAwOo19CajkClzhf9uyiO7ZIL+t8xnGdnHpCCevl
czXxYO7CI9M62/werJ/0XdfOLVUL+CnDlCxLj5iqq+TYMyKKqX8Fh7ZP1CVteEJm6AxDHZ0qOppj
LAWa6uN65mVtdlHpsmmu/0BHL8gZYwQaJPOeUytaxQL6s5HO5QY+i4YgVwOOYnO0bObMmzCPc9Rp
zI7zScNqTvGnEGvmQBlI/uDQVjYYpDQ6Xok/+Ger4gzeriLr0KJsQ+MK+2hjnTTMUyjCDtYEAB74
yBeP+B/EKMCGKkcQzZ0pqJjpmiUBRzfLSv5KsQz4bRkxuZrPjIS0DKgZziIpgZvqwsqhfk/Zc+h+
IBvQ59X6dBDlS+AkeORSaNacnmexTuvszsTZx7QLpVAwRuWd9T8vhaEF2tBhDNsQl72V4PhYhXEc
u9n8VkxCVuyMh+2zXK3S6+8r0vAM8LbKdzi8MUNaf6FwGkiV8PEta1jtw0ExjwvZTlcnw5b45lDm
4XA/xDoat6TD3i43cPeVpnClu+LNkwMQqjcrBIjM3O9QshFzvaN2FoUVAZ0hRCK1tRRXcNCpdPKG
YoWRowg3mcFwtC3IT1LlrB+m+ozNct2n9suB3ytt0aye4H9XxcjElTZsR1CJLnH8Fuvh+62zG0dE
F7t9v9OMsCVj4luqQ9RS6XvA/kDNmv8uDhGIc0lifFaNNNWh0WWW74A4iq2HYskEsPVsAQHH5Poz
rMox7nc1nRpZx2GHProOdk1KTb4Kfy51xDebKSdoCYPHje/5MkxL/WCTU9wqlAvqI+1jPgP7k/Ni
2W0kAKRFjO7Gw8c5cXd/+Fcy0Pspb5hFL+KEAJ++G+kEdxKDNiG6u3QQGg+NWnNa9GYx+g0VOrLW
4tayiiN191VSaVL9IcENFVCrEzSFKu0qjMogcUEohRQMbz0KII/JrQPCe5FHjTKSjITCfIevnVzb
lPNR3yoML0MgNy88ot0QWRMx+bpAKme9hzuMu/gTFenTjepqJTCBkiMaJqlCZL9divNw8TnMqFDG
e5oNlHJXakGa+L/IL7B6Hxf0/IJARm50Cn6uCp2vXQOPcxKqCvveqkeg8wPmeXGc8Mp7BT8AASQr
oEK98xc+SQ1JftRVpCy53ez6yrYDR40E1BBtnfceDlpULAYipAQBnu52Re19oSohazPIi08umgGs
ffwRbNxYiAQFz8hfskmLMQ25ciFWRsi3aVOfo7ia67zLDTybFxlRvHMkS8cvHrklU9+7QluwCcqQ
mgD24aCzH5jXnt5Knn2Q1YihrS/S5MxERzSiiUPZEs6DPbhU/daGMV/KRr85O6U9xz0Q/gzpNMBZ
Bu4p1BuDKJuGF0bJjNeJj2F5VeM6b9Q6V9eC+VtDiigpGHknLljwxYqaN6bNNJZpFK+K2vd5u/Yv
1yWga5JM8gWnUD11bMdZenPPC3qHnvY481vXrQmn4oKVrJu37wnos2KvGwfP+LlZKQ/QSxRAzi9f
PsJfCC2p1eBbfpAZM/c1giP6Iws59TpRyuFUCgOM9OcFHkHuG3Tj+4w6eRhR4nx9VnRHcm57BZgL
8QpX/sCz3E9U88sgEkkR9yxL0iQ1Yd2H0Ph3qVdw7pOPqkEuWnv4ezsRJXslKEWJOf7IGGplJG+O
cvfQreyDebcQKqojtpMVoqf36wki1QdF+teU75V6Eaj6p4NFbBmTR3kIHlXj14hit3nM0SAHpyeL
jTryOIjv5N6IKqU5LYipmtABDpygFIgZa6ljQhNpibnzoldjx1QjPqztT+gLbAntB1+N4+SgUPNG
D0U5u6kAhSRPXI7q9fj/z+tgths0qUbEL4wlBI5O6kwRd7OG3szicJQY91ciT2rCyyBa48K0CC4t
4Q3N3a/ztWBwnLFJ9PwFXQDoqIKllmQ43aDomhkEN9FKjXK2TOilTM4SxvD23o/eyPfdG20eNyTN
oNNnTImfg7Dtyvqceyf88k/2PH6Z/QuykWVYeUlhrbQ5ZdlToarBHiziXcxGrnYVbFFbHIeX8R+R
wDZ7tBMWGjh9vBY26m2JMflxf9s2nqR9LmH+cDSgtKQgzBgO+0Ok2UkZxsD1e5wLUqEeszdYNjKK
tvY3NWP9cEzXgJEhwOIhMK9214N+r9/tuuc/sRvhaxSV4IAo45tmx/WRubcARq+XCX+BlruvdGhX
gmuHBuDnSSdZ6RUIEcJjEOBrYrkWhPVdQ2AOqKW3BM52iVZtixryTuPXUk2Jl79qFzobduXOmVnM
EEemqxclJblxI7KwbZBus2Z4VtOJC1eJfFAPKjNfUan7wvj8ciDCJPeDmFmgSwcK7/gZ9wf/uSXc
RREgXNCk+hgXCitCn96b+WOQ4MZngVKJZTgSvEPzHPlRb3gPWNRhFWKTUqFcP2Tb/P/pW8Gyv6Vt
j/X4H+/VB/XuuFVZdOht32axPzsTnR30qf9OHssWNTxWl41LGB8Fvgdy2kysT7FmzlROg+7rQASx
Nh4yiB/ZEQhFm4hQyszp92CpC1Cf89+Sj+KoW8QVZa5gFMZcFevM2KwuCBOl+73SkkBo5AZYyW2A
rjENpoZDcNe9OMsPiKrQMpkhwdkfIyxCQBDuY4N4Q4uneO5dPJBtE8/ZJ3o9gIXhmXr7fGZrrdzJ
RqdXq9JsicGcc6mOmsFU59QqTQa78icy7kZdHsPN8/wuWtdyiMGynSHLuqdw0zHosjhBtu2zYJeQ
S2DTljx9SmfZrNx/ZXIbUK5yQyqTNLs790/MnvjNCriN1v+sVCqmYdG1u+t0/tUimhxBzDv3LTjq
QXuc+G1NrGbkgGes4KMLXO/KzTGt6siprlLroJzNBBUSFcmKwup0ZExJIARjZYh5atA+6PxucDHQ
BwhvVzr16AFV26MkF9FQA2mu4qLMH3jSBwqiPW97GghFtVz2v7FDk5OCCBlKa1DZKT+ui4qW9Jyb
zdbQWLGOo+SAc9IqfS0eqOC9LU7cxULsqr+HGZtHXGnS6V293qDPfdg6gGJClZ2rvRjt7N5VntIT
63BfeM4M+JeZNI5zYfRHGnIV1J2aN9yW+ya6qwQfTRJXaIf/en3kDVgR59DY7WTWxDdiMlhtahUo
hPMaXRiDSDdzhMrltX1V1TIRtVwAXn/5vpDBi3LEw7ipVTMnAw2z6Zbhu1MAZ334jtaqywVuxcqD
w//Tw3Edq2FFjg4FptswBY0ZaDYLfry549dnK2VcOUHjXSkO3x74Ywdjd54fkKklWdPq6RCx4BoS
/G3aADzBZhFa9l4WmEHcomAGw6FP1aN+8ruBbKzEqCVb/PT09mQ7toUIUGDOOSqw9gmXf1JnjCnt
xOvjtgLSzilwkVrhmwxyBFYtc7rq4NsFB6stj0V/g0lVVeV1XL1jtwN5SY+uPIEcmD56UIE9tlo8
qRWjoW9YrvUAWymMYu54U1cScNNFDffzli8Zsi7D+EvaLyXJ6K3wjDIk49nr/icCOtsSUBiYQjaP
RXGerasbNjNkE0MP9Wuiw/6JNAs0MuRwLLteMMFN9mn/DnfkprgcVTg6tzM021csaKzV3jipsWyN
UViAuDPZbdDo3uVOL3oZeDI4+mspcfVerJcuRzAzbVDmP429Uidfe689VzawuuicqYVcd0KCbkjb
5IXmv+QTYTuqxpR9BJF6AQh9Ygp9JOOpWz5pHD86En8YEJfMSJA1yTWWm6yuvOl9Sf04JJ1KZlPT
2QCg60iqSH/jefOAbn+Jt9dYHnsUY3/k0xLJpWxngk/db0twqqrvB9wJTW+x0JsKX3lrodSsL/XU
RyFoCpuT1r/gISeprfdYlfqvpXG+F6j524CZmmVhY6iO0Gl63mVP4tERvAZIVntthufQjWmgjEWO
vKO+qyVax9TsPdn4P03oCuUf2F4fbvW3BiAgPSFdbR4iuJ/GDPI/MI0YRC0TkilI6nhjGkOYrDWF
JwSzE5XRBvbqND1dhtmDfq30gQLuzPsV58e9RsY27bW3XfR6GW0bsbr/UlYPEsRZV0LBFhbepmLj
ReNP0EwQ3cOBxJZ1oKG5xvgouNIvHFzD3UtG5DeNnL2HDlF4HipnZC4cBy8M62jAIQLRW+ayLkku
TaUmDharbs98HMXnWZmslZPK0gvfAbHVbbH6QG+9WW06GsK/jwtCLRdzwwguFHhWTxSYC2J0isPt
znHqwSl+uMJEvsuHjqgAf+BzppymGpdkAx0lt5U7Jt/vF9M4o15o+2mKTJc8iMlXbNjrLsxjyCG3
eN4aIlUUEUptRHImGq1Z9whnsFmqEptYK2z4gY5ZcRJDue7Q/NPrJ8SuoeLh51gwOCVvfZc7tSlB
NnrOiIPc5WQIob5EBCIgESnfHGi4ssM4Llj66pr2REQGJyjJaYfARe2zxxIBT2FJ77yNUiTeMhn4
p7B/V4IAZTu/PoMPYq56AHycaNKz6Mpl0Wemo8C6xNOBqJQ/MEVVZhT6c6dprA4vHgrOgLOtVw6M
H1Cqsq7XzsfqQH27WXI04Y0whY6AT6jVQwRuSoS7HFlFHO752y5xEUiVM+VniiCQ/qV4n/Yx/Ibc
nuUs3pho/AehXr1ED7jHsrMzdfeb/9xeZbdjVsAc13WmInGQxtLO/aWmpIObm0fV8v5OTRz3OjJx
iM3rbcYqP2xWGMGXTkHEvJbyaMuJeOY7KLOW7jnWCH1g3SwZ0M5fVr8b9H8x705tSlrs54U+dhN0
LsgzfMU932e2VgsnGHQZLobT+PRiSa9V58vYSwd8fb4Uj+eJ4dQ98bKIBbjoJ7tG5c3ry07LJk2t
IlXQll/4YwjMa5k9Jo5YplvYxq6fFTEXVtCZvXh499b1W4l439l/I5ob9Y7+y+laFAHm9VfcWVF3
1maiOQM9hgwdnOUqhyDif103ctlwSquRg2I3040kxv7LDV3/4X/xymFqYkhT5AI5iv6Y9Hwx5L4C
9wI65+vfehgmSocyvjPCBahi1VDhmZ2OoES2rByaVdrtwzzfJj7h8Xytl1pP3FjCdiDOJ9SejQwt
XMJHeJk7FlhWp9qlQxcupbbetNVyMk3NHhm6wHgoz6a6rw+dxLgCGRbPvxqhI+mvR6d8sSvA46FC
Nxk4XyR4qeTsy+97QxC83sNxqbaJArx1VWk41thXwkFowlTZ5h8dM0fMHd8PFIuhIlpY4jCuod0E
l0J3R6Ma5A0rDvVckdnHi2etisSVsd7vf+zOw2co4HOL8HXU2VnLL7zj9JrhjDvVavPFIeckEWr4
mCi1Uwf0SvIO8VtqmDIYPTAHQhNQbUvNmN/eOhfqe4fMuXjN2HS1B3IjYK3+5mCVBGW/cxxkTKJQ
/JNkbLOGR+IOPXMDkJR4VtnlkYdI1dDToS+vwNIvRz8BYL6RbzO86AR1qS2Nax6e7CLakIY/MrPU
kkTXALL/crwVOru5PRjnYcebsYG655QBLkcpcbb/8PDAC37XujvbPNPu7vbH1YUxmTrXwI8Wt4EH
N55rC13YBoGm6xQBm8vLLq09Ou5KyCzKGx67Yi5mCx4viKzzkHdLgkVyeDqJPxcOn1QUVggddJ12
2rIvmrAlaNERHDKMYQUC/GDcEIT9fsqelLNhWeHatrAb4Vhk4ujsZcFJSGZcJtES2Usq1LY0MG5e
5qvjj0ZUsyTkFfwI6Mz4A5LS+g7YVBeHqMnjMdgJyfVEXh7zOty96Fwi6fofnXqrHnHjJ8iMqoDR
01a4yzsbwqooqaXHU3FvwyE6ekBxGLBHY5xqV2wWs20c7DJxTwUbx0UTpBqy9ldYGve3XdtLnXbW
1NO+k3JnIQXSfKLI9zSaQMrk16pt4Vpcn6Zf1kDUVTl00fcwuuBOhZLbAVdCEqZ9vJnOPGhxMas/
Pyg08tFOHzYOiOKvmjOWo4KsrxByfOjnk6JzjYLvPYxsqqGVE8I4VcVo7M3XmOgJIKeR4fmpLnaM
LZ5POAVJvdUo5ACdP2xHPLXRvWUVAJxg1OSGbBEWpmewMBXlue4fiQJmGwB1CFIsDeqSmVeXiYnV
fLiitCCV/uPExqZ+zjCrukGEyL4keeD01R/8f5sRZdZGXXXPN2W1mtxuBxhavSb2EaNIFcryTnzK
hZcEf5MOVK0+SnmJgkkHhbIw/O1LCs1oFwWczq1YMQXC2lI02ycoGCfONMwK5wEUaXLGlqCSdGrM
IoZl/C4c3Gq9tFzTLi6Sld4A5qV+EZvwb8w0o4N2ACiPSISKq4WIl4fO/pF/fddlamDoBsicoBda
vg8wpLf7Mh8vFbNKGI5ipV47MefE6xVyz4d9N/RZJ96e3fIqn7mB4mdO5ApPNzK22c5KECdKBFBS
paCzq0vPYYkUblM26Ojy0YL5rrbkX7LuFRGe0QCDpT5HuCW1a2C5wmiAyASb/KvA4NXPmCN4OyVD
8cB3GY8XHCcahEe71tSZVszEMqCXTFy0S7sMRZl6w5z4DF/85Mz+IUPH2ve+J4oHPwFuG5pdld5l
kOQxKg1MTZrK7cAwp4I1m8ltZ9R8WnL7aAE3K37Su6H11VTE4d9OU34FpxBULxMzXiWdGNTjD1zr
6TxwuG+ZdeU4dhkClbl7EQl5FZWv0d7RXEO6meZ2DcRd9ibk7e5dBjYut68uGliZnTJWuJwjDQ3W
gi4oK8lCZHRDl5fyUkNMJPJ6oBP7mpaKjthWd1Le9qL65rSfDR9DCo1gRp9QLCCVMl+1I3oMMAhx
tCwoCEMlegt6zkYS3haPwzXRVhh+udF+rJiRz0S8+ar7bsNGCgzB6TxLClYy6Fwe2KPlxg3tmR5S
OLpSFjJZbQCBrv8PH9rE7hT3nf0CKABOoP6eWTKk6/jvDYKlSwqodGE/xUu2J3h4uRFyG7rB1oQo
QH4EHlE/twIC92Qr3eETRD3/rLl5tH045lI2Y+rf2xd9LShec8jkDL2avafluzWlIdwLmnfQHe86
73dZGkB9BC6PSWf3yWa1abLdle31Q4srJ7ikSbIw1W1fVPhZ5oKy2j6O2rQJM+Fi5Bh5lDSvUFtp
XupXQJIpUEl85y98M3HCbSsCcQg1eLnX6uQTU+LpyZYOEIbg7HylNcO9y1gRQNl/80/Q6yOCS09R
FmTHYxuoPj0XZS6SfdNuLBFkPL0rqPccFO+1IHXv63xggxtHv96aqdFTijClnTZ2yLqO5eQOjK+W
1Mvq4Oqd2tWEWCOysbhunRjlU92mb1kHjWGr7VukZJJNUWRUQnVast0DmI4CYXGxzHnJGwubsZAu
k17dXjAZTZ9ZLqIQJTF6kFds/sdmvnUtWtFKr54/z3VQWRj+5XN96MA/gE6t9tWxqEdjPCmUY4sx
yxFDYJDN3mkkpPGCM7gcvXbFYCq7NnGB1r0OA2/sklFM19LZ9CJGb3Cy4TtFODDnV/LP+S9flqpN
WADu5+dvtsPTjGtPo4YvvqvXJ6esGWCKrNxrMCgZFem0q5SRDIpQi8qINdLYqisUBnLv2iMTKxOl
UpPx1himFVxjp5SjmHTdwz5oy8eEGSF3/2PiLNTcPcyFyssBLQbfryhk/Tk102pd7GjU591X7rmo
iK6GIppPZAy/8NJs1llKNzoZgphJowBsSxNubhHZPYeAXSdxYlono7ej52NWjvKmKN05lOst+K7P
Y0VEYw1EFWV0uiBwKJy6FoSPYf0PHevwxWP76dhHHWTxZHv1uoBKbVEhpIoP+88ILOe7k0ekQUAl
bKLMgBlUbcxd2/QkvqTveqxv4oc6BDiewYi7bmzWI8cwjum9B+Zon0CyePdx0UiP65PGV3Du5nFT
men0dWRlSO/rFjYcusjAvHViF67MV2V9UVmsAT3vpiWo4TwGMk93pTXQeVE+77lW/jOvvfD2m57V
bsmr66J/TyqShWMYbk5aSjGYaz5wy8TT/U//caPUkNOBKrko0RIKs7DUOn8r+r3w6BIYiCkEGEA0
1drqCWccGG63zuvceTkdcGU/no3qROPKBTq+TtutvkxVlfG7yhU80vh7BzO9eXpgr01U9lgTtYI2
YGmRW/8fR+VEBCxQWKtqdpk0lYql8UmSsXzEj1j25Ddpm+aJNIi6XOdvpgco6o9tlGx8gI+EMOfw
CfQfzkDun8Y0Tth2KCh8Yby8Oec0FT1DbQNYvT9dyFmq+u+nzPsfKsKwXqjWBQQ1hddiQ578jcm1
ilhggLJUeaR8kYvsbQr8PPGT8jeJ3k4DOpclN8uaXnGYfyZ05eNAxgQJMgwr7fcPOeB5JUT31J/p
RuK6BYA0FMv5CtBOxjYkOxW6MGmH7zIHhGNzowu5DviaonBP2Gwoi+A5WeYgbyqtel6cafJzFkt3
cIb7n7FPT6gr4s+Pw+Ro3Cq+SkbS/vFXNPN6t9qYQykVF0wEd552sASRcnYstVaE8UWngTb/5ekE
bXl3Y6zRmvQBlWFSh9gISuYQx26myN5nmb3Pd2qnWZQUyvmhCXrpZrwZk5CLFdtK+EHiMy1hcn4P
b7fV8qTuCYs3ci+Ek4LlrTvU2Qk/lk/JLO0pQ5CBhKsss3v3gQI3fltLth68pBr4AHQeLt9713M4
us7Mib1x+VjkptK0h4VQOs6sOuWkuBGM1vYIv/DyjsY9G+ziurmyG9jDxy2ZmqdqfNkxg/0fHdah
tL9pHgADIm2xjvqWqLUlgYwfLHLGNG2Hhg2sjSOgchU70Q5QPlcfBKjuqe8oSeNtRCqiTwfJarN5
Sott4jXDdfifPFj5wyH8LB4LpVHKrg9NKJX5NECZ1gFhtCHxAVs55EAZN7885gYPeQG9DsbcAnfT
jO47FMfjNhjNy9yiEAJclYYVZNH1D+QUe1AHwy4LrRoRr8B+jjyNf+oCu5F+4y6afSvJeqbiPSHn
vIMwm+qxgSzG1xK7nk1D8xWnCj0TFNDepcq9dt2HqM0v1GMh2ETF6+rJTiDG/6hIj6kchMns9Kzo
rgWIdhbeYl2UGtF8OkfRZUKW26KJVCRZWYpRu2aBet/415TkZJH9u4lUctjBkCEk9oARkyqNFME5
9stjf3zxA3fjckWBdNkWLrQ2fJMVj17HuEf9ofQc1al7E6v9Brg0a/8t8j8WPeiKpmDY40KRoPmj
Rmry7wzsked7pMVtr46jlz0mD/qmNi776tq4FkKBgrgRQyoqbJmEVtvjZkMVbStXViX02YW/Fr+a
f40eB/vQ5IduXDF925zC8ujCy0yi4gYMIEUu03WdoaDhIX7iLme9Wv3bpauFwc3aARNAH6sQsuCl
OUPPvpwZGHFSmAjdJmfn27CTFgiROEGT/7LDYcC+SnAX2KTIOwPzBYWEXt828jtvvOI5b33EmjCT
/tG1N9KV5u1CEcdUjYZ0fYjvarX9TQQjBw0gkpVfc9RB1wFEKUgprRycn4l0lz3gpoahSkdZuFC7
gdDfowPYMZ1Nuwi3x07aPGW5mFlZK4L+WICsrX+vwaEXPhubnIteGIyp7F1mmAgJvb7tXt+a5PJR
Zz+crcKPNmB5l788n00Rh9uoQJt1ozI2N3oztNjEimADq28i4Hi46i/uhcxo0zWlCHyibhcdsX6b
WU/nPrdrnDs+tKoLlJdPtaXm+0mxmvVhrvTXQw8ljRI1zfK9TicmgqJzLdWST/CJeu+/A0YX8sSy
oiJFX9d/rENowPdHwl/giHqKsQT/qj6+6hCcmJLkbl/SNLF4SPpznWJnHCWn7xyhPUlfUByp96Ak
096B90uuHKj4dKdfbqvvsx6VK+2OO700um95A9pfc7oD+MJu46g9MlJ2rJlhaPU++nsHiQFZ+VDv
mtI0ILChQ8oXBuqkJmccGvOd6tMLSSXCY4ecx1TuFN4NPGjaXfYgzicf3xv5rv6DsVgZlBfcoPks
AaKmL2UxhjG8PPbhpYA4mhuV37mj7hJukfhkJY9sUrwFJOgzenmhqyjK7IbFbV2rfMk3QCx/Xpe5
dbEdfcRZVEOEmnDbvBHbtioh7HW3vWWfog+WFGwbkGFB+vZQOEumP8D4wXyzpCqIqlU9m9iFwL2b
eEdBHxge6prJ+CW2QPj8QwqgMeDHJJi9wNOEtg2CsbM/usMNXXKyW4TWYlbaikxsHXky6UAqUbek
jfQRaGmtO8Z3s29gpmseweSMgC41KYy6WmQ4oiEGtETgHfGO23BCLnbt5dVGU60P0+zdsbE/rWzE
K9BlT9YORQ5sURchqAes3ir3HE4ZIOD7nwv1EKr+x2bL7QsPp8IIFQ5mjY8p5LcVvaAMSskR76Vx
qIXPDeMwskQgFLaCIOe3VerrbepoqdkCj6186w/veqM9TzRve/zr3PhAFDRGI6lyuEe2MaKUkxeT
ZVtHJllpRX02U4Ix7e2sxKU3SqL8I8fC90Xnb2YXUwHTBQN3n/PFQHzdRS2psx3fpdKgkyql2VCh
xYfUUX6Xkj3G5eZJFZyKQbPeIUZK7jXJdw4TfStREUwZGbGOFe314TMECl5i7QTFLlDhWpm5R0pD
MYr2F/k0ZJ/IfVItigEE6YOq/nHfxdzWqTcAFPNB5KclH+NhKLtKiQHYsn18kG/SM1yp9HnZQBFO
9jCiRqYZ4WhDHhWOH0vY58c2BHj+qp5KsAAlzbbFLb+WLb6zPLRSilM4XK9WQQizNyO4N1XwieLL
uLXlf41mNL3X5vfrWkHdKGvzm2uT6yez6raskM39yuwETyPmMoqdzNqvJpqBFIPiOwkb5LXzC9tk
JYq4BNoGwDhPOE7NqGhL/8vJW0JMJ7n99PWa8G8/Bp3kh4N6ZJaDiEFq7m9YCnIlJ+ErA2zQEgO9
RRtzZB2ZZnPR0DdMQKx/w6hflr2evPpxRZHGWx3HhMWYqP1WbYeQfRdwulfDpu3qVYcvaY6xZMVb
ZOpTqQlhAUuWhYOvLz/v34qo7CneAecTgUG5Rx/E3ykTe5dVcvswv+wPFT0ZmJy1mbayAUUvkJOF
dcL0Kw96ThQNKD4S7Wk7zX6W5g99Rw9qg5WXKiAkVtNajuicx6zQ9u/mJS76nm2GJN/Qrz/GpL8T
OpGCdEO7DPRZvHWGud2/9jjKtkIP6OtWD6IZCZ/su+EMtAEdyHcW3Qf2RrStKw5R5LeLdmqzvIx4
OYDxdb/Huum9QycvxHWsNTYkMsutVKeh8bPtWgHfewQn488U0446hqRhFT8Ekoz0pcQ+L6jPXDsl
I1yVEqcYhK9zgwwQULD9of+vNg1PjykxHBmdIAVDWgqYuD5QwSGi/xgyfwX13iHRyuinKFEBWUJ3
XXimRDkqgTPNPV0au+dA0Am9Z4OvIw0kvr0UOVYLDg/jdDwHIdB3WQ2rOOwQ98FElEPn7COwzuRf
Jdp+z53DP81KOz4px9gtnyLJiA0eov75OjS6GTAvUb1EI9feujXWQFV6Hq2hXGeW68qrnVRx9M8j
lFijv4QNki0l3Wx0xgA84F8hI3oB+Si746SyEmiM7DXE3I1/AggU/8dj3DsqbfkAkJdBqc54gVSJ
/GO9W3+LCJwdTfyGo3xEJjnKkzePSsJScun9KuI/+F2Q0kRD8GWJzFiurag7lvMipEEv6P+2mn2h
Gimv52NCwIEEZJ+sn5D5dve1XtgBdtQtiGmSmr7KtvL5uLr9TUoaHxF7lySZljQ9gWhkP740LaDK
xmNZFVOi3y4sXR1YJAB/HKGvikAbKOctIcuCxbP3LPmqKnqja1VInT0x2GyZiW9dRI/i2f7CFsyX
3xQA/RrxgwACORXp4AFBett17N8s5eGDyLlHZMULpHjOGqursCiu1E/UbdSBLNFpQCBZiVUe1XUm
r9J7MOczzXSfxv7zzwgqWplK0GFnrsr+dcYsgHdfM4lU887myagKUoQn+z4m6CFxoHesNBT9OJwn
VXoMsT7hTQJWuMdZ6UhMVZsUEY7hkIKwnmJaUv+mtSr4A1zMrR+QirCMOJ0WHJO25wYE4UMiYR7E
PtFhBGNhr+qPFQWFeF/yDB0Z4bjkHk8F8vr08kV+VP8E2OOb2P9sG2l2W0y6bT3tvjmZLATxKQOW
BdEwtNtDSB5GRoFf9KVgwz/NPd5esVRwt5GNQJ3med6P4hSU3p/raQ4SEEBCWEunpFBUsikRXVVB
o0Olb4siznwTakMDo0o8AhREof+bWmzUirIPcJ1Ey9Yw7kJbcX+/fSkXWhqpnhsx2OV5hwPFPZEK
wDCIXjKdXYOnA+a93+GpP7SzZaBSAYYkXjDZ8R1ZQZ0t8yZQDNt5QNd578W/AnoDY/wP01t8Z+xN
J5RNXG/lWQNg4r3ZdfKE1kakspdf/5TE86IxD+7GtGnR2mXVNVIEjKGh8EvZ3Mcgia88gQeE6KhK
Etd9z/hCh7R3/jFhkZKqZgePXNK6pUb1Af+I6Aak1Weaz195OwISO50SZxl2v361IwlDjribK/1k
7ZeGbH7BuJ5uzD6F6mLrSP884gU96WWdNeNbXPKRiJC9vJtGtnzwzZKbI4fuOzVVsWC/ffsM+qiB
gzrXAijpUqA/vWiUbmRBJ/NVAfZjGKgCcPZtmpA2SbqAG33dyfpEeSynXxhTl/FvnhnSJZeP2Pug
Li+Trm/YrD1IiAMqAW8GBJC3h5YZvWoP2RkC9j12gje3OL7iQNmlUnBd9NtNOte3KgSgifJOuX2M
rLyp7uL1F1CFZojIxLuIpfcdu/Ba+aDy3ijgGZm63FaGTY+fWJDtlTMrytiCGilmS3yLibmAbfYx
wsxj9pbtNfzbP3ZRqDs2qgbFlCkfhRNPOvoff3m31tyft69FV0S6Stl34+8ocm/Gm0ISnjieo2DJ
e1N2XTjXm1A5llhGLCXRnR3iZdc923SB7OXkaLpsvI+5M9Ir/MSALVMuj3bE4xkUj1WADe6l49pP
Wv29lbRYmBLTkp+u9gjAuADg9DM3PpV+UxNXRWSePh1tvorznaH3Zsyo4hiGiTRReVlGW/Z1On9N
k2xAV01XCZUmAEwV21eTJqohnx1PZj2d9EiuWBRLqU3J/hrn6iOcU4VSVvo9I3dW94gcZHLZfqWQ
iRzMZJrxWRjOdP13Px+xwwm2HBNG67ryejO+ecqOxWcJ52kKwItilRSp/H+f2AWXgvGuvIZVb6/N
mhJ8UI+kXCWM7uRa93YT7YYqXSFU4wFl4GBijOo0Ops5+GvZwTZ4meMewwFHFlLLhayTr71jozxy
jdjzMNZHnUMp6CbORFZW9ZmA0uiCDfl+VqeLt97zk866HEkGUaGTtmAeqGg+vCbU6C5cbYfj3JEn
O96jVrg4JvmgUdFuX5QozwOE17hWGvUiNMZvaoYaxJlLQC8xzrr+6bM70wL6j9a0eDo8A3v6mYe/
Fi68dQvuUeRuuIiO1Ur3yEHGN8DWuGAjFXzQZ3mT1G+CX0biJVCaStDkPYeDW0rn0JgyS3d08a/1
yfDfhH6848Z9W3af/du+nt3s6F/QVvZpOZbq1NdluVDT9hFR7FhzVm6zHSREkVvrCSW/+X6HHzC7
7y2v4BjHwfI+Xb/V3NdfCyCEWedq7wnaGDqkUTshG9RkcsNhz96X2g+Jef2alQ7Vmt34ihxTZfv6
G64YiewwjAYJlOB03k6GQhy74h9Fb92mmKe6rfRVuZZpdECcUmVQTZOOybcpeKXEmY7TFh7D3IYS
m9X26ntin/grpRemzCD/DO7cO3zGjM6GuPrWjZ/5WCAomS3OAZBZH0oZE6WNsQJlx+taTg3dX4bV
1zKIFiy3uFDoQDws4EkFyTlAuUKioMOjPzaxKpjSi5syjoPpuRVjn3D7HJ6wr4L/+fGM3IrBAXl+
7h++Cvvovtd/4q8/FqRT9fK58xnru09TifmBI81Lzq9RCd7X2Y9db2uAIcJkpbwVMwmvCc5NDjMY
jRfQQTMuWiUdvzJCqCTZ2o7rJCghNUjssVYq2oo/7mpU3Nv3ut0iSZHUZcV9TrZEj4S1jkfQRx4/
O4Y2WmeWzlczGg5mdvXDzkBI59fTZ0GW60MkfA7LChKGgn/loOraRK9l4S2rxLN3SWtrsVRH1U02
8pbrksz6IbhAFnQ6gA7mnx3Bge0k1gSG9BynD7RzqfeedwCmGpSMDhwrly4Jqkc77rvvjMWol2pU
P/CW/61my0eZZkUuFPXlfWi8cDzzLqkcK+LaRb4hPq28RB5LpXWHoTrA8H7GbczSqTp5lfZKeFhA
aQ77YPTvCZwMLxTO5VV2SClAMvU7/b0M4QJwf+4NcIAkZa45lojvEihrfV3ZabFkTNc8qLmMCGdQ
q8TOGdgAXVlEfSPDcl/CIloxGZfOO9DQpqZ/3gsLcZO9eESUFgIfPt3GdjaQbwfBqcVF9iz0cC2x
6la49A1JwTcVeuN5P/U2EKUUaZLI8S1QzJfsHugChkJY46M9k0ptLGHPzUQmaRDP2dsyoH2Sn6sQ
r704w0fAtdGSPEYLiHN6CkOdQG3/T4elwsOasGFfauaB0Wo8h1q/bt2MhZO+GzQka+OCnbdeCi/d
2oz3Lp4OFBTTVo4sWuQKfQGYdut4x+oAvXuQzeyqovd7KbTsduTXPxi2Ic+Mf32g1Fu49iaBpIlb
c3FQDm4kSx2sy3YpxRTHljpFwPW/Q/xw5QMnq/p2qhCc7g0H4ovTierJW/Pt09ADqhbPQghn8CbC
OiR88NlgAJ7/YHbwbOjToV7bL4LKnQ05NFIYN8+lZM5QR3purhlibIZuPkno+f2FSraa7dzrK5JH
CSydcWQVxh6s+JphUGtXe9ehQJpSWJqFIp6U/BzTG6Dpj5S2aAp97W0fGQUj5Whv5Q1IO7/dHxB/
lS4yvivBAXvmR5NP+IFVwUGy7pCUtKbdn5QGhjV2yMUzSTl1xT7KKbqF6Ua+5n/ysfKos3UurbOj
lOEInVP/hGRr/cM3iCk9c+1/oOdE4m1aJVy9Gn6446WFe9IEsJLnnF8wB2vNPyAlWOhkmPW4JVYi
4J5Fj8b0HVvXpO9S4A575GnHKW2Jtfx3dOQFZL8XsUg1ulGBZdDqUpV4zD+ilOnkHxYlH+LhUP/z
wKvTZuspy45QLUdYpj+wG5zQ7zc3CYiyGvgMhwV6yX/Kl3Lex7Gw8WOlvPVOIFwff/FyCWkVDk0G
rDN7HCQQBK/EFJgR3meKpZk/08xpfz8eLS5jq0TvlNaeckoSSrfe9u0Ip5fjc2sZ9fb6bbKoUOt+
Sg9eW3AxQJvlqb4DRwnXQDnkKTo1KNhzoOuXGFfAP2RjwCIMoImy2PBbwMI1Si8y7/+TxsGbIufb
VuCr+VK8YvuXWkn3NnxopyTV/A3x1+W0ZKPpEj4NR0Oi6FoEMuEi08DHqXaGrd6XU5YTe5K1LOUE
CMOxS3O7FT5knprjhtDMJuZWKpzMBmJDluhDYJMXsIVL7yzms2WxgDr8vy5HCETcvZRujiDQaLBH
wzo2B4Hz/9xuHjOqLVEk/PLfnC3WT8RjIQVQeRxkGuz58ZgYNPW90asomU7IrOPGP2XHKs1JZ+Z5
DQI9W0YZySHyDEV8lA+ppLN/DR6fExERU7kzAemMGIdGhLZMIgip4r2JR5XATOdaOxRBfKzysf3r
fdnaTy/4B1xnjPOua5DFRSx9TP2XWer4l1QqCt2gqpO1DKXIDix2XIlh8iGCKItQZQ7CLcKh9En6
zNUffTsicke8ikt/JruVQ95Yi1xLgizE3AI4/jzfSJta4XiyovjCqe4WqTGlaExxQiAzVcLxWTpX
07K1copdQhEwtV9O2NcrKwwfA27gf00898bj/LAXRajLFD3DGa+mRv051WIdMQR5CowEC9kA2jnI
eihLYTMWFtuFvxgePC6QbMa7zI3dwmOhCCIFKQYtkqImuPl6CmF617gu1v0Fw43NWFfYV91pg8vC
Xmgsc3pCJuGe9EyocAGB7NPb8fPu7XvQTcDpkhTUBp6vxeZtr9BMW5DLXP76RjDd4COx0Pnp1WmV
fqG3zFd2fgZEELGipriTcHWfL94WqOTqU6pGHdJytNMkChQfegwukZ8mjjduwugoO56PkZVvmHIN
VALkAVC6Z3LY1jsGVxctRiIYfCU0d5Seodvmp2Pynaw0gb5VjOzfXZw0YC5UsKE/bd4EXt5aNaI6
qKU01+s9qfV5946zllAK2i3RoWtFJ4YFsk6a38OvQOwJwAhfepOs170jWk/+JPZQwxSkoGjlTFvK
nfJrVRJjFgd9cFkBKsx1YOC9lTiZHDbs5R1ak1gWLcFi3KoLe2pUigkxLnHxS/ZelKfi1l8DQzve
Uc6XPx9SwMYs4uwAqz7jHs0DSDTowrmHkMRCAjC1G4Z6w9RjiBbLfQTDK/a/RdsF7b7V8solBAhQ
2ECBoUt7RIOTm76aIH9JfJIZ1gnis3LJ333mwnrYDhPLyKWegZoBnxzPh54n375em008pPl8o2vO
FLP6Dlb3f8aI9m9836sHbbNNq7HUYWE1BguSQpiZun0z1Gg0h0ZNIlenjw8BwV9tjOuMwUna+D2S
+AXBvUiMT6ieiYRtT5lIvs1PtAqgsZ/9CxVJSt3aatgxDLXFA/p83nPsXUYZl+DmgboXoywKCLXy
CgVveIXL9FdwMljW1JEvoP3VDATeQm4L+f7godrtcdbqvD9Ki0DMyfL7BHhkEHTEhjErpGz7LB2v
wBv0Fas2HNluYfJCP7Jy2CHZsVwt1DJkf3yoH3/B9lrYyRbC60TpQnnGpeyZ2O/GeXDKhrHMex0o
rX/uLlAzJ4TUE0V+6cNMbUseq8l6B7LIR85VXbpW/VAsmudjq7XTQHzs5xKn2PdweSjCCxD7s4lL
9Fx+faQPMzzKTL9ZC8isA7nFn7MXJt8KBbR1yOxDTfaa49FZBgdko4QU0RPVugdK423AoCOCXGcB
XsfirN3fppJSW0oOPcTiPHJC5WAD6GU3w30t6d9WmRYOS2wmgumF/XYVNeGixIR0TGzb/pdhqBCE
3DKwfQcExDNeqXhV5UqHQ9yvxH8UW6pwV+T7HvvqDsz0mFZcbuXGtchnODCuabNnOh0kFmBi9Eef
Uv/Pnir9lD9IXZhFPht3rwenpTqmw0yroMXpviX+nDxRZsNMOmIzWUHlFM7eEgx9M0Qa7ohd0K1x
ZNjesxWdv9HBratwo39cNkxG4UInLvHA9jb/OWR5wLcJwAXooE5TsYzY4p6DuCEk5dVdEHjjN8HV
ZNms4BzuRcCDuZ3dp1x+kokgG7pjqFprJyzJBaMwmJStWI0o02dWcMqXErVCrF8iVREn3az8YxDe
MA/UX07ns/P6/20ZPqIQaz0V5oaKP0jVD1rrFpc0qUKGGwpa53pK5Z8qKj/UDrfA820tt0MSnFx+
KnO7y38dCpp+RgfWoX+9F59gAa7LB+F9gdvSZpTD8S5Wk2szs86pTZrf9vGiT39XrV6UHj6OtVyt
iVx+WGTMzUWCT+L/9OVijERggTRPvVC6ZE6tE2AQpKUd1dT7zCHGgZL4z4uV3Iqo8atUlGQ++EVh
fdAnuuQg7ReOPIbzauGiexRsVHzS9TNu2w+l9tXY4HtM1/ueKXM9/kFZKUZnl7krWxmXz7Y/VnXN
VGI+uq+ySo80GwScAWH/1HBeyVPZlJD5/xTCgzKB+FaDqjBR8HMa/bZQ4ZpCVvwvkzkqolqgeJ0b
QILyZiYR+CnLDl4v/rs8TfbfaS00VFWJeFYf0xw/nb7B0dFXZYkqyTfy8TNZnKAbZXFUfIWTd8Mc
hn0c+nqaX1nkLA5gZxaqzRxRa9/Gy/RuK3qM43FoBxrFD1tSowCA34ri8u0eIa+mIpdAzLhfc9oC
8dKqYUu3/1aaQ6VKxz9rfsp4BFtLOudnoOlrowU+P+Nhthp0Uv4Kzboomg1Hb2CU+vB+ks/BvvXl
xT39dxM5/vOPsLbEbNI0eta24yN1fAEd+uKqTwIFo7i9tjrb0NC/wYO4/BtAPyHandlewIyjb9FH
GxKluRQlJgfVYuhsMq2Ex2l/nDIQPiL4vnEIlw+qxZqMERTLH5oNqRr0yAZ+z2Zg2yIH6B/2fogI
adBguuiXNEGbEeX4Z2RSDnAoyH8wY0iTZlrAi/LpqYut8Seu11fj0hfy2jkenufrqrB8G/1Dx57T
1egUndSFbduGa9pvjGhdYOASEpCif5kM3AE3oIEgPvVS4Xr++bINSg3Jp8uTgOAu6dAcCEhE5niw
B/oC4BQRLW2dUn6qnH3wAvdItzud4FFQVsLUxt6LzehBuQeKL6FaQtUFVRPqQ1hFywRlS7WP9rUW
XQ5Glp9riPoztDaE8MPmEp6eDdEWv14rzO27xo+EcfD3sTr+yQMWVJqH4gGdtojmKTbcgU/2jJg9
d6cj1FJHkGevavNBWfULH3XNLERa9JFPmMQd6r5nVGd/LtYWajPpR4QWEclT4jhZ9o0WesOdhmi6
Of6AfNZSRaPxJys9FIbYF8x+JT7CUqFxdlSNVn0kRjvcJJWigqXwbQqRx+ieVrfl8IsaLjky2tfH
yEHpwCkA51ZSgCxmd2rkGuSjcnkI14703hDFjHQrNVe9s5ZnkJirFgJiB5Fn9EE4jsgjXQz1Q4Nm
WhfqjjjXNRxnA2nz5eKRn3A6H909KgbvYbjMcGGgjU4hVkHxkiwYFT4e/NWOVheBnKDnSygyrl0C
eYZ0e90Ob1rQMGEq4UlQ5ROCMpsek0zZv8c+rpmAzBCJNvBWp/n+vJ1X2mrj9A/MresYg/NyxCHb
STngQifFFzjA+B7c3O9XHlysAAwEr5koOt8Fgsq3v8dn7oyncQ5pigR9okx663E1qWb/+aZqqjw8
jp7YcIN//Li//tXDgvSnKwICplZLbwFcwm7rxNflRytmGW/oOE+umNEZFYPANy6pQW/h3L0N/Y2A
y4+FO8e5ZcyDR9Yi7jrM1sc6MSNoqwzPkT+S3y81lwfqX3boR7zOL9IWjlV3TFjahzKm3g758ZfY
HGllwUwYGaynR73r4BcpdG3Mo+ric14taqoTA+E+vtAdMJxSJ1Yw9HJ8eDtyAoDsVmnjd81teKNr
Qhoa3kvs7KRCZmfu6EcTl01P9jQ2DPCbHxfyOUmsJqFQp/ap8GVjW5jcwlQdaZuwY1hlXrU/g6pm
e1Yc0HArxvRZnIalcNsakGdc1VlCAuq1Uve+AUF7oduFjRyKqtcrTOcQrCn4V+VC9qH4YeZv2M86
P273PxXlv/BhlTDiziGwn3rW8c+8obtT8dI4xJevPDQ7RRY3Hkuqubz6cXuu2+wxCrAHWy7T7p4O
LVvMT5bYw7Xim88NoUPMQT4d5M3mjKvcl0SuejYBb1szlXLg3gM5cGZDxfisTUS0xzgddA4XbXTp
xYXWq/EEXV5tBCm54iPd8wVSRnjh56WAMo7EGUF/wLYWfSE9S3lAcwGSPiE2HSV8iIpCue/1mz4T
tdUjmmoYascLa+NTDhSjCb2LGV/UjgRGcsdpsXI9CDAGb1x5nKWVZby786tSoc87jnrPwTfofvIr
r7EJHCHT8NmYe9n2Pm+mb8dCFLMYdJeaUpoOLCOYppw21jYMTJhzjsFPUQZG4lmy2jT6qtOGr+uK
i8dN3iefSqm0NGz/QujGtyCWezzuGr4iMFETTCDxyv9U1yChVzwka8f+7R6hi1DIptLniur+UoUO
aKWytEm6eK81/9FrR7Jq3pq0hnFSqnaJkGCeFPafGJzExtGH+izsbQzhaKx7A614zKkG6Saku8u8
s7reFQ7TKX0Upz/pQm4e1NXVGOA2pXBlRvvtewZdJwbQG4r0gZL6P7ztYwaM32hh/g+7Z/SsY0K9
5Ieb+RZpQBQd8uKhzfJPDAigOocMXRJQnvnGQba9Wz/zkOpFNKQeppNPj6olJLPtO2j+IWgvcYjp
6dXfiZRH/R1clFOz7Y4ypQaetzA0u+qsYqdKxfgam9Tph2AYcsxQJN1PqllAug8Xux7DGe42FimS
d9HbBFy55NuWBFzLNlg5Ti0/EbTGmRhTHlT97JO/Te0PvzWiNY65txjfOSOLVk2a8FDNRCIJcBfV
KkJK/1EUZvdgXh2WTu5ZUUjxHxNb0Q9dQkMwoR82DE178JwTQbRvFZuld4mfsqUJTj3Ppqz4Zdtq
+vrxcHpJln1BwSqBxwDDtvrw5Z8VX4BNme/Z9dSEcriteUXQodCt5LMi80PL1viykjayS/2rfsb7
7CcpUQS5qnDCeXOd30tXzQ9CYMjkXDe2oxmyv7iov0IdDK7BVUSsVvGWxSfnAp+yQaCxrG2L9Nxs
9CLTBUJYp8ohV985iWwpk99SL42XEk/thHfBZ7L0Ix+XJ0dz3Qm4q9LtQ6sTaa+OTlrPm7I0TEEZ
+IuwzW+s4QcucXPWE/He3ubi+5PZfHn+t4kRAXFtufbxeqdjzwo60QSmzQ1e2or7hmVCQpeeH7ua
dUwLVeEThM//Sel/BkdVYBO8UpRPVXAo8PMQdWay/76D9eIFZckuy/QcsAVScg0NygQVr66gbyOH
khf9442CNYNLOssE1t1qFoQK43/q2B0cnQ4XPzT74H5aTOBKJr+L0bHKUFUXikEXGuN248CRzygC
Or4S+oNEcgFVcg5m3A2dEbrL2Ts7AllMHe2+RRBM3kiq4llEzWJGsnpSgadtIxZzUc7TJe95Dcvz
t1rIqPx3FQXs37ohsvny0JxUC3iYIKneMi3dsAvDvVtAiQYOniSSc9mOa4yl7T8ekui4/nojwAYT
HOHXnlul95C3unHLBhq5XYvGzZg2qbBRJQEnVBeqJDrnGTlfesV7kRPGfaO5kNM5hmARsqSgTsRm
3U39a7mFxdQrYah65jR0prMpoIPDn5Vfm1h4tmUmEe6ndyGHQEgGRmeSL3095luSGB+R312bq29n
RVtR+1tCXY6o6JHpkkm8wx7Sv4xV1o9BZ2TCJOvvPlkPrcavVyGBGxFrNExzqRgSAyAlGTApxPbd
WpSfaejUVSrZBObmNTxCLfSCSkcpjF7FOsOwWHa66gkRUF1Qpgs0MxjXCdkwav9/tv/6unwHTVUC
WLbFHZyPkFXpAnu9+Xn+I4FA6p8YynXpyhTlYuUW1eMD1yUCa5Gk37ns8pi76fGF4ajOabF/ZfTv
hgyt3u9HGLYXW20NMzpUrEbJwJwhJCKnr8U0xDzJFsuzS3iicLYoz6mvb6z+AtxeNEbUUdiny5Ea
G6zsPakw64CV3EHKfWHbcBbNyr+8g+xPNVv7xd+7DnbAkMZB85OKSBujnrh1dn5NAV82u08d8ROB
HdP7hbtMJlxK241cEKkxm1UombCNMpS9oVtkLhkewgUz2azS+SmiukbV1QxjWWHdWmxg1NL9XRIN
M1TDrOwGK4Y7DpUqgiaDBuuWtx6U/wfOPvIWVKpj6jgxLjZh3mPoG0nXxoD2kxZp+F9w3w4R6kST
2iYlwvhiGrLqZnFj/69VccWIEwCgeNpIt6YUdvDgeXhcAHA6ecsuj7asc/IHA77Pzi/tINykzUcO
HD5HZO9t3JwyX+SWG8ih98KefzjrXxlhe0iyXFPTFuXCKFzdZzq2B38P6hrO8b10kaPfoTKEzBIL
Eif1OBxZsdphlw78zS3phba7epWsvT0rrpAEm9NEzfxFSdIGX9q64iLbrSC6UxBTpTgW1yEJkgcL
FjbKBSxD9Vu+pOKYsdilpVbA0YK+mIwoOXU4vtMIc5MAnTb18NRnOrH2oBmmUx54+1bvX5LJ1bA5
kMuQOAeYVM4ZnQVlvc1K/QKnx7p1e9tfi1vm67AyqRQ91XYFxXGwmzeelF1/VuveXe2ZWQASgAxh
+pKPeTjigw7twWjs9PzQmq6OSGfn+4DdaXzCoOf4bG21a5uGMYgLwCI1WgYG14utW+/NuGiFleKA
LcA/8w7p2rFucxeomS1pzDwgc5qyaHO3gKwJEJgN0pAubYeufv3X0PnlhDiRt5pH8+pyabGizyCN
kVPG7T/LOyQYErqKjYJbGfWIVEAZp2Lfivzm6rdGPsbyv+h+ey7naGVYA3CdtfHO1hOh10XaJMDM
AEtDxWAISz1QTO8cW3tNjcgV05nzOgr4DwNQsAC7ps5snsy5z1ucDiKvgAKuoIQGIW3SFEbTIIdZ
Ub/53wOV+nFdXX5JEWMGnVt7iqN7i8we6ZO9E0fgxNc1LrZrMl+M6AJS/+1NI6lxV42Hs586M2cX
L83MD4PGnnP6aMO48F1X6x9t9SuHuXrrxgO3lNzBuEOijnQ7HzZQIq8G3menSag5cM/9afKNCb51
BP5LY0UFQtJLNYcjA3H0H07CUuNFae4Wtv2DOSN10sA8tpAxZhxSueVUr5+88DHjK/5JDioDG9W2
CugBpa1j4U5cN7bwAsUJyOpWfIfgfebSy0DjCq8CEVyTeGnfqHWztoMwStxDiSZeKftvBgwSFZiu
WCuwCYGizOhMSS1/+ELlf8phc0wZGK5oAo+zMJ/geOa5y42Nd1xlpQ2V4eDspPs8cHJnBjRonMxF
GbA8DqJwbmUNX2pnvwhKq36CrDdI53obHqJXa0vjZyaedGWMF/tFFElj0P1Z9zOV4sOAqfpZXkBM
bjVn/LT3zz7xGOUqzQrb7MCOORu6HhuT+AL6jaJ/6lnru61v3AO6KcdNHQBcuCybvEepEf3Ub9uT
MVJ71rFR0dCGiIPFG5Vx+8dpLRQAlJn0QKswJP9+HeZDRvlD0miCoy4812CTz/8Z4Ty+jMztpPj8
dwLehUy0z4uIg6JbFiPL9PcCR4QxJTxrPPEvsxYv/GX3ZZT5F7K7nuVpSEoy2uFMKhldcpevi8qJ
9KQxy93Ci37R7luY+WUbzblLoEj18j8TwZTVA7vAiQx7szIbvt7HgGNOhnu94biQd7bKh7ywWZPE
SiCQi4Szzzc1DR+sXgZHFzYkAiwL1abV17hRrWYdBdkwIQgBbtNWBdkZ12K+wCGLDXgzzMYFiOYR
Bes/AX7yK8mFkRMfl7hmAQOTH9g9SBk+ujxIGf+pECcYgTlTtQSTReQs887eYYvyp8xlgMgujma0
/qWxYB2/GqUGpfWOXck806WFhtzMO2q2+J6RZJq7vYeO6Ujohj1JwpX7soZdnxkeNgZWkQOr5O4C
5ycFGrKNpnAgTqNd/IdyRErr3OJOouyfc7XntK6vPWkVYsiv1xIsLTIs7jp+lFxfcVMHu1CRcLmq
pG9cFccRTAWe4QPym0eM/lUDRks5eSRQovtlLygAs/Z9bDere76vK7Eup7EfVVj+xgXdSOY87EDA
ox77c5O3vIsy17fepkmwDWzcJ9gHfHNnpUuzQllktoQRXO7cWLpfEW2Abo8B+CxiAaBuIdFlqetL
XmFBNKpXali/1mc7ldx72NjJyD7xV22TCYOLpPeEJvg69/y33OiKB1w0Ji3uiEd9KHffvGethNtO
a83v3Ea1hazQRr6VwW2/jaZcPlad/qPRxA4SNDlo0Kzg7a6yynJKLPUaPvh8qMfK8gY6XFA0Isgo
FVd8RnB1Gt3VzVgHWQXR3fekSNYLPbjOE0oQiE0oAIuyT11mTSMAFwH40tzDkd2wJKlWEA499aRv
D53T7UvX9FWm+Bxik5Qus3O7ngwIMUs429qz8/XkB45ddhC3C8rxhPJExFH7BJZ0wLUjgi6KSZLH
KDrrtlQQ9krc5lbGWuMjZ9IM4nNK4Zi4wD4jWe5BChzCWKrsa/K+VSqdyRdPUiIEsc1YkAVwOD0c
hPkmN3A7ZhSIEVcIwZaeXbYPwf/5tKBpCG646N9gIingPw7F/mlLYS8iWtOFFBL0Dothl5h1f7wK
ftDgBukcE7usR6z3z7Pn3u8OOTouhWZCOItoEGXTrt2pntwVG+wSen/xCIc7HTNIZLMgjgz05yJ2
Ikvoq4+c6nO12uJxo/X9RsJ5fwRWM850SnCmhXN8sEUYqQBm2dDbF7PHdUbXRpF70ikbEsYS3RgX
H6p7/9rNOxM/jZV0o5TADfS6shTbpwJKboDlvwF1jV+7z0+3E12e+l2MJ7pgB7V+voIMHm1dd2s6
eGmthSto3Kbjtjfk8ufUJb5m0jU4EH2PEcLHqDmZE0FueC2BG5EqtNlyH6GvHiJl9P1ycrnVbx9D
EdEVKsexRDV+0DtLNeM1607fXSxS7IySGGZy9jRkAgCwN2R/k+fkOcpu33NHTYkY+GCkPwhCzLNY
VfPbTXfveXYPePmdwTNYW1GzZ5sFyyAQVH9LP1/5QLqIwqoL/J+82i6gIpwoSn4gagBJwpCh8KGt
5oPtccw64N/2nsDb7RSKcCIF4pmUCb3mxxadWiTbZqo56nEej3nxlMh1Ft0RAuO4KT2+m9e6xlqq
8wmK8ZtcM9ykIjezWwoue98a9/8QK0N/fTuPvtxUIVmy5x5iPN8MmeSnO6f8J7FCVikIECxIVZ6J
mDAZfgU0JyPdvbWLcMk2kEa7OF84RhA+zKJsVVQ9Fjo0bWk4cZm1N88fhwEm25BU2vts6yfAZRSD
alekGU8c0TS/Xy3/Re5RL8laJbfA2Zx5y2zhUN55tLV/B0rRmPek8LVKv+NvuhdZutWvEY9Stzxm
OyNSv3DgOhUTBA3lee+cRqYbUrqwZuBa/EUeG+tizdY3c4Mv2xBlLOGSZ/XnpdzoNcOoYqbW3L89
wtLDxnmL4RAm93YIs3dDQNypI5i3523Uk83oEGLqJIthTu7UBYkPK8mOEtPF4mCHbW4poDvlb0KF
VGyYGSv15RxybZoDPLAUvJrGhOLF/Ahr3Svj106KQnFEM7E8Fl0Q3qCbUm5JiaCxvWhbgkgCJSG6
U4i+6CtZu0RACcoXfzvpRdYGrp50MZyrozjBClqFyuYWWgQYFQNTWJvPoKvAFSePE39+56I1g61E
s78H57fKkGEilfjMelLv/uZLKL+vlLzQYrzYENnEYkEakagD6ypEfi2aqZVCktu7o3Lb4yoZO+iT
P1vfJv3RZjBz9uyW76SLs4Ru1+CW/bE4rM7F0+xtGa39b5nVMiydR8OPhIZbSE1+HFPUzmrjKUWt
oA+ueT61vprHvh77BWjq07VSSiKWKfcRF6WcyY3uN4cyRDmtrCTdzSVW3VdfXNBM+mmnswyyrvMz
qD0SCwqtSRnzLM/eNBzAptYQ8pN5j9/skbpNSn3at99pl0Ji03wFh3FYrcZErVJKkePqyapY4nkQ
aUYM8qqxwTxos+YFNgDwe63fjzpTAKikWj4DWl+5vVW0BQv2n4PzkT+HyZH9TVPIAcLMrjQbEy5r
1CdzE4VF4xOKb5JlG2h1PWTVMZ2OUvLgTZ/cTspwGjS8WjLxwB6RHl+Nw/0GYSDDniEKM/fCmf/w
mBRH70CO1Iu9CDdq2nEvsWE5ApJBi+EutonHhZbgD871oZzgZF3s+bAg3rj9jU4OZcu9raz2ZSEH
GYgqMLNQfRp43RVhApQzTStolR9o6gN7JLZ3Te2p19SbglCfFJinWLdvfCGcUAIJTrRGPxq243lW
/FgnS25Ruv8OPUu4nGJhghvOmOdFFGoibZ2TLtr9sJdk1jvfkj7r2DzuOK1ivjg/v4GhAv35NzU8
0NI+P1wuU0S5w2eA3DZP5O1CRsHqoy1rMt9uoKRzbWZs+4Lu7opY4p8MjT4+SElcJPzvFf5pVRTO
vfZINLkkoF1yT43l5v1+yhH2r0/ZVjKDWXDgiDu/tfbj/J8G1YXlA+6rQ6+QlBqUwRVtKNJxdt3Q
yJLvhmLD+yC27bCoWx45zQkO1F2FXM7OiA0UOLllhzPuN5tc841ANpU3C2MHa6cAQAElipNlkZvA
dnoGLAqie+jzVqzVpJtsRCgnzcLf9/DwYZFdscuNuIJMCnsy41YnCg7yapNzFbloE3D+/prd38Hz
ChonDQYxQn6cJNj2/02PZGdsyDMvTp83iQtthONJas+W+ht0eTl9iTFugMwx8I3Kkx5Rsu+KwwR8
G0RACbCkQj9cVicMjCWVemUhxVi+BOUUSgDK8vFzEGy0gCuN5uteWkIwKgQRJvs5XH+nrSQH77lS
G9LluAoA4YGPCyIf3vpK0JudOf53YKZQzwA+QbMg3wi7P81ziEwcBHwmoEU65XBPvGbbSRNBVj4l
W9Bgh4FqE5XhPBGhdc70yVTht+y2LNZwJIUTVDomS6z4sK6S2NTXUvfKNZwtWdDacuzCGNmnWTiL
NlfHxsbW6wY+6mBLoZImqPwGySAMStD1vFZDmEQ5xbyaR93x0VHxI/qEuTyOsFHsPn+4LtR91JhA
9b7XBL3zO8EchvXqrw8bFVRMBmtGSler7CUWGQKYole0LA7/iLJFHRmzHPBjDxjTm6kRw/dLIaJU
u1AOP/YoJabf1aZnp37b3OqCl8X2xq4b3UB0xez5MtXV6VNUvCG2chnz4RWyjO1ygqAzsmT8uNy8
NTZB+6LiJZHkpkGOlMJWuoIt4XdAl9N2WWIgpFt2PfVnVLpGDxBNDqVtUktnTf0e5dzXGYz6KXGE
pC4ET5PHS37jxBrSuLtESm1ifxG7Zg5aNwNxz5k6qSGmAfQmYNMLpIRd0sCDEHecfsRfR3YHjlXh
1kGuChUaDs9qYwK/bY+ieqYMh89HBq64wVvgN50KpI4yYqc5r2msXGbLeqhbWCWvvhMzCDoF5rNO
ssZ+mr79l+66hc7RDCgRK+aIrjIJkifc0526EI685ax2UlvV20ofUkARlYFo+Rh9yJsEcnQQsSO8
FMk3k6plq9XAngEpp/WrhCMZiidv2JlPxRRCc/DdGlw3M/SI2uJ9Hmfrhg5W2FIdIGuNnFH9QvgQ
uztKeYiGq9D1ug8IQQtr/Iv1VjrbCgza5D9ePB78m8VahouCNRSnoWyycgwtBZACD1fEfueDG+sW
xxOoRcEvbWhMzqneKljo0mU7mxrPQeMVQSmcn/krirwoX0LCgOx6766eaQaMGg0YnCjL9+3EnIT1
BGgZYFBEvH7PWWrZj4SLB77gFIQqBfopBIKqIfJzJpbbhyHsPsTvoFChlR0cDiMNxSTcsyem2VWg
u+O+ekUVhAcMm9o2MFKkOqUjmbjUNdKmsTpXiORdcaTVei0yEJYBf8w3Jnet5bUkTySh8TXasw67
xvnYDn83TFEXGC7kA7XAQaYj8e9qwQ7SE16/gBfMG0i84L7fDIX7kCs3zPtMuy9jkD8auY0vusv+
aoO3BB7QQJAypca4+VGqqB6roX5GA6BS/G25pNJZc3dbBDSEwXpkP72L13JrnbMW+aZGRtb0G5+b
TqiH0HdTUAYIhvqY8SXpUqEFQtvG+PixuBpHaxbbxXts7EPdO+k+vq/WhZm1gfAXoVvdSIt2UqNH
7JL+OG0gVWFIiiQX6WTI86Y6G38UHGuNyY5iFH1wXNVF9QZdBnR4UJFw2abnI898lOsdYOM+VJAJ
VGdm40sFugINnj1o0VUmqxb1nmZXNDXZbywY496U5dOSyY74M8EpWIwkS12eqbca1aV7zCzROx9D
DSIZT8l/WJoJvC252y9xKkva857l2eRS1+lDJq8cCjC9K8LtdiusWEou6VJ6P61tcadEn4mLQJzy
6WceWKjifludPTT5uGXjGYkQXlHf7d9zL2FB0BdDI2lpp5F6F67I9Q+Gt/R0UKsM6QWzDVg3K7G+
qbh/G85aiWkbBpVeu7wAet6Akvs2JIUPALVjGhWpmQp3xbSgv3eUVDGLNmcI87lTr74r+piNfFcd
el0FmPmSxHzasKFSzOzh45M+9cET6v2WmP3xpoxqk0nIpDBCqV2yc1TtPBTg+IXOFQ+MCIut90ka
6eT9AZCSJ9RyP1s4DEVZh4GsOFh1Wf3R3hXaWtUmcgUDxDRHT23GCXO3lSORQKogUcUmrhXhvDhK
eFGDsuQzTACXJAoFHMvxev7MVmqX/GwHK062vT2Gf9iFliXLPD4VQKqOAY4LPdJDEPGzlKFye/Dj
xIDPQICOC0px3F1Fg5JSJ9D6MzgVZamOM2eHrulphAwHIQVAkB9FopwFIeEZBVB5SZXiVFNygVlo
HaD7E6hMsEAo2oCTzUftIgkFdB7yurseTSPbhgBcofXhEGHlyt5mMC8iCQd/OobA/YZ5Gaj++rRu
XksYsoXXUDfHpfo35J0ldRJQLjnoWMvKHdfCib5m0XTTeOIPLcRio9wofMQlUbXLVXoQ4AjkLPWr
8ORLxCk6fvvcmRTQ4lNrzCG/g5WiBhJHBqxv4y7kj92rvdZZBAdp/WaftJj/xCBsAPuZEcbJybQk
ZX71j5qHeZWvadSSKq+ZBIsibQaa5KWF3oDBRRgLV+83K1QrX7r3s9HpoeBM3Lho8UAy3ARFI1Nq
UzRHEjRA0yyG2BCqmpvbv0Cu0m3RWA5dO6IG3qZR647V+NLqc/ueZlBZNxy2vsANylu+v9qPMqTJ
FAmDO17UjNy/Sg2ZpUtd7Nk0XNAhd1tzlW7E9Ic+Mr52L6i8OCGQCEaLb1jEnomfx6jc/dDSRWSM
5D+Se8wYp7k10iT7oR2b5d08SOzOHn7hWhVIb8axvTbsdl5OhwuuueBSWynVQYMBkb5trxBNqvTm
QWEBWuCUY9M9Wp5oglAaHRXN5U7up3ECD8LX+E9qw2+mKeZgMG8ZfT/KdEj17R6K9DPuCFkCAUPZ
G6Nfe9yc0dwUNJBuuu4D/C7QPDvDuDOM4flwCQNJlmUkryBJoBHs0YdvTLDGDs329eEohd3lgNUB
Aa9IvYteR6xLr/ZOMGuBWx+4n41cAF6bElBm10qYkHWalC8ip4jGq66iyT5QgLoEJIqFHrrCu+us
ri7vb9YPz9up1W+AX1d321NW1L2BnPomhhnJcq9qGfzUCdp2SzUDdPoHr+AldOFz+dyQZ1q1hpyf
bQIX6jRL/XIz9bd4xSfLtfa5pMLOq6yTjRRhCK04o2siSuXkaJFAnMgj0B5nYx9DmgmaACzI0V4g
ximtOUbn7YlRiMahnccpgi6b+X/b/f/EbTSeThiy7eQN5uyCg8IL/PdxSghey7fGi0Vzl1JZxuTH
rpJ/Ct5YWQh6E4FIPq3YDgbZ7Heq1mj/0Fw1O+kQWTi88yPtU+GdzXoj1UJve2JvI9Kw4EyzU0y0
+UVz38qVz3SKpmzbcXD16M9GDIPNNKHyXfBL+G34JcGBt0oB4nxUOa9yKSgS/Gw9BthnHt/fStUf
Nrn9o6Ne74ODZACCYyk82jo35gBovYn6Cnrel4LeG36La1QjBmLAR4mM7SKlhdnHGeOmJYMMTvAC
hvSR/Z9yweWUcM24qZFnpvo95e5QgO/cVJu85l789Ho8otSCpAvuSbKDPSXkbXUa+ONQHOHVkPon
E/yx5pUvdt6pNk7sRfWtvl2AM27H42jJJFCzEUX3Ia1cdI7OyZaXxDXfJYApkbEUKfDwjHbltx4Y
uenGN+0L5lT/cCLZ4xbjEXybucGnQgpsck8QJimuxWmnFmSoW9Kd0fPoyx/rItnzaL0/CSB52pCh
DnsRlvWltClW/lKiJ+NBIFI+xrr4FIXiKqJig3qNFHx4QXeSingg3UUd93NGC7IQ0Z6H8d9TcAGd
Wo9527xGEmXpdDepRTbC5xqvLqrKrII3SvSKrbVvQZOO9+SD/7khYI8roHm+Ev2GvbmI3Ow2zq4V
x+nNAfsXxMTLbLjaNZftw2A69lFCWd0YlxAS2QVmxo6dX/KHbsQolWvJyshAo0AK43cWwdP9hG4P
BQewTWR7beCSC78VZCQlo0uow01TayXABfNJbcKPEfvpCwqn9EF0zigtJzxVV3Y+tEiDkZWeICGg
jBO9vsWo+NXl61okJbwppb016+m4VKT2tjKDTNS8jw4lL+w7Kmve3j2qA876cxN6mHCy2lrlobin
U8fCkv0F5pUSB2+Z1xtiv0qpZo1AkzAiB8WP+B2q462ODT1fkTOpaYcGtFln2+mjjvKsD5QegPd5
l0Iv7aY5w1PaaMZgy16fwZvPrJcwwZhNhqmFg6jJS58CXZcBysXer+ZXI6ksOElQX6jZGpOcfuJL
CWCdsu7rCDSYhX1J+VnsplVINW6PNQBJ6au6rMZndZE9HRFtFyx0GB11V36hBFznrrfEawpj7NDy
oiGQZtds2DiUGlXFWPKrGB6ebLGCMCRsHeU4I+O/9i8GmeifJqnADg68M0SkQm9jZVqmeoqEbvXV
gGIomzk3DPFaM8dfSaW8eWKSHQStSTedH9YdzQg+ty8bCiwpaMys7SdaUCSLKeL2I9H/YdOQfGFM
Xi+TdtletF5kuqhvaOOLbPIR1LsBKDJHdpJTnxhjG+fHZZnMlcDDiVcim1xfy5CjEGWm1zxiIZ8S
jmoA5+CJ5iB2HRhSQgg8GpgmNewd77NC6Vouziy7zJiIvg7dH/Nc0YUUMuHRbU13FzLezpJSsqMh
S1GlG/BIdey25IaTAZ4vOqs2TDA9sHWoDv/qYtWUJX15fp+YocegMJqkLjypHHoYRKty8SkCcqZz
NXnYkuN4VpwmboNApvJp3Ud+8/u6M+yOrdStoW9106cApxH4k7rUVZgxizylPUxuGSrESmfh2vFk
2ALzIEsrLtwPR9a6xW2WFV5aEB6Knx+Ak0y4vEF7y1EYz/I6+XaxAR0nXNX2CwSIuDZYfppSF30l
fti6TNW0T4ucY1keyc8cbpJ0MGZuafShonUAYp5XXvDCFwXCXU6/RkJtD5FHHkSjWdkTJ2/pqm2r
JJzYHCelmaSIw8DlBu8A/qfZedKEJeKOd/VFWHbinEwDzlQwXvNHvNacmjgYvpbRZOG97Jyuxsi7
ciEeVxfhJv1i8qQ0jGg5sj9k1vAFViifXSJeySUbcMj0FPN9e24Xn3oYLhmNhUt6mVOlnugAg5Vk
kCmphAyatzmBQP9MMMKo8xp7+SvXTVAPENpMDjJHhqYCoNXtf+tZJwbnu3U1d76mCU9WMYQzTTGS
z0cophl8PPIdA6Du0CIeD1rCfm2E5x0cccKFGrJ5L3pbhTZT9La/zS5pBnNSRAk002PS0iVh80Xs
eZ/bvC1YKRXh73wlE2jMa0WFmyyz9snXFxeO54oH93qBA6Gq1olbEj1Fp86txuFNq4wuIy5FlVA7
MnAv2eWw+p55lXt52wnMvww2l/5pRtwJtq2tc3+eil226WoZkbn3vU/XgBm/Oa71Y3pACzDrSCqm
JLEBTv5xRuCurDciqMLTmqyf4200g0I55BPqL4LxhI8pRFK1n3b/w4ENlBmTACnRdjuc4P/tIieB
YKF0kXuqc/s9Vxq9wC79t6KB9sFW1W00esBneAkPGecbbNr4SjTI046UYGv73lTh1B6dmlkGPNLz
wop5AWtItlxHJdn6b/3AkdPQBhPNdbLplja1M3q2oGgSL6zFMkUdOKJSai9efCHeCYxSzxRDHwlo
CO4pTEF1ZrIofdbgOAr0b2GTwpQaQfg5L5Mt4pBuiubw6uXuEIXVuHzHiiePyZEBbWLk23prD8sg
idsIHo/Si1xQKz9LzjzU6qTLC2njzuxeXfY6u8x1SxjfKGliPE5Mhn/xqsgNZAuyfNEm2/b/bs+v
qzGKlKnHQUJVVv8+lbOe+oFYxMZrbIgVsTNmZAuAPtXH9oR5eps35NmadMLgAUPrJCKLvdKiFCy1
JjY5frl/iWDIXfATTvXg9eoRDhTL+iyZ1VdGjXi4mfS8WZTwgVYe18n2YI/eFqElPg182GT9lFWt
FL0TGzfQ1JmUte+jWjTVDNgKpPi1OpoxbvOvyvd2gC6PpFEFTz3CKKYyCDQgVzxv4A9UiDd7tSbe
UZ9Ge8pGN2WXjR8YdZuZaxYu/RtKXE776ApTGImy4/3w4yiuLd6ksY5+t90YT5Q5legUZepSxOKH
syB0ECq8a8GtXiKJs3q1hxQRPv9Z2c/zSCqzoaUn1olYT019/7X/qMObamW/mZAIf5mtLxCOhpsm
VlXwmyt2ufayH+WpcRtlAare8l2zhS/KN9PIum2uii2/q1NEp/71H01Xa/tIRUZJdevC3S605wkq
2EkCwQaP3gfr88vq0A2muj/PbY2XR/RzR3ApXBank+dxA8zu/eTf4+s1/2clo9yqtxxYkA1pP7rE
Ks5G88bUZkmliAwOxP0vSfcX5vwYQalV99Rw/XBczalnjSUGcQQMp38W/8Ofs50J7x5ozVM00KvJ
1qOGvf+jNd7PK9fPXa1dM6qxVA30sLInntemARBrgWZIz+J6PMOdCx1leHXij9QFeHbzfLYrmqHJ
5p85f1s4m52FWBP944Mwpi5FE1HpfqEvxwIWAq9sm0aD72y5FPTEWxrqeP+VZSBx2ac6THsVXAuR
I9DvV0hGoudEyx+ZkC6NhbbvlpVQ18NgdGiSEdEN5HD/7EFkooZUKi3GZCd50P1bvJtFPbTz7F5U
HAckTwdzccAbX5RCjXIs6fzv1pDg0bjiBFmnWT6pmWKOSQ0qtECZ+55XekXpLUTgy9b7fkrtvjQY
RrfnFpCxEb+nUyp2UFB6EbX25BhNPl3SFgbtIPhKwa1WZh4u+BsinDYfCAu9AsEKAWXRQ45rzS4H
bhRklcM8/VZStx0lYvITVXm142BI/yM2EM+m3fy8K72FpBwzqNviFhaYyWX75CyHFSskfeAqFTVp
V/6/yvzc6U4E9t7u5WGyonghDa92HTqi8qmywfzTCK4TRKn2OkOwzQLhpY4qrVB2hU1QAYls7KOg
2CmrNsC9EfRjbi02orcv6ozJyPlLoe7kYQ0blxwH/PYtIryKFssQzNyMEIGx+owlqO4/BxLtMWRw
lzS3SkLUvxb7x0SHMTQyhg+gaV+zkl+JjMKLi+IqfUaT2I7jEClsJINTwRcYg2F53FrOjPdXKWSC
mNpewiqlyNixuL3HKaqtsb32U4E4KR2F541nER3vk2w6FStnf3cPDqHzCPzxxDIrI9NAnlPN7YbR
Y9/gqnjHuX124TFrTR20e0NvJM42FniV+Da+CjLlKVZertQYEFrujFaOnXOflvL1HedC9DaCgU2U
JTvEzBKVGlC21FhaAeN4pia+g9S46tEtDHTc0uaocOfh93XhLfkhryBwGPY9IvNq13DOiD+nDk+l
Yf4h0ARQ5T1nitn4tXrJSj3GBFw5WDhd0o3c2eexbEBaO3vakie9nXd2FT5GC8aefIxxGpY2HHGa
9f7WhwkhK7nGVsgvkWX3Q4gv5fc9vShuAOw0R0Nov5pEkSThaRQB42T2A+3uz+dc3uXBMnBMG9MJ
HOoY6PzuU6fRPtzDAdEiZ4tEbHpn51wBwqCxGsvH4t/N5l8LclsDqPEom3aZNQplrMxEKNLN/Ylx
7yelBfXHh52qcgSaViNPRETU8bSWtnGnE5zD27rOLUWEGfaAJ8zKCyTnAhpEhRxA65f7bY+wxlAt
d1QsM3t33TOoZTg5VSGxm7Mti1v3ZhCR2KS2wdVDGkZPIcmw8EHnqB9JxUJwJ1mQgJ+/ONAgDPrU
CmNdGFwSZzLmA9qMMeVqVNAFRrNizWU0YBLMTXWzfvDUCqUYhfVMhAxEdw2he0P8p8X8pPmjCZCN
4oN+10RpDwHq4D4ix/KMfdmqWiopCcus84YJLw8coSh1V87R5hJVOvc63kWTQZ+FwLlS3mAk3pSA
mvg5nLozyEXpMX7eZuBnGJZKR9bwC3xnpiDmxO2bcRtkSd04J32OxObPY1Nd2nvjtqggEwbqQ9yB
4lBWt0aIdNoHPx2El/egJjArWL0EfXe/m7/zZFKpri22HMpPC6pYbbZrnuuTVTUwJmcC0GNiBbmK
+D+sRn0T+wFDaqTpOXu8mgfiDMGLIDeecWgC2Ds+qFlvi24tDiDLmObyPuFT5k0Sx2Us5T+zo5SE
4o5DwYW1KAcgrGnlZSQA9IlWWlZKuR2zv+hTRB7tzEPYAtX/CCBDsv7THeqXr5fAE+65+mRrAAfs
4eKqBFy7ojcjpOtT3OsitazuSU+eYaahzQ0WQ3JGrws+6MexDX1R0wxfJce+BqgYnCQbBVj+9zEo
MU1dMFcZTnJxtEjBZTe3mbmEITlvkYCaVfGSzAGaJto+yBT5j6rP7kOeNHrwHw6rxmhWfH7Ch7Mq
RNg8xwiz43SlO8lnYUY/ZCJqD32JaTQ5QqJbjoQu43Rp+Y8KJdftbVY3aUlFgiJT/TSdumIPvPNB
DeM3/laPzwoibbadHrq7wmicOkGM5K5y831xI8bUT30GXBT5t9gu6Vmffcw+9obz5gfn401qTW/v
Y86ph1IHy8GF7i001jhaxltSDj3EtlWIZOmgF3qhCXvYSQvVvsWMgCUFhhp1a1cz+znMUlo70lqT
bnl0kKABDiuTrjvPl6uFoojy2KvPsV5GYbEUl5Rw0zHBBlyt2XvCaFPKnG7feUcWcM3cNLUXrnGY
PzX+L1aNpb/nXLvf0kJmHc8TAqF6xFAQiX4IZvKvRGHBpA7QG4D5+mEZboa9xi+nm5Z5BGjQe5nn
4VwIl2JiprHW9gJw5pkochIPox8WAKD2NXepF1wi1yhZEXgyBmbp8ZeC8IfFemN2SuLcpuCvtzI7
rKrgArpSuig4TJ/mbF7R+LI78HAArXDEovnyhNbDNtAjpy2kzJiCet4+nBPHsdVIiN3rcrTW2y15
mV/LgvIs/YmeR+/4t6taM4R3vtnlBwgoNGovh+QUo2x/ljn/QiZjNE1jDHUoiKJaCbNjLbRO/J4E
h16pXo6Obx8yzoGIjZCZ7bwm+1v9ScvkgNdUJN5y0+XMx0JYCJwXgoIwYMBU6998XS+l9QENzjGT
gukqsMEkGZ56xhP4O462v6x03pByGujQQldX/t34FwQLmrZeLNr7Oi1izJp6pVmWpE0cIKnkFP+D
52VglCOw11Ru0tFAtJRo9hCvpYT+R7jobZkeBNWqHyskQAwLmd2Xbgswg/YCz38uOE4/B25qnKKY
tt4pYXqO0Opm9sNuaQTY2ug8P7CFS+t2MR/SWcEv/VgP43wLA3rE5cTTxzxlZDNvY2Ktu9zpgP3L
lYNGJy/Gux/KnswGbCHcpl2CcTD5WGrYGA1IEqEf9Et3chQGmZfKgtDB+ER4309o8H0EIfPvS79o
r/xighOBtPnvdM5RmC7XQCPq7fET8msa/LafZnti9dfKi5Ak2ZBXk5Z0sy8iNE6uZwfd76k2FphD
MGKWwrTXKw6NWw6l8HKT7Bpj6KpCxLaqAaakBACzq+BGkzw/t2BlXKH2myZ5iljjiVTRGqUz3jjr
us4Aw8SoDMWRX+Hw1qRhhk+NWoGY/KF9T662uSdHhMPdBYtq6MlZQ8jVk6XLvP3efQxe205QjH+b
tk0X1w+peew8ww56XpykomGAFR2gj7ZebTKvsNa7FTEGE6CSZtT2e5fcw/SwH/XIzY09EtPDZ8dg
E9JFFBnP5S1kfDSZhCOIrQ/4uRuX8u9GKeMlec/dx554Xje8xLcxBPixuf9S5KL/j5YK2cUv7yPK
RheHIjy3oQ1wxz1axz6bl+GYk658+nwzRs4hrfNmgdbpJcsF5qS4JsuEq3j2H2wwGlKmjVWDi90m
BjVexrYqtyTfMGl+Re6ayXciluzMkpg2EyseV2zIaKBP+zj6BX1IuFp+mtL9O4FWOd0tmxM5kTtH
GWUhLa/rXIaS6miJw5D51gerMkbKRSfrHaeDhgzL9Gxs+gOZ8ucPhESrhx2bUHLNT50TX7+1yiwK
vQASf7Dhu/MbL+ORaS2q8HIjAdLrS42Z//2zkxx+sCrzOzlYkVX+NNHL0fHJbqPYwO91SXxwV9A8
on27UjBa1d1pm4hkjjbyZ31+ApFW9xb1+jrmgbnUMmjn99ht6tt87Ky0T56stfpx98Du7kKXqc4K
EpkPYcFFHxS0tAY8Wm16r9zefARGqieV1otRveJf6waz1K6wtwqQWnOZJasWIpKJ5AsVaNlQYPqB
aTcDrNVcOBWsnwYHYfLz5/mznTBlzxQJkzIS7DgHv/VxfSA7PrKi8/rqPFUBR4AFIValUIdmlevJ
O+BZF5FkzGms7FX6Q0gl2av4dfh05EEWdc9Kic4MjJtNuUED+I0RXcQk2X1N5nY5F6o7NGl7AFCX
DXVJViF6H6qbhpQft0gZmhOQkg0GxQj0o6p+5vqhJ9WA5elNlxf/0r5O4VgTsRuSx78gbAC9BaB4
D9AGK/v+nuqWilBf3GZwMH0hEVxf1Ye0md340HzmPosO5SMIlprmBNp1N/ID8GPp+vzD1SKl94SG
fgUKtk67cm/QCSXU9GuuZJ5WMn5ZgE7zxmacprhm20FG3OM0VCq749ul6gdVPnGdVSAYIlKJq9lc
s8pYnmJyYyBcan7so2TjwhTa4+VmXOivimiUWAZIvUx9wJGIRjMn3iR8blEtNEDpuqge+FeylEeq
eOVT0rEupjXJIp9BQ592w+SbXlfza1jqHM7jyjhJ8BXIaGsXRRPjr347yASyip7DCoHgbOWW/6fa
gpb0lcMBMtYHJsTSZBUwDUf/YiYjkBNJwVZbNEW7Z3BV2eHkE2iH0CP37O91jwjG0LJ43c+stBHa
zzEDKbS6kSDdUwC5wUoR+3m6to11Nnx0yGj5XAJY59ALRNaBxRL7F/gcXw0YYvVcJLEpQN2VNSkC
UaxKx+YwtmVIh6/+QucAZVT1x7dsMNipTYAUdUCrL55zhS/+DMlUbzwAUK6TF+zX4kSvxXTqnjCn
SQxRbSRyif6mVU0BgEwUDu9sceKyGjN0Ak2HtBXy34+xgagiGiB66f+I5ZxdmPtnsKG6LaNv3cfN
sNiVFqMtLBocopE3EqgO5V9/0Lrm2MFG5UCF5I8i8P0xZwfcI++NkcXvp6LhQR4eVKSdQQksyOCU
K+Qm0i0RR2XkVfazgfo2Q+DHcCdu2a7lraB93JYFJKUVWkqX79FQbJxP+6yUoVdMhxkHOZWoiQZq
oW2OK1zB5PY2grRcXYGueACoRLmBou3JjhS8+0sYOZ6DA516e585Dsdt/uiPVm/GSIqKKuLHN4ci
9KhmRErPKmyHqDAv6+rrvy08SS/mrXr1VMjMNoD1SWbkP3cpYGkIK54zQYTTVhPXt/BkP3mQlIZ6
7dl0vV3xynerIamN7w98ItZbhRI+XWxCZGWEJX9u6Q2fKkWpK7FOgeDxbQ+VEya3qX9+drIjRJvV
YVvo2+pFVbG6dTxNRusa+VGB6M13aFK2vA+wNatjDC6C0eu12iYEkMNAQKii2UJE3KLbjaMoTnyi
QX4WY76tEAAS6R5kvV4DncMyAzUr5w+Su+a0ZtwaEpnpMzlMhqjYjBSCzDAk7lOXYP1GPpYmopVv
6Q4+DPTb+YIxxmmpvjwhHPN63b5cwk26+lCxuUf7Ql325+CbMYmlXw+5EZe2tffWffMHLDO5eOa5
naP3k0tJSacQ4NGCR8GmuGxEf8no4Oj4NiUnkl+JniqeeE0iGbWBwVSPhL2izGWfKz4Xbgk6Vq/t
gZwcFAtHbTL33k1aoQqSQpZwmw3qDMyn6tJ+Hf2uzbFQW5AcXaWXdeTyj1ko3dkDgxe/iMXBLf/7
jSDEMhINCi4DdNAkhAXkLRnUOil4OFIwm1hRhjVXHDM4arHFRuWR1GXPPUxHBGMx/ZPFt7s1UTyN
WQH5BngcfRgz/dkIdm+MRtkVlIbKVx98SpOQCPN6UzsUoldsx0Lltu3Fgq7vB2iF1uuljWbgc1dO
03SdBVribcIv5/mq7HzL7KTKdWLgVFj6mg23fegMQ01SPSGbWYWZYfpSXK7hou3dulIz3rCaphm+
mnSotgYqjNmKDp+29pypsRX8YDuJhK/JH5DrFZSouGhbMWWnlHlJLF/KCw/bNOFsGjkXQV8POzCD
2vv5dGLW4268apMy8eBxJFLNuUSn2M1ejmAqiWse7WR8FTEwZgeff4fN5BWAnv2uIsZp1FN2w0Rt
G/O75p93dTT76BfQ7CLY6UINB/JMRv/s1U0dXnBVfgdZ/yEYiGPD4ESyjjSUDhoYacyF3SGfh3kX
rGiwyUH745m1IysMRtauxZvpqg4YdOZSId7yTM43aWCqQyXkllwPBdX1On6swT0BZ1U51oFZpLXZ
AkHyAZpehpUJ66mdUijqR4ScC5KOZ5rSkOXWmoV2AQPzoZhx2/Nbc9+wgXIuLBany4FoI+2AUZWz
gKPMRLYkWcG12wDbZoNI0QmQ9RUzAlmq1giFPPbu5Y1BGCq/32AQjHgedv5arUHNOljCsrxaCp4O
3lK0XqAPQqfEHfjV9Uyeui+YzhLDEdiX4VL+YN12YfT41sVm7jIEenCRqTSDthoOgcbTD4hc4USS
lEb+5HDfOGArg0qzhW+zg1i+R7ettBmxlmhNweKDMWmGbnyjS7cNeSp6TWoSYVO7XODealloD+cl
MjSSxX8+9I8x7zjJDmi2Y+vxoERI9V2ilSazzHOwDbV9OGUTqXC9dJN3s08+4tZg3kRKKI2jZf+O
bg5qL2dessRgpNnkbm6CG0Zx9EW9ctGB6tgZUZ/yaikyFavAKV8doezGRvtxNQM+Bk78iXfwdG6O
uG5olCwz3SgNlcGdFhQSlkCDb/ZtAul/AHUIwEfYNyfCHduJ6t/HaefvyX9WtwVRm4RsV2C4Ou61
JC2iQF3ii83ln3ceQDyLUGCaT2azqwpK2GEwiFpuUw3hwJ5Hz/shHr4nen5/IEYRMSb3LfuUJyfH
XLGp9StAdqaXCJFWJv00z871yGT9hB74IB6KHkyhH23vyX6vHVmxFqksNuOe+zDRYHx/Tx5/Yapj
gptuhO5ijiRCVRFYwGRKF8HZG3X0oJwAWzQorry+V0hVwQ/H9Xz8knAleth5YIWc+XldOtkpGvmi
MDCEOU+iXsHcNQseAbinSWn11wv1gYZuBCoBQI894MNZO65Pr2Ekg2XyopHOFdTFhp9hB9tCkOP9
i2qBIomXis1ROfaRHD7vsQ/0KxXomEjlM3OgtdGS+GyV3xCJ6Mud7PePnDSj3y+621ML96747m2+
kPUV0Lw5fFnultJJkijsL6v2+p0cXOBxzJa6kkqB1+XFJflByOVnX9D1++yDt5wCpKpDeFwiwfYJ
l/fy4McAkE/EQxcLAJ52qyRyJ1aq4E6swPKhIv1cLzzkXQGsvF+nWj2qziJEwWhLNcwJ8cJNruNk
LR4MNHu/6CyVhaDhUeUZXy9d60kys0jqGeUQG5Z2td84WvxvRO2Gg3+jKKADNm/t/mjhbX/AQtlQ
r1PPlNoMcZSKg5JOY5SdPfGyZMeXZDAYJu3MqcNBUy+ZbYydjFv5Q0aYV4vzFuDfDrq9Vft7VArJ
24AVxpYwrZqI3D36Tulgtu8p34Ca10qWF2hpQGJwC3SRB850km90pgR+goMoe4s3kiwoSE+69F+d
7FxkcBNwbXRqcxwdk55TZFTFiuMEnA8kw7DaakEmrGBbFAnA8xEXguarQkHSOQKY3y3fH7ZVfsyU
6uGshpx2H42noYSeBFDwH2HkifIkFgCXSeSrffPLly0/V7VgWWCTVamtrlVm4HUx5yfe1KQKrjnP
i/RNN/wB/FJm9x9oyA2ov0+ANLWP8WubsJYmM2aiEx3Fby4yCLIOQm26hY8efm1WJRqVa5AyegLn
BJJIlgh6NaPZYAXKVs2Z/y8eqpCgmtL5Vh7mIILObD4f7ykz5b5W6mVBJt9aI3zQsnbP7a1gLRZh
UQ6pr1/1G8NJPXbGlgyoaIZ45TfKc5dg54G4rJmw6tk9uSwal6GrwVlmg0+m+D37jKE0qgYuWB5S
kol+9du3UzPTMRJVGWa9mIzODCeowRHyNRMwn8YZ0DHFUFL/BY63b0oIcQy0S9ijWK48cOz1pR5c
vR2/x9YtkNIfvHJKwQ1FvyyLKHel5pHafHXJ3MLpkhTFbN6uBiDNVSFp90eQmqJa6pi6XlJXOB3p
Dsv0lW2TiHkO/vrkIQKH9b8JiYOz8fxHPXsqDSWamku3CwLrp0SfflllQlIp3nlipUsCBLJ2+M7t
RjcKjsUj35S4DSLpKu5mkMnKARDhkw06qBL66UkSou9eU7HNhsx+JD+eIDsHihW0nxZjEwmpRO4i
DvUAddKEBSLm9QI2hYqnK2S/9yKTE3LQIVt8mDxzZ37srLCuSuSwZMObI8Sy3szP2UFI2RFSJdN7
78JTWWpGCQUvi6oAQ52VU2yxdeQvF6YM+uVUOzB9EbrsKaAb3TEZMP6fyw6jJzg4cYEoQfwizM8p
GG9jrD0BUJ/Ne5MfHDGeSjHsaxVjbL0g47pQ5OQfUtLYm7blVgpu6tbSHqc2N7/wuzH2UtxAdaD/
eN8bQ/N+jfHR1vNbnrplZauTGF5Is1x8TFcgBfZJamzh0MkCcwg25UNJjTOOVtMGThD0ymxr+uEw
pUeqRGxKJeG6a5Z64fzU0l5ysAR16YwGU03GjVhozUeGjP3CVJSH1mXkfn6jd8tA7Sol90frHj4u
z+HeqClXUmp0S3OIyuIkIW1HDLpdhjzWBU25lZgmZl/wQR6MDJ3w1aRce8brG+0uJO7ExrGhJLka
zA76yXZSWrcYpEi7E5/D/qFj06mc37Quhv/tETTbhLQeu7N38lt8k1Rm+J3m+eibjY84p1YI9imQ
PiIIwWxxjUoDTORZ17hLOrP5hkrNb6etmq0Z2XrZIeknSh+8BdAxTnFBZ5LGwM6BwH/7kTZEr3lD
3iUjiGv/OIPsUhYQz6Vf7FLynBGJyrYFFRwx7RQU23ifzil46F3W8K7GzAI2ql5M36BplfCe96WN
IqX60Nlyt5Now4EbZvMehg/ngsSNc3A0ps+mPu1epBaNXRyCL3rb88fy1SlVfP+bUkRxH9JElJX8
WktdrJKfk5A0PTDFX3k7MBRuqC49Yl63Ablz+YgRZk/lzGUyc83XAU7al5OKcYW3oOK/oMG5mPK+
2X2Gd8P09zLFxNMgxmlDLqoXJXMcLsXLdZtfn66lAKAfiDLJm+ZDzk70lJF5P2TNytG2UY96kbUy
CLGxj5/xHNm/CvwmDzOH4uXEsbj0pGSPIOqIhyEpuqGq0a3gj0Q1oAbBX4bjp6XpPWa2YyRjftSq
5gWyplzBwo0rYVcot6Kq9zQmL/36q0hFB7Sl90DGKVE0dLZ8AiJrGm4CcWat3TZOTDvkUfj8hi0n
s/jjInJSBfw/s3R/nrd4UWXHa8SeOwQqYwsNv5WsqGItvOaK4QUJzJhQPrhSeFRe06Wt4FhgwL42
ElDNzuLchzcdDsEk66VS/gK1kHhoXGGvCZb+2i+n+zOzzOTNwVqkkWD6xhLJ6Tcp94oumbtwvlu+
ya/5Dkl8GgL49lWejHU6SthC4r9Hr5paaX7//wpQqD+LNE/C7Ynp8mOFQ5Qd5RTIYVvCpphT7zbp
TRm4zdVzwDxye8Cjd6S2gkC+ZstfWPriZjYgB/qy1j4JgEfijvHuTIh1X4+mdPOEwBeJ8fEVb5Xy
bAtQByAkC8gt2bzr9iHUv5SLD6bEWZzZDgX9k7t/AbwAjc9kdZuX8v9+qnslIFGxR0N1VypUDDf1
P8uhmrVb8Gy72v/FVpsObp0sZ1OyYQ==
`protect end_protected
