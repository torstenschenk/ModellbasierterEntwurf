`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j+npTEkrOuoAYyMX9/wRnMYX5goQTEisG66YW+i1AlzpOzLle1lXgu4EgeH5FLw294DViS5wgySE
5m4qv4CG/g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gUZcfjlaOFMdX4kb0TbR60nJXJPsPe1GyqlMGQubcZlG9I4tJ/ZhHd1EMxwWjzpXAI7Q26CbWB5d
M0N6EdylvFtjmg1EUNKbV6Du+MfiD40m8//+pZe9DGyPJfpmuD4+Zj3hF5SrXabgZ6C1Xp1icJbQ
L5r4LZJ7J0joZtYvw4s=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m5BR7gQYyud1p/OTN3ItnmfZf+MrbBm5KEryxpppgQ4iwUC0k6E0EmeGOhQnOMR89C/Uz4vDj5vP
kR/7K+K3yLfHLs+S12FpPBZ3NyuY74QU5rOfBxCPg1sdBKjM7iwVGn/Ecb4QkpmrleGslFvuCXCG
V1QSO28mdm007Vi1l3E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B4L9p7tgqm98VIH/YFg16sVSk71xEJ5QzzMkqAXSOWwulHN1TAbp/Anvm0mHWyNUaf7zrkLBC1E3
DyXIIdN8sGBbSREiq3gWYd0NIbQUfdJZZYvs3uJPPU2+ALQYTUwHJ5s3WX/NzIzGuAAOCxw/hePs
QWaSntCuSjeJws9v8g1EGOV7yq5Osdtd8x2LUU5JN2WFDJuVRSHIv/ompQlok9q1EkqQ7S7sQz+i
a0PnTbVY7uVeCYr+SXmQ0ogUGteEgW6M1VHjoHTsYDuZz4WbwB51Vlt9WJ1soaYWFGDCJlDxH59G
F3endzqkQitpYnFk4ShPiMODHQv12VpfJYbHRg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hwYr4TS/aBHf+wunP3cLIe0CYKkGOTJ5Jld+NMc8xGN3F8TLtDkRxbVMutpF4XfSBJhLcHSU4iQL
iFpWN0M+yLVcuPEGASE+OmR037wzVwI4JbEmc01MfjDNWHEY5ss30fwhsdWHpqgsyV3rfWe51mO/
8TIpFsSC0FG+zpoqHyDwegAf/Lmf4zKpgFLLo+3OtJAc3YmnzL6aNZ5o46AbwYzVu/XN7Ak3E8lI
/q6Y4ANFXbA7iDszKKZ71HKX3ByW0rvpUTg5gri77obs5l7sIyfp4En11ig6Opv8IgX7A29qw9SP
SM2VCK7D7eVxqxbxDEPCIbcxsa+cEizeFb3ajA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fLcMKoU95J0rpQurE7HrpDJ+JK9crolX2l3JMVmKcpL0dY4KtTMeR9YZVRrUm6v6lYXi1gKv9VGR
rJoz1MY0q0spfAy5jHcnDVY24WoZRTIRmr1rwKTVmYW99Be9KcesnhPZ4WuQur2Sv45IkqlI47hK
jnLtqX84PKzW0ap4HnvRWci/sP2vA5n5UU1zybiOUtlCnJBxpHY65IfbMy3yrF80TfTrR26jC/co
4alM2f8ErqkNMnUr0tMjzecZ/pjdWFH5wg5jNvR9C2o/vcUC0kr2fnXRwsQXgxT9vAbEitKz9+8m
p1Mwc+il16beY7eojdApx4J9ojOFXIxI8G/fSg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 65376)
`protect data_block
VNYkwl0rEcKPMuF52+DMTiwkVE0PXKjdmKTZm9hzBJ0M61xQHprx2DyMkMRez7fXqwm0u7OwJmom
NOYL9CVwl3VoX+biZLOHa0mNCMD1XxkrGnkpWsrdZ2cCTSIMPWr1x4yW68NmqBJ0UP9woQJyqHkm
Yd84zOcj+z3yOD0ZLfN+JCcItkzxjmlNoeP2vZUMPB5LTL1Ca03cysncGUqCGVysI8TJCkzlSP/B
9JSoo3kY6JiYEtpbuT7+LebhYU05qHBQHLoVWR7IQCZbU3/iGQZ2sOdQ9V27L+1xUQmhFTh6xdGQ
w5Yu2hasqBfxusAMuGXR6PP+EWS/T8Olv8aaVFPwhKN3tKIPYybzdOZIKfRul92efHBqEzN2GAS8
ZcPAxf9m+m2Mba4uGvt5LEWu6dRg0vSBRIdBrLc4DeJN7CdSC2rY0BdvIUmy7ZqRQdfEWLMZuncW
V0IyqPfQBW98VlKTK4LLS4gdXZxf+roBLcQYD7RMRhV0VoazE7ET94NsnLB6jYsLbOx1Elgh89ID
yy7snqxqgLzd3c5QJDiyhN5di1s9QJlv9Wz3MIyNtrQZy2iX27eqVJ489FkSaMIT69UBMyhk1CiG
8JqIGRVL3uQj7yjS5AW7gK1pSXMNjcvr4Pjq3+gH07FDmsQ9jHY+MLNuun/4yjejy2PeMdA8cu+X
0YCGBQd7jeXcQW4jvqgLJmFLPKsA2/r7uKfUPrbo85V49cY2xyxjQd8SeEs56RSmNZ+C8qfsLuZD
3gnk0Nw8HM0DumlSuP1vSeDTA66++eeyNmDkCHVSKOGfEm18RMtmwn0a9ja410WMSF/ZKQKJ4kzv
hT67f6xjCTfEqiInZLeiXTq82+HQhwhWnta2qNWf3Uu62goMQ+j07cOsOcDcnN/Dn9wvLbFezW2A
K/JgWZuLZ8S47TCC2Ba0N6DeLJ37YW/lmsZy6wvuvi75YrZFvtFUT9wQWr0itJ5ZwtL+YeswyKGP
TKMJ7y/z5TTOXW1sUN1r2JSUosv2jy3bJWSpU2KV7+k6GPYjd3Kf+5yGNLZFO1+9ayR1QsXNSKyk
WYmE9YnRBQnjznCKCD5zF8E4pTudCs5X0g0siInYato17+AAUM1X8Ydwy/jptZkcGhDv3kDuhPVl
A4EwIXuu3rHVFToNq3muOchI37/7bZI92n5LnWIAEmxtkA3BNgbTde8R5s/g95V4rt+ykvYTyHHM
xf8/yjMZpsCFemKxlRR4jB1SSIh8n31GHslRWL1qlpmDGTrAaqfZ5fzZPKSIWwTHO0juJFtVjwEi
IyE7fNf729xw6nSvI1lldyRMqcrKQ09iIErR40nmzJakJxaqfmzqEVxUKTfyQdAn43ijTycjyD+e
zi0JBTTVvAfwuPBMjb88F73L+jPfeWU3IK0r6o0CKFdeNFJv9Avq3E2koMrxwowphBqGRUIZuagB
yhmBJ1B4qjIFV/fGhHDfV9Uvk6PywkTWkJkZGPIsQ2Aviaq40TJYnfvZQ6k/iaZBu5GX6p0PI6OJ
cqiDXlxfVdHqPtggF7kQgcBjCk1+Ak88L65uiiAJ6aJXq89IY74bApE2Eoq0SieRqGbmHIbJoida
nWRkxJ2wme3CWqe2z562gYYtfKpSEXWJvFqfQb0CL9AxyZ7++Wm2TMajoVlZR34xOH2pROAz37Nx
YSLbX0irCnUDX+uiYsUsyjPSHxcB2t8pscw2sowzUCHpKNI/9C8tR9m1q3iKWh/2hbAFjttb2n+H
YscvcjS8q/nWw2yfH55gtluy+0cPrHwSMnrPwSFLZs3Wz2FscgZP+lt+tfFibS8xXPNl+SFqAAEm
/zPqy86nbqc8b+/Yzt5BiBioOZ0A+4bKxvEfFv4WXWl3wm3qFqUm2eh/5vvsVpS0MK5MxIp59bLf
DvPtdWhyhWUFOv69uIZLTPG+EQu0gGUugBVWudnek0hStm7hg3cSx/GETrButiR6Rucd75FQ0QBT
Nu3aHcaseo7FJXsoMjVwduA0pijhGnBLTqJE3vbp0Hl3+3/sglJsmVRX/fxwSjiD3A1k02V135jq
70YvFEFthQV3OMjdIRo2wa05P/0P+PsZMaomFw8vkCEgBGdm88dCMZi/VHw9QcXU3CD2zqDd/KxL
yGMr8ge6zWzWV7xsud4Rj5mu+si/DwTAmimZH9mJC6GUA2R7NRGx8gEW5LZA1X3WVec5JGoB7moV
w4W9yulVtBHBqb9e44jaiCiWSb/DmNxgNaFMnXgazzadj4cePo6Pa801aWroR70wurNOtyu/FZid
t1CVX0mdMa1nH96rbUSh3V+zERSTdTdTw5y4qQTrjfnDUAU2eSUHscBG9/okw7xnyiGqXX0GMzbU
ANjJRemQhjgGBXJXQDD+aRaOuY9LuyJYOqEvluDvhdsweoZP/W2SAjL/z2t/Xerj9xN6zNVbWZ1H
UoxtX0Znt5aCFykKT4pcTeOfPiNLRXsc1yg/dXz2TE2MAfo/dOUooK4AY4w/ZFUf0o786hteO+MC
VEdODRC91Czq+Mnnb64dS+g3NiAST7ulP+dO6wcGBlXZDX824G8VEvkLeg/f6kq9g/RkurdZNCzS
0/RlpH6tsEdYjzEISxFwvwwlOPZ2t3W8hOzO3GmJN9oa+x65yT289qrH9wYHxani0tPPfudFEFLX
++UMzfe4BwpfojmO2p1NATVmItkkxn15EQ15nrCbn4mMUj3WoNe/Zi6dD9OzPnPPzhezA4aQpPXy
pwuQgXugMKOcSybDltX0SsKNk8ix4aFRbI+BdlAw2lF0vMUVs6SEDM44j8nQm6Xa4sYcBsEh9UGu
yLIhN4qFYjT8iS6C71VCnA3Eq6NzmflEPa98jODHW4WW2Y4hn6mAEn47HXt7WgGTSdOFE9ynoIOA
E6J+dGiNXVf46clFr/clzUSQEyk5MBpTxug3HfN3tw8ikNkbBbZkeiRnuBwVLHW9OaO2kz5Cb3bH
crbBdP6tbEL6EymBDJDmuCyD5lwANYBBfnJxqGQhR0qWcekZXODfDiCsLHmIQAuCE9B7RTMxYOgV
0ULDnr89X5RoNPaaQs6ebijs1TjJhDOI1lTCZlnP7hmTNrJQX1j5cfR3OX+GA/wCgqOIFd4c66Cj
9zBYdDRY94lpb94ZJgTGPCT8HSILIbP/7LSAdt+ouuApuEjgucV3XiGuC/0ebfQ9t53qqiGaCA43
i+ow0YTmw9J1pwRdKqpSUD4xUBnr/T5evGDAxle1io1DPPoPxdE1ySJ/CVFDrHzOPhtP3/rD/fHJ
SvXl8syflOdovnoszE2S4npESf14kMJ4wMR3wd1XwHK7mQTRLmyAexbb9g1VJ44KnAqiubX0v8Sd
ZXc+1NGkBNMq6k89djruXERWGDbRhxE2Ct/X62e0lddaJiZlgw+HuqmXQsH9VwEpg6TkFIQf4Ver
XQ7cddbJ3I8cybyTuGw/shEmV7iT01UfdxvFxIoEFAjzEwNPPaYJmvooxmVWDOqOJJXXJgF65t+m
ijmlgayz7cNfIo/3xZFyNgULeJ4wNwd6iCH7pKeRAjnluX5N7qFs+frrqaxe8SWRbe8InIo/Zk6j
y+m7GpwY5crl5LsTCg9EkNnthxZFWQETjFu6P8NFmaehnXkuC+kcW6FOhatCmZY5484y/QvGvL1S
WvmvjeU9iJQwaCYiwcm+MerP61N7CZD30BwjNaqkjbKEfo70XxRFHUSdc903u98oa/yetLc+mfWw
Wtl8WqztDVbaN9sz4ok8FOn/kasNNvRgnsPZGwVn5hGoSUTjfjCqC623EPuukzvvcHIZ3RCtOCSk
/hYlEWz95e8ssrd7/DOdu8c+yn8V0kaz47xzkjACx6MZ2R81JIOnvZI3qrLJkkch4eUPjdcl0IGi
5A4/fkt2n/WMr4hEtWbTsPsGFZOh7TfQFHiWrzzzXaHcrj/HvtwzgWA146SmGjDidF1MRktLYWmP
3OtEiHK0pyDvDJbvvuT/SLoG2vvWg9RpyIpCV+uluseAVwyaEosvAJsDDx4vzSIE9DpJjUCkCeJo
k2lhZ05DqjlaIhcbCt8j6zRPkAJ0CzRGPH96eWfWePE9v1v5aJR3hr/UYTasSOLuE7fBtXZBwOmx
WsxWmz31fqqlmkk95wBKG7fkH6cZg6Awh4cxUW+Uh3nwJR4ZJuXKiQlJfhGvYV3XY3xMDDKVKdHB
H4VJEHfpbbUV0hz2eh+rjTuxxvyaLMwl1o4bZUy2hc5IrVQ/t9FeJn5gyT+elvNW3Chre/Ejp+sS
QQwYJBk/lnXDHZEP6DMkrq8wEKjbaUkHMOspoVEq0G+rjOTgevtLv1U3ZcDWwKlDNnkvgkYxhq91
eAZn0cyvKs+nsAWw3e+aRcczWeX8fuDdXgksQev5MUDDl2SlqYCjc+Vb+pHAsdh7AJG0vwqtmlNg
XMZntkiAKfVDS/nNoq4cWkJ6GoVhPtfMDLI5ZYs3KwOBKucr4ulSA2+ES4D3OqE8BJ5R3xLfkBND
DL72ltJkLyUmecsi/NuDKn4sNAJEMTaEMgu73M6XAyd7qaG/hqcggxNoLZHy5flmbqYNqlRwoIm/
njikayxIoKw1XQBChhBGXPVXX/wbVBNBl8YlMfbRXMPpjXoieZH4CfDcv6bfLmnM8RzLMe1uXzj/
HZ8DjSQpRN6ezsEKTmbmRCYqZHtPmXydwgSL2tL1eeOkVQuxAA8/Y8shZwu79wzdN15GQOqe2xUI
9F6GGyIOn8ggr8WGAXDLhtJiot9toA7VXGN7sXZjaUALa/YcA+e6zB4BfqRuiou0LBCR5XzjiSEX
8sqL9aaMiAssCgJ0GbP8YpRgamVU0Qb1G0m+W8PAnt7s+7UyRzTXTwhgwfYB+pxokhVEueTOUqm9
7Azx/J5do35dBAyGG5J1AnzpmHp7ZpoXz/jBXgygT8TcCteF0o7opqchghiXDZKZrTVnBHWI3Ka0
oTHIYMJqOtrzXDU+vZ8Ur4jmq/sesVp6he54m9IA1W7fppoE/JW3K62A7dt7Qe9NggCnkroGKmIl
nKJEgiHYIiAGTjh5zoyAt3m8j8u1P8t3LUiB6QwcZvOCvC/6a9lpxya6XdwRK6q0Z6KEv1g7eq4n
qZgUSG6OqC5Wr79nU2dSwon2ABtuzDsdZ9xH0cnu0rlMB2z495DnGRlEYWgj4Uogihj+8WWM88/U
32/N/Y9VMTs+a1MzeaGMVtEPgzegAPRSSFVr6JOibGvligAB9+7Tc00UQYibXXghaqOYyoJzOyu4
qT0Fsugf8bkOMH8ATt/dRZutxHWlycPRoGdQvKl31mKRkvrjP6dqi7ikqwR7krHoLIUZe6hzW0rC
R242Mc9NF3vqC1o5m2MvbuSVzIuVFtIDEjyegLGBjXdCejggHvLazes+NPMKhS1P4Xkr5zFDla2F
2hgyrZJtfJajwQliqXUsI6onHUnyCg+uGwckqP+NcucX+l85y2s5jfCPSyws9MCyRykSoecM5UBq
vVQX3Apm05t9fIUV5t0bDg/0AkzrBLxw+sZ2h32zKwjirYRq4Z4VMJxlrnKH5OeL4I6ZB7WTKNKX
CaZf54vgrqd9rW2wlUhDzlbmW58D91JaY0FLkFOF73DaVxjUB8XheoUSH2EGcBbReH7Vjfon8UQn
BcNDCGJs+0BSqsuXSI6WhOZk1RShCWRlpl35UgGgIuUH2WMKDi9LqgvDJxnnos3gClvTI6gD4nWd
rTSeOGR5u6fiw0OG2M1POT3zwyC4XDenMSa4O9mbLggSgEgtDLLhXFmsGesJEEARZ/fFLaK7FzWP
bbSMuNgEEY/rKJ/bU/PW7Oc7EyDWzHZJF5T1w/2UjJusX1coJILF0pjKnTAnw0AVZX2K3a4NtfZY
SFLHyGG6DklTeT2ScvjSJPCUPBDfZBm/pnDHq6ZpdYeWb8BgN8qj2WmN4W5e+16X2m52328IhC/P
RPXUldS6rqyfdpQh/zHa8rG487CoXZLUpCxCVAMfWraevGXcMnGjgIL8HkMul/9YuH/YjjeIPrTS
sKyqzn6Cn02AhRXHn2kbV9OJ+7GAywPzOBrlo1Jlx3ovq9jpWumOHvafrSfni/b4o+F7/1KGhHRj
rK+HJ7likGtb4G4CJmqVpFJMGw9o0B8NWKV5FNgwDncwjkcge7C7QHTNJvXuBiY00R5e6z14g+xV
WTIqcoSqyYBRkk/gN7kSiOf7q30q3SZvMc3SM4u+uFUip/8n9KIgJXU1bVycWOd1uCKvnsWU5yrt
CWqzjkvR6oddBQGN106YiwAqmBoiJMmg+B8oNJi7hmLXTPn3j84PArzbA369xl9EaHLhTDTuaYhK
WHiWxUjk2pXm6Tk0XmqPug0HEGzSA+0USMU1d9Y6EpFe6eQCeQCWglqz9JOm9pVt+42uv8sWtpcq
qGR/gFOLbUhEwiayUlM9+rocbSw9x8JUJeAjAXDSOmWwdAyUSF29A0vm6H0JA3ddG6EZHkhgotVq
0BcgHhq39j0tcNK4AvHIJcY0dlO1ST2tI10IedczA/CIGUdchACjyVnK0C97NqAi4H66BbSke+7Z
DzG0Q7rd9wl+H3DdYvxomnhnq1bqGCzdM18d871hikfovGm0XJul/S6fv7yfjhz8CDDQV640C9Ad
/R/XAfCGms1WL/a6JOVkbww31psqAdk7ZkoCFEG1x/CKrbJZDSG+Lq1sQ3dVK1glf0gqCVc8wCtu
ZrkhN1EJ6f+UzAd97PMjM1DADoKOqIOLuiodxMJI/RMDkeq9DYgiNpcUasYU5dF1E7q0OWqdXEv7
jKC8adDx5ESo6Mio13pue1eu9U38BNucAqJOszzkL2ihiNjgSlZ+cU7gcU9nvX4i8/AZCxQvl8iw
Bd95g28N6zo/WgvIFUngVMEwsXHYjqNox10faPF1/BJirSZ/quJMbD770HqshaL5UHfF9hcZWGU/
wahLrVk2NMBfxNsRMigtcO5AVr4yJ+vt29yvab8NAdLIyUHTMVqQ1iRr/U7Q3JCGCQiBWFKmN3tk
ICeGpphX2P5ydaCe/KZd7t2rZKEXa1WY36hBW2BApPUx+Q3FfCaqHCZt60l+heAI04+WvEb3fWrC
A2qUk1XxjKyN2sNfpaxVLH16R/1vH15RVRFTr7UifQAAykayjVqoi7RtEYOB5oLYwuRr+mj7136N
6DQwdObTfp+Sukd0G4vVYaMsmYg9U50i07VK2esCOKjOR3W1JYe/VIVtYC8VsnGbpS6fkMBsKqOG
ixtwaNdHnYDC1rq4p4sPvXMFYBLBkjJghL8jm8OAwhSOoQeNiEPZstrXm5/zbNQxOm934eS75liG
IogDY6/QuDXpfQmjaGOa1q5ztBqYifI7TDBt0ZwWtEv1kg6ZZU2jZiYhtyzBxMVFgG2JTHN3p+6V
6mV3M8uYpYJgFrq4iHuC2Gpb5N6a/9osvLMs2UfHudOIXHznFhDb8w+QWR8J5h0H2McTEtItFpJ3
/2rt6g/ld6hQ2I0zwBc9vXF2PRR0sbmTYc2x/tZiXkl4OQP1gzwoLNx68neodd6YLiWDE05jyBzJ
SptLpYbSl/HPUkA1fRiwl8h0MLmwpwiq07ycZrD+3UuCQ7GM+quPhGFflLleEnUgNYaIUxZTl+OI
KbQuQbk/e9Z4jDw3nMdkD24Pk4ta5qu0jpLG1RCDhMTB0EwW2RnGmcOPsb9gmxL5apscAGoIhmEs
oHa2K5q2rgC2QUhkB3OalTcq+J9sJvMMROLvoq5ldAqL0BTJw+GfIiVEGCshOAb2inEkyHc4+9Zf
sdNZYRi1nC13JuIQZs3lRP7KGQ9K+utUeZwMYJYTUu1z8lAuQdBpR7gxKIpPwUbhJBSZzmIPdnJg
6OcnV1/xLRkZ0rEeVrpQ1a1ggcepUfL8AjyID6eBSrJWMgYwh7FjFru58xklp77NlwZQquIZ+Uk8
y0eYKdNgfX50HXpF8GRS+cAAh5L9BTLxLilTFxuqywfegd1hQe5BJB9xbvkQIi2pnyqGj15Y2egi
ZMs9uRwC+iV9shiEwpzoGRbAVJ8uu6tAaQVg+iZBwNyALBugRmiIs1mYSEb7G5G/4MR+w6B0tSlp
y5DHuFEI6KSeTaK7R99Hk+9nkr4FHyJ40I6Z9Fl7BQ3+fg1rE+STtL5J6q5O5VEKog1xYzAsrXkp
xxqDZ8P1PTnwBa6g33SoUqlz5s/gOVZOMcQulgP7tp93rWg36sll6U1c+Wm7+r0JOSSzig1NPntX
GIWJf/r9rXE5aFhMRzsFhBRd4fV7mWD57vSOCe7zk7jnDqihR+t9CIgetqlWHt8f/5j7L1m1rzBd
dGIFM4LVYawD1yWTM+gLbaF4ySGbzQJbIGqjQ9awZxkDeB+XpYDkL1cCapiXpY89PjmWZ3DhNLeo
k2wg8ZbJcr2kaU17XzDZkbJGKmnNi1WarQ6CAp/2uM66VEfTM1wmIbb6SJE9+wdBVmHAJiI54RWN
Gls0DqjHPVAHK3N8WDzsbtc+IVPC0zjgvt4sPUM0y2u/HTgcU+HAsYqGQlt5cTZiRlzjKTbO/P50
LJfkYsOdtXIAWYFD5G0FjEPLLKqJV4FK0gTBI7n9kXyZVVjxceBG3jUx7K4kcJpoThbJzDsm92Fy
JQh2mnnsdRLZvZ4xowxQt+CZtFqCk78yYRA2eR6qUz+AAoSy5s1BicKicifS7CWV+iUiLIsPn2TI
gVHmvsjDnvm67WDJBc0lyI1dCWjJPHEvK06n0OLNIGcsb10RmCgn3CUyGSfdZxV2YAc0d5BZ1ZFV
CgE6000V3WHoBW/hGoaSde0kbkoxi1pAlCBBJgQfGLiqHCM1BsTd13v7d8YEhoFzXrNQlpUKLluR
msRMck9DiPieEyR0ZiOjARvYEHOLA/qZwUSN7bZaayqNrRKCGH9OOMu5FeM3CGV8LfzMBHHFnPPw
EA18X6rUGbRth9Li2zEKfczh0+ZoREi+gHKSNoRMVGlSfn5WRdpqkJ1n6X3W/Ejttm+4ekUVDwGX
rQ6HUB8eRq1N81hh912oJLygIFUb2dN/AG5XvKCvxL5rarH+4UFjyaU4rnnAsF0QQ8S+M7TNgjL3
0QdeQOJYhR+eur+g60tSAPhGjbFvTmF6KsUSlIkaxT1Y3VI15CrAgTHlJa/LRzatd/MbxcaqymkA
MhPO+aL4Notkiy6ueARv/LbSCRWdIPNl+g1xaJyOoLG4k3yuZwTG6vO3svpcy0Nk6ltMz59uyCdS
7D68Bw+9smsxks9S3UQiZku6M/toF//JnOADObsHYyHcedA+apxH1pfBFlNvKK9qEma9C5LVvUZm
Pm7GRCRYA56pk745FaZJX7s3Qqm7lkugFdlwfYchzC6s+nH3acFiJG4N+VOrcu3OSGEezXG3cmiM
hzwmNe0Lzj6pf3xGSTCy5pFhoNbxEEt/xIb6ziLqR5xYbqnvYkqYdZekvda6A+XeVaHUedXC7hvJ
SmgnufZvUVr4l8EnU/kasQ+7L5AdVypR+HSyXZUSUTZMAxKUm2yIrgLKwMQlK8uI//+wTCxwQqe1
FtTjoULxgUriLJrBq1niPbjPsrgMldCG64CYsceTzzCqef5jN93H8dPQOQOBHYPnOepMekuwr8sk
9ObkLr+ha/od34ddn5r3Kk5aSq+qOVXQwI0tqfa8QFDb1NtaRZz/XT2CSp0O2MdSkk8L3iwH3QCg
vopVqI17Wz3FYq/YhZV0QZfE2JkB/L53YOL5mmJjl14Hwo1Rme7tBS1Irg3gQamhSPbR9y0HN6M8
99OsQv0avlMkblz4b9it+6gzI5vQJMWpVVpOF9y2K6zcFl5udAN1yK27Z29mdwnjBqPMCkwBK9TT
s7/fg2m8WRfN61beYD1KsZhJa9Do+tM41NxTi+6OOmm9n71iDxqo5vf73rCAYJJQb9kmbRi/Bx6K
MOfUXZOd6H8qwBERKEvdWUZy8jgjNz6iPwFzfWMX8LGUfJyW4jr899XRviGmWHAEM6jL76IxiX0d
ZEGfuzsi8snvhYqninjVBwxtsiElGCmLmo6VWWild+NyrN6z7MnVeS+OhsNRbQMWR3hCNbjPS5IF
b4eBQ7yv/KM0mDIDwdzE1LowMuVPXB/63b1gBGNRlVJh5JZ2aS2rSOR5KJO+N/uVhEkDZnD7TnU+
SmvN4JejtQV5WEncua+0lZ2Lw+X1ohkpsjA8owmaskAsddCZwWKOIQigz91OdM/WjxUH6kCLpceH
VbEIqBKbt22WKfrAbt4p3zEPsk9ig1wpn+mY2X1NaSYEnmsgWiClEl7npQwDXRkyp+Nfd5nexRvJ
IvTQVeAiiwr7OWccHMa75vNYMiKv3XuoeW7nxK/yj+Ov+nTDdgs+MmzPAjdjqW8nmpNK7bax2gBw
o7ySUnhEjNTemlKMdUv4qIMAP0c0C0qwzcKmVU2bvYaj2ArCt7eyRuU0+fahmNQPgJXl0E+nS7rU
8RZi+rMorIq8VZuia6K0sVER6z3bfHaR+273fjab+L/XcWJrLU7meP9UROrMI9jSKyg7wxcgWfYO
xcdUGnC4HikGHfaqO12kMBM1xPrF/y4mdj3BB/kbcr/2cFe/x3Zoalf2pAVjJi1UJwZ9xDSHn7pD
n42BQh3eMNSGRmgNrUR67BhCRRBPX64p4YSnR9CmBEum0zmmy+QrThIafQNofd5amE/jAVb16XNB
glWbtGbs8aBPvjF0MW54iQE4r3B31SCU7BMafWeSuL6YW+L2zHzuYa68zDFeczdpGzUZXeE2NaAs
Ok6Orqr9eDou3pO6WBgBYNNzX7CvD2tJVTjCRYM4R3chNyN3c9IcEFKeq7zEHyb0EltbqW6NB9TA
ixYTvEuCSIMflXDX2r+ThvAhzvGma5Q3yQn6ww1bykAdt9g0MOf2msalv6NoUrb8T6QFb4qsgvmk
maHEv3pLX2fLltZW+lsri9AuF3xo0Lhq7XGcAabMyiT4Ba8Nir1JUni0rzsA4xTT0DIvFmLf3Iaz
r9in0pwLbHUfSnWZxJXnKxlGpomMK6+z7gvZNy5S5ata0jopue4WXs82OjXimX/FaPwa1Vn0tUS0
FpYl/yrFtFtrV6KmB4tKIZRfe89lAe5EagVVkdMraX4xuOn9A0HBsOeqiHaxLbrD/S5/2+2RLkYQ
tUFhJ04qRugCQmLhl1LJftgRGmCi/yuNDAEUcBtF/Bf7KTZ9R1lTEOY+VAEpIm3jHE8UPn4EywpO
sj8esj2mhkdAZp3bYeE7HvFXk1/vh8wdAQcDA0BT52G2VmKNXn80w1hn5qAECjbW25LZqzVK0ZKp
o5YGu+LO4ge/bcdpcfbG3+H73iJ9bBQP6q9kOY4TB6ws8St6mLUEAo5ekg0sCCKHvr/ePfyugacW
x8nJOxFmR5sX5GNttF4Z/u3WWuA1ERmz15VQ3tPWwqUGZD/Pp2iANs9JefhNn3DKWxX5+vs0iPFD
imXNv7iNNwnHlYhP94kKn4wee4v9QrM9MWOtPF4p2WX0ksd30nIobQu0ncF3c/E30dRnb8YBar/W
BsMxwn9SfAI3JNzHVkppnz6bSAPNRtqFmonyVmu3d9JeYRGcv7T6Pq0blDQXGMqbhowWMtqd9yEb
wp1CBuxHsd2DEvQ3Rlv3rT8bBdkobikTaK0jS3wBozFgR+U32eJhPq41TtcEoAX0JZoyrhLPtJl0
I/Sdv+f/MpxegB9EchruiTO6P6kzlB+kDs44SeKlVlgSGC8gYMWi47lUSiGHv+ScKDTNSjATYcEx
n2Fd8dJGC31oliQv89No9i5hdibHKS9oWYEjiRfZxNZPNMmplFuFMny9zh4u7MayehMtlVD7qgoK
RjBBVbumGGmadUkPu/czWAIgrepk1leDpp437NepYX9ICEesa5K0/lQ/XIQ4f3t2/IJnh7OcSeeu
15iborrlT3+xbssfj3a3XTkpT6tG3vLblDlv8KhReEQ/R22xweN4LBFHo5DTvWyX7O7LTDeYkv1A
k/piIdFMcAGD95hGZTa9D6hZ3FUk/zHydkfEOncnwP/l4yhLGrnV9CaWSdMm/dbgOD0cdtoc5P2h
w0yGkLqvUB6HiiMiUoXaOCFI7HY15sUIZ69tW/KNflLeqZdYERxgjCd3c59u8N4vXdCi2UBEe1wS
aNeocqdVSHdaPNYInR7K8WBHowhY0CAgYPHmJ+cqvj4jcKObRCl5ZqbBktQWL5ukoceO6WDnMoLL
KeyqIdc9cyCxmHgXm64wDOlpyZau1xlodXagDd2R/daffoD+zx9v/Bq7Ud2aSLTAXT5poFPlmq1w
341nLyAd56F4jjIlUl3CRIE5VB3/D8HlXtkSbShOJzI+gPI7+B5LakMihVClZZgpO3WEPrGLbgC0
dKSomJPno+EyIMUzFxWzbA+GHoSLGCEom2nicP9MjR3H83KXALNTIlzvGnas9KzuhGSj8C0WWx2Q
wn6nGTGXUV1ZarOqcZsmzOE+DXjYbykJa8O835BflP9H3vv9vBUGKNxpX7tWTAUoGnH6bx9/KuBZ
NfIB2mZ9hy/+Xdc+NE3ZDWXIj+uXLbpF3Ou/FLJ/elsVHYsCDM9X4Vm9gWqqtBVWpPDim32T4tWC
5oshprJ3uVO6dIDcYo1PUaDjDIWPcWRAVHiH8Acca20yG+WmcT9liPb7x3D7f5Ee1runrradwElH
Y28FMtzkFQHWZDJRIgX2OM+6vTzj2uHZQ0YArybNkvTCdVIHvnKiJ/Tw+0ORmw59MxiecVt5mjx/
p+trqmAXsT6Wjx9I4zNr6rXzRfT2QF6hqnc+LPV8v4sFz9Svu/38Y783EG3m4ufsnqoVdX6yHVtQ
5Zb8houDwxozpaH29mworjiAuOUe06+dq+zYC1ktxpfR/UufXHdRbplS+aipGXaI4LuHUYFSsMf6
K46rIKY9YaE4lSr/E2xvOnTxerLYxr0jMwst+1ofi4Fz0S6lWLTfJa5xVEp/a0GQm76eGkPgE5y+
EIMMKdOQ1zCUXQJJ/+9vYTGCsLaed8ft46tn0WVec1qeP87lAU+wpG99DhgXReCoJlKjtpNbjbi4
u4BJ+0NGph+H3lodR0u2nwbP6grXbyFxqP0MQZQdRlWnQRRQn8dfDuqPmczSFJp1yjX0WnVbsAP1
yOmwDyx/ZQUUPtsYK9HYC689VXE9vbnUadT0yBEfFxePRqFKBkyJb8bEOTPw5xSc56srOcg+Q4sT
GjpuX9gtYG4lh2KsJRPXj/2ekVyLAXmxukzwyxNvtqdyLhavVdv2Bi6lpC2o28vfVB3pkphzu5JF
m3rr28jL9pkB0STKlQsP62IGdTmMDvQ5BVl7Dnbt9Ags3jbXLrpM9fdv0Q4gBMlQ7uMwNGDG2MfC
B2oqWMV0UPsIg5mISIuTlAvY7Lhi8YtT7lwY5EkimaK4qski2bSb6ksQ3ytabIWyu4CsaLjRjdco
IPrwwmcZeZKi6hl24HseNNILBNOR5eS7j330oDBne1DJ1e3vaBns+CVo/cKS0CrY1aDJKdY+B6aC
8/rV9Aq9QGcoMpwCsVsGUanCCxGf/zrOsPfafEo03ZQhr7gA0nfDacL1pplJMg1aE3soSQJxVVkf
in/zweIpiWyMi1TpvEBeocrsgi6Us6OX4JaxMs3ncxez5oj7BFW9xFCeK17sShuDlxk2MoGiRcuP
o4Ec41EOVGXZZE9Kbq2tHlp169YZ6WMDe/OGby+5ORun++hsOFOV3JUH3AFgb4jghGGwyPS29q41
SFkzK1QfN04cbAuzrrOhdH+EcQZiRBqdDQW0AlR0EgnQbmEQwJx11AilENEwgGn8HY1yBpvJhjq8
wu93KeUCaFoAQ2XUQGYJ2eIDZ5ufs+1CA+1bW3U1XuBknnHLl7K+x53vPCMkM+HZPYf22UQONKX6
gclM0TMkANBkYZr+iK8Yvbw9Nr6DFOjLau+YyAP+GDVh5ZNmrmt3ra015umwwCAsA20GRCf/O6O9
zmJkaT8qX5uxEMDNaUFVuSK/svbaPHGTK/lOacdq2kR5uytp0JX5ioHkWjSci83oROLhAkHwNxuk
IL63bfepa3ORt1Oze2RFP0z10GZAE+Yb3b8SL07HRk08FH0HYzc8x3QSBtnW4iKW4PobUgfZBcnV
qDIo90ZFrglNQK6WttXOGnLdqNoorwBs6mdigRWmb9xtygb4rEUwWkzDPfRTs/I3GdBXm/iodVIu
c421oDQtRfjKmrZ8vBiHnNKWb8C5gep7xf0y7W8z+DlM/2a8sxUQEXdDEh7C8TOUJSt6zzOGIe4o
nCLY3K5fb8M5zlUus+tZMabCmlq3+NOS1C02yW9SAxckCmyOTc2Oysed4Whu4gKhhxOcodYuvcGP
41JVKJY7h4Yvi3UDszJIrCDcCRYxV4DebXUGkkL7hfX0MXUaXNTJRmZRb++m1+YinMlw9R/HTMJl
6Vvs8jQNBnWQ8bIHm9DvoHKrf/oHHwaYjfE+2vNU+ivj8T7OWQ1XxTWfa9MiVZEHi5ycf+mEDwAS
8AG6tiPi7O3m5e5MntqLd/V8zxjDtjI3prqNrg4rcaWLiYzg5CVUA+YKlv94uSFOeKalBSy2Vu4h
PJZl0E+NkNHo9R9YydyMLpX4h7JRPn1FQcBBw3yyRZVL5dFW86+9sExvvep/Uo/NuVso2gOSdoB7
yLb+UOZbH5YAPIz7tK8dqYsQZ9yNnvAzagRKHn0Vw85ne6H+tL4FLOcb5TVLhZoXVf4qjfxrP2Gi
88n7s1KrxAhAAPspZDXERXjgydT5Se1mubjbR4Nq71MBdIoSr1cKbGctJj9ON836Z+svNyWKw/hx
8eqrEzf8tUg0/9puluESQZ0aAT0MX8zX8tY92Xi/irhdqlqk69ku4s0SU++CuBKIJhK6vRRWyZlD
L4zQx2y7p3V5kaQrHR6gJlg+cVWvLsQn0lmr5tDS4QcugjX7K3CX0aZZwpaWyzBrk20aagxrY/6z
enteS3TCJ4AaDhSeGTxpzAPFMDhMqE0Lse1okq3TepWcnHB7E3orrsbh9/OuP11NHOMK7Jg9Z4U9
pLcFZMAQKKMBx4NSPZDA3x/nIyRbNhMQktWd83/syQhmlFxQPiLUMTM7y6nnDQu9mulTD4H/psWg
NVFNmNZLxfJ0EU4lIubjEA/BOsQuJ18fxehnpB/CcCtU5Q5Z5udYuX7UFF6elbsVhYBOGuPcMlvP
BRsSDEVf3z9G26zKVflXFUdmzPKHv73ONMujVI7TdKzMTRfXEFxzAnEI/4jXZvUCz8k3FuQvurLG
f5iATQRPVRXyEzzN2YMbDcBCLzHtgC7yMTE8JOiwtuQgeLGGj0Y9dFJLSXypHfaWiXBfHdGMGYcE
FY9sQcTUsR6imgDpitRwAAEWZlnhyXEM+K2WutgnJU3tFtIr0qjVqWXmUyNTPZ8Qg1v1d6LjTW3t
IwliOrxU0BCOnt9r3QG+gAP3Z4zuUtAg0BhLrQXYdFdcKhWxG+qnUOCELYJUUDzpOFzDsgdy5ErO
IXr4f3QC5yC7m+P07r+3fHlONweYK/InpJwCQ86BL4EoD0ZoWK0NgTPOKntDHbChzp5vrxDLXfEH
e5Zttx96G9G4OVtYFJzxW3HMqmZmpZjgQ+K+/IYOye9VNFwkgc9f76dJngQ9qFlhePtRyFAGW45Z
Y0/dhs1X67bCGhYGV6v1p74Jjd+1pqBkNnDie6nzb4fR2IzJ9mRnHLfBdz7DJiT5VYFEece+h830
v+R0va+ha6d55M6+UI3WthgQEC81u//SrOrbXaLhSNhyLcQbTXdTlKarbedLlbZk4p99K52ZCAtO
5Pn4mBtorEFu4C24eUUx3SMBA6ACv8vEIhm3PEQtIRGje1VPPaBcdQNCuMifNBUs+w72cM5RKM6F
18ypQR0DXa7LZ8MF9/m1Bc3AKWJQ60lJETl6wwAeM9vr/jEeQuteRtfbT2yvAY5FKJm1CMPy+KE4
ZIuDFOSb+L61V1yvpB4IzdZ+lYT/DSMUSd/s/BhV2ct6xM7fAe+5FiVJ/BbUSoAiHnAbFLPzHg2S
VcpGkQvrOyUd7ERRiCZ0qUfbAu6LJTpUbNKdKZBz/8+CEhxP/lnTFB7ytdgnvebMcbv3R2g8oWAr
hgxvlEcBaEWyXOGv5LgrbrAmLSPyRGWpnxVuU2x0soSAvpF3zmrJzEbkP7MnMzn5Ifu1CYTS0lch
MaPHX3JW/2sGkgaP2eSmP6CWOQsXpG3wpsbxfLtVDUrrtrMu4N90ESwSVRie7gD2vp5rEcoYa/KW
4TunJTxy/8G81twQi0957Gg6bT3+EHHkd/imUN+2VyXdvjgTILov5PCjnzA21b5oCHKFw39P8SBJ
AQ2qL+6sWUmfE/80UzypPUhXs2rzR5DxJYSOkcKVQ6NthAo6YyuLMBnHRbWAZfOGPHQ+bJNwqmx4
Ft4yu7W1dnztB3FC0B9mVnWK+/MXuQ2xysrhdgmhYJxsL0/VAjTC6DsF2YTX2TEM9VkA9GoJaXjO
nrn42zmzxzp254MPtxsz/nKdfiCMM9Yz97frNlq5Q1LNXglLaMFVeeo7RzwkYyIRwpapiQHLDV8s
rPIogK2whZQ14/YTe8dQevVLYmwbiD7nnGZDsBmfU5l2YacqkOyvWl9lLnJdnz2h17X1EhvfkGAp
BlXCmuqF9qKMjyXKLRjhHpdMYs7f13MD+CRg1eFH3V+URhadMYSMY4AwXmueHIfTgQki5HjJGWd0
qHgG3iZXjLnVFn+i24OMcWZITnidiZ3Asxwliwwd6J2PN46HP2mOOsTH2wN335pzu2JS6460UtG3
l8qwr18FOhZ5rOxKQYCIp0STB4eWa6CN0h8qrFNgXXrFB9os2tw/10LhzSOwZLZTgT26fuOzTVpG
rsMg1Gvj3kWp8YQuAcOr+CglnHlPwvYsqK0OZ0TUMYWCVuYCMo8MeDhhTmMfypIP/NOuI8QMV3AX
c2ATCnT8bT/rInzAsY8ibHalta7YeFpYTc6Bx/iWyuL18u9oZv6Laep2++R1umsRtA/G+3XYiNxs
S9JXg18GabiM6eKQhYu0BSw5JYYMPaa2Kz40UJJFt0vue9kUJ9gVBbcdwzWQ4Zi5WFVM3/FKgSmg
0ifVKrVtt+QkpSjG5fZEShaUJpNEEqxH/K6U1LBSxpmIXMTcX/HcWSdM9OmyqbSXg6PhCd3iMqKn
71bdStKpgWYRGbOOCaICWczDwP4q3pPX3M2JMHR751BHr7h1D1nzdTGxRK6uLT9HvChaEHPrE/xV
p38Hu7YjcLRLcll2o2GHKltL8gUKGGV/PsFM03q+yQMXB1OyC+2Qgn15me5ZPgspKA8XKTDuocHC
J7e5Uu+Rrss1DmFz+0CynzMVycMelH0oTgCP82Mb+BTRjw2gCT+2f/dltRY9zPLwlFsG0y21XV95
3zu+ttaZobhY9utmcKKvhv5z7rx7w0acc1XQx/4XohBS9vgjxb+ys5os5sjC75J0ep5fUjQCCVP4
YtQVWf9FY6aaPJ0XwHBDHrkp3+RvCr9dxfX9UXBpNgk0tnT1VnWh1EMP1iyNh/6yJ5usUP+Dgij+
yvdyB5AhUG/YvNhjErfkwjyXni89Ujbemp/absWusVWzfH7UdTHOMDcGpPttOMrKocaZDjtiWcEO
0i+2a6EUqHAkarWwzxQMiKdzO46QVe8YEZJuoRMP1ybnDQivHO8gfUSepuvhQ33rn1IwxlaFSnXq
Ok1JNtWuw8719S5YYqZewrA90qlxFl3dwE937Kt1L7YEzHl71G3Q223rVuXVIr1O3s9Fu8lQfXxM
8+yXZF/4DkxozvzpPhNIt4ByKWNmuOdJPQjw/L2BgrI6+18ICGtrlnJnxYyLrAenMMwrNEBtQinz
F6w3Nb1kL2izDTU2qhPHPjajsGlgai5pfMfUUABydp5yJ2wDzFwA8FdY8NfEjyfJKd6iu25tzf7G
F7wAXLGP/NBMzzN7QDa+0KrcD6QywxNueeqYUW5IeKcyfysC0FMxwqVbV9v2CeFu/uQIc//GE1i+
dEZEdGTUiT0krrjOFwR1MI/hUGhB9F550b7wPa9Y3YN7OUxXzMdyUUAf9TsWqeQN54ml7VsbReBp
OHbvMzg9EXOBhNLmQRxjFJHo545WgrLQ6c8TLLBRiBFZTDENF11yXxa0M/3kfs9Huih5XhqzcWvL
jOjwEeM40PxI6jkItklW09haI/TK4YfeExZ7jxvJHGEfWmUBC+y1beQP8PbxanBelECXjIkNlO5d
mV7lWYA6gcPfl5YXkVWS1NI+MvpaBuyAv5ojDGq1TmBkcVJYpG1/86G0t8EwaVHj0CRga0JENdyy
I3k9IH/Mt846M0fiSKWWcqg8++i8P5vzEj2Irz/rCAouCUrG6JkmExsRLFb0SK12QQDp+f2TjIl7
r1EGH38ATLYsMTT+w5z7K2H6esXJ2lp97rZivGFOUrS14/Gx5g/XwugehfVTevL6RQkX7OZT7IS1
1OmlsS89xO0FgnT/EZX4CtsA8M1HIogKvU523n40NbAvpBUtCwdraOTPVQEOL6g7F76YztTuURnr
NOYRIK4pi9nkWMpRSDYCPajFgmD6a41Aik8IxYpDBB+n1pBsU6q8uObLN7Z5GDSAVNOcsbVyw3PZ
CR8NcOsJ2Juu1t1LaBEahJ11oa7Fpr4AHuEFxR7aQ58oVDnA7cVWJAHgZ1x7cD6V5lWnrZUMPmbw
X+M55TJ3WsYbxCyVHetYFoZnvnbpfcC4y++FM/Hm38Sff4unFpe4xWTq6Bv6A5uxNEhZbCkzt4Lj
oqYmozBqO/glCrU9dP31bRiVMqx/9rDouO3tVjOSdQt/tk+aAit85Oc2hgr/P6rE03j/5cb2Hi/O
dnZv5XVMurrWE2YkatLd4sVkuiEQoNxKfDe7IF2cnYltU46wt4pILC+bDEBXwYQFqFsMYgtQuDGP
mLZaqPphSrGy261hdffdzkWYqdGc+JPwIYKtfcqs8OAj1hlgnAkRw+kTSYTfEnSZIIZsCiCvspIZ
biedC3+bzuTG9E5ELUheo4xj14sxlLRpMB9vFCd1wA5h88e/lg1nNgVXtxoDqfOJrauKaYhw1xK6
u06rd1Caf9W+gdCCKuh4/f9EFvyvUDLW7A6BnJIjM8nKK9s+n28NdXQ0qFg8DajeVnLurldv0Qin
hs3hhYbt+y346UgL6wSNxcuCfwHw4ORTCuaSKmCnLmeSBu72Dalh9U0IjiwTuUM/11WDLELvq9sx
zxvKoFifVyKBuKdMDp/OPYB7/7ieV/3zjTXlWx2eHTz9FK1UzVyOZONZmb5moJ/eYEQrMlC3hMiI
jnPqaOkWQqqFE4cG7Eh1oRNh0Cmys9PGE5X5aM7EytfqcjtEfPTMGVWAJ8wkDPM2TqPyp9P0wAk5
68feubg4PCHzWOapMNdIPdQhqqfVxKENoH92ldwfzfAAaNS+QDQLGvDPHggE/R/js+12xIeb3iOf
vR0n0R6X5cZdQ3V8NxYudtNR6Afoiyl5GF8URMeZEKAZTaRKqg1m+KG/qqKUxkBsIdq3FK7IbnnO
2InW0drfmRI7HQ0+e/7r59VYu7QrMR5kJ6F/xLbICC+pws180yr7kJqcWtNCuTl+k4ENYXwJCo5S
YZHAN3vowiQslxNwe/SPN8A9sPJbSED6bJfkg29HWtphIajCEnCFMspDcSLmVWGo2G1u72u2teSr
fDvVnQdnYRNlzoTvzvSqzTk8Ngc/hANeTC/6eK+4Pl+lVEw8e0BNFW2yjELK9VJ3PWUcP/H39bvR
SZCgaAwHz3sb8m7OyNZGOqhHgkJm3GI2e69+AKDNyCgsIREfQp1VNnjgrtqZFT+QDPi2iFNbmCtT
61wQ7ZxfQl84DUv8f1eTHy/vQa/omF11Ho42Y1XSQKm95vVk3M5fD5hO0gs0hpwUyBiYHtiGP3MA
euAL5nD+Dbl6beJZRvxVvTk0Lh8TTR3thDqIMEJ2jl01LkvV7aGLbAkl+1wKRccep4G2MrqVZ3qM
nAeGFKsTayBnS8FXlxRiksOHi3YLIbXKc6NdJkuDsUd0Lwr8/mDop1vFkH8R31LJSKEdPJ68zk1V
b0IGesvqIbdD82VuZr8v4N+FG86HWrH4s7Jv34PkH6Od3sDVqPBaGJ78rZGV51cZ5WxBArt7vl4O
qj2z43c5z7XyzOQ/lPFbfAf2N6QHfwMgxJ3VG2H4MLMOEXBpCBv0GqZfHBFJzvm/hRmaYBNM6CXV
Vf78F1DVegz0DGXU5sH3xPtPNuqiKV1nNiv1Adi0MDJKQy4ewpLLj9uAH+eJyVx3fSWjkkqQGvR9
lBMNO4h6QjnaLxb9YQo7tmdx8Ro/7m9QdOMjXHP+6h2fw47Ka6gY7I4kshxGANGNGbzHZIUlDpv8
mpFU/e0PidYhnM5u7+GqSPhXXAcCoX/V2gslhR1T8mVZPQlgKXVa5DQJh3NyZfh8DTD3gmBFjuut
PacmPavQrlr8y4CGzCm/PgMJ0qLIba7aopd8yakuxBPNv15F4/CR4Mv/f79Wi7sWadPQx/V1SNea
pEiNaUcZIjUmGOOJO532Jgv84Tr7F8oQZTKIZ4ZSn3IuL6dn8skiE0SyIiPd9ozTnpIGEvpfF9w9
ZhCh0SNOHxVUA7c+s34jwhPRrm1tCH2LSUSKWl25VFKI1hhp5qCm91QIleM5zMjGsTg1qLCJqLTN
t1D5Qhqviho8A37flFgA1D8vZgZ1pcruxCHlPc97M/+qPlMPiWhR7R7Q6zLnMVypX7lwMP34CqEO
lHxII7qe4myBm8B0dkF7xnDhJ/d2VbIjsl9n6ruwU7qJBkpPxBVSSfofJtXQ9ov2iHfqkzYIzsgb
e2LTlU4R6wboPCCVaGlqJqDM0aWitBKm7gol8dgNkBI62JC5J2KzqwU6oqf+mJC/yI2Luwss1PCe
Cq6LuGojlvXFOjTtLm9dB2R2ro2dIwTLqyR9RmBU2THP+iq9gc0DmCmSBxhkEtWCCEVFEFIH5DT1
gAYCrE5TgN7zpR87+nFdoIzTejekcLDHitHxnia6tN5+qrkpA3q+YQZ9cm2WrK7FCzef01FYfaM7
vSuSN5v9/Cjxq3ZWHHgCM1bt2tWbukWrfFu0+PXnSLnw9woIbIdWZi7SK5VQX7gt6/HNm500KG/5
EU49JcA6OhL6/GbifE/olIxc3VoNO9HFLpB+l6g67RSaTSmjtHAZS3UPv9YDRycxMVWHVHXs3icI
eXbCTv+44VnR+igQsgxbDNMbKt/NYzsifI0cVhwJqdt0g2JAIMa8MEoMfrv5LxXtFhDOTxEF0APJ
ifQ6oqLuKqhh77CjE2i5wnrMoWze5q6F8eV5wC83y+rqrUJ9+gf8OhLM6tgQBpZtbsO6lWVXm40/
7sTqw0NcfyzW/su8DRxIjvWcSfpx8f1Gxe66zp1LW+GQDweXMLLfRGwcP6CJopWmYfzCT2/M13B3
V7IlQIU/piKlUHsrE/cu3XVqEfo2hf4LIoQjnW4aP6+KaJZj8d2Q5/7rixnsc549G50dZqIb8FTN
lmYBg4Y8d7fpH4gBwffWHNxCv1L3o3e7ps7FRx2v3rITfBE2BG1kude8y0UoEv2o5/R33WMB8Ev5
yXHI40rx2o+IN8/TJJZhcil1klJt37Y6VTrBm2S2e/5ssJmI+fwW8KkS26iEM2OYuFR62f/CprmS
ZDfPHjTFXUabKobQlchnCGCIUak+/QYDSrlXhRDtVEOuy99TFPc4k3pvmPlHr6bDf14e6z6XjumG
JBL7i4nV1kCK8LaZYcIfXwrTrPALntQHBDi9uRZlbJPLxtcAyul0DgAIhVTK++StphoeGBMUV9UA
T+To1c/Q0UyPfa92FqWZscyMbY5Hwr+0ZGzdjC/9cG1F9f7br6qUcP2d7L73tKp8yIAIKYy9cpu1
T3Noe2oCP2ChbKAGwKHxVdKuwKM6Xd3rVE9qRS9m5V9Sn21TIemj5SZeiOdhSx8Um2oU+JrzTNlN
sl7S4+kPW0X5EdIZYOLY8juokJRw0E04Z82WWF979APWq4hhc0iMqafQkpXzKB1n3PO1RcLuv/+O
tj1oZDDYDp0ksdHvb8hsDUeNk6J8GrVv47b9lz0eNkHE2Jktzg1LLZDjLPrKT2iGlO5iGjM9pmPC
IyeaQmyKN2aILPkYwDdFDjRD/4mQo5pTpK3RARE/KOlsmA5N+zBM6lSBCKtlOx2umYcTSOE1a+1w
7qKSlGTRylahwo4NmreJJCMPaUdY2x1jC1UFyZN3937ULBiNOnmalKutiKsjM2UJXgzfzcbPjcDO
6kGf0O1r10X6eP48lWSxAplEk/ZcjceqTsmzQlXbYJinFGPGNjcltDLrBwq604tK+5t5Xju2Dq8G
4A4X1FvryHyjHJC5e9eEXzI1F0+1T9+zH1aNke+WdQliuueAvKrvDmNALENcg9UX14XiMOUMAc67
qAZScnN1tq3dOacJF6ASgdHUDhAcHkhACOTiOd1NnDH/MYzLbiOXKhWv0muM7G0h2bBEnfr3I9ip
gCe0/pysPjDDEPR76qQaKxoFdBax16tXMCo1+NWfxHUz7yOnEuDWkQBzPbByDXRIIHKl/+fGT6sW
+ooNi46Udx1pEW2VK8ySMmzYscmJrnNH/3qwmXs7b0MBJ8aiea06mWSVdSAigPN75V90Eg1sAgW5
3qNihVo6NtqwGHWkc9471t8wxHNFQswxr0jmLUzoIbUnVZNMifbpP35jtz4clv0mobl8FoixAcc6
2z+4fzca7cStXduNfj/W521vYoZUhYO91w3as17Cx1Da/GoLSTlTB5WShtO2C16x0ebz/y7TMA1g
ze6IJUV3aMbUoap5nAX7PJ9hI+zRzmVNj1lSrerDe88cl0jZk7zOa6TMJDHyhmdcpBYHh7MIld9x
BZp1GigBvNzWZIRsy9fCdxySo0n5tkhqgQt31ezGPxi5lsMql6RVkRANYESaDgRH0L3nUi+/N/Ga
kAlhUfmdcAe27DFeHHVPA5OmONYsW6dzcjM5otud6mf6c7eVAoX3i1cBET2BykwdnMr1JF6gSXry
6YxkQht/Ny1tezNti51FQIE5+v9oh9nms+5J6rUX+1Uw23i1x7zOKaJ4LQxVWaFM/okndfex1wkK
uFZPjUki3tLvxKLIUbLaFY45j+NsGEbPah20cuYe1Ev2LJ84cJ4SB6ozZj5ij+EjvMfW3jnRQo3z
Bc+wwFY4PnuCmynQhuBFXzXYvEQvd5zc3VgH+PxT6z07fNMlYAqh0XpMhmA4MDJxbTQ/+yGxroI9
E6I/pX4MiQypbMDWdKvtjp7Xl+F054JeRwjOmYtP/n9L7fc0qSpw7PEfl/1zixlCdh8aw4oYUCPr
DJ4pUV5xgPa0wFiKV2ZDjskhSMQEa2wBZh5WpLAPjU1uOkoxvVx8C7YPRa93KWuCmJk3UdUDpEDH
pZGhv6oijODQ+Dh/GAILugBpH4zflPfT6886UBXJ9O18dKAVxPIQyrkHnTYkaIu2OAU+f4bUNPJZ
oGpS6tsNMqm/nvqhmickk2lpX99xlFqok5RpSAbRf+Jk2ped9AxOqwtNfejG7OjL0OTCeSJZYTun
CqfA7HZkXADoSQXydMzPS3xlpjctFY+nTASf3t7oln4s8KPecc432KNL0rvvzk8Fpd19lC6TCrUu
Obh//cR5oUhI/h7kCnu5QhbS36L6VKHQLNY7NeDmltm4+h4e6ZgAis1SvxaUQK3y1LfO5hkpAs+O
6imubzSG4TNZaKVvSnk3GNPfk5u522wiQ5Et0OnjmjAxLFVsZzgFFcqHunfRhKzLTROk6DN8XBAg
emQDY61UJNlnxuzQhpaMmDh81S/Qy3UOA0udYVSc0IEU3Ba65ru6beRunYvnlkav8fdbTLDtCPfG
FXDT8sbtTFxvVVEfkVw7W1qJH/tvojvqrrMxV9BjJ0vo4gGZJB1C1j5iKdGAXb2pQPWlkvwMIp3H
1Fajta6do+EKDN9fazM3VppK5geeDSznn0BLDw6kRx3bLr2UpNm4IfjftuQprR7pvom4JumBTNB9
K6K+eh/yaU1f3VrYHj99Of3nyCnxGgxvPKl2oWBW+SOPLcwkglsox1H2mBFV5055pOHgebrSeWzI
xKV7wcHkznhdMoBFCanW1GQfh/jAjJav7+Y/67b0+jXSiP7yOyX7Ifr/jWESIlcpe6F2Zqs5Z3hL
/6FkNBLcWSMRs6RnRWEvnJo3Z1bMuwl4CPp9WibZaQToUnywtzmnNjySgUnAMnKBH+mBamB3aWAG
28ll58SYKyuiQP0xQ0FkD7U3ftyFAfdsck77GQtTZAOgf3insVTeKHfJb3/EhX5VtfZIgmDo1bF3
R06QmeckVNdLwoH7fD+MyOKqO5sehJkuOXoNTD33ChkiVXx9cOh1U6yRZlANofkKVFISSSTYZNN4
lemBCqHaC/FVNPExZxCXAWReyMhTLGftOIyT+Oon8GdVdkQsa22UZOMFllWuxFMHqjCF56xBK1Zi
3xX0a3ZYdf3wBRD21Ew3jvIwn4sHPapSt7JydIkg3+dYdKrUqqpxtdPaD66mVBU8Vk9rRpfII5Jw
iH6V05kQdWFfWOp7wDMeSFtRup8DZpd3TB9rYyliIrebgX/7Q7b+JRwauMI4/rpmzIzp/Lkt8cDy
EQFL+yPm0iN2tZkvsuv/aXxEpb34vVsVe1En0htTQDccRGQaCqNYW0n5AR9ZigY/A4mkn5DWnIva
x8l722hWvVv3JYMiKG3vA1BtKbOgq2qgabiXTnCrDzRUMPb8Zj1IhCSswodHbinaGkI+vdHzjQS9
U8hT/3AXPz0lPqhSlEWtfnqfox1U2/yW3aCeEwwVNNtymeSTQikqtcJWlHVQkUiruHl9mrjj0OzP
lOpOnLYrSnpSNZeJW5tOPoB7jQfW3TmgQfZPQ3Y0ltWy5mSKZ6RGAg+uBsuvhlxVm3LZc66ZGh+G
X7UJqosaEIrc5EsYsNZel2OoejkgBm4wh6EJ+TK5YlkPurnMYR9N9UOEqRaUiU5GVEP2GVqN1jhs
f2eSaT2Ks4so2Yyq0TQZkXBwzNL7MooPyy4BT6Vc/vwjaZqMFOKl1eX9iyUqWBsypnouxD/2idTO
sFTZNw8Xms04yxDAYgY2ElLBzb83vqm+3+JpkIShBj6nyfCSgQadX6P7vG2fWVLnUngdiuXinaWp
Oa9qRb3kgxdTy/lIxsQ/iAhywuVLFxgvdPL9OlSAqW84hO/wBpKKLx8xdy696uBjZffel2MCi81u
9aRmrGDvhC7uaC59zcxdW7eWnKLBJETjYsr+GH3rg+6Yp5l8vjaOnA0zekIS2DqiKZ5QYGRDPMXf
FfI+DD/ff3VGemdgAQ/n5Z+O+16J8AGnUE/yfH3eHgxuijDJGl9SiAtpN5egAsWDhVlor5Mx9lLK
Ay80SKbbs0MT+jqXsWpm4QOYXk09V6wNjbtgVoV1h568Hn57V6vudnv1D/TRnLj+VBk3UkG87L5V
TDOHTLCTvpJ2UJ1kuOLf36fYFNK81/ubj0AKFyYVCMrk1+BdcGNngsc7gea812lv8W7R4ZsDhqeL
BRHrjmtTMryYhgwe+1GnM+KioIBYcEHzL+rqSjfOH6zDEzaKbaQk8vB2T3lgNh5EcyB5nCOlAVgU
p8TQzV3jrobAeCPvE1aDIJYODJ0l9G/3uUwppK2jEU9Oh5hFhJC0/iEnN5RSx+OSyJT9KHbnMVFX
D6u04vCkxzEuDYmBshVBGhuxjtSkhK3uDT2/p7LlIXTmaRV+iokqGdiniM57H3EZPCiqXndDdN1H
7If0Y6SV2+L51GCy+F0fhUD/PmVfWibmPHOWw1gyP/oXgcJkk+WDOa1rpd7dKTMVhjuwPfIjUOkA
c7fpp4nuM1eFqOelN5VZDS2aeA1oPIqTNxo9LbAFiIUdWtiISumy6Un6mvvl1m/1oOY1j1bsxXhO
Sz/E0LHDSAfhJIkDj/u7drUlokBh14Fm5dsUQkoAy+us6yVrX4gUDdTHKyHbV60+k8RXg6C9PE4B
jPO7SeBBTLV+t75tM50ARkQF52cv1Ugr6clsX8juSI/zy40jr1Jp7KlFTDwrfPqmDNyEU64an7+H
DZrCpFfIPuZ/y43btSpG7Z5j4CWbH1+I9wbM243amL9CEk1FylpPU6fImDCxztaF78a7aMvZYIgR
V9YnsINwZSkQ0T7mWf9rX2hQCd6GP3vB0vQEoPGd4n5ODFvWpsdKoH8pYmH/O91MUguhJ/flt9Fk
SUY7/dm1tws+tLRkJ9VLjjDuHdcJEMdbvLfwBi3b3HZ21wZFZU97qUkpCW8iY2HGZ/ASFLKBHb1t
bUh87zgo8k4DFUmgsj7iBpxdEkFWxUvUG6YNoqiplap/lfYbZxfTurfIiNKbIEUVEInm7g208DSo
FpqufG9OkecDnd7Wi93KDYMjFBBR39oZcu8BlJX0jaeSyrcpOiwvsAfp+jmnt43noYpSZ3nereij
9NzYXczhdJj64ee0vwsbnPBpFIkfrMa8m8YYnd4Cd081lc4xtnuo1hVzWRnoaMGiUL7RSZkEMQ8+
39V7bBQCoy/nGpH3KP/toftPnpPYZJZ629WlM4RZ0jzlGLcBX0BlKyH7XWfZ/xo9SDdv9tUlABvk
BFKDEdquB1+bYszTwi/11ss+FebvofANavRbAPYEI+ze2Q10YOzaARwuc3f4bIJMV3shhRSwdBh9
cdRC0TG7lExtvAoTOX7rSMkSUo7nnsSMFxDEBSaOLhFKUDmZlEGT5yMpx+5vThK5CRmlZgPkusgX
mCEbPUmJvqtAalsSg95t0xKTYODOrW8h5pzyz5hFnkUrZaGFcUTeGkLWX02psycUavGp4Nv1o3nU
UWl3ZYstgqxyvD78Y2M1xhbxUXhBeyUxhGH/MNl7qW20B3V1NLmlXleXw+HGJidqgfLM1kITF3Od
xD/IXS5GE5u0GV6z4YPFhQSXPEb+18hrlkemVGt1GQB/6h2CYwCi8FwFGWJlD1wrKXPIsyX2mYbK
RmAzIsSZrPDDsA742V8pCSMDQpN2uJR5pWNOygXiYs/MbzMj6MVm/qrChNNLqjtt8Dm566BBgfnz
63Wah9zEGL0rxmZ0PiuDMKECp/A5ITi8KRorS8k1yUbZqpcPlYZKtdqvX0ZOuuY7F+nv/5hCs5Pd
pMlgdfP9stzFJFhgy+HABzfHKia0GGb0zP9i9JTbALyHbjtFwlGFbAr2fYJi5tPEBtqKJDbsGtP1
v0PutROSW6dfDmDAaFF6WfqMepqdwlQMkcop5GG3brmX6yBiEOOMdo9ZuIUe7V8qhAEign9KRfmu
Q7irb5nAbqKgzfUdQ37+KHitutOuRPEgROxRUPfNzvOufFGtOZeAFH5brvqsdgqePOOIA3vHC1FV
unM34duS6TK2y7LS0boU1bAKPnABXc/65XD5zYol+RLYNYwFJUyMAxjA7uwnWC+fTNpyU0jokE2o
NX8srpBlPQCk+gLAsn4lIK/z+RV9rJu3Y5b049wp84rBAugSXEj2UA7QmRobjHxQ5OQ2prZ7+/Lp
Vpx1cJJNkt6APkzP6sCLapN6w2O8NiLoBnNQoSH8RTjAcx3W3TIAdgNuPhMh3tlJWHcgqX1Lv8/g
1J07lZT6Rp6yS3p+wcI2RfjFduVNTLeJpyVQCMqNFDvY/gNaKpbEc+4ImVLSHSV06FD50u38w47f
eQ7Rp1p8H+XjKQ+9h9S2q5NQ9ag46wKtVKLlEdb0Ijo75T6DwzWCegYsgn2yFj8iV6r/d8Nh0tnz
G7j+cn5dRkwRf5tBcg5GugbGcOSGz+Kabl6x0YeDaRshLK4ccftUHE9Kl7jiJOh8/Eqgoc7dbVfu
iVkjPKf2DrsUVBawJoWk+o7YjRKYTI0RBWmQHlBqW84HdoksPR51qCaet/f5G6VHNBESyAVFETma
82JoMb9fiYJDZXxv4n3R9MvXHRk7x1f6ZGJl4HN+E2IHeQXbHpIM7rb+3fnCZZOJpFUf78jeNwO3
MaPeHJBahwjzYBAz4MAUGo2QIFy97K3lTZLX1IKxCWlyvw8NkfdVjY4r7gwyIwKjhIJoEkJP2jI4
bsk9hX+a6JBuqti28NTW1xAt95/TuURWbEe38iSfQxV2rq7YTk1NCViV8XuVlHPOr+kaged9g/A6
yu4wDhzr0CkqbPQNx/VC8AQe2HUw+RDvf1P3oPSPxKV02tVKijq9v7uJvwgje/FUBhqOMrbnI6Ff
BvpXFVXlNK3q/lx9odA+zRHZBU3YUjzVjslTLeEvSr7UwZ4SQhZTKCBeFZeFJwqqhHbeR4MY9lF9
uaJaJEx25jFo2YIfMKgrkUgl+g+QP7IUmlC/6C2nF82Ksuvw7LF+dbzagBhS8I/T8xaerOa2rgLa
a2zq6RlSKjVYe0Omrx8EY6YpNEaYTShqX+67CkSJCXVMqt1rvDcre+TFun6zCGC4XCcQClOnT3UT
ap+LieywOIsG5F4dFL1qYkDaYxvqRQgMhaZtUcFJD+Sxwl3ED9/cgR19ylIzr+5C8r1HmGwuUh9K
maHkDfHjV/CnP2TT6zV0t+tQG5WuPMJkZoCwgi4dLmk+CLl83UwjwrxwU4lRCxn2MPMYoqqQNIP2
CeceHr0VQuUXEjxFjPYwOJKP8sfGVFUx8wu+R0K1NYy1VlbCWdZO05zBMGKVXaY8zZ+8RzhMPfLU
w6ilW7prHCAdgSgzzzILOtFJ2KRFVE+ECyBFeDoGHjTO46hDG3D7HBtRmANfvRSgQU1bcVbZ0MtK
2dcR9z9B+Tyy+0Qo/dtdCMMCe0mZ3P9l5vR3/CGJx4+6oZ1Ip1G5/xE57LdvyI53mYHuYnMjVWmo
0DLsKyihfPep9vMDnyBBK4IxkhRD6EA3DK3nHsCkYaKGhpCjCO8MX/6O2my0GNrKBc19GUt9qUvU
JeQySDi4xy1taklCYZRnfXuguTTJD41gki/P/ELVy1PrrQbYjbv8qk0vF9UW8wpfo7VxMa8g0+UJ
/C28dCbB5UaQFuvnykSz2e4r/AIyahylAeoCQYU6ZMaS7Ok6ahptEzn4yJ0wBniIJx8eYPuJWopM
dFjHaxJHMuUudqquHGPzmuBSxn814cIbo5oDetREiD8KfBSTpoP0o+T2vkawg9X9+6TWKbysssab
9366EGO0E4Mye9GaK+PM1dKsSTYqPjV1Uc0rq/Y+O3Fe1hMfaAHUA8SD4c73sS/VqKKPuIw1SJvz
SZsKcAvgSZMVQc/GxA7xVruOfOkthH+D/VpuLBVjRmquUxsg6YVzVfMyThZlcBazjYjt6IgeZgc9
y2XYC5Q5yRotzLPHkHNMDh4ueS2GMxaQQHHhwhp4qsiKioourizfREKpszXjuLFTDVVsLBu+YIpE
v2ax3qnPUlewoQNyJQnZ8urhMD9b6nUlhj5iI9iI9zu1SMmMbRm6WC9mkgKf04KmP1IH7NmpWyfl
CmgQ4DQbZIGztp0RAiiJxg7NojIHmvoesgcgM+vV+AbsmSIcy3fYb7PL5omuiwh3hSIoRgbg87Ox
oH3V9kG4Luh7JqcK4tf7qdkAhit2On/OmNs9CoE168YmqoNbbUOx0SnxQITfQDADUcDMgac0+TBM
aA9lPpLpaBrPkwh0sNolcQAUR1EdbgUERGB4I/jdv/g1J+v0ka3FFYx5qK01wobxcsmMgJtE4ZDs
wtMgOyZu8uMR3iT+VUIpUhqDq1D1Tp0ICZl2TYDi0b8F7DrQLEKXcsImVnu2SjpvaemYpx8nqCah
L57Yn97VQEc4985TXvEV93IeIiQYWts9qjkvM+CVUgZhwu13YOmQxgvY3nDFEYFkYSFA//DdQn4w
g9iRKMG9KU8jyt2wQCOk5x97oQMY0hrs9gqo7FV8+lZhAa4GkPts7YteQhAUHrpIikzErukktmGK
dpixokbIkuoJ0uxP6BtcT8I8wBZ0xU3cKYsDl3dsm+v3f8iXcXK8c5LF0+U6jcMjD4V4ELy3GcVL
NqYSs3+IPAuuqPRG54lPiYiwDJLUKRO08RD9ktlJwsSxHICaic3ldxWuNYtC8/9F2ySYkjPO5IN6
aReZ7TFNne9wOUfVk6AtDJeRtx4AJW24O2EbEZyJa6b6zuhl7+m0A4PKDxOeXzOJ+P6cOqvsMIjP
4NfPbwTHCu9HpiTSx18ZVGQWXY8IG8sDgfTZfbddk1JIqmySd5s8sYzqgY8CpfagvzMTVHwX/d6W
1VF3kClW2aotNDJuPFeYDiu23mU4dnkwM/g/VfGF+JbOiItLgWwjSb97xSznejg5hXmYEFO4fw18
fY2cCOQ4nbvqvKZZ4S4L1Dlc6WeQFJd/YdaMw+CQKeOamCsgtE4KrASx8Rs0wZ7xGTCYLRpPYT0/
x02TxaAQFOwQOdQaNUuPWyz/ReIII1lBb+G94JThkq2oR1SuTMcvTN2FQOQt/BR3uykMqLVlWG3w
7+OnBwHxiJRoPozRXIoChK2BUkLF9llRFXwiNOD5qqwzEqm41jHuNTEoc2JW1GPVY2mx4482BdlA
hznIJzND4Q1G+Y2aRMVxiGgJJLSZaKcrTQTZD7WmDd/W5QFppcYV9guqRGsPoNj8lmtdgV1C9tSk
iuROJnqnC2m8V7VmkBcAlTF4yHnBFXELKsn0zvaCYSHc+VZ7j2lfjqY0d0HiBbszrMAO/qY0+7Ww
RL4LBDtnB2tFLK9H1sCX3IJHXGA211U8inadbqgy47iQVJluZTLrzqwjFJqevJLRRViGHyJALedt
3/FGwFe2jB10CS3jt7ykasY9phbqkI7hbZGyDPI2JkDm+lj9mJ1Erk/JSZbpMyK4plDCc60tc7Mo
xoXt0uqLLn/r5++43xUCMsqrZGW6ZJQuL1MVJ8R/dwCnlHt7w77Isclbv2dhyrI+zf3DCL7PXLqH
Nqgv0f0oeyU1JoM4U0RwF7Jm3W3otBaicIMUSaQyK3kKMF26b3UMtalhKaSd+O1/te8x9lyNaCvQ
2tDbxeF05DkK5Ct9hIv/Gb/o9Pey1LhUjYepBBT8XkooJ+TE9hD6bMuns40H3TL+RJVX7AglIdfO
H2vO1gvRRTCnrOICwdFwy7FG4P/OmVkjdM8iP8LQ1M4Dh0zFwXlWbjkFJwnhNnkZNnA60ZFvTzH9
BzF4o0ar6xHsNf7rngn9/Cnhada3ySTaCnbDxQgPyj6phyl72SE4RQBZwo5/OvELNLEsRtx3qLYx
fVnsShoxEjU7DbDZ+OjnSDiaZxrzyyPaYJ9wfF58XCP9EgpOkCtS/BvORymISPkK/J3Y4XuFIjhg
fKYSfzbsj4JFd0DhXL0OZwOFtRitDLaYEFIhLxax9SoQzi78JfLez82NGBAMvYS0+94u9NOIantB
IT6MxPhiHdhjCjrNqQdEhB50kRamz+2DqXNOympqcM1D0bmA5fhNTVDzlKj0w4HbncFglOD5KYSa
NTol/KT3tuIkNK2pLA6U70fLT26Sl2E7gANSQy5RIUcwSjbmAcvclwV0whWKE5c0oOi0dWDJPWZ5
SDnOOoj9dfgav9sd22GjCCeVJ0H3J4c8u4qLBoEIzLml7gTppmxWpqiOLFMtf+wBZreIJojeOQ5z
luvvzFWCIKkqanFmy0l8uE+eLE/7n4aF/FzoCvlkoHFB+64ZvkhkZA9eDoCeLnnT8bqxdO5z9fzg
wdCsz74+f7JCQA25bt7laUwgrVrz3YYxHAHfnE7fJUgFiTRFGa6ZbzQmKIVqoJ0LqMSl7Q8Rg51U
z17uXe4yzDgY8feYzKbryKk2ycOkCQlsuYaqOp5qWMlZMX4araQ3OQBJb2lU9WCLpADIVEMvru1t
/2X8q4m7kDSDl4mFDBlDnuUAutqmwM8V8+y9pJemmWYf35mdkK/3srRLqyGYaog8V57p7pDGL2yJ
TgBkSwLclk4iFLW5j15DLop+4206NcuFYh+uFf8mA7QxQ8telgz586ibTkN95gh9K/UPRbGKZ9Nt
TLpv4y0NLlJpOIF0IPhlxcXNJMyWxtjLZcDTjO9+LmjNyGe8cwRlPQKjh6tD5LyDMrPAYiQxvqbK
wcobdQ5oy5jhuS0s9FwmfR8wGinvpjBrj/cDGkcKOdT3M9VcGqx/i7wuciwj/+QJaasZvoMR/ERs
Jn3aBCJwBuVZv/X4SZ/wHiszRVYJQkKZXqkApNt6KkrBR4GDLLAGUEeBd1tfsg8GlMFL156MfNJr
CF/VJZVn7a0hNgpFklepj9HM5YOPfbcOQ0wfvJIUsoonP0zP29H38J443+nRYHo5cwde/qPM0hgu
dJzbdJtDcmI9lJgpCCHZvPBgf6iQGti2ph5ZZkMEpNMjguFw17YxpLZ4akxH8KaHyweIC93eS0G1
RMOs1PhYPFM2bfWgi5Y2USAMu9N+y5g5ddf5mjAzxpHOwywNcACts8REgvOYzod79eBWyYo/fT2l
qWn1q0ZRpG+PUt7xUz0fepDXy2mBjLJfL5SnmYoi5qineEW3gfyZyP7PsxHnkFhCN8GzfwIWCMhN
7S/O5hQxH5okTzHcC+GQox+kulcJENXa6ysLytFF5M7BJO5n2x3VW72fkv/u71qvsousxTxwQUSe
uTbx/H85B2a5NlmMEwVxv+7o3UPiB35+wRVNcJYB9epKaGwDQavkaOXGFXEAlIuuj6Cr39reAUv5
NsDIA5MmgHkBGErGwcc+R8aWFvgOTh/6kYLFtYa45ZZij1V2yQteiybJwKUnTiYDvfxkY+Sl0L8i
NYNDPruBOFU04qFcceyiWC9ldZr/6YBARsoxR4j4WqqWIRUFOap9qgnCvOiRF8Xz1WQjv48hFgU4
UacIC9s0y/pYTmOTKJk67AxwMPFbLrpFZ62q5AzkQ0ZRGcx8xeeHuyswOrNVB/rNL0IeHxaXt1sn
Ff/3dhO31sjxoghelbIpP8q69jBNF5g0LkPQ3F507Ou/ahM0LPFp8qqCs69e7FS5PJTB0srxjsAf
TLWGGzDusArdAnDqv/9NioSFjSocliwSavMKR2Jt4ALuy6nrj0/FSDay7kaMyC0zShCLhIEFAgTL
ubZZYp+1mA3Cckx7aJjE05CsylQl/KMYVlEvWJZKrpOqsCc4y4+qa/PmZEuQwC8bhiNwshbZu6nk
BQeDfA8P7Wz40frjjKb2jwojKzDTX67G71tMqT/XkRvSSLE95nUA6NJY/gK81dr3lrG5wr4VWDRo
Nk4QJdr5aJbqWPvCYJv/R7CnoM9b3cadpea35etTrnKTvJe+zNyuhMWlZbXDxqBlFlqs2PcVG0Id
5d1mSUV47+ea0/vj7bng50XIyf/g/IGYDfATIt2oEDzp0LJnFpkpGFfr8FXbXdbW3jjq/XoNdw/2
EHqNPXEAG8fx0Jkh089YiF15UbuMc9QjmW5KNXbiOoJpddEZeiTo588BOZksc1A8xsevFDyTUJPH
Lps++LcKD0kkQGpqbFUnL7367o/fcRbSpTqTFJklZr6JVpZO4xRiNxuhYb7+HTmCegJmZ2HWQuqj
Bn0hOfmRxZxHRowU6Z2ojwBrH1vM26Zw9bW0LpgBBaEL8pwckTyPXO3KthqecSQ2oSfn//46PwDl
pyJ3w9SVlycx28Du2vdmjWqcebPlsdZJa1gHZiseXOuW3eFXeF8ss2hdgGgVdA0TUyiHtv5zM5+q
GfmVr9lpjwAKnnNo+mMmcYcm6Gz1dABOV56Ely+iPDpyBEenkVIZgROdWJ5qk0ZKcmOWVz7upRTH
G9FbLd1bOxR12cQ+tJp7YuAuiPKAmgBgqUn8sxsh83iXaIEI6wop3TO4Q8r7bDCX0pnxkCpio1s5
uJUqCJdGh0NUY6YXHvossFTP/2fL4cE6F/W3UN+vbdB2dT0Hcq42l1vMuCzqydoO9zsKDE/1uUod
bk1AcFVR78JBkfrN9eokDLtA7x7BH+bVDIf5R2RQ+dLQ5W1H7nju7dFUCc33Tu6UZnGGBaRCz9FU
2P2LuqztQLP76s8aWpNmqwoFUZDbcjEpfa/gzoyVDaIbS0l6vW+3qfbOIDNDjfFkEhBO9q/yG+sS
944M4mZxbASs1ZkRnAwQP2cy1zPA16vyzXnAsagX6jCB0EIW5WVCXY6JH2vRw20y9iUOkr32o4ch
Bsa/szSnD0hf1ndG/6poDRMj3UjqUOMZlksBsP3eeh5SneOdJb06pqxYg2YEzSvsL8T9Z6Waa+ul
qnr9zImd8h9KBkvkBn+oltwQ3V084KRi03QpZwc8Lc6MhYL2NGx/ipKC4s1ZPZ6W6fmYmYO1PwWx
vUvYkrRkKs/iQi6NN3FQ/0zloBGqmgpEa5oiFBO/dN4IXihuExT3igXipLPahBiPEkmQcl+LeMgy
n0RHSd4oCTxoSxMfEfa6QZhelXCX2zVYV07L82/dHJoOmB/vxnRpYLheySK6JzdUdPwHFoiptwFo
XqgITqx08Kj3EuWaVtDqCMtmAYlWllTtRpkRMtCUuiUnODtKsJuBnaSf9g4D/rGq5Zl6kIbONe4b
m1/jTSCtDf0TFVrfYz7fBO973d23bFV6cfFE/dTNRd+WgJQo9ee3z9D3+ne5cpLztJcq1+gm3tF6
Z6EoS+KHa2qK9grHfp8lGaWdbiw1TGBrbjjPwMAcVS10xFWTEF3V6sOPAF+FPbLZELz+7/QmJEL9
bh8GETsL2N5Y4LfTxdhMy9EdnFtRZ3a7bHcC5R07TtrBoKjv2xmdVCncBckByS19hvXomAaEvgbR
sLUVGNPmWcTpE2VFG1yHhRZJ5et6Snt7fH2LnDrCE7xmQ122iy/Ofz03YmvqKbdbBwAOpiqNgjIA
GpS0LI0zEuOqTdama68Jc0xIVlaPChQhaHJrlMVaFjugWSa8JGUwwwQ1NgmPCcr36rgHhEvItSNs
JRdoHVevKfE//ahCuWsds0GXdjhV9OIlv2d7ZfGj7aHZqmEG9xMYknD0yO0qNYDzdon0eL0+SKXv
JX2YzEWiHXRwB9iqamwgnx4YjRRFFagfLIH5+zEHcURSetkieFFXkJ5O3J7HxaP1zNA684OLzp+P
m6KBRZB+qC9iTdzL3kL8mWQsy8Y2cLO1aKDD1T+WuRvbZuWPEbTy6ugEDsi9iTHwBjLXiDTs+hU7
tNh4yEvEJrDBRYBtnzDC0EHvxax1HpWiKpv+KXPjaG9GU2We+9XCJhyDM7DLICZMFz+D9tVW/NED
Eg4M2sG3jmL7Rn9tQzgt70So7AjqnnlnFq2cTV7fU+DPM/dAsEKNQMPhBUPwoBRVp0s9Kb5HFOz0
+TjqlbyxxBxVVD4LuctVokzSphLtwpDs9dkWfAZqV7+T1jh4eS4UuhxxnGykazuXxzZwMkJIcDb4
Xr40qqiYb2rU4Uwk6ytm73xQHdbASokoaLVsrjPlxz988bcGSJBnGJj9+BsXNSfKNjCLVsLIrL0e
L/mBLfjrDSx9H5HZOiue7OyO18G/oEVH5tfoRgEvBF07iO0LhEtghZCmfYs8lHz/Fnv1Iu60jDrV
baOyxV5mhUk3K3CyJrnSfm83T3TOVbXqLmEZgjSz9veXeNmIW8oopVVB6477FAZbwFySMvHL3/kS
7Agi3Svinl+Ml6vZksHtv2zFzrMMTtPuNF6/M5J+sWdWVpuseckFlIeIOF1pIdCVDufBOyJmX9vq
7wcJxbrUkkY5EtT3QDnPnK49NwqK8cynyz0EJOwQP7GTbyuHPBnNS2wACezWYEdBWkV1/sVVeBWM
W1GRUnAZYMHDsOGiRG5cg3XlqHOkgE2v/C9hB1sYIMI/W7Yst4pUL1FKp3AcdYkbaDuG9TyjTSRd
w9tMoSVYBkHxpkgHsn8XC/izvjF0af552vIGDR9U2C3CmbAV0EArQ90T43QA1HHRvkkPm0ghAj3m
Exba44g1/PCRKraA7MHM2pQBMDlh1ftHDSRg2y4gbLaha2b0Gns+aZS1WijucxsWddL9e98NQc05
P9AX7mC7qBPifBYN2dln1ynyNCYcbWPnLbdc/m4qf5NAX9QDRhqcRm30AIS655dPLXDwJJiV0lRT
OEO0msMdWesP785cmhe+WWfk32+iA874F8QP+xX6X18OWIVlCkT6rtvFve33XvivGxEZA64HUT7U
jvIEyJg5EVk8t1iKp6ytOKj9VDrXEwM6XrO89KnpldO761EImQ7Dpq9rjcVZXrMecP3N+IINe0eD
IB3SbhMhCWtYXG5Jnc2ddBekeVkQfYnQrT9cbIyyqtyFYuyLZ92zGzfZCcicme3aWueZ0Gwa/xj1
JdF6lyV1lGb5EjHAlhdQ71KygL6j0xOxknKbt3/mef7dUfZZYdUHbbI17dt/jTzDqkD5n48wIZAU
0qCTMm+13MNlfU5ahyTSIDGRqyj44Cb4sVe9LxCBMMnPwwTspnYXyA8OMoVxuueCsRfo31QxF7DU
qiqTROjLBe2fO8R+lLCpAb2SEnQXPhKvnXTsFo5/aKywHpxhjEzNQwMVea8s5GztMIC0C6/sMXxW
o9spXIi/CO45CD3DjipcITWTb4wxvxyWbqnWg5Pp9g1ozpr2txdjfHVr9omVkbj/E86kHEM29U/X
Gb4CDgnVWZoWoHFQ1VXA5FHuUu76rQ99f9McxC7lFYqdGSEKIdoSO9aFeLrIPEVMiNNZt/wRiplm
+abypO68GFZqira+5EBQggpDg/7vYqTBY8YZMqVQG5k4peTVXNi4QVviBf9OT2FLJvzgu3KKhyit
uNblrFYLSs5e01dWm0R70f8k+Q+HcHxBbfubDhnD6cQCQpaRqqooQ2mAHPleuiztK8+TjZWpmUOd
OJ7wDt2zOdirYqPuZdzDrav+gcQwgPG0pE8gbGxR2u92ab6pOPk0LHGr9H6A3lpKU3iOZA/djsjA
EAfpdzqnSnP0VXtTYmpQun4k/EDjZZJMtmzJTuwICeP6y0VwZZuflItvCSdrWsNwFVJi6r9Tg/x+
3tVaY/VdhLjhsx6xQA4Ushw8KDX9gAtyccWJhhLZsOa6WchcEo2YdDjCXu66GWVUISxUKPM/ln5P
wONpzcOihzX5dFwCrLQtOY58GJ/FJB1ytioLwxMsHLWkhNRQxpOfgDuArbPRfMqx47ox6I00KYmQ
bfEXU9HEOjDcNU7JhG7+yGhhGNyTX9nXevmY6dNlsArMhey4LmGUPWpIoWCtNS7Iyxl8uxWvx2eq
JYLgkCi2/uh6CFXMQjLCVShNpMTgn71fOzuLmcRVo79bNcjaexafoKXTmX3bKNAfrj9y6VcJHYUN
IShhKOK/Nt6+VN4NwyLlhtIB08uB9dQipmkUcIMoSna/6BmAixQLO3mUtQLd5ylvrWsBNh5p9qfh
L1GpGB1s++/pKfBuH0h370cH/BVyrRwRNzzIv7wq7mqDPwH3RxoptUZDOH744y+rHwuM9yrh+uPB
fjT4V12rCCRtErL2fHF0XGjj1DXNQ8rfST9Z+e0vQ4b8vbyVVNTZazHcyz2L0sycCpCrddnr3nF8
WU/kV6dUFn5gZnOecWV/w4NGI02t4pK1pzRg3NpnQXSxbEPT/m9/1rjBQtri3z/CZAlMzmA1SoxZ
KwlKrboOEEIL+iOAAlPxX8b8+JmlfXrWl7zBoYqUV5MFs+ghvW8IkIg0mmNGl/QVrLySWfrgPrmt
am4csgOD7q8LAWssTUMcUzfSt8eXrKjkMLa7NcRhnkk0e7GfEYlRGtkshPe9GCDm8kNlZSOKBxcQ
q28gMTH8uaaRrypEnsK1mgPQ5RFEncVkOH3Q8G5aP53SSa4+VU1nAFEOgBaVSR6y5OoVTsEm10yJ
oJ2PUcRmV2KodS44FpeYVWQrIGy5pABEQtlWV09PjEX12Uua2qjQik9rP/+B8v3FxoIwJkvfBY9b
Y6Nk1UiuFIHFhfcMJQi2LtQVr7pos5U1R2fd87aB2N88hL/3cqK8FlM9tLNxN7ed21LyqrXQp9eK
MvHX1rR39T+DVFqu1S5OpwPJvzMB0Po2BvpAVpZISxPhq8XzSFfGXdhE2lkjjnSOY2pacgc1R5IL
naeLcEdEVWJWVupnZUoX60ruhGm/XNkc8Ds9MK1BSo+FCi+diZR40/PMU5+M6HB5VoFanrkAURyL
WF1wYWwGB5ZxSgsHDc64vyvadPIqyFCnOYmuw1Nky1oGCBO6T8zUOrkJc4GLk/pN4Vv8CmXx4NQf
LKPH1cgwyy/dy7EXa/BAoNqCtfyXjpyGBFnvUSlnrFFkA8HyRGGAVhG0h6wM5HhR83kfo1TzHvjf
3wPsjXGUbEnyW9BJYW5b6e7urx3arEDdxQj8q5mfjFVPX/leQ6z7DR5LSkOJ67rQjMXCItp/Xbqt
jPNgwyVmEmTfv1UGRjXGtz8NULnL+mnd3e06X2SG05u54NSUmvYRTd84Gq8WbnA8SGpB80oKbF9u
AnBxb5GPDn+b9v7fFKnx8YYPrrZ0BjsyaVrpDMqG8+ahmEV9LrvMQP4xP2zi777AnMHnF7CUtG8n
0wJ0V8hqtJlenSEFgYf8eLyh9RNI6eqlUbtFjo2t3uUJMAjRoo3GvYCauRLymqY5mc2+mUfa+DNw
i1UOV290EQE3xJNX/3qOvAGHqr7953lRZUShJ/eIG/uLtnDPcXCZwzL1TfmMbq+MQtR9o3+QOeMW
e8el/CCbM9cvWHc5VjLd4167uQHmxqV4YAZOl2T142RjQOC1lzm8xK87bww6P3Kpfyn+a/6exdDh
+Hs3lfxRhYDdDUJuLUG9+6OWAH2Ap+iH/rl+558hDtHFu7JAUMw8rge+Q+eGkZsy0YHkpBJEa26r
64RSDnXHmK5JSRMs/xWKnESjjTiX0DQU7CE8YlwaUfcvLgveMvAM2XtsdGMCksfK6ggRKEvOjYyp
M00HIIu0f3GY8bt2i3W9UdZI+c2JNTD//HcAnHBi+qqy+Gl068YV6ymx/UhxnlTChs6u0roB4hhD
g2bGnUmrRAYSbv5SOwThYk3KUG/M4GCVlx2QCWAlkWfYPgZTBWGbTbew/LWo9+B9hBJ5OkWNaZ/w
bABgY1wrzOhqRyKcqwhljzXUO9AYGKOpZKSzGaodXOKe+5XjwFg4u3I0uJPEizTY3v9cbXj3DDOx
C0pefYPMsDGA36BJtdeZfkG2JAJTbA7aAwsvSyaRnBhtHfUasikKD5Cd4Ta0VeH05SXLy3paRXyz
cDuDjJKDkm2pVFxBYg9aGSqW9AhJ1B1M7aVFhv6Oiuqhj22VhMl3dHiyGhuPDUAeJRaUNZRT9qHr
dFHB0yFOsEYHLI5WxEhki/f3jwseQx3K7wnAXgdedJLzyxYjS9WH0AsBri5h20Xrm9XBfcsFWaIP
s85Mbi3BWjJSiUArx1XCAgN5kqRW91km163IDk26/4cBTlBpw3aVPkcoTZzudXKhv5eLi8O6HOwI
rs+w3yOiNIm11GdZPK1cpAiIwTHIKOcd2yehNTnW7XWcQdSOcuzR4rvuzyA8IDzxuafnZ/22OTLA
wqkT3/1uU5Kamp9uHj/JTGIdhMYfeDnt+At2zO/Iwe4DjlsztBvKO5MU4Wuig5F1YBq0OBpwbsfX
pJET00srLVAlYOg8G0NFr19Yzij8ugi4rMrHHGpTGxESahaShBKlHTnAFto5g4dmBJl++70Xlzm1
kLP+tImYRxpF+yUakZ558Mapmk1kqI1T4zlkMV4u+jR2YLTEfOxYanIkVqwpedhBjyWM6oVeG7Q/
4aNna0kMh9lqO/M/rwies8NSlSOuHn2YV9RcQ5U1IDINDO6Mh+l9ebkjzZ6f7KdAL3ImJgRvM+Zc
bYSxnepyaoOuyjUMvJebvfXeieB35umRS9+SuRkEvBxzgQKioFyxlLa3du3Fn3sLRwSps6EPF70P
H8odShJKkTaXYn4oX4KvQ2qTdAWk2bViw8Q+AqcZ57kOIcbJk6ain/bBZHr2UfYzY4eOlMlzHRIB
S0xcGKEvYRQGZbizbH0IbH1GJP1UIMHatBQN5Xu6iic3GAsfdUQEB3cgoq0MJHwmsOwp/r/0KA3r
AwqI/ignA64gvK0z2QD/YqF/1vQB2tg+5xIZ7tjjvYRM2eA723uNXXzxisyK7AYzygPH7yoVIfpX
S0nK039oI/vzv3txW7VWppo+hGOrvYAivVHXSCt+2Jutg3R44C5AXCluFU7JhdVk74Z5qbTa7GA/
YjZnCRTKhuzmDxhjZdvTtCcfgyBZZko46jU1HW3jUrvaJEgpx13AeoYb/7wl8UEbPma+98WudHTf
Yio1qYd6Tp8B67vW/VmCGPe0KQ2YdK6aaGnoSHuEOxkK5eNMZ5KPLf9ySCK0xfr+/fSXLVh0HVaT
lhKoHMqEGZ00wZz0Zb+tJnZAJenK/jmKtmD5h5XM5MHNCDtGfRaeGT5gGnCRxMq+U+hwvl0fvaxu
0MC6IJltnd3Eq7rUk7mwgwxeP7OlClOkyCM1gsuX4n9ZIEpmJl6VzXfJjynrjH5FhUWcIZJfX2Yi
yyKaDK56U+xOJvup0GsOeC9iysek1zM5G/mrWlT34zlkk/u+x3F3IIzmGkvAUI+M7UFx36OFQWrr
703HAW9ASmqi3fgl7VOlziAInHTUqc5LARr2QHYR14fjGJdfr0rIvKVLtGXJFdADXeZDQYw4w5t0
musmfu9HnaDAutEV/+UL74vzJbwp0WhwpvlPPSPUnUtWkx9h2n6V/T7BmZshVMqtG2Tk/HijG7KK
pAvxbDobNJwQ2ZicdVixlVrBJSTCyWYk6ZFWaQYnwfjIRH00xgR0Xu71CwrQEZdf4ExXy5qEb+ut
jxgR8fD3TzPUCWY3jVV2ddtlkBXbYaqrsqVwO8uAMwUnp4c625J/QsgrhawWNuQw5qdh1p8fPmLb
YTi0++hnHwC2YKb9gnUmtm78pCI2vB+Uy/5oqlvcXgDSlqAqUsB7omHpCwXlyF3bicBc+jvzb5mp
6Vev6C1jcSIMTY0zno4uYYR8Ie9xag1EcPfvJSclvc0QpwAsypB38Y6Vk2X0c3QnE/r7WPu6fPp+
0hsPq/M16RY96+OycCOg3JLShkz4AHavQXXytv2Td7MPZ08bXYow7mUOxuUidsIDNwaq52YwudAY
ob8ZR4ID2QxvoseD5/kDN7i9Fhbl01MIk0U7N04XvNT2ZRejkIT1J0M+AQUW5MS8XeDn7JhsvHJw
5y//yixMLdXJfX39Pw44gSf1Dhdydg9QsMX+6wCujqwLi9H9t37lVxJebHcFG5scylTKyUcd2feM
UFzsWAuc6Da3e3RepE7447ZzMJll9pwyhr2aancg/2kS9EwyThXOH5sAGvkpP4Q8sNx7E4zpMPXf
LtSNV/2ngjDYWMPu0+rLUMhH0xJnXcPIg/0qkUuEzlSDOLmpO8TRpXJ8kL6RfdrpTTLYe31C0REl
e8n0VhUcvcPPTJaSduhuJGxCpRJ761/IKhOW6mwzvUwrIjT6fGMfXJWYOaQBZ9ldmbldqbzepDjR
bTc0hnTK5/UeR6ymX8Jk9WemEPpTxSwbRO2oxsRHvoYuzufZNPgYWnMT2EnuUEHpfmLF8/4uruCX
mUQ6VshSoFuvTrM9Ye61wvdtsR4kXeX3Zn/z8muZkTU1NMIrzT03hhsVIuK/yP7rdVbF8LjBJ6HC
KpY1BqlwZiqYOCYMAKyKU+TrJnO9OW5ic1iEQgL1NceZDb4Lek0tANhi3c4NHLOqyCsA7TkAtHny
V6bTNDp+G3CCUeViaj9PeqvmTWHHiHP1UbfRproM1ujhunylcDtVFO8ChPbV+FWXVAlIcmQvcJIv
Ti6TuksVz9T2rFwAFqmsehgBOIpHbg35hZmEshy4Ri0k8kvcxuZNteAtBGdHU9WKunPq1zuDDnZ9
9TUNvHiBVntjDSuNEB1fUmwlwBuEPjf7fTvvSSA3Lcrh3KzIBi/F0poOLId1gJkGEFHSpIiIDAWT
59+dhmez+d7X47Fr0v7Z6dDdVrwZiyLgONlda97YqMjbM2m0C3Uq1h5VM5kRcsR2Jp9aAj47T1k+
UheXQfqrLPxoNLrwYkdNdMCSzLE26VmVtK3uUGeUf1m8fXj3i70ocSZo7VJI05Uf0gewv0+Z/E7I
ZLGstOE7ZYkzoWi1bcVIDgVVEk/d2+Uf/JMgtuMbAThIyl5/rZs2d5JPJY3lTxDrfQXhTTHLitAs
YJ9steDQXntnrdYCbfshkt+133IwYhzoHHOnX6g3zAHIKsPjVq1h6jOVIaMV5jIW2wHYaQgHvYr+
99XFJTZImFGO9aHTWMz/lFBUEQzQzS/EHVT/gLTJ42GFPLkflBGw4cZ00fYYthz8HkbWmq6oWg1t
Y2yOYaZhaL+lVf9DB1Dzq9oP4tgVxnPSs7BubkQVoUCfMuwjHYQIxF8RCOVPnBoaXkr5EBIMQqTb
wAAzbBY029JcPtAmY9iRAjZCqqO6cMflW2SBE0Txvkg1i/JgmHZ05LfohCK2+TOjL31Dr7lfrLkZ
Ih0RmAGzMg+lRsUE1PEssm+CdcbgK3DkDLKPNqB0Np2sIh3juUfJCepHi2qyip63qAA3ttN28i7k
8eDcCwpsAUP1dfmh6ryYeOc92zelnCu/THHnZuV4dqvq3qKvRJz3eqgNHcwAmkxOhnidgRaijAVr
jNN7EVsDGCGRfiSPia2K1SaSTq7wBygj66gP5yWBmiAcVRgXIwB2weNOwOfNIWt1hI+5HK4KOx8G
/JyEME3+urjRU17P3XcgbXA9ej8x9A2CKvgyCZivdT4FXOczdNA/gdh8WvbEqUV79SHJ7c3IpSIt
teozzdU+bKpbR8mnLQu+FMpL3eNdpTJodQehDcihOKM0BoZtP2evoVNQocdd+glwokFnLMY8QXwg
9KS7Vk2UhpcCl8BSY6NyZk4Q+hZL6k2HE7gHTiKsBWz9n4m+Ljui5yDQysOOn/DpqOs2qRcGabwi
1wwzZkEvZHUIlpR3E4l3Gou4tTkDV6Mkkjdws2SZUsGq/rGEQXFysZqTVWDq6HOutuaimTUY4grV
y+iu6dgeFz0pp1AIsOaGdQTZYf9eFemrAl+v21MEcoBloUJChj7Kk1Tf3VJEpGEojibwZGljGQP2
JTXHSBeR7ra7VayPJmbmNVQcaVlSJx/0bkx+5PfXyBavT5718By7qyowYb/zQhkvy34uDl2g+csJ
PIJGHAytsO4sDNhJmhsKPzHvogIM/Vq2kJRLoNw4CqNbn95t4F5jN2FbX8vrH2JB97N+EK/ycFUn
VdexExgXPJ+mISH5AvRCZnIxMzsnp8b8J90ggdsfwCi7EM0d9ossujpAFErHtZ2aWne9xFocIcwQ
WUXH1SlSYTYtcTiU7E7APh7IXE5AqAuabSmYj1mINdUw8DL06w7YzGc3wPqf5utZ1tmTs5p0fch6
KD+3ES0OgbcSfqC+TXjzuP9or/zmQy6W4hnuzRsiTXHutvQgXjFjXW02HR1EhauafUu3aOw9hn5A
dknOLIIB7Ku4Zd5En059gJv68TB7Vo6+hg91O/EkXZa6SZJ9dgidEafnLm9fot8x0Vh5pTZjFzx0
O0GTj5Hm/MriUkp5eiMrQyRq/AYNe0BzUWpXO6tbyWDbllwdGc6cvfF6Zz3KReNrNdloGgXWKiCU
Lsw3j+pf94FdAt2UWW1NjxMB02otuE9gi9EbatnaO8dlt/iu6VFtpOHjqdUCcSMN0p+XLmf5g/sn
smE1RH13o9RPUdPTKU1BErejGMVJMJJ/cD+VvZD4onrEXHv+kYCCBIpk6SrhuZP5jTIzi39QtDCb
e6HvW4TbtVneibkcXHHruqpjtCIuEoF/ik4z3JmX30q+22jR4x+D2InoM/VM/hYmJeQpp7G0V0G5
zhlapnI76nmCv0gMRKwbfDlTaXfPba+jFJ2LSbUkfl05arFXScyfUl9vKjo0CxhR9DDvWA+qsBDj
esTXDxD/XuwZAFC7l8FrdV9Shu35Re2UNry7MGNzzyw4banNqVfhHtR5c1MMARuK/djqgvfSMl9A
4kzl9pChzsdPHM96869h3L9dmji/sOwX/C211D0DWRTtpb1HpByhFK3MhFP0X1JT7IMTRA+HYGuX
9hEco0iQkNLNoj6yv8LYe2i+Wm7mjL8PciWGTFYMDpD2wAEuB7acwtR9KBhLGwCTyxWobX2c/s5i
RcLqD6DhxSMCyNcmBFyZL3lwIO//mpyDGkjTDrsPQYaSxsVSX7qE7kh6zqZMAP1IwgObKEuDvm/B
ZfKJJwixdyyjNWyxO+XTQ66tBrLcR4EY/GjI27EE51p4itYSzDFxRGhUXOcQs7rC6euYPqLOuhVw
aPDQRZTpS7Iio/WqF9HxLp1AvWP9D8DoJAQ7v8TAKGltID4M5aPljOALKyorhB9kcLbuJJx1B4LF
Vxy9mfAoD3nd33EiXnygrEx/xzU+KaYxHOOHnefbsxcc053IeWtI8H1NK4PoDDYx6WVHXDjBtetH
p0//ZDEX1X4bDv/jFgIG/A8peP5HvEam51ic3IfoVKpMnqsB2ryO+enaWTMwF17kEyR8N5ZS826g
YBvVNzv167QMUvCac1+sIg+8p7rC2051eXbU0vdlfs+sF1WbV2KTCrWE/VZzGCFUafj7+6EnGsTR
TJdFiurygtHh5LWxITzvDuge+V8jOaHUJKtv+AMjTERsaaJIh4B8PeDUeUGwxziaMHmYSI9nWx43
0N10I8AMoYdGX1pJLk1eAvK+Q8yaRhhuLnAjwvWcofSMMyRuWJKdh6MNjjKEv1oaIEZ81iOBjN7z
eg/THr5TnxotecPZ67GwMSnVISfUj0sXSE9U0XOTCEcEdhohRuryxf5ObtSShDkp1hHj/Y5In1u1
3kWwyLP29mOW54YzG2wlmmTj01KA4bWF+Kub/NHbvCmPiM/gLUmE1EMJDwpxjGrBOxCp/gwPXO/N
C/r7mq9w/+5BXdHyTxCpXytJ9i82o80vpNaXMaMhYjp2eDKXlzwy7KAjNQ8W/tRRY8f5AB/dE9zn
r3eq9zS3n5vkp4aNSduOGFE194lGA7Zw5SKbsuMr28b+sdjwfWRmlLQuLttMTW890YWJkmOI08Ev
2FyPDIj+5T1jcEq/jERsHqaQ8GumI78Oj/LhBfn3KkZpMMw/bY0WzM7lx48ZwBkDuR4XPWcN7U26
Vge25QP7RfgeTeHeTV2U1IioWG9kvjdxxMTc1UHGwdVL8qngz5S8Py+6rSN4cn+nou5T4T3r/4Be
pLBRMon0dUf/JF2ljQttyJD4qvrpFbfjdljuUKLBOjIQ3kDZID9hUIIYz+sQAahHAyXP2MmMY7JI
RGhim95Fr9ybHJScGBN8Ar8bSP52eqfKeT9BZ7+hyDyMIBBT978Bd7bDwKSjXPge3b6rvZ0CnBCe
K9YBCvSXqX9hDVGhmN2EmUMhswQvChQYFzpeg3FJK7jvv/vtdYr1Ek5b2lImjym/JX07V5LDhUhd
wK5oPHxjnyomEGmqdchYzFJlBc4wEDF84wT2RGRLBKz7RX1Wn98KawoY+Nj8jQQ7gLJPx9yjXWP+
9yi5nt0rFqnOqWFgpUazqeJ5zBWSDwCRrLKCmFebzvkuM8V7Xwz/mjMAOBJzuIcoC/WLZlMWkkgq
B8g2cVo1hahuDfZsCbazkfPh0Dyx3zvjk6wdU5GbN4T6IoyWEaY5IQ73Skug06gIlMaJh21beNNZ
NhfbLb1cD4ZNXdJGs/ozZxT98zuNSbos5n/cXqEeAfRe5O19aeR4Icd8ozgrASNrJPT3/KTJV1iN
3suOuupFSDfBG5k/zWVveN83p3ng9z4S8LUAGj0BFQHB1uygdekuzl1GU+WApqAZPvMJ9k9Aw6M+
cUbFPxBr1EzHJyluieaMyYggITKIEm70qyHF0GysVDIrCxo9f3Dzn4bvrqgnUjYQnn3+m9a7JvT7
WlrdTfOs1pVRbt9y3jHgn7lMS9tpe5ObK90xfRG5WqAiMNLMhDPQ2tMiAcrXBn6ID5n+9rJ/921/
1S7JpgEOsB5zRVcG/6O/2WN+mPAAIII1NJnHUaUmNkrXsRGt+iJSnQ+Hn4WK29eQJ7xhD2149XyA
uRkReWfOvJIv0NNeysT5cNplOd7Ns5daUpOHqIRgzfDHZ5bMLvS50qyr9GxTZWLnyTknLcff/x70
XdHXHpvy632WhsO3pDiF8WGTXvURyPE8mf0/Z0S6GSPeG/gBPTulFPrGCRsJUlqBRCOyVlquwRJb
a1hwGfUOXMSQmSl9QYcKDHT69+G0NU6qR03DImx5nSBQ8PlEcEstrMpIvKPOejyAeWnanIwKFFMf
cKYAItXMn2VwUvry/QBI7XzjnxtNjmCdcTmeDNj0qsJVL7xeaZKZ14kwVGb3VRiULI8YHZQlT9oX
B5Gg0a744O4DW5NJakU2Jd9Wp5bdB0AN2fJCWwWCCBmtLM6vrE0ELuwe+OR8JE1FJr7Urs/LeRWX
gLGpPRtCo7yNhgw9GVUKJBeNFZ3F38MhYwyHpqvdE0eHVfCGPOj7g/o8onTlA8ZtCR5NCJ67XAex
TlnpmH5KgvnMBUH8lCl/u9YZb0KHKMkFQ8F0yXPjO1MhZtuWnbqCrrWiM8BuLM3PCfNpphPmw/C1
vf5yKKrz23zJwCpWkdSW9VrIfsLsSgTI3bRi2S7KJ5o+JHbSyjhI2a4lcbwuorJgf4HCJHDBSp3F
Mdaec0MTjIplGvm7hj+p9+eyNCCfERJfSPkYSm+sU6BLk3gJtpqMGYaQatwZK64mEv7SdUox8OCz
cS0QKycEFNjhIHovKAI5OcL47hrUvbZsWG2dpzC0GKQgdznEIWVNJQyBKLP/I5SSWQnRORFnbxwj
lO6mb2r7cdn1Z79swhgSR+Gyrm0eTwrAco/80GdSGVeZ+3osCp1+AFbBkAKtXlchPQ7kABCTIA6C
2d7tKMbaZKqUIr4sf/Xgt/0JIVV+rYZv3Hw3D2xITeBlyU11u56c/Eaufkh4+XJbdPz0BjyazEVA
c0PgZIPXOnYm0jvHTjF7Nql43uVhECXuJvCamlkpBcuMaKanYiSOqVO9O5LeNejxPz4fZAvdisjN
jUjZsMcdiXh+bHT0M2LXk3Arjt0Kqg5qfnRZiDDn+4O9XBvhDemfjZxkNFhuTPhl/8y6i7wKUSK8
NtNCAVcaeXKUEy5vgy/5gUaqbARKXLcOA0VgxhxCWvIYD5WgTUxRrYUu3n7NzGSK4UqKIFGX4ep1
E9vGwEBSnEHxIMdUpICzQDMX3fkmYlbys40VmkG/6IsrD5a2ds87F3jaTncFXgOFcAYBzHS4wa2s
EXBV7zjMlMd7wflXADcTbpI22GUHr1Kp8oWPzypojtQa+APD2oS5Z417cCCixstLXh/0ebhe6MH7
vvPDZvftT1F3gfCw+Q+vFtt0G+02eaczBqDtgKtPXzTdl+QoltpSl1yoyD+YufFkWY18YeLkWnyX
qqiW0JAvZ1Gask/i2NbJrLZl7IRw87YsA5qauf9/NgAACDSOD1WC6f2qkqpSsNNj8EV7AbBaxdb9
wNoQGWafYVmmfTgxfLRMum5qiUaJvnX5Bz8Vm/4N/K5y82XRaSwXvVG7bWj23Jgv+GiX1a5bLk19
1c8irZLuYKOa5y68Y/v5TIH0NgKgCmA0uodJD/Nzwv+GLtMVPhbb1kOW2uSCJR32joMU48iG3C8P
m9PvySrU6xRzVP/psSM0qT7QRqUkgEumo5p6TqFmKD0SKto4v9c0WH8SBG6Kwq6v0ioy2840H7Ai
jz+1Kr/TWKHvAaru94ImnIBgHHGJGuLlzqaWZIC36VF2pckaZcOSD4WrQDN/Fau52Hg5mLoOTkzG
O/ptw6gCEHkVmmwxoKrjV8lnow2NIxJvsdNPndEzKCjgG339gXk/PWHMvMOohVBvs5CBZpn2VTs0
8OwXyVtRa4zkwvM48Q0KMcBxswS1nv49Ko8sIU4BqEWY+iDgG+w9eRSibdksmq4bLsGHnzA4f2Yz
dqlWyjVhY/+0SQRPlm45PibMX7Q4hMxuTUWuumYi8/FO2wR66LSqFszlQvNiueLaWlRIigrS/mls
l1Ulo9Hz5QcpJ8nc8lg6hNY5jTSf3jonuXKk42qU8ClLW19ZW9egXW9tqS2Cc2CX6YYerwyWOidr
8g4DvH9RtDHds8txvGQjP+C5s1fp9b8i/d/xGnckyyrnWBQ42wHusj6TYT70NaDYKpqq2QQo1EZ6
b9A1EwORe7eMaLdQWLJyV/5Y5hopmBoAIdrDFXGK1EvP/QL/HMjgZKbwYA9rPW5iVD4ViuCgYuMg
TS94ksNHtCoGGNUXlA8tB9DfOFvHspr7ubn/oyxSwk/GFO9FR60ax6XMa6WIbPwuczNHEMA7goBU
0mRun05mWf5UPfZqWLNc4PXcZ2yw9ycTTcZGjRoRVNn27kC6AKN4Xt/j3JIjRmG1KD+SOBmYKxdU
UeVAgn2MrMbZNvI7vK60XosTp4RmLQ1JYV+bIXBaIuTAp+ycVj5OqTlmYPt5vNi/Q7d5h7y3/JIv
0kD8ozR/QrXkJyiJJHkPq0gXD3wqsRX0dCh2jH663sW53kImhMXgdPkCHeJSIMHyqqeKU/TLGU6X
3kx9e15IR0V2Ni/uNqN0KKvtbNZwAl1l00hNs9liPz/dzEMXvb5TED+ekO4Vg8D+wlAuBbXpT6OH
3c/Y6J4Y7LOaSTB78Kku+/VWO52bVFVvgmaYTigIS/ixhSNr23X8lnIVv6KXuEzMSPoCZm5m5OLh
QHsViYNmzDgk71OhOCHloygjZER7Qg5ewrfow5Mtr+iUSoHBLixqk3sDT8RylkdvsFyEBcaFIYk0
jUW8BvOjTpWfH+ANaEPcP1e5u94xoH2HEpFgxX2qFIdSNit5qHaPUWFQiEIxg2IGiN2YQ1jiKPFl
L4A6PaX9fCZeAO2eIr1l0RwsLNEZUanVuqsxsdyjgqpOIE7y3a1d1C6/R9/x3Zr+WJU25miNEOGV
QRTZKxFx3ykjohpMW0zwc7eDOufW09f7vvjvsKJmtCVH0cpu3L4fTUSUEm3IcOKqYY/VX503tvNa
BkwRT9FtoHwxh53K93OhE8CDoF/G7/WYIyG5b0ffhOdSxq0CtHOiJZUSe4paQZIAGIVRdoVQoEUR
7HSnVFc6U5cjE1C8HrrlDryhthEUxL966Pi7zhm/DWiUtQI9VX5JSf5vxr2QPcD89tepMt8sqNT/
xQRqmOlDmEDnLydyeAYCHGAqa3/PaBF1V+7bTU5EUVjcXVBUA0dQxU2nz3ovY5DS4Di6KR0Xvb1v
nNboGwSrkzzo1A39IBbI0RkpOjYGRNFelpkW29SrL+KuGatGTT43hw9hsKh8WbzdU8rp5jYMoQWO
ZQIdRqjggYINhRZJ49r5+6la0JXLUZkHyYCQGUtSGeDHos9lN/I7BBeuzWFsXc46iCasUcx1bpoZ
jslULZKwfT5uo4U0U8Dc+tdyG7Xkd+yR6SY4w0tXB07VDsZkXuSUNAmsll6WtRIHYiWobpjVrCjP
5vwGmve2Hcvt9prFYWLUhstvbfklIZRDjqgPdjS2hBpQ/ZnT7I7ovUXeASA8HyAWdpzSvkoyQyEv
gR3Qr8BTbM1lUmyxH2kl5AAWB/SvfeVIcicDrGy++D12DmJG+nGn3/4Uf1mMYFb3P/ZVjtJ0eppG
MTm85MvzQ27n48neRxhOo3CnnVMAm06xMAcxCb5fM1uAcRKOvgjwe0XO+q2ErFDSEm8JtiYXuLI2
R6IGHlOxE8ORNaIUp3siFYAcnHjPtXEkuQ24dDNtFXXcfDnrOnwDqKwtOqH7StR/FsNBcLhjnxeg
oMn6tz6vIfiqDwlBmMRpGq6lHPT2ZPJZD3MKUr/jMmpSBePTAW3bZY3M7CdA/ewwCVu5iuviia+1
o5f8vHOK/kIDFrVL6KgylyPDw3ZxdnF26uPO5glsj8W5P0rsOwY/ET7kXvqUhTZP4t9ewlNXHnMp
h3jKPw6Fp00X8LFmQ6BzIoIeRUOQRHSSoinmTV1mKP841w/kaeGC69cpCe70Ea5BF4e/eubagxCJ
7MMntxgxTVvgABAey/aYp8zBwFp6+ZaEFk4kY2HSDbQNHN0ggxmmcii4XLZAkWE2M6eGXQTq9yyb
219HQtYZwbUhQrpaWUJOrRmFQqCdMHy6+bUsm2zL4yjio4X/V1wQQE2RFWh92+X0UIeoNFY757n7
KD4dFce/pbWBSFwUe5i7JwaFRrqoyb296/I9x+gzpYgWJ253b9DQw1Ig54K/PiBQf+OgqH+jWoZp
CbK2dlR03YsKcqUTwT5hCDgGCgy/NvEIwml/BuvgUEQz1Mngq3TRcBLSdVgF6ei95ul3IBjul91o
jXjuwfW8tMGyfjP+8c2BqMRRpUwIbb+Zusa+XGGdbJJ9i5TJN9X0Jb/rTc31QIoVrp7nagwXn0xZ
zS3CrbpVw6KMO3fuKdMJVUAUiXetFdIld/IW1IlMV6tDVqz89b9qbxy50ZyP6+sk0DEqY6Wtx7ay
bKvU8OKV4Abk9H21/FpTrAyB6AEdrVr8xi/oOsDPArsfUjYBEoBLNSO5xDR8i59mrkCDXmw+wkuQ
v+sGvlcwt+Qu88G7ajZ/U0G/INCaNddewEdhDrI34+JkgISwU4KLgbesDkEGZxK3vDtpS15NE5J9
fwFtOW21hh7vn27+uUzQEjlJILorvpWDDDwxp1sUk+4nK5EiNkOYDGaQU0KG9EPIdbE1QHwykbO6
24Tibi/TawZlmYgnqQaQoQAddCUSUeqvDKwiJByd2+WmkIvFZIrbiEGHu6rw6wxX/MLR4LAM4Jw+
EUW28VDOvzdkF2+PC/L33XBwEUVH+opfP6Im4u10Aw0Xiipc1Dq4KUx/VawYzxdobPGZB1Je2LMK
M5u3oBtMU0kY9rNL6Itx/NobThTKPUjR7qP6aIR907fHUh2WGgYIx8SQ6Qk5lbBqsOsvtGFdQtrX
8Y/GGUbDhWGQFaYdLsgXBKevePjvNxBgbStMCUI/1rIkpfqyvO4OGYSIJGLYy91FuFlmGX8a8jp/
8a25j/ITQxfqzadw4BiHy1Y9oGiopLCJrteYJYQLq+f8EhaKgbvYkSk43cdDgjwVVe19s+8FJK3Y
MqKZOtojUifNYUUPmcN13ofwUZ4Z3ncX9E2ttyVbnCZuPaPV/R4yvbb+grU7AHXWhQuDOrtibbvu
XU1ncGeTTJwpyJ5NTKdGXn/IMtE/KzyCyPsn7VQViKEhW7cgWTKAva5YNhM1oEmpZ4KH8ECZJ5F6
Vs96e8rriobXw0NTMwKKm7TTDJYVEQnzXYfBSE5H70qtWAbXq8yY+gLWauh9EMyl1iQ0YCwD1VTJ
XGxm5C0y71vrU3jFEVQEqpRzBfs28B6TCLDGzO3AnMPHNl0m0S4Vgp4ts4b7B9Eqs8R4JwViAnfB
BCyd6ecOlKDcuYADO9whwWI3REuxOVLvkP13DNowpUNiQ/F2mYWa2fu/kXMvdtkoPG4yVr+12O6V
d2XLNeOz48LURJsuqcloOBjMQewSMwp6I30XcP3J2Yz9OGa61NsDPF1o+M258ox1LqlTtWIkAExU
XL6Fy08T8P+3I6mK9mKqWuO2WV9XmbMgZcCn7qtzz1wg98V1Xwk3vjDxw6LAY1cl32rnddJdEWev
D60CWuezn+Ek3Dpmq7qnYgXKpDIYrfXFMC3pTGATt47N1ViZVZxy7L1e+bu43JatzI0fL94PNtrR
gy+uWM0I+PoGh6qQHxBxJLehFSYocfNK5ZReQUjihnuxkwAwQ6qs+k4bL8luxIN2eI/yMokXuySa
UMfWvWh4lqkFpHzlP9Grcd+wkIchys17em8ZJeZoGwR81SYbyBoBlc37JhjTUjCdbf3byUwVQZu3
N2aVUxRFIeWHZcDmfNbKffiUEw3MBp6CHBg/GKfZJA6Wy9N3qRdJSrzy6zAllDC6Bz92bS7UY8T4
GyYjudrMrgkKFmDgDIlAo+lBbtJ0TFej7VZJ16I6t64JUxgIIU0fBq5HIiMrwwY5tjxNr2itI5fN
BvjJQshhoMhdaGqyU0RQ2yTmdn+x7Q0h5qNXOP8SxCwsaq/v88i2EAmr7g4BsFb1Y2BE/HsEYtdS
vA7u93XlohXMxsrCY0wZRkwmEK8h2e0/AHprOBP5/vQpko+Lz4cRIqzBNfwQHTZdES29C/iBcbnD
7bmDIjjezKhnTzK088ivtrHEpTiG84U4pSOgJChRLXNtZS8MNKMXqR0N6av9rpfkJMh5R7VqPybo
qSbs8h1pkE1KEilBcsb6SIubz7LvdW/PoQyL/7oRz021exJct8r/iAr9kK4WXJGP01ufZDNfDhfP
OQDFap1fhK75yyvp92tpTfll+nuXrspiQM6VrxBIpUHJjn3S+SOIFGNi/9u7R4C3yr08aWVN2CDA
nSiCciKA7BJld05fpMyKnKZ/oouVNl52hr77AugdauRT6KCuRmXT8qtH9smj3PaRgXfm53A/Rjhn
qIXAx5Othq2j0c401NK0DqWhh7txnl/4ZejqhUP1MwFOhy4hovtil2SXoPmzqB8zrN85bzjqmcKd
JspNzbw8nWh8ytTI0Xq0MukEGBZdh26gIGOBjkPPv1IH/9Ob3kUdKTMXCD7I4vlC+l46nTZUytpE
5WA1/2AP6JME9DGhlGexvvkY5R/SffK1o8YCSFK1mdOjfnjUuXa89vdgF5E+pgmrZpOSFBqhzZrs
ak8G8MYA5gWVHurCEobr2cJvd1heJT6OsDZbAvLE1RwBIb7K61keN11PAxlT9VmdX/RncbhcpgJ4
S/BKp/BGab17cggWgYB1FKl8dBBD2g8p5v1aPJYkdHzMd2bcWkekuHwPozguvxll1ELccPBqKTxn
3wjanO6dSOvR35PXmMnZOOVTkArFJveVH6/+AVVkmkM6rahu3ElgsrMgXfEnWMmprAZ++Ml5uxvv
1k4TKgXkCpv7j2zbHWy51PY3Zb1+z0yZ+h0K7A2BNpxpmwAeswieufbwYUyx2ogQjyiu4d5Kz7bO
3F+KBonZt4wC94IMlf/KLv3FzAQtzE+rBu4ef0aZGdqH5J1FqIsF5mmHTJOh9R72L2MobccAtFou
79rxLmM5XxWJcral5m9CWRRUggBYgKpTNJl6fy+e8xMoyUFIib429C8aY9sjIUSCDk9oHtSF83Xr
0Nmi3QPxwB2kwZgj8ajtZVHtxEY4QxdFxhfZP4KvDeAMW4bqj5nS9HYJ5ZSQ6aNNK8yQJuIXAiZ7
lkPpzDYGCVyXd0z2VjutnVjgsIKfB/hlCfZtPmSYBCXoyBg+USwZuvQeItZ+lprERUpiuIqkm6kI
HqsJ/22U9FlWFTHaMnoamzZisrcLTuLhZVESEY1sjxEuGstax6JxpaA6tB+dB+RkPPv1gQ2xszFy
pj5CgkHpgGyIiPLIWdSug465C5atrlK0GYMH/MR4hC2DLcocEtlMs1O7yXHCxIk1WPyksJkJrpBK
6foAZC+4Nsw1fNLTrIphzlxOZopPNisnqQR20yCiOSS0KZJhRw69dHMNxROOAo0tfd8iuMJzlwYp
z7NfiG8eEYlMWf6DmpkbF8veDO5LN+9OGy/54Mi8YJufRiX5eO4vLHLsBmKlOqPyMkchuLWcUYzn
1dLEJrNu1ZDNaKN7eV9Qqxsl/QfX366gfyvzZRHcQz+8TPmEjP5kok8E6ydPwd/kDHxNb7PtkRmT
0mxu3sPqriRyfRy0YXo+GqKaOKxZAbytzsFCAcKcc7Tc7I/6LxiSkMY/dZyUiNag1bHUNQj0Q27z
/5vva7m8cReKj7ptqYpOITlBODLV8N3dy084dwlSosaZjdLjt9fbM3wcWIFbXt83V6UEqCtizs07
Lwhabq3FJlc4jco5raH/DHax33glBOkapZSbqP2Bv/OnrpFKLg7IopEkMBLXlu3XJAAEqF3UilOg
hBf89/hR63DeeTJDdtsJd1sWjKxRCcc9vFPgXKZy6IZ/UCL85qcVR2FgMdS1z3fzjO4VJdUAycEP
/bzlu20aIcYXzJ6KPVNaahSooNp9T5Kj4hs6/P9YFlLvOp9maTJVaYy/8WkK3YGHL7tHMIRBvoVB
HlEQpCkpZaqrL3nzdPN7uqOs/Z6xRGOnoDltu277gZ9SJuKDW4XcwW2MXGoAsgT9qKI/NTVVWZVA
NnaKkXLMKiVRvV4iK1sYPxccmzspgUaVrU7kkUsnE80ZHI6qk/kMzUPzVyG3/mr40tzm0XJ/+w2N
f/jHPmeOjtiwZk8Eps3zBiJwqz4MAbq4bvij507giv7CCd9OjEiS1yaCnwzvhlkpIlIo9WiDXHhZ
OOrOlImnuCHnT1fyN4vNS/uvt9/rzozM8zzZzMkD/ucodRGhA1WJQ1q9pUyqBeqJK7EXF86x6kDB
l5r+RTjVTLbKromxNr4Pd04ne4c5HO9c+VRQ/ZhvrKN56H71T2pmT7sDY/jEORm2YJm3us4m57Au
aSe/yvBTgWuPOJqcFPubxKraM855G04FDSCj6lCDP9G+1+8As3ITYlnYhJlIXOWugqGmlWm2ECff
Xm0ENNr9L5vsTx9Fo9TQ1kk5s1xB3PygRovV74yD8MZqhl8FHK1w/OfoO1uOjpSfFewnbBv8aHx7
XHsNPZtpB+EKIzbzCJgrZldb19/3Cekw2tqW3lPYVKnrAv13h15bzDL0lBAlAbhEzZRJbDGPU6k/
lmFdQ3zNqCFSjNJV80WMaiaKth2MyJ79n6S6xd96thhKLCoTE0cS3OZAwX5W7sq1mq3r4yZhJd+Y
pg6q03SUWPrpLxqaaaRgSL93ISIa+O3sdsiDzrDBV6cI0xQaJ12mGCym3HgZaAlHQI3WaGltIERb
kPdZSCnDr+uAbJGWiFMwXZhOTJSdk74V2uAEvOTFyOOJ/bByc3Bdvl8BoDd0F/nwzi0T8g94M5tz
skbTlkkl6ankTLKmO3In1v0tt7oiu6K3IkpvghwmyWs5mRr4qtg/5zL1nMCGDYtJTNuHG7F8q8r+
U04P5BJkwjMkV2T6giDZ1WLl1pmCyxO2cp+/xteg48VVX/Un/f9AF/P4xs5WC3+Qn1Q4hCv2tmmE
0Cd6ZQclL0CTGsMM0fTGmpi6X2MPRyD0SibuE8Q3DhUuFoWpi8LpUT0QSjGYR08lmorFMP3dzS/k
pB7hK0TBBg+btuUXR4w1PR7PmayXNzEYLGaU+ryWiJa+DKiQAJoNtjglov5ELHuOe5k5BuZp4g+4
klXuSjtGh+PyCukG2dYtotlflRo2mmN0CmsyI3C61d7DoaAQTGQaC+x02xUd6d55n2+42soyh3lu
Hjlu8i9dK3cGx9H3osLjYB2L8WhqJ66Eo6xNTCpXjKsZibTKMC7NXCLWTKEnG2EtznU3HqKt6y+1
j8Xxk0RLx4n70AwFaXxA9b4Bvc1t7Rw8wRZaYg16Nc5XZhHNy1dnqkQn/PLPWIeWhK1ABGfRbjTN
+jOowRNH2TFCMSO54Mmh9twfvnqqDE+JPYQmJuWC1kK5b6fLFZ+wH4nsXh2QKKOGkk3p7B4skkDZ
GSifWZdfI0tajI/kUYrN6rfNWPsL15G01SMgFWS1JbkAiJpzvp3xcy+IysUVNtJi+reNTmhQlzS3
sY4X8TIDKCdFLqx6S/wR8Cvks9Up5GcR/W2Bpja/lNxnuYMbja9f6rQVlcSXZBfeKPKZewTsFlhP
YPC091t0fIkdgoU5Xjph298Dv9Fe9QCSOiMhWTFoEs0i/9waghOCCwwfNZw5oFHVZoRY/YPJ/OIW
FBITMYkWHz1p3DWe7UjgMUZMJoV9MLWhsdXiY/uTn3sKea1SfptsSbwPyDT8bKDSw2DBIC20dC/x
I3pskJ7k3Qgp9JfI60kN6hpcd0P7VyUH+Bf8dn/4YMSGmzyB0APhxki1EqUxLVwpVKmwpImhhEAP
p5l73j2wzvT5Z22+BsniE809uG0paYzQsmUFP+oNpn0A+ConzecmE8Xv3FIWsbWQGL9CHD/hBr58
SRFn1jhVDZjv9uUnCc9Qg0aBx2uOUA7zojo9rIpu0Rs283FNpPyFcClREX6rLdTibpOdM4ZSFi8x
Zhc6YVcrvyQkgCqS24ZnzxCzTbDWddlzqcS7paAs8IyKDDnHgdrALI4EBF4wB/0WlgamPQBK+vN7
iLc0X14hR+Qd+rvpVUiaOoNqDcZECdADzFxVePJpMT+6n7ehqzhq+DuYHh5GkhZeI5+LVcKesqjo
r7bzWBJL9x8dwfT/iWMpPMdxO/0SlNVh42kyg7k5IUsjdkfII2nvf4EH+Ksya1DzMElmVku9C5/K
OojKvzBhWX9ejSnjo25EzzGicdYWdzdhq0NFfj4Qvmo9jX9P4xFyax9/9hgdvAoLl6lYyOdepL55
73/i7GKdpkMC064UHRUnO83TyiHf8OcB6DoZzX5RhRswrAulIhA+wfUjOCDLJoH/Dr7f67fH/4Oo
xgsVRMMb8MWVCHKDf4zaZkENVM3ZW2YJ+vR15BX5WLPWIeAr4KzDGQKBwUXyhqsolFiDYgFEs/eD
IdrHnlzEAIOEAjneeoxuAn085xAJlpRBk/dYlQ6PiOF7g47x9vNVLG/nvZJxaVRD3nbndpSV1+bK
T4uWST5pATOZn2ijs9NA0VSV078XPv7sldDxGbbegpkWDZ2n2UKE5NiBfjoveCfwg6ny7jG33e5j
fCHIA6qRTHXxumsKzWZPoM06HSlD3pvpR/JH2yxdFImCEZHG1bf8XZo8MvWbDoLxnTOczWbR5U8a
UVg69KhvlqCtJqxIA+fkEnxx05agzm9LxChjy9mFvzyCqquYw/jHIOZKM4ZxEafLwL7W2XK/QoDx
VGZ/69aHjbvDxBuDCFV37+kBhYmJ5+ogvZaBL/Ot6ljeDHFdL12Br3xb4AJPAxOvr3YXyY5GtCLy
zkF/eqxSR0J7QT97Sy/bjelYyV/gdZuIbpNH4quLBw5aSUcTNVXMZvY9dSIhwHBQUOccZgGW3s0U
kU6sQdgJWUWz5h/0+croj4Fm05WQBH9/XSb+nHxZrrnjQ5CmrVSSifW4VNBbOnE4qsjMVNahkyAG
2UIJTdX2qp7GaqKe9HP4hra6eX5kr3eukJC44wkb+unLhmPISvyGscAeFV2CxjVPBRzAmIblTSyx
JvnCffn+cd6ObbiYgpXOECUNsjpCDpTJbWKAXVCtf1WV0q1rI3G4hELPRcq6VMYxP2kXxyiZDawp
bD89FqxfKPjpY9cVUplaOUYTej0InkoVpw0PjlZR/pdU1SgEfAok0NzZq4WKN6tg9PSMzsCO+YdF
2nYsfJ4S70jpTzLIQwvpuxm33Rg7jaafFjgSpkKhk07r9vk7ooBOk747nSFEvQKntc7XzcxkJB5y
/pJS6EqMWPP9QWSK+tFsRA0K/myaR4SSUhwS2R3cB44PsrC5Wsc8TiiFD6ojXbhJJFxeq/R0exka
IZXOZfM1XuT6YfSgGRkv4t82v9RG3ZrEWRrvqiQ1TqFs1BIwslshNUxUzu5w6jI8Tfb0RNs3Xf8v
gJM+6HXqqCP5oBT/KPiXk2bw+Jdt4tdxkx+nEEP0vCmj8iSKc1N8ciUrmVnNhZSajhOB3rkjfLZS
gHkl7UuHL08Y96a99dFqf43vgKf0d73OCBmkcUwVnfdVAKOWiZ8Gupf8digbV1kKIE98fFmhd6EL
ml++xQeevas3WiDlkddK3UzZAve4Zn32TT67YSOaFU8Q69eL69LN5DA2Y90lKdf9aAps1A1Cp+FJ
nzrU4imbTicfJjLwPEG0nqrnLEf8jccyNk2Blb1NvkCaxaZXJYdmLrVLozRjjHA0koFjnC+XuPQw
sSEKALGH44u620l4zPJ9NagZpx7VLbHx3TJvE2SChH4r5J/u2qLfrCBUuNo5kEEdg/RTxkkwwcnf
EJx7btoQgUmOg4/qpzm/TvimzqpSQS/tIK7NjtuRrSU1xnceR7h5HWEOUV0wBQo0vqlzSX3iDg37
QmDxOnm2/ipmXyNBSbTpAl2zUAtxr/0T32AEIwonQAJ47UKS09Dj3y/iIE2+2M+zGEAY05qiWOvG
5aLNMIwHOmnmn9u7rUayGfxBd06kERa0r9aFykheg5yPYudE9EiUUEIu5KIFUFU553iefqAI04z3
DH/+E3A+I30Jo4HbjZQ/ab7Tb8HV4OpDMnvreA373fg6tuW6gdYptm0I5oytM7mTs/kY+N1GDinu
Cnh+SSMGtuxKGfku1kPH7eMRyrohxRWvHEY3837YjtBx4XLto+5lKihOi+1P9U7ZOfPsZ4xnYCbq
SXUwdlW1XUY7iBHm45HPjaSVmCO8uPSS9Ca8b90XjrX3WMaI4/28t1AqMq5ABmTFvnucHzidXdD6
KViK4vo1VZa0cS/AtjKSF17t6NZaqt19sMegQHuSw6Bw8R/lwBYU/Oo5ABF1zPc4nKhG4UwCHjF9
8p1fdVVSvfVDQq7+HMzrLiJ3NWKmAwAglMrOXe9KEAVNKFqMVOz5J2Gn24aOeW6Qetnw5NGljTxt
XkRvXjphrIA6E4ZXBTwheDa15jJ9giQiUTJTgyArqu/URZxs/qMJ6eqe+cVuOqw/D554DhGEhVI3
+91Y6T8WnPwgp5MoZYC4zJO7B9CP0sg2fWH7otRun9obra8ehWhmE1b2Xt7fOogNfkc8KQbc2Yw4
CYoKugb/9S66DDKtI6+RKtpbyG4CMwFrMyBiQcbeHvZu29wtpTnyu21PlpCZJr5a8SzErPQQojHm
/Asc0r6TQjiWn74vVfzEArw2JTWKfyYHXxvt4AB/Ltm0dGaU2OAXY5TQfpaIDvrjiJS+tqDZej9W
MclsL6ppSx0nc+gnY9suCFgp7geq4QP/R+d4dylSyPIgk2tLVOigyyywYRe1VZfseOvxzUBhga4W
qj60c+VtrFq6OS61xdTy3C+pcN5q6lO09LtNXtv946M9Fd++Tl60K00r9hO5vYQW5XbKrw/0yH8G
qB0tmV8JegExGD8j7zNELiMJjZiKxoJvmpX0CUIwQpoaaQAEuIEWs4Ndu06+nN1fdUf4eIK3E+tJ
iPbNEgKFkdCtY38agU6ifI3zM0068MRsyuISFhvu/DPJPDSe7E19dIz6ojBX4RUdlwlh5u0n6tSX
xh848kHxQS0CHLa2/kqvtxjmGiUaQbbK9HZ3bP1QniEM2DIVmvTeWLfE6uGdWvOeU43OOBgY3Vk/
Nf+dXqhpCIYNlpcGXXE8QBm4PTXaJV2m6UKqhb4t3Mf5ksGL+CtVB8CZaq8lgftuxPRaGUV76pR0
fhVfgcgM7ohd7PlOufL4QMYM03ReGd6jA0NSYGNPjDolW6IrQUOFfS3QJVMV+FevAfKBbdkkmeEW
BIbGVe3qFaknDBoMTuW5pZkIDWXOTSuJHBN20mkNdY/e8rWWJbrf4fJNqtFKQGnadsaJzgy11mZB
r7qPYEqS4ryCmTzk86wFnY/CRrUsZGxIL9R3ExqzCaskqC7kuBiFM5azjRfRBk1xs3I63ARFDXzu
9BlLflGL0TQA63DfkX62A5FLADi8L+kI0Et7UlCULlZpxyQv4XEHazfXaGWRnTDlbm3eJR02iOQb
sHeRWuYrsOwtJk17F4iZswmlmZOaJRw8aHRVLYhDDJOPqL/b20dd3i+4s5dcOzPf3VzoSxii0JhI
8dVYnKck0x8eICc1df4/Aml0DVzsxxdizq2KB0cYae9AN+jrU+EST5zwCp2Gl9VVuH7eGToGLmSn
XmjMEXx6IGXEDj0jS3uZtLJuxd49vYsKW3cEadJ7jOyZF8r2LXHWO8cldglMo4Ka1MBD4H2yQKZz
WitwK1m/taI8zyAoGEEM0ZtQvCRwL1EoCyulR5T87WqyhLM/7Khb/B8T2676y86q363U5Slh36wM
1mUPQItwXXdgU8jSJMGEX/No5RgvWzi/C+avgvSXT4BP5pVpa+KfzPv428NqRioKtzD/dNXcRiyo
Vw92VM5So8UchzJ9REfRoBvyatvLiU+Tzg9vaOF4X72rCYEIzDuk/JGCXnXDdM4rolgwBjwmZZCu
UUO3oo1krZrrr2AEAoCaquXYttn1H52rpD8TMlwY5mp7d0o2uEf7w+XSCJA038YYTqD3xv2O6Zza
xC2bT3l/AiZFgGvXvy5HBiHaANYo/Cz9XwphDYjzp3CyyEgVSGq3gSy9U0+0W/gOHJxf66ZADfFr
LAegmxbkmJuK2RZpn8Oa/hBcLfTNr9ByCB6272AXfaFuBOhoviccmxi0JpmRQvXHWGGP+8l2oqBi
9U2mycsVaxr8y0LoaBDppvPbOawqkDmYWl6gVquIsoTDG5d1QV0seEIcd3xgJjp8lI5AfDkruPfE
7wlbiRVc0DYBna0XuXF5Fg1F8TjNcmzWbVcawPPKJ1pDhTAH+tGdIbhA5SPNJKNn+hy+cLLcTaEU
kge8CdXJItyZ3GuzQgjl1/+BIv0Mh+Rs/pGM1Aa6ahdJQsyJIW+DDsgvG/TIl4qiRJlCa/nCK3+J
6MFqBgvo51WgIpmUrM7urD+ePYYucJpuuM4OyJLx1tDq9OL6xDCCrPWbmJay/vcrgoDKBuEITwYa
IRrgk4n2DwfCXuEbJjJLvC/wF2q0xeDjgdEz1c+q7oXp71OvgvfOoZ/55UJ9j5B84NSnILuJz3qN
roek2yAwS8B/xoAMDV6g5pTUvqN3OzLEO4qsvhYgNfth4kQfM6gt4B+lROqfAo7oc8yprvoFAH3K
wgfgLYTZGCT0nEvKUMjQv1NSSFvrZHWDk+A8EiDZWH3MsTZ91foENSHkHwdqc7CA5e+0LY/nLkYB
bqYPz88xsWojbnVBJ7wpenFcaHNh5wnS7UUTxY+Y1Per16rS85GezTQkHvHT9AgKS6wlW9C0x9pC
kc0vfr1pKeUZ01XAaBwDKmfsgxVLrktOeV838dEG2K2Ctxep47zsivCXuZg9PihvLMOzm4lbMeer
xb9a5bOSMX6d2oR+E6L97vFC9e4E2twL9JxgPe8hovmUivp91R4Hil6uxe3JYHpqSS8cWNTyiaVa
UiREzcn5HbDnEArXsvPy9CBPOfpOtMiRHfOl2Ur0K5mZ2BfaPFLqMjbUk+sgCULmLfv3hXKWCW5n
hdpU9IsXEt9b4/SY8Ojwsx7I1Rkg+c1YK7945aqTtxouLlZMpYzc211+4mmIv0MB5oHoWziA6nT8
Xrfi94TfOCqY5Xw9TYmmcAtebxUgZWb0jyOhfNUN8YSmK8mR6PxDRI637ZZ1cCNVTIsURWJphKH2
tk1SpmmZAnq209xJ/N+fUOB/DUrf2x1YtlTOqOStpMFggrel5eZDtveq+wGzX6YCfSOMjZaMxA9U
0k46BcVWCzyENZSdkoM2NmCgMlPKp74bWv0PXnDORqs5fSAPB3R5i/at21ptLvcUWAR/iwc5m4NF
rKhF8Dgz8j8wJI5eiT+Kq6PrBgT1vN03k/5a2Xl/TC/UL5CCo/4QFMIKTr/5xSWzj2NAGWgQKFUF
xwTk0rYfoYjzVsJLaWxzzhRuRZiCt9nv+MJK9W5b3Ea49HqProSBo6pWVMxHB9K4zQHq1lfTXzlZ
7uqd98yz/vD4NktvCljfyfbtOAuOdbAfzoYxY5dUZ6Fx45E9KD3b9TKDWTjxm61Gv+CCf2p9CAvv
nBN++v+6q1UVw6DEhOJYPmNgUNr6rRQt+uQjhBKC+RL7GBY3ncD2rF04NfpUgTw4dgmrn+PRwTYu
eOWgdx9/+TLfz3AWKMJVEa4+HM7DZUZBFiLwyTFJWp61fZWSFp1UfoQgWzRXJGSe/p4OV3gTQcIl
VPN5DaIo0BthxTw21CFouUdBZJm6xGgNqIU7pr94rl49XlKMvQGrK0oBzycpzOWGMfkKX/U2vGYl
T9/nWlPU4UpVUVRiMcFFdcvULgSVhCDjtYskSK/8m6ccFmAxZdcYkO+0Eqele8JYw22ee6jVhrn0
kIGXA0W+kxI1jNlRk3w3dxczRzmUymhF9juei+GIcvfnE9vLDgSLF46O3X4COxDaDCI9WS9EdrSL
tkznEoxVj7nhyzD5CaXGV6NFREkQnv8WKkIiXHamQaajVj8mRwMKofzLCh45Hwc0/7GTbD0zZgMg
GJA8hjyvAXJSrk0m+jB40wqKH1Ot9KLstNpLS5VfWo1GsHsXts4u2AzI0aP25nEHWeyZ3O/7GkLV
90gmcVEyHnRwXsyoTQYlnfxVCCgsDIU/ICi6HgO234e0B4pb1XsXp0w/Q1sm35CzxzwVolgQexNZ
us/81ChQcrRrirsjlU1IzsaqqUEWpHzpkKegpq0MlhgbWUUnhUAb7UK7P+JoiTkpLdBNvf9+Je/i
ISbQKkhrTlZjO6cFUdxzKn9727ZctEkaZxf2XLl8bIHj+f7IYyGJmyl1fcTDCbCw95xD0l9HHHn8
ZlKfTp+cw1Trsvx03OXCw7VrpiN+bZUdOW0aN3e3Pd80yG7SEQSx74/yTsd9TcjE4qAAfO3sAAb6
i1YOrPw+17vKxUIKR9IA+pkUn60GYWq69FdOL6HsHy/bb8D+Q59kTMaTUMV57kil31r3s3ruERV4
MY6uiLxoYvm51r+tHPzQCm9VvG6JWZaSUO0TmHbOLNUifldJr0m4gpoDxbA1u2BN6Jswg12VtXri
T6B1qYFb5n156SO4K1PJZNx9vQT1i184DEDZqFQ89a7bHvBUipMysUQa6tNbsVqd+Nl9i2CKMNEp
SIe68/Bj7FnCjQmAr4/g8J8dAyVXRFqIxPigJixWtwXRerbBANPgra5QGO6jk2zj3Lo7fDjP4PAC
EHBdWzRyFnAMgId2q43VyztkHcbQO3Wq4IeEwEah6Cuf1C8BVfu9FD3eJXkE335XsvKhhSjVD3OQ
57AvlzAzBSwyZE4jfdjOhLR5/A0eGvzlZarGLZgtVgZDss1R0ZikzNw6LHhHJGcXzgG1ZfkDlAcx
MN086tBM6wRTwOTz4ENPBZUHnWRz/PpEZ0h2zcdH+NtBDKQXRFbnQkdq8uCSDmcYkVIp3ZBOMa1T
+R50ez8yhhyg6Q1rqsvwzrK3Jtqu+pF+qTUNQPo1wO9UHNOHf2nLi3iH+QGZsd5DLeaQrOaZV3SC
VWAaVK/8BsAbTvivs0pcp43qjctZ/GBddP33xgBStUXraPeutfE3LhmXcvF+p5oxiMqa93x+KbTo
gyZl/PviVsqsForiZ16Uu32+xV2KMli/jDeMUGxqetHBCOTpHD70TEsmtr+d7qvVkzzCRZBrqInK
tk7CZrs0IZIoI/DG5CJK1w83w2JJa2fQx3CLfnxUGhRX6nz9VB2FfJniXD+rPea7aQEzYmnLXvVi
aLstp2OkjBpMiX11e/HzpTf4jFTu5b2+kdI9Wm2otoKUEie7IOflZ3jkBiCkI7Y6tpK9HybM2pUn
HLKNeAxaeyTrRwVo5aAPScrLIPkycRjqkaLeygA1e0eHbtoAWyk1YXUcYCfEOsRWzJ7o4At11pa5
HKHreGkzxRx4ErzoyVr8Qr734Gv7H30CqvopOeajtu9drzAyFfh7/fGNm9zAALfy30M9bsvuR+Jb
8dwGS2ASDPrUcSpS1zzySIukxIBjQj1FDxzOp1lcdxN0gxYDSTmw4Csg7vKet/MsBvYiHG+tN3ET
Jvw60z3k51YlP5MR0oSr6Kc2WjB7SVbbXCcxkK2jEINWEjysEhZdvpolf7lhwbSCfkvp3uSEcuEd
pxAw7g73C0Ako/rJ7fqxebp6HnpZd6ggoEpM7BMc4KoEKF4XOosGn8gaLVJjStnUxKaHkLhZLhno
hOaXfVkXCC5DZu4uikZGxVeHO1wUb5HSvgLmfdRaf97DcaCVqXtWtRouK67XiW1xLnNV2UStItG7
keiWuxbnHWIHw6Pakv60d9grvPED7rCfcXnWryxMKlbPhCCOkc1/CLjzDthLN3gfagrzmYrcaom2
PErqProl4yKzEA+YKVmVADcxeFoguJvBryDj+9VMsal8crmJWr0yH4WFy/gaCUgrVZ/RPadDrAiz
3/6y74ZJv6/UGOQSqfE/fFsfyXoZsm2WoU0IFQDwKx96gUuyA9mMWM6AhYcxoXRAovKAizOdfEAR
DXbQ0x6r21JdpWOwPo+xXA/FRbboYaCs9n09XcXm/yPvjbjS/V1+JsCm3p/TS7jp1yHOQwZA1Ett
tWIoMl20PTV7OYHeuGtSgZTPC9ai4xo6XbWhMhIdZaUalZQMMftH0LA7vdJMVZKntZtq6sVxfBPR
hjm0A7QYbiYWS6/rAAFLjpUyO2Fu9Yauj/HtvNOUSogb58j0zE/yzBFLo+RKy5TL8X1X8blyyPts
R/g1VqLRpR7SoMDfAOuykBsLDa57cPVroczzUj8Dl/rTntgqsIrJRfEs4CGmTXiqVdGZi7MiLNcb
xdJatKZnvKKlzi87hjW/JGXSmC3IAQkHJHQ98r2GzbtEHWVPwE9PfWlM4p+zDn7BldB1Ln2171pT
tHbjEMMOtKj/pwGttKYkjClwLn4JEz09UBB7ZHaPdvNL0XLlNM+kobbTCPM9LzBEypDwNIdXYhHq
TXWE8BjNMRFbNK9l2G4KgB0AxHZjdUqJxA7PFtOlfTnvQ7wezQaZZ4Qmv8nIq70MYhxjajb7Nc5p
9gBso1DhagW4E+wG4yN6MLdLbC+4YbL6nA7xjWm+Z3twiXLYoQ9P4EzMPJFiwyiStMLCksfc1c10
94L/T9HXiBExCLQ4FzJtqvIRZUwLxHFKxJ2v7F1CsP/ljJpV4zta/IV+mz9T0rvlNZf+OzKQHNwh
fSnLpRhv+O+dIvssb8tYuZTNcGgfeQ7T58lj63OOZrM4RUdqHui3kh/KU8zdQCGIDVFApcOHb96X
sfTiQyV7uMWYwrCCZf+Vnz7pSxa8zDjrt5qoW88U3PfhzQBiWJhbqhwny9FLih7KcMEk3G53ld/8
7PawsEGcX/PdxWuKqmzWDFlyMTD9luwB0j9GljTLyHL4IR1vllswF5kC6Hv1GrDGPg4RR0lWrSqK
1sKA/V+amcHt/DyGHu2G/AGen1arrMZbhnUthuGdQ6Pp3Sdg6Wu8NViUMO53uYef/EXe+ntZHkwl
hDKTH93oKQ6AnmhCDcuyBzoxjkMZUneJnP6XvftfcdYEwYeAVsNHjbvVkfqPk/9tgc3TnGyIiAfI
pjNDR216W6X7yc5kubhM2nwb2S/Gvzoj3FepCRiDxD6psOYw9wePpVqGg5EbxyX9hi3X2OLXBV1t
6wAMreuJxJy8hct8ULtwF4M4CI93TqGRIMg5S0kmLtmcJO0GqYYziahrrPv28I2fh7komPyE7Twf
QPsTglNSOmOikx7n65l7xqhc+drQZCM6+f0DHVqH2meqWAHQhqWzToVPtzQbSwlSXY3AnHGJwD7c
VT8CJ4dB01KRTG6oM9F47m4W6hAulcqyJBTWmiM5StK889pHTgJgHpjiqUxa6Y06jKQjVDs1tJ4Z
dEYAUiZPhlQne24VDTbKUsXoX4sj1C2AQ/qRrcBw5dQl3JWd0WA9nZKiRwwrSDxNZTvtGAtxMo5x
Pqwk2ylipl9y+BDZpS7Ac8J9lkUTnhRyfujmFdiK3wWNbuZVJr9xahEb8K8OgTC7RvwPvifKndhq
MmlGd2qd5ijq+BDqueKrfHIiiLqK4jPEjsS5dF6vPWf4PAl/q4rKhCLY03Ef/3KWtNIJpvIokAsn
r/O+U9EEIWZggAnYqq1l9LGqyaO6WYEhMDcld0V/EIiLmqTPXoYiuCEe6VHlHuGEP4Cj/YeeLpr3
2qsYEhoJRDdIGXO7pcjENX0ME8B29rOLZO5BS0KfnHsZI4tnATqV4MUm/3ItAqzQM3i8s6aUXbvf
TknK/bdgbo1p8JHAlrA/9hu35mq7CMDgfqwngVQQImaKvHNai/Usrl485zTc3S1axJeMk93m7xdw
+STSEJ8Do8g/2LvAVpz3Ms0VcKz9iBFRhJPJEPLuahT/FIke/mP5dPT+8FkflRoGJIveJG4XGHtu
l1EEe+clMaO9xze/1jbIJs6OeKypqliWzyT2KNfjuY6nHKRBVDqKzvRCOBf1rnRLUR/wgjNqLchZ
XVtuR5OVBMCLjYWFDRuZI9tXZwxECIzWXqSf3VEkEPz5uj4ROuOx7TexE5Fg/JkQzE/Uerv8HZuU
OvHY0sTZG1T9/6vtV3VRS1tQ2uwwai3iBsM3DdDdZixfHLWQfNyEuBndfhqWieu+We5Ggvxbn2d5
QOSzLuZamTTQRe7oPsWhA1/Vo84njwrDnNY91Ssdsm1NrRTlPWcpr7+owsIH7wP+3SBx3qnYJ8Wx
ayCiDExcUyNSh9OKn+RTFvsYE4ucCgk1UE7dg3zYePlt103a0dVB/2OnCH0j6jn2av6IidrvZ7OY
IA2WKpJulxFWXJ2zBXGt65E9JHXXTyWbh5FTapKx5GiIHV5ETb/8FrrciWwT4qYXVPIoGDIzGVmh
6t19HYmPidlKRCPf65Y809MHFDKwIgbn/2nb513XBM8MPl6Y7XaHmeCAnYR+Smt23kKH4PzO/nWx
QeYURRUfYZczrtJnGhiF6xe9d56ZW1i8Uqv0BlwkYbZ4rSIw7Pa6ZgANlJp8sG9qj6S96hm/3WWa
8gKCB25kQzGicuBpjHVzo7uttTZYHEqFsPftW+ohE1WWY6IKc/7KTArCEfOA1NeEMdQaPUObtKFn
rYRM/LvoBFy8fRIRSg3QAy8W45vJDNjBh1n9ZANam26FVUVzQRlk/4L3xZiZ2vC5JWTMoxcBEB4y
fhStUN1BJQF4H7ROW9cJbaVKuA/w/zQzSRsa9T09fmMl44bBxMlBoEb5Mk0i3SYuzW62YakpqbKK
H8KZ2H45j5FZ67zLa9neE92BNFUd/r0AWHggOmJ3OqvehPFY8qsc60Hwas0+ZIhRTTSs/ieLX0j0
v0DFZHigsOl4tHn28qbkoGlA/8A5Hw6BP0KQsytMBCdEBjOfB/luoWMBf8r+wbmxlkjmQ58kU/xt
3stmH6ctewzPVREVvkGV/51Ikz/9KXuJVGfiCf8Z5eaCNcIxA3X3u6R6/X8/eNabb+vZpHITPdFb
VgE+kqAYNKnY3Ll38ZhrM47KSEDjQTKsw1yG53i/TLCJ+6Nxt/4EeSZfELAjwa1cRkQmTM39+teT
2Tuj+d/P88afjR+DFb2WcqxF7WHer29pv5PEqh10jsIDOsRZkZmm6uevqKJOYmZ6cRBfGqJpVKRp
8dGs4D+6GzraHSeKv2dEcdhWvEnEK9+kG8GzBNavFIGLwkq6EJMDlpR4jaPDLqvrcqg4sdI2yNSK
fevg+VgRDcPM83nSTNtsQQeDvOGctv+dN8BxttT3RquB5lcq3ztXg05sv4/9mfKmRGt4UuaCLFDN
7fJNBHxIvMp098QXfJe7KPCefqGI324xgeDaVdWUnsr97BwJKSaZlSh//SPKCFaAYclzLTmRP4Pd
02ERaH8SuS2A1p/Tex/4ZqTA6+VrpgzoYzOcteX5NcadRQ8e3mjEM2CojHdz0iAl4Z0B7EckgOfU
VEZjl4lqYo67gf76EuEVd6VrxpL56hN3PCSUMpKvc4RhoKh0Vp0Yr+9EoseSMCsVmBVSBB6zwWI0
QBhff6Gu6mafZlp4b7ccu/0I42u4RwMPfi1V0xj7XxU3Ch58nwocYVvwrg3anCTLtikp/Ega054r
rAfkkgs2XQo/usME1y4d+lwvEjDs2Um7Y5/GwcVa5xkBYhP1RZ5Tps2PkuLXWfidit33E+PYBc8v
pCh+eVVuHSCKAn4HgaaKSUhpEOaTEWoiHkzyFfDXqXWSYVGDQfze5L2/q+Qryn9l3pjsJV80fFRb
vF9rUtWV9ne2ICJ4XbPq16+dmzIEYR8Lb5G2oMwc2HqM74ouhYx/90d1LoGcxpUi4ul4SJ+5iE01
Re+Fw+kpIP/0kfayxN+4w/MTWS6kP/GT0+dHXbZ4/HQEH6xq/is8zYS2b0xj89MSEPKUg2Nr0HsS
ZVbP3k0hta4azGkNUWFHBsCfXwUtIQlgvF42GHpGgWX0Tj6BKwQdNXubERSdb+VjDJcU4cdA3ssH
MCHyrcUmbZ/J9ouBKzd9hSsll4t6jSVAA+69xd3FILWrwmgvbALErW5q/jQ5/t+p9VOd8Waf5Ddm
tYQGBDaFZqzTIzarztiyi+x/QNDBcCoIwi+tgHKI6rQGz+jNtcVIzqbCtnozQhEnSZu8OwKql/sE
ajeAZr/tbfHOyp3Lu50FC7BsPb+0kolQtH+EFSpDgiISeP+wjWkJE/gMcP+Stou8ZCOlI/DH0FfQ
htB7dEyqxsYCGOCRlU7nNc8TgiPv3o64FNkvbxZi2QXeD55L+TQXd7/PBHVwIebJUiyNJUtBD8KY
DIecVAC569fDLHR6NMdsn3YIhB5HOqxIAzSQYztBDqwN+1Ztfqv9Zu90XDf0tSW3VD1vh1R+0IL4
6/1suBpMtMYkpOWoiAMaKZaKmbFHVVOZ92JwQT6Zsyx4LgV27HdJ775/V4mufmWjHfw5jEvPNOSX
ojtVffYV9MHwu4al7MiZBqgNlNq3lxkERdGiXpQpWflzUsPuvxBhocUUI5dZSfAKjbl2hBDfGKpK
P8Fj0HPWUuPh6ukfeSX/m3hNZasZHa04vEx76uO6KMrQ+iA3V1I964j/MyxHdjiQOgmsr5fPATv6
ae3z36xehJp76v/uRIxOhWtiU2gqDitPCaTpdyo4XPpk63BuavP3atf12p2fPLLr4NskiKJJLeut
40jMLV8HbKzYFPnI2oNfWToE2zhCzscMVtj4yA6YSdwE7l8H615+K8RvKNHgZvOWhlu6zfqRGxyE
7SIqdrQWLc5F3GAxUvikS1pC18GEyGLWq8JwKwt5mqotIU42t1/wgJW+7rfpQ8xSkLsTR/DO360s
OZEKUrflNlKZ5p+qQ/R6B5ZRoyg9O+W8wqGMmWy4nWzdMZwZjp5GR3wqjH2dmWh00FrRcVVFL253
HVQKvFmxrNlpwuKL+xHlMXL+jH+YJKBUGD0F1VihOLsTssndDMNYJzA2s8Ag0LVKhbs2CuD730Y1
jK8k4izlTmt9MNUgIat/uRQPSM58HZAa1uYCXYqrlJtHTkW8OIoiHfBjDR4pEEuRebC/JoXIJrdo
bnsA160tBPD7etVt0hS8dPOMJ1N2OLiffKFYR7Og8QK1mq9GBK3av6ZKNarIa402Lq/iLtlwlcrQ
dvzWGaHc03cvz/20zLZ81+5DpM5B1H5jLiOHz+KR8gM5+QH2ius3D4C+j3F98dXqGoqka0dXTEx3
nX8pjUH2X/ny1qwklZrpsKHhwo1RXAs1crP/4AipD9TwV3+Ucti60QRI/0Kr73aUs3Kv1mWuHiis
tr3ypzsCaWR4YAjhYgSF/nkmazugdnH+X18p81T14kpWkGjFElSIODeO8E9On+g7sdOEv/QASPap
BDUZw8q+CMVXcAT/tJ7Q8DqyBLQRp5hn+1xdnD9Mp4V3LQmTB2Y7tQ+C2W+/sH0xmbD+RAj/bHt4
WXR0JL/TL0vAw529YWgAcIWxN3+grCEWv+dcm/DzCSlmh5DxkoP6aMw9gSS19d/Jp8O2zc21vO1A
dtWPyPNvFnB8S710gnmopZcpDV0aAFij1oYVEeLVfX+BnNgOyDdnQgdjJlea3aZiT9X8C0ju3/p0
73138x7ENhdQFtblck1rgKCO/9v5GdXADCyyjIll1vhf5HKC9NgF3X0YtGzqIfkpx8q/3QpaG5Kg
CsyhLKZZaxl11iBT7AUVSGI/Zhd/B4MQnPSu4ShinLBTMWlWkQ46qKPai/hNjLSic0pE4+9Zkr8c
O41WBA7BjxMsrobv5XxR89pcALYqgnaXl4VqFM8oNrqGXIc6tPk5adPmz5QWoedSbuxmodyua9De
yyeYEgRf41r+Yz7GbLJ7Zq98J9/xJfjm3r8CLETCTKF9KyfJpS2orRzxRF6R49k9NiHldp2CB+Ga
Payx4BDvo6zCQHmgEduF1otmv88OsPtnQ9yLucGuYA2Ed2h3uEdwP71USMJIYFuK526kMeYnn75K
DO3B+se5PXOcOJn34GFKSM4Kz4u62/+4i96enmTpkak6yky3SEuFl19ZuUYOajs1sFJlAtFJ9Ls0
HpYaLUH+7Jp/xrBWjVsY+n0fx0srgeUXM5d+9J4dch4a7agWbltlStmM3GSy0EJtWOqJmMoLyRjk
zmIzAIMHpLQcsusP0LR7s/v3WOzdghTQwzrDEIBBgoY2L7faZkM6UrgOceAJo5WlqDdK5HZF8t3I
Q9lI2HkunFnsOLVWaKt+TXe8Kg+gBLTAYM5u3wDDFz2sWIa/04YS5aoAvXRz4zIIw6sspxLEIoCM
54IMsZt7tz8nt/uFP1yow/7sV2q16lfXU13h42+UtbUMm6fz4/jMkhnAmpsboQOM7ul/0mPI2YEf
snPfhHOpETKphPiFpPmm+Hdu08CWdueMpDiEpwA87uBfa9i4V1JGKUtgxQZJXDZxQnOIbRNzsYRE
zY1rhDACkbE9cRN1cROAFBJg1cfqc4CHvnVCIeqVxJFBKl8FkzfuhsBoTiG2xuEFNsVBkONEICDp
KRTMAV2+Tyltr69zmQkBbAXfnj42XWhkEFKtEAxEBHroIOJ1LLVVE/weHlLBbsgGzxs1SU0d5BZS
DuOFVIjSE5WZkqPxpekmCIAVc613i5wFU5ybUgm+iiooWHFzZKH2TDLZDt91Qj/mlPQElri20jEc
15hFzq4xAFuzBLAS5hhN8avJrjryWvC7AN70uz9EHTSFG7S0fNfEl8OV00GMBxMXsqH8MKinkPrS
MYqj+BLvXCL8CZui2409XcacSIzhxYa6bVLmZafuj3u5lOp0+82M2xAhhBqqIil9YfX/9+qQr6vz
UWZGQ9l4yrNrzfXEOwRmkJTI0H/h5IWMT7XHY+G3bq5Y/evydum2U37Y+CN/wAvf0O3MtXNEBzpD
Aya756NlEO6rBgO74US2I9Eww13ldqGeGS03UPS2t9xwBGrCQRUV6nMLSYwr9JRlQq0Vg6JVD5Kz
pWR/tTykSTZzwYIWt/9awYVRhRk+5LiyQC/xFREjwUgXCYvz25XhZPGiMaOuSiWXzpqUmAt9Ta0M
Fb4v2mrkfldItCXAaiz8zees73VpBffjTmeTgmfrduvvbZ2vQi79W92B5AyhVyJBBIYR2CuIPbNv
zNe8n109hrGdVImuj2E//4bM9riE93S9cSq81zcpS/7W5bn63U8IdQOehZQCCw4pDo6I3SEywWxh
ZD+1x6M1jJgZNaF2NgxXqOyVo5o2RMVGEmHjVsEVEaHwDPWkkStZkEmr4bJttjUYd1mOBWgFcrQx
WfFVGUBjGWZ8zSEsmWXSvvpIPorkPekjb1uZZ0sIOfFEgDA/j15mkw2mRDEmN6Wna1j71bHsWWxL
K2h1uvcPc4eKcKX9GfoRUok3KhiGZ5LFdnKeZtfezf8BD6KvY2prZGj9iYPAWa4F9gLlhmJ5G8D5
Z2xJqhY47bow5dCdhQMsNKSvSOXBTRzfx6UKVDmcbOce/tW6vRUxOp59IGEBXMEWpzqY/oFYSo7U
u27OjNwexFUDHT+BbFDOVBr/yy7MfgLpf+tCfqVyKOR34x8KtaYFfxkBXLnEQsxhzIUiBHIIWctP
Xf+EvoUlw6Q0O+Cv93CJ43J7uKNQFzdTgBOWNrA7hBTDewiUK3SH1IPfMqKxQWfWSwkTe+KhdrXI
Z4uUlOGmc2L94BmZo/Vl7EAI4xf9XeLUxqG62HzzEwr0MX9t+or4oZfnC/Gk/MqtOLAU3K1A5Qom
oC/v9KryQojN/3l05qx/qv7OqBw4Y+4sQk6eMomJnrpzGlT3xyt7knsslXN6rFTvxm9hVnAbuA/d
wX5mo77XsMVf7FGZJu8b4ybWdMHQ8qIF/bRgG4ZwrOdLTbBEertT438nkvIkqK+/8U2d8IoyA4yM
BYGhcLAmcCW7ARABrGYYs15+LgO2RiwwH8zoMkIle7+XNbP3FepwwqGFZBxOT/SbqZdZ/3SdSq8X
Xu03wFPOiiJ7xfmTjnUWMntPxl9Mhj7FQV3EeDREJU/Z8TsdbagfV90un/vc0XJMCQpyCWM6S4Mb
918N/FNlbE88lBAnA2mjUpCHVadIqX5bT75mw9ip7aTOpzPjULiumZ2j3Heo3LGNCigWgQaRnEtp
2lqnTQ9/X3kLWpVfjVzRdJ2FXJO17pPR+w+gJLMhWsOun+DVqxmFeeR9MVg5wbo0bz5Cx4QOlHzp
J/1CMutLwmzZ6zN7IKYzNyLGygWODlSVZtx6Rf5zTTMKRQdi2op7r9+1jTOHDxSH1JGaT0rsTD8G
GccDeD16aLiwzBkH1WDtCdDaioimfTpQ9FwAKfn7fp1F0DTdCGbcF1wQR7+WArx+JVBTYwoHVDT6
hPxb01XXUWEljQWOJu95/oVINn0UWKVELDzxptD2JxE1h92UA3HFmDxJpmCKU2av5H0v7wwiJ/2C
W3SIzT6iIRg3MS3P7FLlymnaeYNnvUkoW4Bdcr9rWFq2PqtMIp+eMdVNqVXW7LSLgO5UVGAiIm0N
i/mRqKYH3Zm+4r3N2Jek5H4tZI0eCy+a8iEuKYE11ksEDKzzpCwAzCCYSBMVwn/Kc9WdnXWaNuDa
6XR80xmj8HQWMzy/PcKRia12ptX82DYPHMuYdLQ+3X743ngkJBX3EH1oQ3LP5dLWgd/295CpLHSq
tAi2Y0h57S1eyxKMkzXZdlUI+baHzuNeu9Y9aUfflscvQeru005W24xjqN9maVXVAI5/mu/T4QdP
dDn/cpzrar3lhwCi3V78JE678jsQLB7OKdVpDgY6ctugxE0TQMVsIJl/I9XWCDmpwe2Wtuv/KOcQ
R8Keyt30ks/xeeAFz3uXc5OBh1D0apE0h66rziDQ+YeUMJ2bGCIJopCHQ2M+p2dT5muwPMT2StG8
VJxxKnmWJunh/mW+rKc3EsgYK4w4IYMIb3ScJ/xS30MsytnW1eABWRihMW0OThNwhZ3Qpg1jYr9Y
uk4oMC7+Hsv4i6amplb8HIvo4Y+6VPm8xr7uCXQvSWY8loUqYZqDEE8ZgsN1A7OdXja65jgsraEI
fG3b2G7KTefh7rx0iR89GlqMq/vNoNSrSmhuuyBzK+tYRMUn6ByN3gp0rSWi5RoNXoonb/nHwgS1
6uHCXfeYDIVxu8kWTkYRveGcuz8aPsz1vQSXeq4AArjGeft9NxtvMrW95aaYgXgqdmx9NmWwxQ1M
D4iLH3SiGnosu5cNq73kVbvMOoN65QWa4jhPC4V/4QDbviFebMDmVCLlUKc0XD+ZIRJjk7bXX01T
yAmvrCwEq5kk/oPZ/mmkLVWN4ciUFX1BHzVRNlWLfneEgZC6/Fl0G6vI8yHlwiIKxzHKDx+88Au0
5vF52mHUUK8oChbg3gb+jWR7ut5xhXDMBza6Ys7GT1bzu+5bx4D0zw9BFl9ZBXlwyQIGAygorM8Y
LGYDsVyFdXrb4f7PFNljz9ZFN+jqkr7szfS9GHhFd2LmOCowf/IQPO8LLQz4Z1zNLwudRhnYZ2ha
AF96rz1AgM+ci6p+dGoB1sYtKCVM62crzv5u9esRM6s8QkXdS2xoLl3Nv43h8Bv8hcOblp2WbhPg
pctvV8RBRNxjZ6WjxQ/sL4cv88XqdxmjUbICYmq8IPJtkqWvnQz+0WnQHjmwjwWnOkfkUqDX31uD
tNSfzU2JBC0CpJF410ffoxuEYYH2fqpunaedaDI/YUO2Q6MpEHApUqQRT7LXxzBou9T32WVfBDNd
+3cO9YQ35Fy3vx+Cg1tb4+Io/GwGxMGmXl2HcVncIYU6knqCSQ9Rnxbo8kEMAik1B1iXMqJdw55o
SO6Noh0RYjfuMd0wBz9H5BHg0NbgGkVIZWCFrrwIrC910II+ieWuAqVjn4Tqdf80uGAy/Gfcepzf
jkb84gQXnMIzbLPvLxBMAUceoE8AGM1rPxXl55m8BFDoDMn7zj9utb2SxcwAn7PtLBSFM6sICsoT
9/AmZGI1G7YfuMu6stQ4NpSexcZOKsv0KCapeXwShdJM9WQlRyQhpX7wbcucuAVpSR+Ra9RY/WiI
oUmGdali7rKiji/d9ceko1SbugAfnPpbWXdd9HmnDoDuwfSg5vbj/mi510T6nH570+I49b3qqjBd
27Fcp/GwqlNoQEx+w3TAFtKhn8npk4/8SlFTgyqPnVM6RfDiKad9zEJkHgBN9yFDGD/RVuEckU2P
iAS8pEY1uXMvwHfSlsDy54+PY9lEKFd2uiujLthXEr9pbiQfjQGONHMqnSjlfSf+zxv/0yeHAsNr
Z5j1zFM0DrUVEtMoHel0pFkHrosLIs1cmqNPRXzyPPauyc0Q/AmxuepwSFCsVuC8dt2wJbhcBtEl
x4CXj3csjUvxtae4mR8kWffuHwm3KI46Oqrg5mftNOVwl9yB780Jp7UcEWfhutpl4YDbDKSR5q+Z
37qUnUaAVwB7nop/8kvY8kUJvg/Q0fiy1bGfclQaMWNcfwcFBZCPn2Y6jY8uXYHmQG31tYl6QZb7
NysCUhB4G8epg1VGhTm8Rwk5KaPUikXPIRgNaQgh+L9jUwS+CIYlX7P3bW00seES4mbhBzXHCmek
5stR8AtfaF5G6dUWeY6VW/d/A7VGiCeZlNAVmAhDzWOugVakfHQNMwvlMwlmAXzDBrWPlOTdB/9L
BP/ab3t3XoYnlsqJW5CF5x5iGqoXa5EXiz+BVQNcheRsGTPKFa3xKobPcoJvyfe2G3JdSaJESLif
J7KMXP3pm5a1k29+pZf48Brg+iKmAHOTTfmebdjAlqSBKep8SfXY0UOcCIX218zOD/4MKVRbzs/c
zNtT7oE3N0fyY5SwyRbGAymS6YggCYde20uYjkbqxS2WWglYa8+xEaMK/X/Ezwrjyk3KqetYOtiQ
rQqaJ+oBisD8RbuNdLlY4acuQhr2emkF/Fpdv5A0tfqReYOdg8qY2yMYtpS2dozXz//O2/pNsCfD
/spCP4vc3PdjQvBJHgOyOWk+LRShagnquaBkjlnbowK6sQRn0dDPzx5z6fFwLRznzDZe/e+C6g6l
jVneHxHXST1fHhiJJ3AGKd4Q/D4hQe/jNP7lZ24Ly6tuWfmNeScs9ddcE0lD0dh4mKYiLO9yP2kF
uftDvr3gacwh2/d/DKchaiR+qiX1ESzFgoaCdpol85DyMYNXRIbsAf+dHGrGLVjVDwxxpe8+2iN4
uX1E7eWV4hPsjOt3kvInGLpaTfGsXYsoLyEDFrZnwcff1kl+AUOnAQVYAuV+pAP3IeF1MWtA7JVG
nMDHYY2RN2kb7ixzMQW7utLQfxd0bZ7HpsYhZUvsyZFDIlLR2GlY6yJQ7orhMFwFgunZmt1bSQtw
uTf9jomX+1xO1xK62pUVel5rG/yu4kJfFwkta6OMNqlRL4sAeISTX1B8B80qaye56aFxPOFuAsgf
KyogiIE8CvBMxWqY+vu2AZogNrlM23q6fjUqvg8twm7tGa3n5/U9BwUiwcqzlJ1PRyPWvrLcgq3a
U9EYzt7dZ/IH/q3KXQ66bFyWnW4+1AwX4CbhK3JLThzYH7GU5L5WEeZ42ROrljKMP5Ir7RpiT/ib
eWHxi14Im4PPEnoZAPvzvkbezF97Vlk19Q9Zqkb+GImcPthCx2Nk4HnMmztOLVhQUtBnBU6WVhIz
KZnXwMtf7ldNMAJHgjWNaVepOgJLykz8QXt3U94q4xv3Q6Zn89ztQVyMPyfdtGnzJyukTLpHlhxO
BlUN3XxO5w6gzd6LD6WUnlp4kqyymGIyitkSkZsWgnEb0Mm/4J3xVE4QWFNy4OddWuOKvV5+VQ46
KEyUcKajGJsSNUW8/oYH+DvWhxt+5Of6uhtQHYkxYrmSpIOt3vRfcQhFURglLKQSnBWe60mbjbhm
nyYRMG9DBgJldM9m0QFUjClzdJ7/E1Nd/S7bQ1BMLnmmP1DAbUwrpoVrCO7hpSJBbQavWMH4hCz4
DLEdkjpx9y9CF6TjjD9pf8ilBSmLK7q4Q2wOZLOYfuPa9GrLT0D/3CN1o7GXuzjECOevzv5Ld9l9
qltdiHz/DxDQe6/rhJMRq1o82HHhtJpVYrPuv+GEuBkGVZ3j0y2VIp6FdU/BXCM7Bk8xGKEQrvdK
F84S7keXYyVSZX5VRm324+WSwdm9MtO0292m6wNXfh0sKiVxkX2ZMGJCPTrGXZR46KN2zVEqAg68
qVCzEa5UkZvMHP5pqFfmW315h7qLZLZarBlEopQwFxs10WJw1yWesDPI2Gxok+W47t0RYvf/urdr
Onz8Emu9ftGBHUmv6F6Oz6O+Jxaauz4LjihLsdpIkMJk3g10D4RoAqHd0VmIQkgN32BTXbdA1UVp
JZGxnvtCC5ypfvCY9i1opgupLh4w4SlJbwMzzsjsqSTn0QflDFw9rTUJDbqbNP1U+q1s3qly90UX
FwB0tonKt4Hd8upoFwatF8POHRphDPJan03E1oqL2rKuxia+Y+Kyvv7mI5jBTsbpkFq9oNuhUXt6
qkcj7pQUvGl5U6hDNrwsKN2PIheFeTUQBRIyHzUcOdN8bihifOp59zILA3y7KXS+zpTL56XNdyMy
ZqH2PaMfz/CeAhrMVnOXnS7XUURSbVLH9Va4/xfDkQTJCVIoumYcqyjtgIRTJ5p4MmlakHOjp0cX
FtqxxdaTKLu1mu7ETjVIreS9k7eOYRx5+4MTDx18jxg3MnN1uR9Y/sstQgxXOvRKdkgjwAbJtW1I
hHya3JF6Pi6dKOicupavKBXyTRcXXIu3UN9s5U6KQUbo3lGhsKaMby83dKFeLYBjPB8K57XYEsrT
fq3dNLiNq3SOoRV82qEfoyYtsRtWYTki0vBIcrzwqHmDvovc+ZulO/CL18StFbasV68XGnOLenFU
L1jXs9ybbJlwazvkOT87FWjnekaoQGB7vsUlBjIIzMTpxAxwClNiR3TDcJJ8wytBC9COIkK/Iu1R
OaRRPBueYTlVaMwgQ3WYccw4EXYmVQDs0PI1Ntn/icUZNbfbr5ql85RTAk+Np5U13eONAtwbwv8L
IbY+2gE22xvThc5ROPMQBTBMj+Jgxx2phr2mnsYlJ8lS7PGl7eNyVKO07GQwg6pCvQuw32qZ8bkS
OmDwIdisQgPzUCmYdO0KxJZ8h0YWyWe/nNvImfmIDP+rPpAnZceDeshFZRa6xeI3UecwbV3HT+ga
4aYKj00hsNpuFYMOHzcbvrDzv7kRomkJvo8BBksZ83HA7u6BtptdvzGIt5Kvg7Z3zBddjxwhpb3M
eL9ZHulABj0b8gvYCvdYYxwqWSjnpxiKjZvKwyLbpXsAiwAM/2C4mYPBI2luySFOej8/vKniAhKR
szmLnDykdtWDOM26q9p33Isg3Lbct/7iRAm7LOQym1Gij6t+B5rlAAUvNFDKBgYBZ09+4Th2tEsl
ysKA/RBw2q13XtZnZPnsyMQtJ7z2o3JetmX+EHh5C2DQlj1amQHnwrvvvCMDImShf2SnPUjnWrXX
0kanjo2ri5EPsERc7BxViM2gOJ5SYYFeGhqv0W/q7reZRcMMDLUS2Sg2HH2t/xAVn9Miwkyc02AG
h3XVtCbka/v8z6UIsHR5u0PfwsWlAqoQFqjgnqWHNvfouWzzBFdHEhcCBvi9KlohL1V/X7VhcNCF
7maThPO3w2PgvhBusPo3y3yWTqFtGkcOblF2/mM45r8vTqwBpGScN3zDJbegAR2TkXxfH9QdxupJ
RItsZXP+VIkwLrRXU7CWj9U82g/SlHKtup+2aji0nmXDuvzh8yOCCSBjTbeqarTBV9cptROpMcZH
X1A3kt6OukDqicIwDzGGx8hLVOVKvuNJ5pyogo99ZMVvnxiC5edRL84O2PM8uxiVDpyH5H3buyZl
zY6ZA+PiG7SmOw4/QRtEjaEVrGniwoVPAMa6bpsqK1QMCo4voofYOH0QstfGDPTwQ/D0WlmXE+wg
L0dE5DERnxAhVIuv174YTSBxxF/ZP4S4zifMQD8WDOZVY6C9pjEs4V7+D+ZlD2AfBhRYfppHgqxI
gX5ZRm2PO4L67jux/opqo/+JQQtLb8c6bfekiiiWM9z6l1BdjTLvNIO8ZYUZwhApd1EkeXIZaIaN
MV3oWW1OPIcx5d3ZzLX34VYALpu91fJFfegEnorh+SB2RTacJyVI7F02OPrC1i/THE5hRfhfoTAi
QnEvQf+BJHILdMAi3HfZVo9p74DIOE/2vP4jmUiyZDtgOVwNRB9W0P3OjvQUujkBxBdTLpZjyz46
vLPtrJREeYVOWZ5Fa7cksM2f/EDTTOV02LY4V1VBD8dUiASFT5xVtJ6lWXUnPVLNCQbHekMq1Q3V
xZws3IJ7qXzzXG6XoOpbs776NYr6o/u1x1huxYsuikUCU1drMbOlfu7Jzjs00SnIW6qSzrgnS4nl
uCQ+8yZ7hahK7Tne80Tkf62XCpCGDArU2dlszMonDPvOYXnwxON7lIZGPsm6ZvEY9V7P8U+8Ldc1
Ac9Pcdklbu7EwSm2lY0vN0OimKLWsTExDdZpcfh4Uf7PTYoW2N7WH9/8Rbx/RW4ZysS86mPvDNGe
6YbyW+SFtvJEZdqj3NuYcSFz022Z9K8ZhlWGsdDOnavA+jEzzTiyehp8WO0NVu+EslkcPPJ2lt9r
pd4yooydNZ+I9WOvkThf80b6FXP2ywwIUpQlVmuAcO7PU88TMLwxtegGvng4WbFBZIjqmcpzFIj4
7nBop6FvuHAIvX7lqFREP4ptIAjtUwhD23MF65yiYnLDWK6AgrHt3SOFwS7mMW9S1dC+gr760itQ
8W9WElC6uSf0F/oVulbmv3UmExsEIZlb3TdJsiAdgxBS4ilPpwN9ewBC2J+daBbejWttSyRowBak
1ZJRXf2hxQQLLSNo/VStMro8fri6O05KrwsxHoTNaCtacgOhH4Pzxx28wDFch4bIrEJQydQdxEWk
b8z7K/q5AZQ1wfWPu7mgFSeKzV7U39SbbQl8PS/wwu5VQXO+Z8TCZqEh+c0vqjh+SpicWXEuGSsF
dZwV1sCxezWov0qITrIXEzrGZNiSe5H9OuuPf8KIOr5ivp3sycP7qhJEvrzPBPiugWLL5F95TuTs
0z5AGxiWSpBCwYxIPIlEniBCG1SFemwrUnffcq4/zLl/2D26fMolP07vKclyJvmPF0Yvc9X5BWl4
KI/9YwrFoGgIt5zakPkKrgiZvlmj+xPalQJVUKmh5jYTL4H/fNx5ksP4AApE75DiCvbnbz9TsyMT
/Nn9MiVayH6tPmiiXN+uZMdjV+6TVXZxdlkTqnhZ5elTn6JOUa3hbTJQ1SMmPAAYCmoyqDY5uGsM
jk+ZFEd0oMqWB/aDRRkqHSy5xCcYxB7QEhe4i47e32To7zAFK+ZInYh5igGpu0qhfsIj6ZqwyxK4
msGE4PXQU9jqbruWpZ0rnMVJFDuM0nMPbv3qmLxAGxAsO9GCRTNaCbk6na0LZyLsITPvj0hC//Zn
LyZAeE0Kk1WOlN1XYqRZBubvxj5Q5a9PnoGtlrQQZWl0JoWxF++XhmuDhEqq2W94z8lJXHtp5Kfl
IBMZdY9radUUr2lgnOo1hTCu3bJbGL5qA9MrCd5nx0EgcM9MBFhs4/c7baD90OawbR5NTnD97L/0
IjGD9tdeJsT/q5laGEqOab3f2x+Wk4yD7r9QV+AorJB13ar5uPlXK0cbTUnR8ZPnXUvSQSFwC6cT
TIbhy0eORRVPgroqxaXk14ioUr14jFSzJDNzA58HJ67R2BWo8K7w05jlA9pSK11CVlKLTuw/b+ZO
Grzsn8FKckajxzr89EL+inD5vRqA85BK0TsX6AF6b2jlTZgli8JBp9DN8my3ldfgbuFXdKAvnYpz
qXBO/0qr3OfJND22X3ebOvCXT+IRWaQ4F2WB9fUmm8wXUgGEXSaibblWDII+Ig9cUeGHjKJ321nJ
BUSuiXNA8IiFsPsbzS4jsyRuaOki8QJ9rBwniQthtBmNzXkKfQRiNHQdqmKTOKngJqm9Tjwpx63q
pMyBqzNsq/ObNdMhzrBnuOkyjaeu/5bHq/KNtIHRkb9G9yuvBnCKyDJ0kj6gUXR/M2vly7y6WAtc
8qyHiFEY2GweLtzZ5WeDP9lX0K/0wStBj/9iRwQAZYgXDo0FxKF0/OUJ0JlnAfOLsdx77oXyL6nZ
s3WDZ0R+GHInmbJAbbQExOdHpJuvaFxBekOnG2UstSCIwUVqbB3LuKQYOfsMO2SNqORgXVg1Td5F
UQky581SVZwvW4jJ2PIrwnfIT0S4riN3M75SJXmvfN6gWSEBUSp3aEWSOXB3aWoPoiAYQcxMV7aD
mNSxiVZmKaCP8LKg6rOu9w0bHus1Ld7r0Qa830IHmPrGyO+nCPbnvEda8tiEm9Alok9MwpnV9r1x
+xCyqvfcrnP9mUsVPkuT5wDvDCxDXKsRNG+2gNZO3AZseWJzCxzbqMg9D9l5nW+OwaLkhTDitji8
0oWvSMd1A+XfrjyTHNWKRSnKeBAICNo6x2Sd8L7OoTAvtB3/o+M7rcZhu6/q5sPDzIBoTjiMhtv4
2C3PVzJSLH/fCQfWg702p3Hq9dqW2pnQjMgleJtrfhY7tE4W/2LbDLQpzPW6oR4MgcWybg+Hnsqi
+TB172DrW4dq6Ve9s/R7Q7q591iw9/raFEWIDasGyQzV26RzCFknq+9xExBjxqUs9gdjDlyDstnl
a3mvvU4ApVTSjVSJK5GvfVuiYa/mBk0sWLJ1xHahyzzuI93bQMCF6ub/57tBmAOURAFHDG+bfuN3
nWIselAMzpPd/wxbXauyT6SnXyEiydU9neNSm4i9dvLy5cS+aT/w+yGUGs2xYOYdRet/BEffDszq
GrGYGaU+uXu+LYCggmr/0f6g7yi9ol4LLGq+am7jP/KmtavvKAWA6Psy1OIBUMsTRHimTsVop2X4
XknIzRdIYIQev32tgTCRoCN+ePa6SPI2zfwCdmVFESs448Bngr/02EekuSLC+RPBuM+PGq6zIz2I
i9UJ2d1lOx3FdSLofOLj8NK2t+r4CFhUcnyyXaZoH7ZJkUEGMtRx1l7RCnxJENm4bkd6EOm1VF6r
uzLhfLyHtuTHwq8UR5Go9pz6+uw++MN/6BY2lee/2X4ugeBbumvd1nvfuPUIYmK/LMKNJOVp+zky
y0VY0MSmVQG67rXTBmgZYQH2Ogve4guQCQWmLftzf3ZDeP3u7HH3g3scglfCh7XYzXI/cHzae4CG
+FZNwN8q6qHbRiWoWxLZ7Od3uxR6ZICU2Kj9dJxrxx2W2fZNdoTnLmD7zTM7stQmkxkj+XAw8+68
H3+++MaS4UNtcLpllV+9w26G4Hw2khcKbRaUvcRv5NoxOgGZKKLyZLx479UWODeuLSJLYqglt83v
38fB0njc2XC2bMibdlke7Wrxnk98MYS00Z9yz0urWuwS6pP7+V9rwvCVC+hB0dOAuLYlCZIkxzbt
f2yfD27v3r0sOBiwrHOL+rlblFBXdmKucEElhrV3kNSaxGiTSLegpWKvN2hYPIom5tWhcvNqTS3n
t/aQ1ExiYEdq19CMaC3aaw+6VTVOy9e9zFyBelq/fjnF9J1ICQgJJpEUqa3d1KOrn45nXbRtx+q+
Jm6aS6B7pUonWH5LJnuVwYB1PkKJC4KuNAXtuoyjAVj6/1qGd7HPgrrfImqpD/KDlWPkfknbceSU
0Y8gg8wudGeia396jKOZFLHaKwaOv7hHbzT/7M8askthInxMbKUaieY2Ykst3vZsVSaRDRteXNp5
mZwQMVCGh+6d5O7qykeBhZfUibGOn6xOtJCuwhSUDPd1/NPvs2ZOIilkt5TtcO+auWE7PmYvOCke
amFWHk6IDtza0q7kVrGZSVhPK+/vubmNr/IXReqavChKHNgvQoXxI1T/hTeLgVbYiMY20kWyxXxn
Mu2l1ssizMvMB40mEszsGKnK+WcyuI1sone/34hM/dlHjAG4r8iAeB5A4kFRCSZsr50kknnm2x5B
y+KwL0uEr96yxKi1eCLhf769sBizte+w8WvOF3YjhWbTd/PAZ3uah4I4osSzL9j0DRmn3SQdewGT
MEnpSAX+9Q7KHfZABlEvSzZISPHGIzQc/m7ggTwFEOESZNBGHiY8371EP6o8m9tTXgYYdmsvcsxm
4dQd+kEgrFGA4elayDjfI+R4XoJVY+6Bke0mdhJRG8QtJIofaT6GqB5POwME4pUq88q7YZqf8YvW
wJcZNwKaTMqt/rkqqGZPdg0QNF4YSttfYed5hmJcRERzS7RS3TlGeJopOQJYZw8VuTMJ9HqeEg+Y
3NQTLyJdZH+ZOHz3NzwXlCmgWKeEkw+sjvyiGUdpyRFAmiSg90ClwjqfRrplTyfd3h+nEZz0NmZc
Y95UVml6PI2h4m6d/tA6x4zOUDGATIuLMq8igEmyW0voi+Co/eij8QvMteiXxylQrMzz9hjecLyE
ffDJIxQIcoq0puhKiYVLoEYup4UKb1PG5aA5e3Og781hx+BK5sE0zR5r3LPfWFlCDyMDVnfwkQOx
BuhCfGz6jV7jduzZbiV0xevNha4RbTn8VUxigC0QtWcf2urMs7IYJ5Uiac5Uk2dbZdmBSSX0GD4U
POiatD3UtWhplE61KNBnxkQ8ahEgaUJfiv2R7nBy5vi6NNwz3NzxqF1fyj+lCgG6GgkfSI9NHZTd
Ejwoke5qC/u24oU1NLF2BM6VI2fi1H4nDM1rVURtkiA77404hqwI5Ph/q+w6L8WkfXgPL7iSiA8E
+tJ6yJtmFzXHcewzgs4b5kmaiu3jwVntFujhzRi4HctUGExKIG9pxpX15mPfPy8BCu+Spr8g6jar
PN+z79ORYAR5fnTwQge2z+TY8MW7D5Lluq29u3WLiTBK2e/8BngASlZ7GX5t0T5R3IeOuMrsfPuN
0eKgkojjH4iRUcbThga1vBHOfKsRFQc5f9Oz+BRdlcogwpM/PMC0G7YjGvomtTPcVrWnEsCHugWy
miYtc/a+Hz31ZL5AuAXR+8o9VDx8jqPu7j9Esljia0IsJc+Rjh0qssI+IlHhtDaiOOWKABSzn+UT
/0n1swM37vDzG+Cnr26nE9reSVsx66SqEI4yR34PcZmCf6HyN9g5rt6V4BoA16Zq7aOV+e+FYN91
o8hjWFz2pu5U2uN6DtiNmrP5zZsxyhYQIoVsqO+5ZXuycKArB4x/WU7/owpHDCBNYoogGHycVlXL
K+VFeBGDWV+3xBitUM/BlfeM2z1oGZ3CwYchSD11DecrfGvUlKa2emDR6/g7ddlTn2yINUtS7FDh
GfefWv60gwIjabfyQ6EnfKQLFQCV29yv/p27c+6s9gSuZPLg1ZaNrae4X3Sum2U/NFnIY0aR9JKd
8SwMuJqk/2y0HVwONKRL9EY81/kuauR5cABViq+Ktrj581ubrZLkcg9HXKPYiO/hbLDoasxQ/Z41
JypGidLHybuBWBT/p5UgesjOLVbtXAcwVrAHdqC9NqMvolyYvWF0IWjAc3IAJCROdh17ao/QDv9W
TVriig65E7b+8yyVsJb/ZMtK77WlZ5yhjPA0ATx+OaqZ9xwDlxpy0RvuG28xA+UpDGcz9v2jzRkl
iPvK5XsUFDrhmCP97H7XkrwSKh0Y1+atVa5D4VyPrD7IyrBn6Y0ueDde/+fuZmxLFEw4eyL+m8yb
3kbWKa5e/RNtw0EnIuRAbnkMsqTJEvqp1e7q2AhnE2iUHUES5ynrWcM4uehBA70mzwcNBm/0Lg4x
d4MrG1SJgkWbcyi6Y8JK6XMfBH+NeHigPzTkqxdcnPHdprTIzfpVz/ds/wWo5tjxmZsx8ZrfkoUs
osZgi8l65oP7r39TisCYdYR0m1To2wfTyYDfwCA1LlhyZxkYvrL+1+Ub+liNdi2IglSGkxyJQz/A
/KxPspf+Rp8Nd8YP0TIyqlnrcXow0jp9WmybmTlCB7NxOfjgeuGqdqXDvBpnWu8DCpcrSxlBRNgv
bwBMbZeqihKLlqutII7c2Oksbyjn8vrWqN2zsbLDtks3q9VzTVa3pfBAGI5pLZpZi79ikhEAB62t
S1Yp1llh7bCr3WmkRNpeedDCMsRib4SAaMk/NoRk5MGVLYhjahaHclQj4eqpXhDesQH4XEBsn/Z0
aHEn5qbw4ZYi74lNp0RKu3Ens5yy8I9CYUWUnPYWRSsANcldEs81HMlUA9DMw1vbXdGtrmgeLjwr
ZGXfgYS6u6B0BbrCGV46wWEcLKHD5a12PArFXwEKdPMW4P+CrlsNWtzgzgP1K5ZyQygsdQJDMoCT
llAgwMz2bPhgL6XEaQkQ4qp8Zmgz+cQd0CMItC4Orld4oMczZZEUtjw7M58ef286/SFJzdj6jBJk
bdgppab+q8umEkjy063z0YxQUSQrWo0+wFN3IBnTdzXZvGNq8xw3wkd8lEwg5jheJX7zOcDZ+u6c
AelDvZ6FvlOR9lzW6zoJQtaAtWWT/mSk43+5XeFLgFZWO3BKDBUBuDdkrOoe+nwpzNuVRRcBbZ2r
ZQPABqkIF686xgs5XqhBSrTe5eZEtEFXPwhpkkRqz3zUqr9VFcWE6QfhArndRaIYvI2TYXtEJE9e
L6sQSeJGg0Eyp1kZhFNh29G+TF4noiPEdvpviZLmyPQpndOd0PWB/UuXrzWkx/iS8IVkojkLW1/J
T6cDolpEWO0pb36GEBqPUpHbddTudOnDJdvnDfksQa5Am6EwWnHL7f7M5WcBbNwH4Z3MKnEO+ZVm
BFiBC7gLMcPIfgrF3HxkEkgbKLsSL3NrHlckaPxbMeO8vjdCs7+rIRmNKOxWAZNXiKQPyhYX1734
LcWQZot1yTINFGjasK8uqKTatFSO8sjCtN2dLt1fJX42ctrjDy4U8PSnDAcK/Piu60j5ShDVvbRT
rVFrfgQxu7AM55zu+QehVxwzT9lJBNf+CPJaDPtfDiJSr5hACaHEGZpBo8RI2unoNe845pssy3Xs
Ve8aeXhOtCwi0RbWD/4KQJsUT2PEo7cX4rc07d6l2p6IeKKm3YXk81f/TtpiSDHgdyYOakJpqr2f
YPC01VvWZ66MQ7bdONIncft5ztHNVRhFQZSvUN7A1GwTvKLf5tGapbsKCM/T1NoUOk56bSZtiXdK
LuwzimZwLAeNTC1BoJDH6VKIUJTNP4OEipVvYj6EfiXloeNkGWewpiKCFXtJKfCVy++FiJoiPcX6
ipE+l8HDsP4lskDVlMQIkvS8Hiy02BfFJtEU45amQibX7NH0SxJS56SC6BuVpzOH5nGWoNpX4ibO
Mz0qSpf+HQwcWI6zFooW25StuJGy+UZ5p7iPADAWQynQwIVjDDNtv+WaLYQ6tPcY4Z3ujdDKOIRz
x3BM9SJwikQNxlOWK/x50odEMzCEQIjcrN3nS6M0NBplUpja7Zo2EhVZsNRyfM0PN0p/WsDS/u1m
4RwjitLfDB2JjcqgkMXFqDx7PFlLLCmMUynmDE3wtbIyy1ymPoh9aKJUgQZtz3u97T0uQ13uCS24
TZ2w6vRu3C+9hBIf5dxjpmqOsBe2bn6u2GHu0tSinCek9fv/X0UiQGC2P8wX0PjwrPPN9DYZ+Cl4
wl1OCN5aCFJOVJ+HxqG2MKMRKbTlHZDjzGhEVvIFi7GKL73QGJen2nl+WCfWroLSEFyvqKtf1dae
4qsi7PPrhV4FFeEmCjbaC+gJ1GEimFwTWrR9QAnqrOFSEF0MxTbsPUOiEs09jYCOpkhS9kgWuPor
7QSMour3Ln7i4pP75n0oZ9/xb48XQmkScLEgV3dbh+fOobirUNYvmbN2eeVoJSsgVGSRzCnjhmad
Q1pRxlovxRvR9waJzfAxGCnHlmCeb/6SNA2N407OCWalI+W63oOgyj8uFp8qstbB+j9mKP8VXrCn
LDQCO3ZpfNFCwJ5msxmw3VmyLddo7D3Yqd/74HLrebCk6xXDBR8LVwsDF44N0l6aPl+/s9x/nOfJ
T953lQzYbtvjFmcCcoTd366q1ZIOIARp2AnJtKQzYY0yAvac/Rjeb1mPwrA0EChbgKbe79bKDgrV
rt+Htx3ZGMkUO4ppMwpNq4b6CofAlkQd57AcAM0u2oa4Xc0pE3m/9/BHn/iALc3lLEm1xplGV2Xp
IYSO5FeyPcYhMEiMzgKln07aXNuiePrRrGnq3QDANcii9dxzIMGowrzWTr1nGFHG3s13y/bgIBX9
RbiuO5SvHn9X7CRwDR8z0FB0GLZuXG0ET0Rwz8ZhBcLyIWOqTbDHkrkxX60pLkDIEGiakR7/dV8Y
aE44BESbY8d2a2pF7LXQxsYrZihdPQghNbblqpgEibuEzORBZ2lJgubOmUkMocyX5xanafh64kCd
ZbbkB1GOM2UjegATAgbWwK42GlbXyvi7igK1AtapGYmQ3f6pProjzGDILIVv5SxvJzupm8Ccd6uq
RU8YSqIplQsU4lNjxHAyVXNr4e9O0bfXK4/PcsS3ey0l9lv8VaYcfXnIAmF32P+KQERLLffSNUSv
FrNGS6VlC42w7sFqKLWesCO7TwbJPg3pt7xuKnddTwQWx9VAZLpzd5QNGPi+/U9fBxtqfXvHENB/
AsBMZFmcC08hfB9nBk3PmfGyBFMpnhk0d+aUOaGLbzQizMVe9Zj4TE5cq1vpsz5uFVMRLOTgQy3Q
dKMW6eXz6WUDrKJwBhdZ8XPziJx6NKl3LDY3LYSsQPMvR22YByDm2NXl3as2F1qFyAs+Y4yJenEJ
vqbjhGmaCQCQlj3/cdA17UEqej3jGAfJazgpUgW34hddE0xsMdJpBDfq6ciJukhB2hJdOdWbPiGj
+3WmC5vArNIRUeJ7w+rcIzunt8j9t29aB8/wDeZ5pFUna8+oPQwg069DS5Ry4AkM3RpzJtKpIYXi
G0gwpVl8kk7UpuDzNYAJv/OdD/wnr3Yldg9hEuZSt/OcOYdcycTbRhOCAN863x7w1DAPfeM1cJUK
jXkmm9QXM6F16vTdfiZQz6BAvFZiGU/SqhPNvhL69S48/m2YcBy5kqF08cbEEcj5K3aUiNKed5LV
Hi4UX8wnlINMw/WNIReBzFUz8nOOG1VTXVIaf+V8tLw8Kk2vXnGmteH4C03tMohiUf3VGE0mNiAP
jow/nasfaJLhdSYqwXfYl0140Clou3m57Nuv9cYAA8kvyRFsiCL+rhZ3RucpMq9+zeQiin+gBdLs
xckGt0tr2RYyotwiuMOBBxJczO3Jj/Rn/xSyp9ScxCc5T3kLcUGukD6FQWLpaA0qlQ93aYw9qHVV
oaWDrn0r7mkg4t4uLjSct4DAQy5yuWyCzvmlk3h1hrHohRvaYgwOad4UOhakGKXAwS8Z2BlFQ+mS
Q2adxoRDb5bWKZ5jK4qcG+MfnSR9ibOv3EqqiAhFCbY+y2A0Zo/9Z073cGAC8vj8GcGZZEAWq887
ubLaEIuW1tlqsbEXLtWVBoKpNTw5MX8bL3+rTKkUSlzV5Pc4auOCwS8JzFBxj5O4QzWnNyvp7eTy
bV4owWM+bsdytmWJ0Rqn6jm1ZlRgAO6P6l3dHRrDz7zBczwyxVjjYBoM0lQIJt5SUvaE79z0
`protect end_protected
