`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
j+npTEkrOuoAYyMX9/wRnMYX5goQTEisG66YW+i1AlzpOzLle1lXgu4EgeH5FLw294DViS5wgySE
5m4qv4CG/g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
gUZcfjlaOFMdX4kb0TbR60nJXJPsPe1GyqlMGQubcZlG9I4tJ/ZhHd1EMxwWjzpXAI7Q26CbWB5d
M0N6EdylvFtjmg1EUNKbV6Du+MfiD40m8//+pZe9DGyPJfpmuD4+Zj3hF5SrXabgZ6C1Xp1icJbQ
L5r4LZJ7J0joZtYvw4s=

`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
m5BR7gQYyud1p/OTN3ItnmfZf+MrbBm5KEryxpppgQ4iwUC0k6E0EmeGOhQnOMR89C/Uz4vDj5vP
kR/7K+K3yLfHLs+S12FpPBZ3NyuY74QU5rOfBxCPg1sdBKjM7iwVGn/Ecb4QkpmrleGslFvuCXCG
V1QSO28mdm007Vi1l3E=

`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
B4L9p7tgqm98VIH/YFg16sVSk71xEJ5QzzMkqAXSOWwulHN1TAbp/Anvm0mHWyNUaf7zrkLBC1E3
DyXIIdN8sGBbSREiq3gWYd0NIbQUfdJZZYvs3uJPPU2+ALQYTUwHJ5s3WX/NzIzGuAAOCxw/hePs
QWaSntCuSjeJws9v8g1EGOV7yq5Osdtd8x2LUU5JN2WFDJuVRSHIv/ompQlok9q1EkqQ7S7sQz+i
a0PnTbVY7uVeCYr+SXmQ0ogUGteEgW6M1VHjoHTsYDuZz4WbwB51Vlt9WJ1soaYWFGDCJlDxH59G
F3endzqkQitpYnFk4ShPiMODHQv12VpfJYbHRg==

`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hwYr4TS/aBHf+wunP3cLIe0CYKkGOTJ5Jld+NMc8xGN3F8TLtDkRxbVMutpF4XfSBJhLcHSU4iQL
iFpWN0M+yLVcuPEGASE+OmR037wzVwI4JbEmc01MfjDNWHEY5ss30fwhsdWHpqgsyV3rfWe51mO/
8TIpFsSC0FG+zpoqHyDwegAf/Lmf4zKpgFLLo+3OtJAc3YmnzL6aNZ5o46AbwYzVu/XN7Ak3E8lI
/q6Y4ANFXbA7iDszKKZ71HKX3ByW0rvpUTg5gri77obs5l7sIyfp4En11ig6Opv8IgX7A29qw9SP
SM2VCK7D7eVxqxbxDEPCIbcxsa+cEizeFb3ajA==

`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2015_12", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fLcMKoU95J0rpQurE7HrpDJ+JK9crolX2l3JMVmKcpL0dY4KtTMeR9YZVRrUm6v6lYXi1gKv9VGR
rJoz1MY0q0spfAy5jHcnDVY24WoZRTIRmr1rwKTVmYW99Be9KcesnhPZ4WuQur2Sv45IkqlI47hK
jnLtqX84PKzW0ap4HnvRWci/sP2vA5n5UU1zybiOUtlCnJBxpHY65IfbMy3yrF80TfTrR26jC/co
4alM2f8ErqkNMnUr0tMjzecZ/pjdWFH5wg5jNvR9C2o/vcUC0kr2fnXRwsQXgxT9vAbEitKz9+8m
p1Mwc+il16beY7eojdApx4J9ojOFXIxI8G/fSg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1032656)
`protect data_block
VNYkwl0rEcKPMuF52+DMTsHR6VK3mFUVlRavY+1qMoEJd6RSiKV9iv+7wZi4qu/mtmdxWhWs69aM
tlQ+O1GubAIaI5VIDbUp99jEG13mVRFGqe/Bbtuc/vIDOwgv2SggkNsfbmbqOoKaK17awzcAh6jU
0qoJxdAzek1gXMw8FQAxKt+aD1HcpTF3wlB0jrzsc2nH4zkROYDGqroyE4zRLu8ZuQ8CqZ2G86EQ
8W4ptV1ZJbqWRuDcM+8x+0ishDPpwg03BFj78V14232FpWZB1ynMPYEFK52gjfAakIAI53D8FBig
Fc220JG1uT6DW3hxNgQuCp2RbkwB7Z+s7U9AC2/IW29diqCK6+BvopOWdJIsLUogSMw7fqqQ4IFU
ubtJ2OiQ9q0tqA5O/CQTXl2x2l3/Eeb/HwSWG5tGI+eFn8XhUgdSI4YZk4xGarJgdGThA1i3+cO8
VaB3Q4B/bBX+193Y7E0gLWwh8gKC+C5TKdY99+qAt5vjE8Tn+5DSnQzojKa5VAiuGZ4iNzfboAq6
ZpIY9OzDM55EGobnUYRxLOkNyMhaNRben9i3fJDac60dEQB1a1SJD11sFVs785zaXKCk9YBjiGLT
NxP1Nc8/VRMLgVaqTlVw+SHB8eObmp9mpz//z9kJd8FYh11lSZUz+qnM3o6ilMh/Poa/S6lVDHYz
MRZoJTimQfbxNN+/izG6zNVmrDdD8oi6QD7mF/0vIvAEoAhxh7rrxj0wvwYPD7AabaAO/URCJaZ0
4MvSY/lBNmdOWfyGXr8NCqARNMJaCJnw0RrqILSxQWZBqVZBaJRPsUFF/oFwK/QXQqskGEOgD11H
E5RswR8Iiz/3Nje4Ygv3RyTOURSiaOiAEvWlJ2xdlD1oofoKTGIDJr+gCwQdQ1hSI0m2oW3Q3+C3
wUjnPraDHCUdYuoZm+L1x2zpXClv3Tzdw0SpcdSkOpde8fQX81UrFC0osCOZ5o0vaibVIUkc/4CJ
A8iRMcUp1ImFsf2eJd8LAy0txsT0uEY4g/IOrHVh/c/rznijW7Um0UMxQwlzoEpVX/kfvT/crPoe
JNMmUXYlWgb1dw8GMW8xEyQ9nrEoM+ESDiNkx1pHjlpb9U72RX6yrFt9uYC06koYogmCrkT+GI/v
zFV8GXWHwRFQSB9pqf9F9JetP9ls+BAggKEEg41qwkNhRYgaTL4hxHpn1AaoF+f8nMhyc6/ygsV8
OSneO/JZu7zOS/PybaYejsl1I0jQvOr/bOEnW0upvG7RwMaf2FuGr2fNgX/geN7GG650etM8bmQh
OXt0ik4UFl6mUzUyOHuRI5DbBctKahNzZPjVlU3JHB9TNeUdJ/SfCWz5Xt15xbKSQfjm4YhxJqBd
ZuUfjSBLNw7j9QiEpFfi5b/d3l5yGIhbxqgjt04rhKQ1LEVGp/ghGSMzoY0yQ69kHH7UuTbuA6Ct
QpOq8EikujPIA5EcUzxFtpeKtGTunEihDckMNUK5AVv4bYcS2yemwbDeN9SRO2vuD6xsPNMa5+lE
SupunKxVDpLmB4aQpzCv4dDn0jHFGpXkp5/tZQhsTBRinDtDiaZh6LlYr1MoE/0jSx+qV7OknRVV
lEVjVoh9oaUeMAM3tJU6XHP1uuskBvUBylVLuP8yfDeEHoC8inS9d4m2hRQGCBKIEz8AgLZ29Fqx
of3PZ7CtCxOxBJ2d9z/iIo/3F2ocemaoN/61DBqJsrIG5rYk4sLRqBH8M8leKWspRn289yXhxN0k
GppzI92AZDP52wLCEJqPj/ZIi+edxsi+QVUpoRwo/mSACJRFq9LUCUdt4Kf4nf0X50ShwekXQiK+
UgitZVZY8OSDkmQ+qr5y9mIFN6YzM+vTDzNek//m8UlzE5U6Y02Lb3GY9rCH0qysgOideBhqLrui
I8mh7NFXf48ysyi+M3m8GfDsmVaowyLFT1AIhUIOyxtMhPEgjW6bClGfhSWQYHzzIyeyHFlM21gc
9WxtIZqsrb8Ps5hABaaeWvKdJLjgf8Vs4YN+wr1+GjGqJGn4TNAi3wqfORvmfuHPPBQmlwOWvDJe
JcmMsu8XlVEbpKQDD7YqgISC9Tws+ULJCkTZOeLWyRKxb4VrfbxfEntLylnXdD7NVuDJUCfUnr1k
/3JYdGfFahJSMFM59+FZ5ndT3kuvj3B6Jca0NcF5twppje67+z9A51NX7L9OBrKuaB9tHmyrNqdK
awDxV7mhI+8uLqltZaWgrbaTBpoXDNBWc7jb3tQOw3meJdpuAwnO5jFlihvZqHFN/+xOfHl8HTpP
CuxXJGWU6pfTjIJhPboWO1hdCxWKwbtvBiFu6thptZHPaB4+8gdXBrNm7JLVjA0qkPYUtSEbk5vJ
VnUoUeli0pxivkONDpbjiq3aGGvuUuf3+R3bmxYwLL9lyZtdKjlzduwJkpX1bmeYr8D5b/1APp28
yQCjH4O+XCt6ooMzf6iHRcuCQuMAESXY12oNLBp3iVFKgk6TuiildR1DmQr1Yy6FCrgOeC9R89hR
PFTyL2zGZeGbtELSZ+OauwTU9km2nC1WNHBGPw4j9Wt9QtaF5Trw1MpWxsRDHFmLg77q0vaknGQJ
0e8vomyhnwMv6P0itVs6Euxe1n5hb5knYdj+CN08d9R9rQTYGdaiHGS+Uu1+nRII7l6yJ0D1cThZ
Huo1rSN9J69sCelYx6VPOwIeneATO3WVtXYnm/adV4P/PT5QvWPHx/oTUa3qZrDeMLrBT7wQEhPK
/xkSvvNb3KUfgo4BkhQ0t2q6AIsM+SdOeY1IlQaPIZTzdwvfEaub9lw59kW7afBvc1sRYwQQhBJH
RsIywfmU4wLWczN9OL/xXFp5Gm0+72jQEJf9/3xab8mbUiKLGegksxcnqlFE1yhJOZ8yy/Tqe358
otctZUmy8rtRSbILS4pypzd1aEOf2JMjkqZfwDQPJADrCrL0Qqr2dMybn6dz+LagdDauMmkLC3CU
WwlI5vWMPxyHdJlo+g1XZWkAJNZkL2RBQHWm4GZoI9YpCcYNaMI+CNlh5MlYFthmP6lJJBtX23gz
zUJxHY4CWuWV9FQFUPD91+FRcBzQHvQWnEvNXTFm2BiiA7LPYp41UoYkEsGepD89OquNuMeu0D5+
4KhUFaRD6h1qgnhJRjpGI8ntcapsL8zfNuJ+ICjTk7RP13NwBd76Dj6ub2KAGC4TbcnCoWL9FF0l
Y0VDnioMpknUc1AgE/g4VR/+JyKuVjo6R9oYMc7hQPhOH3t+J8r3yuWyDfhSS7usxE5Ih2YSRxfy
wqBMVXunVAppcRJoNVyZpe1O7YE+MkuZE/PpXOa5IvIb4cv6R0ne1KrV86UAUwCDS7u3yPSGOrx5
Fvx66SptCn2bwodRk8tIg+GSCYrvtt07mZ/RiMqS0lN/DPA+YlB0vH2q1pOlMYf7x9iknUn6T3xh
Pd0JtLGNl/LlMmQaTKUEnJuEenGzromK3ntTJHcTdECxu6a+QcvOtoaPyW3+Hq9m5b1RY4gew/3H
caS2P6F7BsMTmlOTKfEnVP2zQuBakefYso8e1e7JJMQX8ZnO/put9UNR4vw4yWKu8BGlDGn6pBoE
I91nBRSZHBQlDU3usNQ3RWUHrNBMhwVkOZHfmxpx2P8skOvt2b2bn2OCpDq6U+k+5jkpxeaMrudN
KDQXhBfgOsdjpmTaoZFNCg3H/goaxAhb/eE1qxZsFXEOfNf9Q8ctLz7jnJrjZwCdsyIkJUtAEg7A
OwvEBjZ/DBlK9eDip/imR3Lv/B7G8cQVHQ83Ooq4EdOyhlGavpJUvxY5PecMcnvdTYQlz/9PcgDN
whKxjKfbqIoEQMTVUe1w3a08NCCUkOHiFvsCox3N/5D3mxkDEeAKiw033rztgBdkLBHaHHAKExsB
a0nymZn2AFcEWLYzsV7wpJOmkxyUHDNGBHiM0YnVMGIZOrsVe+/0YMN4ppb+9vtxvOHLK7b98ILP
sZCDngnuMPzFaz6x/kPpYTznEUp4BH06vRBF2WyO6WGbJxWL72Ed7bB0aKcT0WKkynCkGYSR1j4i
1DdT16a10Mj5y5llki6LoCWdQAgmnELM+xnq4UQbRc4I4vCJ5N0hq9xcORJLExtZ+7FYKP/dDYzb
ZOht4ruqBGxPeGXqg/9p0YegHNlFS+OQXmMmNmaWstCUy5RPkns9y9f+pF6v40dBihccFORWE5BW
FtUkBTkCggjT9GrBkWC2kyGSeVG+JdPYRYjD55Hl6eZgyQIHFLctQGiV/ZXYcAjHPRgEgVqdhKrm
SF+YXPKXDMDIiusLrD578BYCA1j0fQ0wuzWsy1gVC3RnJ6rTTjwi4i8IO2lcSLWiE5yEQbZlIhHa
0Eca9CmJmQeP0ffVnRE9HBXz+N0vONtomWx4ZF6wNGwwnntr1Vy0SgO0k2HMz3GqpWa+PK0JeyFN
tiwqOPtFH1HeVkil4JKDO4Gwhj9xfGBdio//CU/Uzwg+1QPBJBfpBlEzm9ZQLBRTJ6pLsbuiJOcN
NQfzRshm2Chg6mHnFujwaSENu3m7Gpwf7vhe4tEAFnMphCFCEvZIbvlkRsxWoKx+Sm8KlKu/EeHK
SDF8JaOH75DORCIKVts5nkmLu5JbELm/vTMw5bCQDtaYRGNi4Ajswcf2PClhnA7jQp3CZrqcWFZ4
6CVX4zpexuvv5jKXq/BpVx7kmI/E065XI5btYlmSGWK0YeMBD+y3T7NlAqpyn30ifO6kLGd/pHAb
AHQCREywh35rI6YwUYnB/uhbjH3RBtPRi9TbjY+T0HHjmI/yFv22Fh5M8DPJAk8f7KN6FXCUVcmv
NNfaPUyKjj2AOjpNgSzreYinq4f0T1mUWuhEvd8jfBrGJqXXcsu0PqHe4HlrN3ffGs+D0bXBFc5H
B3AN8HN9/UyWCA3dpYyIt8/wxkU4MRKmZWZJMY1HERRVl4nCQD0MWjmbCq+nVac/bwFOYq0HSbhu
EnCJuv5ri8JQ1AAsMJDgvsD+CIdIFK16AOHPEi1OT52bo7xyft1oiwTyxZwNhEIRDc2ui5aSpdEJ
eSXkhrwAIBcp8VsnefMc4nbsVKYQTupMTK49zs55dH2Se/2m+pqPxH95SgQOd0q8ONw/0eFa1pAi
ZWrn9hyIlt54JgvnG4lsKs/ydZyBYWrbSMVQoj24MrxyNTWted2N6g1hSx3NTy0BGJljqvNuOzng
UniuRvUCx1DtTogDHXpxHSOv6AVBu7ugp7CkgPDGZB1bSNi+rRbiju4TqR/7hJQjZ89mTQy/jcyR
X2mO9z+sjb0CNrcHs03+p2i8YClX1eub+1AZAVCcrXVzxLMZ/uGjJ1C7KKwZtifLiDiSCBbzlFFH
XfZqjtJUeP0j5EjatbCbgdwvl2J2trKGVRDx1XlPDKDFjrbtXJyGNvojEhXbuDXReMe+Dm+PsSAr
uXvLR3hOnvNLhtzvmsp8nC/PgRVx2rFSpSiaiSozteNhUrJ+BcE5KljqWBtRSnQqPZwB58qFSEyh
3kntaRbv/Nrc/wyCm6cyXVf86nZ6m9eYDhLY/tKTDr1PYLFWtDl33p2JnRb9zrKdRABt50XJRcGd
axHMxfSjOrj66HEAE6a7LmEs2mcI+FivNMU89CUIHNo6zAkGNocDpj5mXdtyYu8K2WbjBLLvUSH+
4+VOdh0r1dwBQ56CCiE2cd1FMUluJu5TG0Sq41rrccEG5FVOoCrcNdRYc8izKeF5n672fPK9HytU
pqfEyT2q+0xkN/vcWPiD3etgnZLZXgO/yUNJMGxWMEb6xrVxF3iHbmL9nlFzS0oVtdX5vXWvc+Y/
jyhA3tqhPo0acK0BqJ/EaPv5g+w4PSlhUtIT/qhixlNnjxw1otKh7GfKHFsu+0V5o1Zc6UFcfurd
9qhrhPLVvjclX9GEm+cdpQNrVVNG0MyfyZGIfWguqIy1+fsyPnxMlh348bChcTgOHpUC0ZDQz3+q
+7pAGEmuqamSOE9q2LTe2BpbvL1xo/FKUoxDWXUdgjLKd+ko1/MUtSd9OUN0v4ul11T15/iGq2/K
utIKdlsb/tpnJ1LSWRSGvjgZ/J/pmMgB6F03mzwsvGFJUsl/pLqKv7tdP/wy6CwPGzRg2ciKmP0s
A2+NNYe3zVXCcsl8yNN1EWtjeASj2hLKBEc1Jsof1SHJCj2T4o69CsxGoJYj0ncic/i6Stn5i9PV
TGSqKxWm80v48N5oLKxnvmr1bCKYq41CEYnKfcAMZAfcQoybzyxMI/od4V+Op2hwWD+9GyRb7855
fYFe/ChgWorgd/u2qsPtFo417pS1wmgo6VcX6ujOU6XEt93tDYLBkHeWv+T8B/X/QXQJ8iAwnXhf
DeN1SQwarjzM9di5EXzDI5eYNT//InDbaI5EZ4b0BRxJTHaeA1Av8UuR2aJK5rguRxIwmb15C+8/
lwuDwg249WWXNWzeNZW/h+xKV4IF6/FhCr2CY5+LaI1YtWxZDxKGuo/+DZ3VWsl6Jav0UYTMEjPm
ssRKkKCwBci5SPM+pSZHiYyUBC27W3+jcEp+S2zaLrnN0t5QDPKKxV6E+uSoMh/jvFPN+BXwXaNG
1hc46hUILPJLa/yGkWm50gSiWwcZFV6CANECa+3R9QA48RB1b5rjrlDEw8pJGe0WzYlsN5M+Ujho
S4B6b+xNh8aRUHMxThvnI+uXXBh2IUuHHqxH7/vBjcJraPjPIwAVGfQR7aZowWKf3/rJmZMJHTBR
kwECvll5mGthXxVdLPly7k0Yn8GawHfxEBqaoH5t/tQdA1Uab5ydKHs9/eCq3x0d2Xy7IF429D9c
mh967BAqyACNr3iczbI4DWFDM760+t8HF94vkx5PIvictip4awtL2E1yrNtfgh0UTyoaAbH9ekQC
TGSdcJfCzFwy60S9OE6LMbNicMoAXPaWv8eJTTT0b4nPVmUlu/+JufWpk1ezFpMFSwmeglRNC57p
QWq39l2WZYKm/S0EVdgYSUmL/lPRWLpejfium2ATcddvLjZQH1Y+cj8D8XNRbsdouCtHuFtOtx0d
tsRBnfRJCYn/eYW5sa5b2feFvKCum98Uwy1VnT5qLywL5vG8CINgKnVxDQXe60niDxeeYPDKB7XR
cdRDtaaoiJAMxbXaWmy565JGc3Yf8c/MZKdmLyltO5W7wCQ8tL5qPGzwMJ2XFqoZ7ohCOSctgTrg
C8dUG0d6+DXO3LpLY8lty6w9y2i3JrmeDykljziMLhuyNTr22ZhVav/Hll3AZsP8nM9pCJz1pGWE
P/QfstkLYy08Ts7LpGrUyYC4z9ivYK57bALD0ZQkVbnKhoNgALy2Zw+vyja8/l52d9AQQFeN5CMy
C05NE+kFnM3XOKHFhmKagf7KoQxVoBxRaWM8nhkxFReGWMAbuNRJfi09JpSY6sHQXARZ5bYE5FtA
2mXbDqRP8gwDHE4AbgtYF0+ONG5kOcsBSES6PRb+RBk0ad9Aown0pvqWcjd0c0hRJytwAc5St6J7
jIzNhfM2osA+7wUS60fvN28HoA38/m5VaPllH2ZlGpr5uKYDWdn5h1Xlq6SfvpV505vzmuE3mAqK
zQuU1P26j5wYSCEwGhnHmCF7mACQhG7PVJ0zsxpX4OSJI8K0xwqTGGD6IN8dwHW+I9SgwcV9RHga
a/v/qbG0etOUBsVPrqaG+oztYUheG4J4LlGDKM/uAr1S79lOi6Ra/rQy4Hnq+L1XVQ4seJw20fQJ
eqpUt9/9tUqpN1FGc8FgH+k+omiH4jqxLAaPzwgZ49xmIrZawGez/OUJo4kpElOy9u4ayIm5P+ea
ogzfuCK0WhTJgNxK4prJtYvhA7WlG9S6L0oJpS/6y88xRMk1j0rCJ9mbAPbbMpu3LI3n2PHlcIhk
BQ7HjGVK+4fdzoHWDGrPOUh/srbpaqGYvpGwt2D8t3TTmsi1ki0AE9B9r6l+PWTBWOU+YUYdstkm
DFtkT5a7MbxFncQoEPrxQDovt40dtD5twD0DvwdwN/xNfV8PsIOEg1l+PoFH0xozKLptZ9TO8MXQ
x2N8dLa6wPsxbYaTAPME3aCZbnl7Vy0nFo9Z5LZqvxL0wR9HaxhbRe16TeAdBfluK6hTvfcL/s6L
wphwiHRQt8rwFKxL+m3Or/F52Kh0fXlyMJkJrt02eIqn3gPw0QgwCgR5gU+N4LgFU6EvpUjTxtMA
9cMs5EOgq/IqcLfp2nuG/3OYxGiQtqe7Yk3tLTCbcUt3/QJE7sSlircvTnq568ltkfmIdxoJv+Cj
Ck/K/w2Onm72CNuE41zfct1Yvvb7R3SqtnUzPTYAMfUVkGi2a/fsgitFVZBsOTV/xHaf5UfxPwrN
NV2HBHRxWniuGETqru6/Cul1WPz7cUJvftB/3JxL09cw9283W4ykHNsNorBNrPMjXK09DYwqYmk4
nj/dcRJ2ARNFdpoFHbtSqmJmWQ8ZNMVoa+13KCfndmbe8RCHrKJ0C9v/anSdzi8rVv78C/CF2il1
w/FTnixzZfetwjSh4jeD5KX4yOzlIzCsE7hbJFpVUcRjTRcPP2InKlM0gAPwaj7r5PBFdMlS3qmC
PeRlWV+KkxTjMjohMGuUBPBm/2d0tScIYjjXJtrwR1LtZRFMYUFM+IFSQszHSKt29p983VSjddEG
bXkDZJ/H5VPYJxo7lX9q1HDmvfJ8xQznlTfTWJEF0ilhtYT04ffO3so4zN/DvbbqBM6k6QRgJX9g
IYgc+NP4divzu4PBPchpkbQLlN0uZMxguR6Ao04rZC4jSNkm+UIcpg3rCDZnyNY8H5FibzQ5G8ZS
e+39y1H1f0CdkmRStkMLU9DA0P/JwZanxzEFt67peeEvUzEdJ7kFDGfY2JbnSscK0RWQmDsBwDvu
OnPwsmH0zinRp6ry9fQOsRwoX4WFQJSlsC5F33BsYUyEqQhvflojUoV59guI5RhwPgFedOp7kHxW
LUw8ur9wrfPefkDap9FVZuhBE6Lz3ReM+FE04D2PLE0BHQsH+MPRE00AeqUme1OMH8xtoDrwmx/J
f3iBaYugjEbsj2Gh0PyGf2Bu6vmz9mFHlwJLQoIPFqkN0VGxFWUxvDRAkbgmpjYMIFBDedIFv1yj
aJtxSj3f8AD6/nI6HxHbTqkrJENFAch1A2dlGTcEYGIRj0IkpJxVn+DLcXNsQff/cTxbfgdOdHnz
IHJYgwQaITXC5UlhSMHx8UHca19OsSoPi97pymInbDJ3TrasT0/Ddh5+UNqut2MDDG0dT7033qjr
kpEfSBTj/8xclAUOuYpRksDM0DRAHBIR2BM1WEbYp9DsV7FPByTsAqUOpkTSMIy+L5ELo2cxUzzv
mojXF3wKswM5JEupK6R7DtlkVfAfq4XbfhNDS2O9fFNfaTRRqw/UiScRHyEhiOptY8fEsaKl/20Y
YFMtxJ6QJWReGPouq9ZiLq9Yxnq16JXVXqkeNQ37J4lhBz695pgvz69HJ2672smr1p/dCmMYNQxU
wnGw73CMKL0KfiYm6VO0nwMLYdVvrZKSM7T4jwuXcNzf/4eAMKM92xkfAOpR9OcSqs7RKETdKhD5
U5e9YagprZxFX+r31orFMHT4p8r7Ke4rZyKM6l9MvZ4Wd1XaICLlVPs+i2AhYPAuzvZ09Drr4+LP
9OaFHu0u76AaYXRUqo+lAToGFE9548DHudLMag9diyaz1ntFCKw1T8/hlIgJRu7tDM+IUQREokEn
/Xw0kfZZ6JPNc1XmMV1GsEoDN4njMjPZ41kfsHmegVbmcNmDxYu8Xq04xBo0jjfzzF8RApWItTTf
55Bo0BDYRmOERlQGO8AkPa85cDiDEbqhqunzRWRchNWAtVgbjWXCNvo6POW4Jpb8gzZTq3K/R8QU
YQzTuF8MHiMp484N3Hyii87+sMacIYYi0+SJE5WiR8fZdSs1UPQWlk8qD79lZ8QyHxXLM25/DMX8
IKPLKBxipzFsUy6owfgK5d6qkfFUeCnmP1pskyDB2ZhYIok5nvsPypjV22FM91wiocKWNVWs6Z2F
0Uw8XT0MunkNXlucI8WWKaysNuHlICFHJ+KmNf2vWcXBJuxbmr9sguwguif4rOsjCsDCqAyIMUyu
o0zyxjhGcOFYwC3VELXv+gNxyd3ZJb9oJAK61e1dlDz/QfRLo+1SZEjMVhcuijmaEFNVekDqCYWg
2BFt5UXgiT6E75SpSeIpTaVEKBrKGIsJsmfsIZ5PTuBlWJrSiwew6+PrBEPSJqM8IIa3TeqKma2Q
/pcZxgDxYMYPTAWh98eDgYYaAOMcu/uh4ZTX6PmdOR3EDGvR0eg9p73UDuUbN2oNEAE+JBmgE5ce
m9TS+LkDub6+nuU2vN6PmcdUcD1QkXn+nsbRfOazbuHHw8rKgSvZptoiSCqh/FIyJhfr1hnEcQjl
RbiKZYiMdzezhFqRikS3hHa0GElKl4n0Ls4JrmYrIx/rRjV+Q1OVAhnM3+QTLwWpzcATqKy49g3O
UHEKrDJRKnk28AhgzcXU9sWBJ8Qj5teY0fRL+RynP6clM3auRiXv0W20wkF3zwuItWD6hAz7MQFh
Wv+nESlK3boofatzEGkZlYRv+8f+nf4/qSOtLAzdbPcH4h5Ey06mGeAb+N5nExXOnpwreN18S+AE
YYsUcEoePS2c3iR7nrusXL31VZdJfhGJBRpDgUY3VRi/Cn4FhVUBF4QDiysiU2E/n8dCpYxNRKwF
mS1y7lj9xe9g7qc6XU3RCarLWEHGGHEyNcpfFxhBr103sLRwYFwYwIo5oOJSeBtR72WgGjxlKb4R
95ohCaiqHqujZKV+kvx46Y5uPbGX46Qm5cr3lSS+m5uzJIP61JD+RdGF+goP5j8gHaufKIZ1fyCw
GyI9Kw9zJ9xUDTFPpIqWwVzDUWv1gyZ95+luhZig2nrOMc5U1hn0u8RbuZ/2Uh2zZqdBp1rBVlsC
yz7v6TWEo/IFy1I5TVHbRIXowXeXpOr5eUl2JGq0/5ANL9Y7GrJJoc33HzwAI5fqoMQWrlGkMWJg
kIB4UgPmXAlcBV6O+tk1WxrN2ayvzF8TC/RX4R2h3pFV24mwazp3MnP+d91rnwGh/9bdiDp/1boC
ut3FMPWOYUiQfGVaeDSNWmXpINjbkvg6vzJw0WYViybItLw5JnVs2oXSXViUuUKrF2eWcVRIhIqI
9yByXIzeN70DiwFsJdl56y0r9A+1IleIyALrZPecYLz0SLz01sHEpiglWpTGTwFZ3kxeEZHh7/cN
a9sCtY0Uieh/agu4ZLy0DnP1xautrXHVqFbbqW60LUmd9Ddx8kFXSD8vlFfD42Xpx7NPv4mNWxGm
TtUitAEUhuq1ssXVFc0cjT9Ti35Qvsk8cHUp9eMyTxsHlm5go5rKxwqFMqBMGbSZo7r9KajVGrch
lrEPc4DFxH0QsVJBNoEclCsSZjgbwCoSnwFAFeKnEgHLCZfkmVCesAMPnoRQiVfXROsOCoNPrJ+4
EhtpSgWYZQfbaO9yVyjF8tvC8HKvFXrHhg/B2cDNlK87MuIK3OCvT4kJOwMCMrq/3Imo/w+KUXmB
lsZFsvHFoE4AMtOiWRr+YM/7K7Gvl1LDDLO//p5tqnX1NOxKvy2kgtOlqTentfrQXOCnhQtWk+di
h7hxCviRyOo2pcAfxlVejg19JGzykvM4lZSMWDCy36uR17r0aVGirx/G13vQPgx1yPXOSCZrQSnW
2bzvzVgnEkvfqArTR+GAKtI3O0oLWuITmJdAvri9FpWpAmeTxhnse1/rFpDtRh7FWzb3474VcIk8
J4FEde0sUgNpuJmhfmSk/WX/AxZ+gD4JmKdmPsqSUQruMMkMmcwucFKUDYVJkSXoDL3yjHbPwJcj
c0JdhnH0frtpWoIwPRyMs8CtB68RdSYiJanTO3uBT+6z2yjRWCzoKw9kEiqvU4qZapLqV33N00Q0
/R983Q1JeWm9VL3lq2lZJ9SSfVVxtlUpWKdkPVVA1XiRWGmeBmbFZVM7YkmCKkHZ127ItprhD9Rc
71TNrbL78YzxIg4WO07yTyOBZg8lRReQsk3eOqSyVSV0YTCFOL7MdtgIftre4nsia/Jqy4AK39g5
bI2RgMcgTLu1oMf/n0TJo0GxWLN1wdTCjA7OFwds5FOo/nfSJ1oxgK3TPdBK1f90/T67f6foJ7pF
gkpL2YYt6phatoolOiXwB1T4uf27B/RWQwUHJbVppD7Zu4PYgkvp0ejpDixfSqt2a/lA21061KQS
1KFNiA8VdxvYfRdur/WiPhiQJzN9erWd6WrtQjwUhDpAPBXacDdHLDTBRIzUA6D9tfRIKo4JIibC
1ZBXhhTX42tJh5x5hwCvEYY0T/jutqJZspX/wGwxhtp/Myjc1nIATBXaDhY9dthXQaMqlnl4Olde
dZvvtvAzcREjaFCzTqt0rzKUk4QOxma0rDJOIFXCFStTPqfesEtOCZhmsk9UuSQ21eQsEe9qE5Kp
MEqU2RpEIh6vd13IzrxpVUy/Qm75ZvktBCpwSUxp23lilt9K2wg8hX9a1GINVUhaIohRcGx4/Nvd
vKFMYx+x2kd5AOQCRZ+bZePH8ZcPMrDI0tHX8Uo2+zbXL83hHmUWBeh8/9GI+tN0hi2ZaESgV7Sm
YxYh/JeHsf/8BYmOvDlG/wMe2Q7BiyODvo5tR6plN9vjG8f40kyYjWyq//1O70PRyM1tqJOEyfgF
p4mS1uoVtBCa+c0GeT5/au7lCYVdyWaComgsOuRxE3QD4vudBg4zoTSFSqFTxJ+5lBOnhWD3y1on
CxBAi1qVkmMx89wGQok13UtNkio5kJORPHSnPyKRkX0bcTXxzL9gxjx+9pU9TPAUEnFNhN5a5Q86
aI2Y4H+afH7/YyJ3bTuM0xFXj1touxa9JVuJX62ziPfN0lnBzVIe/WOR5A1y4LQxfaV4Wu5Z1RcF
fm3xppNMxFTUWfeinAPbpl9ze9XVynZG7wHFBFthbDoEi334SYXe7NiSz366ZNxKPLI6zPupyL8f
op+vKOerlJ5uZV5zaUl6cLTP5Zd/db/EFIlkq89gn5QEiRo5L0bQWtK2yYozKODwKbwBA7MKHo13
2/kg3DYpxbFpXTjJ4JaOzXhaiVP2WfXkL9TcwQZ7uY0Ejs/x1hprtALzjD55GN0F/lC11SAAfPfL
e35DUNdzrwVcncRNxqsXUud89T6eXw5TVP3XkVJsAsH+mCCSI+PaFNr0rGr/azpMzvuWqy8YDBBx
ybei5ISo3PoKfw2o7ZLWrqWbHu1J4OvCLPwue55pgQ2uZxJ4qrc3fvQbHHVYdoEcYWQBxMv5L7Se
r69gU0JOVjrWhFawOOrGCjHSXbiE2mIlOmoeO5PCjYYg5Jafkecya3J9JWhKGKM7gO56+gyZ6Nft
Mm19mNOHO/00LTkz8eCDuehMSzNzMG0MpEXwSsUGpL+HO/t4EuPbGfARVL7HFIv9iU7CFL2+wLF9
TOyrqCNM1Zzv6OuufwS95Ox/HlW4D9GRTi4s+CTi+cP8caWonla4ZHfMzx2pHZzCcDVe7yiMKr0u
QWdjgwkDJsbVaoJiEs7l4aJfWmmiE695TrFkDmOHeuZAbLqWqOkLpX4ielbk2ltfiDQqFCHFFZOf
L89iCZEDsqnbR9Kj0EsKEKF+WusBok0EcC80yOyUdSC7SXOVov+pWO++HUgWL0pYtLbGA51kM1a5
yKHZn1gykGAcapHDHJBPW5Y68fX/Oh5OZWXyjnTzyroUWjdYNNS+QclnFQzc3TDxPnSHg2aAW0kp
ebIQQZ4PxlcnJnp1n/j9TQo1aDemCLWh5qEo1ooQXEqgAHkv4Mux/G+pizWc+bcH+JRrE60YWnTK
t4j2HEbVmQUadK8SUyXNaxZEIxxamnPP4k7b6ghCiVJ1/of4+MFO2oHQAFLSvm2MODyHtlsFQW0N
u4jLqWFYSX8FFP5QXtktB7/zzVQC38pl1663qfEQQIUDZcd8nkjS7qZ/H3JXoP1mc8ZUSBXNLZ6D
l4SCF3qrIDKu4ghWyeQt9EQGFcSxzt4P0KU1ChPuKVLcK/x4gKqSI+y9uzHUzpnYz4RF3KFMULAC
ANHtzeLXIkPU7OFW6RXDcnSFuJFXsDLgiMyzAqqA26FidC73DBIfPbS7DaxbvhDGIsqjH2JDo8yQ
yZc8vnwAglhDLgbUgKDcWJcueuwngPYXyOg+/UXDUtZRf5y8gv1gHO2Wuh59m4vvvFaC3Y45PcDz
BASfWSILBSyqu7j8Fs/+6anTaNYo7V6VpbJSt+NGFjC6sqpAnNewBfK1f9mdC9mmDOWDLfEJNKgJ
ueyVEXlniGNk2UMvtyUO5LYh5aaHNtVXV86MYGqdxnYFh5kAbuhjbXlfz9L5xkXdD4v+yxfVSuGw
mVIgx8fJYXt4LvzI32Yc8vEIeOp8dQnufZYuXrEyYaXYX2GzLfyd+XOmD00sawnFRUKaAtgoEQjH
agzQ0VMrIrCaDqbBfra9zWipkdWTwfsenbiM1ra3Vpxo33fftifFLTTpGnSrDposjvY/n8TUkP1X
xRWkYI89J7JqWY5ekKusgmXC/pfQmrTkpNPzkRARiVzcMd9ZWyKMB6yAg4I5Z1SIVDYTA9Gyk8eN
1vsWVGmuO/VYPfk3BFH/0XBbqrDWPpC6ceywkTXDo35MAVjtjfSklnc8HDvucpSYkiwPFmuJHknH
jTa1PMLrVJ12DeFLrvjUt99xr3p1KPrVsyt74FSQgDdy/h9QtWraNLI0Q+oSAcKKmcR33aGv5QlM
Q7P8opzRLUU5RFK8ueYCk3On49bjhjL4Z7gLAX2ngqsbPASJFHBxL/MGKwLJspHFV9n0ymQs1PJ9
li7KCc/4a+s8m6hyMM+Vpu9P0fb+GmHciYA3Ok1KNspM/3lcyR9wBSJphLGeFQ8Vc4oQF/XifCdD
CpLhGf7m1EKJEQDMVZNg83ENC3LD7HWZfdsWUEjWT2dQbh9y6IynOPVn716fn6DLAoSt8gIiAhqU
rwRRJlJsA7x7gMmLlIo9HpdkUpttTHbw84rUAVkSP3Vf2ghxGF6uXbxDVsoI2bnPVr92wrj6OtCU
tX1miZgrMlagA19PnGCWCprohq2FiYjBcbzWoPMY9dztOVWG2Qay6BIl4DRtyQC6VTmQS175VLcO
dbOYgxftJRJUIHe+B9sDvrtmOYMtwXdoO0Gqc3SVc3Hhq0acyYvMh1bWyQ5H5JPqo0GGFkUvQfN4
U0tKcjTi0JHqNZclkgnHEm/+tFdteUiD2ImtA22kiq3Y4pfwmzSfoEigH7TixHPwa/EGmIM++acT
MqFAeiMBAzpb2ImN6FiFHC6DCbt1F7wX6lE1HgjFmTuJhKp+NeN8mDgqDikSyu4VD/+gVen9oNW5
i0f5AJ1FbeMP5tQAbLFnrBdVzXjbISa5SvbqdlggDsImO8T2cQMkIBzunZFXl9kpRnO+AmHP2hWb
rhvf4NrwHe9oZUyHsF/M8ksL+zJovhdXDfro5JYwZn0tNSwgVnu9EUjU3RzWZyM8XE+IBVinobKK
XQMnbPHGr2MWd/ryd5yLyOI+ghnhB20p9YMWpOqkzgY0NbszZlH2xHUy7YTHLRCBt7xfwRpoMENg
esarb2Pr0w4HzedKgA8VX1ooM7+LBaoAhcTDARP0nn3YbumB9PS/dG8hY8o/t9dB2bmRgRGSUtmQ
Ozj5HKpgPuV+dnYmvJ/Mei2KYMBGtPxO6rU2iS6Ook6S3IA5RgFw4hOla6qflgpH8PVDHsJqbTdT
ZXlottgQPqMzAEjSTfgvMeqYyUOxWsfYRJweFxnfxi4ewhgQUZ0cQsY/9yJuaKWp7PP02XF/9bjz
TVROwjfU4RwGIAvNasXoC3HngRD9XDV81SL/ms3kdcJY5dyKNGyFw5+wnz5zEuUg9VtTLxQugxOe
sOF9Og38px/oR20aZDLa7UsSZSYfD5XkQ1vfjVXvZg1HqJ5DdY1etwRRpxUOnIt7DKyD1qxXDPpn
Qt++tyz25PwM2H3gJ6UCESux1px0qWU1s6uVLcQ354Y+yfOTSZXZoLDTnzU4Gw6NfoKOcoOrI4w7
WFNLODdmBMOBrl1hgIeOQcaACSBHKRIYsdYGx2yiABYK8sUIManhkyWyz5iMD6IiOiRYW/+dziAm
VGIJARoi1jaOcNzgXdpQZEx43i+f13E3QZ/28WEgYkH1y/n/tgFrRkqWyAinJRADU5kNGh48ZBN5
D4X1cQwbXOHE6S5TduVqhwqR/hZpR4xCP/tcl6G4PMAdiAy5ScJqEImtKZGSkXkzi+9Cs3lrYpH9
94E3jA/697bd60Qq3XF21kNmsSxQTG+iAHUQffe8i23RY2FrTh5p/xXiFwS4JFiumzx+ki9p1nIs
5yW5Rfi5kfyobMJHJTaq5RStcRj+9i+p9p1ftYFFf1/4vOxjiQb5bqK/9kshsPWC3Xfk1bluanHJ
3Dx/ImLziXBe9hAqa56oHl6h5fQces7ycd0wWWsxMAJBNtuEWpe4+AvSfRIHCMI0vxPBHW8AJ2U7
1Tf+/0iaRmMvO8gLwjwtHcl0WSAFOU5DkSyC0OgOY5Jew/kXHWj/6l9stpO5ZLJP6pLoFqQqKGOT
W/igAgqov4kabf7yS5TzmhcY8ccktQLITtrylgQigPgyV71Ky4qtXdUcRxDsC1j9w+dN4VLm5SzA
8VEMnB9vvsHKphaWMqb0EAYE+dKcQeaX3H0On/NgOkA67FubPSgMgIOyKuoVuK+C0rgnoBx/PgHz
UpEc/AluimHHZDUw6JIoFUgjmzFvYHMvDrbwB3rB17/ckfXa2zcnt6bGcjndxVzXFOMC7tP9x6sK
lMA0m+B8RXdO4DI4jxf3z4GP7djSo6ix0Y1cdZ3e2G1N5kLf4SmXXplePaIZhL/oZXvLsa+sX8Jk
6U2JBV3GwFNrLF7RhHTQYUusa/QmomBXsBio0s0bDogpT8+a5q2GlNd7hDbNXML4MB7nDtiqnC2q
tmiVoiiKxFByOrdfG98lk+ySEyhuoyVamho8PtUAU1tBb9mkh8nMqGkOrbh1vs3Nx54KhMHL+DSc
U/mjcpXW6Mk/+QzWmjJcB20oDLpGwvxvq4JdSZrWtHLHoLwR+h255dqt6cS3se5mtRlTD7rrom3Y
GVfMxBFs1cxWkHx5qkfQFtRbzEbpUwhxzAzeJF+j6xWnRXdS20UnwC5PXMcobaKjdO0JoJiHYg0h
dTGOn6xgdDjukN8TPgPOlhj+Bwm7pd6/QIGmJrGk36pSvBi5Cne8WckcD7DzQWSqzvros5cOXRrb
RVYP2TXC34p3D7BYRB1HEpwVxvH4xoYN9o+8TSFWUZjfFXK1utEGxuXbpwMReSztxaLmKEidfxZd
ANKU8gNlsj8VeIDk5ywthmJ9cIGbQ0VkpbqESuQiq+ClDwniDone5mAWiTq0oSv+9uPjqCxwHQi4
xL07FSwkUWN3nPjWh/8qcf/IjRVMWnDm919A8M+tnJeGP7Tg2tme2ROjCbvysNNCkO1KZxcUYmCZ
CQWQz3NcE2WNLZ3HCZ/zUG5VDKZlYqaiEswNfnQbWUo92eX4FuT3zzWoU17I4sNnz/TrMbV1uEO2
/BzHCcEsaKE5coVUfwoBbXCm0voqUsH3q9kPfzlFK0m3+o8A/I8lEj58Keg0Yr3XezLdbzVQzd/h
w0KCimc5WfHQ6e77rhaaDFfhSs6/WwdAzMQG6HN9BO7QxQWc8ZNnt66QBMZlwjlIdyssWfqsZYJF
6pGpy7+HOBqp0m8z3cOVrUhh12lAHWkNJo1LDTYQI6j/Xk3SWjmypexud+UvMruGtWtr9JJNiYad
/Xd4ilwK5YVgYVVEQuNvz9UzgjBb4kwWRrD0FRPFkoIUjtlBGda2rOlJ0j+PcX+3+HSBeDxgp8VO
RBBwZWt6Us9u8fepbVtQUhVXzXUIyNFqU89oJmvcUgxHxjvDt8OK583y8N8vw7edxEzhHpsLbN29
3M6LSDQ6CxAq7Px7//zJ1GEmWu1xq9SBfxsNlni2yNs5omG4zNt1PR0VmYeA3BZq4w4zPwWQTxgF
kHuFbzcjD5XGkWcBnEFiA5bs+5pOhxwYTwon1MWr0LWp2bt3A/jl5TI9Gjm9GdIALgZ2beLkfB8G
e6q7z8Axu2xTto7CdODm5xOSXs+UQgUiSzwC2M6+c6M+vMnPcmR3ROmYgLtfccm35071Qop96LCD
QtxVdB6FgHscCorXFfKB4bMRTjOYGNAbRX4KF2p65rRpWEUfpPExhLQx3kHd+JwH55+W2mqV9AN6
StI+PVMeSnOSbAf2vMusIU9ubEUQgZgnOsXjgSE0UX+bGm9l9Rp8iUfBoYZbEKWF7cOPa7JnVxGK
ML43lbqutHLCQGpxzaBpwa3v/DvNy8GPeqGn6s2+NBrOlfaEr6WVoXDcB0StS6Ht45wgfynyENNU
ogVQkOkNpXKohLOP5rPbfLlydYtVfoy6h/9KlhNE6RATQfEE8mi6VaL1NLSj04DGnPORjBhZjzoF
LOt5WhOf3/d5PFVhPlvNFvXkKsPzNA03hJHkCyw3hR18FxrUfYSXZoJ+oA7R4SnW8jzO1hM3e4YS
96AXcNrWkWOkZmdVzTeHxFEja6gHkVgLoZ+9C/rRSKdfjmjlPK8OR3qa4G5OryDf/yB78k+sDZLj
v0/a5OwmZdVWin/ifJVSraDfuJsLsPSyr84cfEvEqo/foDPb03sE7HeXkl/0unBIHIoVqISC8oLa
WLef6kAWCLEgnZi5IT1IIPHAaW+d2cKBD55xsnLXcsPuaSEhAxOfPRhurFn0EAAMdF1l7auSWqgv
1PqMw3sJpAEh03+ocISz7a72dWupEFnrMM3A1A4d18h/4UiA5qfegwBpyvEbNMZM3yPziWSE2lKq
ckWDOh/0FhnyMakPRuizKlnT9x/2Z5IyFNGlpRgerJXM8orkkENMrOS2+o2a+zMsLVHsvQDfbOSh
OPEBD4/n3hwynD1Jprgw0kqK2IHpmdAnVoccjs5k2erY5K6hxoWPT+okKeA0SYxEkbyLgioJiHxm
99d5I1TjEj3OpJbVXKu54xuWJDtj1pjl0ituzmSzhz3V7lE6qfkf5gAJoaXIteMSzKk7U6QJVwJt
FRqw48GuFWrSkVh4DY2UJljVWujzUBbsu86fMN6IDE6TmMw3EjtzOKBY0yk9AJeFnpLXgrNuBkXM
sHbVLn4A1C6jSsBRJIv6VbBGPVgCl8wWMT3bx3MzDKy1bzE1BHHt4IiTExX4nF/RYcu4sqUoq/Ri
Hhegos/G0EFtKVHPh8nZVRvzHcu+Fk+gXRinH18H1fm0nGFa/SIULdOLHpB+10gNaHG4/C/QCZO9
pAQ6gP6jGbS1hRMdjXj5ctTRKFYPW+gn3XEIlc83/7vmpVmnCKhqieFQr48hqAG4mKSJ7Xj3Nohw
tWmu/v9gZhHNbgBGBKEjQAcbomkmuHg7SQ6j0j1uayXrAJHGA2a/QZaXl7VT7eHjxBWXJ6vH5qGw
+IjeGbV68cPRdfKV/JkbEsduKceus7UHbt4FA0l8iCqtrMU2DHhZHUah4bq1naniQK/ggw6OV3rB
EguOfSMZmsn605L2mbow4r45SWKlbxriNkSBVyRR39b9cP/PR3GP0MVoeq8NNgNuzgjmk10QB2Mb
AtUh7pFt+6MuqyhfWZfA5PLOBBMAvpyCy+Agcj1gMq+0Nxxa5eVquJEmurEcV5U5gyztDJARgLti
+IlNRc+dDR+rOTb3d0q7sHpsRncQ44K7cWC8YKU1qJ4fuEjOwgLKsBPjGVvCLJ9dGB59G5UluU0z
IheJcOOSndzY3XgMFGmhs0I2cH4YUzX0AtkGBOkmDmA8ngHN8jcSUh41Z8W6qUfELoJgqKtOYA2G
iIEKprcxtoRyUO1yTjV3t98Vh3b+0mLffnYIs8TpIbCFLBIF/iPgPljd/zjqH2Y2g12kJrO8+ijg
uUsACy3WOuOvG504cFBIl3uO1sZYmm2d8AoGFLaSSsgtMjOHNIB9gvXEwsQgYU3oRsNgBcFTAaq6
KweuDe3upJpwP1/LWRIw0GHl73nsRmdv0bP+zeG7lZBsJTcLqETYCuub2KE3bPazmScHNaux0pVk
WZd3IJsyuVP7DcBc9ieR96zrt9lE2ls0J/rBPHtcJ9kRRXhn8sKPmleIf0MaAsOWBezOVvJa6c8f
eC3Gy4ShVO5+GYw7j2vapTIKG9jE9RdIDEzQYGdu1zFmPK553/12pTKEyFdsDizMn7vFBVGBsms5
LhaTO4I5RADa4hYkPGzQg7QRT/iUVDpMyvAVbmySpXedd4o2wEIxCfmRNNcqpy6VBAlJvvRqFppa
2vKGhKO5qg8RqW2vHMak+9lc1dA+xyc2117i6NXcqaP3bwFgIvRRWXPil0cxuGC9Dbb4eTOUZbRy
6s+nmjF3FtiN+swxnOsZUj6DdYNpmzO5FCBeebbsZU/uBpiQpPPj/d3DxTMBeegI3bDO2RmgdrnS
13IegEoLYsLhGqtqb/iTo+on8V79Z9lN9NbcZ99Yp5R/31tOO50ZsGyUR/YW1ziIpA7UC0wTywjL
ezkw4w/s5Io8bbk6qUYnc3cXk8Xbsef/ayIqfTag0JOzXpXtor4BSYgd8ePU0yZsoLbUkdDJabuC
k+3CjSEIoYeB4JtDbAIWILMbn95Kq4EZ9L1pA4VJpLK2J872k01UWIN7PpvoaWJCOv26ih2i5T2z
4UpdvZaY8CgFf6A7BUFa6/bsDJBJfJrLI2t94rJBvCS2JqcJnR7xWSD277aRHXZjMZR7HI3v6tBX
JznfHPPhAYJ8n5JYNHV0ZnFam5YE56kL3zjilgvRe9ZePKEEOkcDw+25yEkCj4pzM2orxoKlD2ef
/54MHFHcA6ZrUjavUCFrrJuPhSuza4WsDyWHSqYcJ8ABk+3ooI8Uf4f78ENlQriZ0BTzCy86gXnH
/Z54zpstnndjgrtKNBKwsVrt+xfeybRLdUUxvLTBAkG2JChRGTHRAunq0bQFh6ZwIyxA1SWLNmKW
SIR3NaJ9eAUOfyWnbxKQhs+T4rlLqaxU/cXreFJ6fsljTKw3blLPFQNkby1LWehi18ejy0Rl+TnZ
h1lATjtYk8BNMzIaMwHt5t1SUxfpp9Wd7Nf6gZlvIT1PWm8Fyg8ahpfgycMzzOF8JePhKVvbxdX1
f0K8TLKnjPTn/L7zcTf72FC86N02Dx0RrqVQpDo9gn48L7ilDGDlqkyQi+zSqLlwcm3whsJ4bGOR
Nz25ISow5SuvwW/UlrBVoSqWFuUTJ58072ORGyzXiJqgdC3B7FEl09KNPvA9scTA15RPGNASjJzN
KWhKE8mGITWuUTJhISvLUrYBLYM19OaHkHbM5jAr/k+TSdBshpYF2Wg/EDvwNzwBzTcex+Jm2wZG
IYaH4qi55XPd855BZyfjxZZZUuSXBvuJcAlFSdNBrr+A1Mi9zomCW5pGJZQcU9Cpo4Gqwp+s6O0B
GY6DVUJiboEbgprg+L4PkSPsUGtlPMTKLYGpuZc1IJdT0SQ6VVpoRXcyfCfRfy+Id2tFRxm1BmHc
272SsAlkGyamM+TkQzXD4E9zFTWqrRFTdJJrs894Oabtn6jLWP4Y1B1q+7NJTsdXjSIc5X5zHqK7
nUCpnN9mivj99MuEkLl/bwFyJxZR8PxRZ3Km4VdVFbiE+FBzC/knApw9ICvAivQctnLIeSGMTRwz
bNghvC5ExetjpD+c9YH/pl8Um+FrOeUPbjhTxnU2M4n0lUnsSPxBPJN5rQaHJhs73F8+gjTEE8i0
CGm4ufDMUFJjcY9uoOtg1e6MFtBUX/46uRK3iHwhyaP64EmBa72b6q1XDD+hFe/gPigeuAfVIJuO
wYrH1CMhH3LzNWsu3+rNV69xLtTi6WIK7WbFQprOXrVrYQaC3y5bxgreaciGyJ8yRqGrwlNoUcoQ
s1fTTW6YfNExatQuontOlIGtC0dUyhZeIBXq1Qv/h+kazFKFJrWWXlrRKWomeUXQfby7mKrzIBhb
4XtDh7L2idbcq7D3T4ZwORW1OG5IOwnDteR9JunxkA5PryMBhathG88Y2KdZbKQ8OQKAVMhKj0oK
/pj7a5kNFJfyfkPZJi69qxJcx6rJg2q7AGAKOKUkNEcrK5f45Lh78pM4TGvmmtdU8N5xaFWzkNok
OkhP3MYVwL48/FCuxC83QQIPU2Koi+kvlTlrk/Dcz0XbvJDXclywI8k275fVNSf6YTxfmnXXlvxM
US8Ju7VIGquEN5q7FjN7mKdZr9VOVYgpsueKf4sowxJxyuO5imDNF88g5FwfOnciAe4Vmwvmnpcr
bFBiYpo1jYpt5UNm9EBVDuYwuA1ogBQxQgNEnV5sxOsOV8PIsudvQAfe3o4jUrZYv3X/8DDLqENU
9dLBYJ+0M68V+DJjuRyJFjtnu6haw3UQ9PVtBKgPrX6qWidWFuk8yvRQf+PGqDKBDtNfevZWRoQB
JGJLQEHBM1VEMQHZvKXMc2gJhQzlK1yWSyNMpsZfQOzP+a2NO+yFKnbsuaSkfb6qJATv1LaPmC0P
QQEpX7n0mE13QVJShKN7bxjg1tttEcgeDOwm2ro2Cmm/Ep13p7/vh9jZyGIarrx8WXb91oeteU5I
8UmbsqNa/DZdYaZsyWE5Jr+yDz7RqtgCg2z3kBqCLkUJoURtsDNxc8TqfPxTBSIZnfuzetdg5qsm
5Am+7UTUGFPTd6YQKj37mBw3IuoBVQYz6ca9jefuxHklWHc2q1O4LvX6h5vGfTtCrFRUukXNsZ/w
hn1iaLho4raDJJR//xtLMzUTt75N9dtvTe4YtldUAYI3nJibNYLGap18Qn/k844AF98SJvYzCpzR
4e/th4v4i8VyLHBJpGtSXrAyR13Cu8uf9O2a+OatltjzExQE3g33pekC7fa/aCCfzQG5t4D0N9S+
hiM9s4/RVsJ36ctx1CYwZ4CCLMuSbSuMCtFeBoEmfFEio6Y88fu7++N9izNFJqVUJ6FrBx8axGXf
RGIiKysIyisIpFmMnV1YpTyTOicWUSOQObAkQXdHU5lVpF1/DYbtzBD4ETlhsanQCT+1juPsSRgi
YNHGd6osbkghzq3Ky7M61vkbwKpK60cjqt0uHonLFrwdLl488iFBq2IgiCYgjvKsKRKrPd6NlMeH
vnPTYnU9LGUQlnvvkjqILEAYAyV9GPo9vZ40hah2JRkn6+0Jf4/rt2FCAdXZdbbTEAzBhmadl8T0
NweslHmV9ACAVF4a84CDcFztA7KsL20XvMzTr1lVEYAGgXMdd0XnBBU2gR7kgE6BU2AMb0XOLATx
CjJiKMQa3TIeGnGeKbLkIbFI8msICFlWlYRzLmREgd5+pYQhXYCU+snOfxQJ925Zu+HP/eFfKRYS
egJKX2W+WF4niHcFZmiwEZ7tdwv0pESS+rxa7Qqt6cW46/JVfoxiW+LDc1aGT/ingcJTpK5Cuq+S
Cxx/FIZ2QsXHcQa19fwblmx4ubCVlwnGINjx4QWsCG8j+R4YVMaHSE1nk3qj5FX/yU4DvAc/Zkjk
OduN9iamIykhtLZ7TCEiC+oRu3PhB0gb8yLtyLfg76Ao1Ng9qeiQtiwTPSO7FiacjMz9XbMw35Vz
Zso7Fg7RlrqfHTVkBYudOLuIBIfktk7C+e3nv/7ep9FCzW/IA0f/i0W0sXkEKQWup31D2irkYyrw
z+vl+EzAcoaaIBWbvjrPWh6TAT8KZdSwK+7nTk7k7MhSEZDh39k4wl04raev3S46QTOBpbeQARXS
bktarjAclQGw31uZt+3e4AFpS/IrSyTnbU6QipEiH52aL1xwK9He0bwYIdJ8QQ5lPZY6Ji41J8Vm
QzeIOs3AqdirF6cqAtRN/mx1vqGl0lWYgP2mQUGqZ7OwdN6xJYG0uLVrtcIMmF4v2nt2DoGQuQxP
neFCsEnL1zNpvFDeABpGDxhXw8nnJ5QYeYoNOVhJrpk/xtbD0By7rKDeELeGdskADtPOC1L1FzT2
WpAxPH0tbJlPNrRwDhpPrR1LXN/QFiqZvScJaVMb+xXjHnG5B9zZRwt1ENI4RhtTWhpCYpCeW+RE
KBDxoN1x5IKooO5UapK85IpEubB6cqtEZ+NMVBhXzFhr2kz3gYZQuhmbg8UxoBJcOexlr4ZZwfuz
Ey2jgtFiZNH+dPNVovACPDVWGZWRtB9s3BV/GTFELpvTg6G2rjo7tu2zs91vmb+X76wI/3QLdjeu
PzhbsqVd5yRqOwYDJQNl6jV90cH7HFTHfqXCy4ucGcmC445Pq1SgzUjX8NA07HsZ4dgXuis5MA7i
JY7JWacVazYCW1lIiV+C7Ewic2H6Sm3R7H27YG20igpNiyS/cEdvdsRACYc2NnHUtVi/DDg7Y8qQ
JLyunDU2sL55bK6YeC9eaeWIbsRNdBKjAhk9R44a/2ipFHm1UJ3Fe0UamXZMW69d1Z6oa+atEFUN
71Rc3UIRRdh373TEG1BXlAdwuLiqH3o89oyPWsPu+x1IlYsSF5YOma4YleF69v9KQKW5PiD8TwFF
Z0qqrJfk/v4/AuUidCq8jUhG3zuNsAa4Iq4U7cNBEecy4busc0zDgsMETFSaWXBAGRQf+f65/3GS
U6Zgs/UazJgqVyOQZqsbRN+WrngIn3dlUwgXHswhUxATjGDPle+ouCvXAzYrwSDOhc3xkxTrM/lr
+VVV/r5mfoMTBikeBHqvEJuaI7QrjPIjVhKGKhNeqLYhNHIa65i9+k3YtzfDJIb+jTMB9cn55Fq+
e6i9oqMJpP4h4ax4IEJVHr1Pwerh9sxilYSV7yEXuXv37SSIf6tr/eqsLuib7EqjK2W55pJ8mmmw
n2Tw8v3V4Sew7h4OAOjqV/NN0TxmtPBQ9re2uQNDp+D/fMy6aDGRzsBTC0i+WtdVacXaKeGVrM8O
WxtNt8Ypr/giMLe/1A41pax8SpnlAjum226w35EwlsEfUX/VG/Z5ZRDaGjhPp4vozKelL9DWfZ1S
RreImNtk8OZckHnxLs4M1jPbP8cbBrq+KFp8Pe0dgb7oS4wYvobcrP7JQP40DKNJzXLhK9VSWvbH
6RXt41uJhr2xSQAfekL0rr2idv2MKylpjF3IsCR/55OlDkbEjtqMNIPEuRcCu7uKkaPYUueHsl20
amVFZTeiztL4hUqxsywUDfrae+Hu8iGGA/cdr4sxxkGrgbtRw7hdHPCKS29KaLOFUHpYqvsOwMHi
hmv9urQTVrJ4bGY81Vdml5+qzJwcROwdvUwevnwzKQF3JLlQW/uLJfQ3Up2QYCndZ1fWHZgCrujs
hTpmgPMMpXOqgxbhZG59OyKR4zBlxkb5PqUNQdOUH/KLaWW3iuofJNwtZnogtAK49m1ke4SuHm/z
ZhTY3vBT6xr0d6ALovtuamPgcgw3vxpbJ0f65uPfA/DQV0eyJ4D3iy6lzvRk5PNL9sI7wTa7YTwQ
bl+iAKa5gNJE7H2nZ3tQiiJgIK4anRI45uchms945QrjE1nw47JbB+ClnnKnqkRjOhbFgV30xLh6
861Kf+UVE7UcP/lUyDAKPllBc3aCBcYCx75YDA74peFDfIJQ/1yYtKh65gmT5uiNPm9zn/4wyOL0
fS3acwRQcOzvETeZEEDdsX5sHd4sDfKVhnqIOYtSOTqAcMTy0nYrkgjcYjGc+6ZiAqNHl/QeqBGK
blTaWFXg2Che2U7Fxny7nfXfeft9aVXsH8oMgV1T6Fjiq6G+6htUqaFH6i8CwT/ItUZRodUnkjXw
/xiA+gepco8fPSoJ9+GHsfWsBblTkjqyogkixXW2cSZE8BFVvyQzt1JlL+qPeiqQauTqCHvDhtBx
HH+C5Btd81Mf5nC+1LSpOpVUrqSbwHFi8w0z4ewmshc/5eSIH+bHslOLnGJTiRQy0TYMJ20Mc96U
4ip8tJoWIk1xTZJ1u+tuXbW5SQAVTbPTM0nAJq7HpnUCpOihn4SRv7V5v1kAeexYy7dzh2hNXO7N
BlVnWE0tO05Xa03POUyHQrM5zOSaVsYiA9M8C7VNzSG/YvNF/mt6KN6d32Ld8PmE1cklSyXQrXzT
8BJ2tJRu2SmwOCwYiwg36WRmACoucy477Stn2Kuf7usq/NtHmo8+1dixLevYnda2i50/4JqD7Un5
UAL7Puq/rMJV05o6lwzkVS1hzWYKOl63yws5vedDGUi5Xum1sXtU5RIyLkBPlo4JB38k+SaZIkXt
IO+3ZlXeElunZp+ja+zXNMDjYiuWXxIa1+2hdGVfQv3Y8Lf6NGXKTCnE7nUhRcZ1laf0kTkdEvzm
uk1KxJGnOCebGz8d3kYhnAF56TSbfDG0H3z0z5dXIc1JWyCOvGprQuMS3scgfRX5/8Yv+F8w9d2b
8OI/GpE8QYssWsffKK6wNW7h4hnmhELlnmb41Rr73yop9Y2P7lELTWF7lmgNeRyvkOQ+pEvS+ZSu
ynAxRRE0aPOBRhqyWVSlnxdrC+wRRkiwd4JqTm+PhnD6sI+7csVGz1iGvwQ9LEWtALo7OJLCj0FU
a/DHMqMXSrFYdaUhWfLbbP/BJg47FzGITKA8xrENgLU3S1y+S+bSxH/IjIhgVwzGdeYCCQIF9DFe
jXmt60oIWJtnlXZ1I/lw05ee05M5Qgr6E25Ws1NWZYB8QIOmrsvflXphL3PBt5R06lydxt4CnV4N
zaWe8gQdq4nyxKZ+n8Z1f4TG8T3GRb8uB97jcRNzGjXej6G8m+LnRekq+WCFaXQAXM29LZifxzNh
Mj9fstBn4wZaSnXJium9JzqownljuoLJa/QQu2kZqxbYfMGRfM456vXX9Unm3tMgnzNFxRDsnVOe
7nV+H13P5jXywYxNQAPm7bxh4Gl34cCmY9uuv1pYT8Kd5Q0X86II26EdfIb5ao80niOMgXL39rCf
MraJcOEc3Qx1KYg7bV6GrQqDsSjo1Jpm7o2KT1HS27sOYFdkAUjxkFbl4ywUOKqBTlnt8FnVouXE
hHtQjtzoKHaPqjaGe2DRDyMKvZpLDSB5yaw/54SQ6nbr+hkt4VXIiKAzPJq00WZwyc9DvzymO0Rg
4/2R56AW4FaX5S81mWfnF/xsb5pmSv7tJgo4Ylglqwmlv/y0ouDAGV1DXNkLTrhYsu97bNupDfMT
JTMSHwGCPL6INXaR6/yS36s3GlXTrZTamjc64YyfNmJXFMEagRZnfgCPYWdYvKdszONexavdFseS
lt290naxP6SU+WA/GF8rQUB0l3OMWUlmy0t4xfNaQIUxDYYGN8sXLu09S+wr2ea3fClevzPOO4/B
r6n9vQEaBBfxuqd56x9bz8t77SsfG3nPyElhPtjXOk/G05aYQjW/MvtRh/hvYQwRlYHZEufq5lhG
JGKWD1TrGFRh5ySZu/sDpOkXb4SWYqKDCnrjDsf9LRzY0OAUHFcit5+N8HMbKizG0TuIOKbNiPUb
NB5xvomySf6Bf4QBORXcihf2PX2/zCU2vFRnh/y4YiKqM8XrUBxFXaZzw9wjzWR83E8n5Bf8LYah
4tl0lYjnQX4znCuc4XAagzQp1xAdrqiBxYgm0pV17rodCVQHsdn3QTquPb14qgWhDMBgEi3akiot
+e4HlPrp1rxcjIlRLv9d/035ffALJ1D1B4JCvEIaC78X3tqpIg9LMta/cfLE+O8tOnIIcn51C36Z
yeVfWVxNGeIzzWQbig4vKXB0lCDJkK+R5ElHtME0qVa4gIpmHMyYMb1wrJtjydH8lu2ks6TL1PRH
iyAtnh+B6OY3opl1MtF3wqcmVjPY6qHhjWOy5XVFL9DpD7nacX35fqEPycJUTS3W4dG36bNjy/dr
RsgFehbUWHzrLP9Ufq7Drl8YoyPboo8WLwaj4XK3fii4U8RKWVNZkXQFQ3jesMWKUjElnxj4SMgf
3N2aWMD3joMoDtfpm7Sdna1352CI3cFi/DZq+5eBgZlhIYHdxRkJleCuBoQ26m/pdojqGMZdiPx3
O0t2dCtbSIEvDoZJcjVJELvK8KH+9Xjjbu6L2l/EFV6ztdF0Im/6xlaXGFu2wwFBwodgN0N8f3Mc
nvDdd1aOkTpdDTIkEAIkqQf9OSNZNi8V1lDF9pNRsETV4LNBzjeiK7z1nbXOhfFfVDCl4kusOdEh
kTXWy1SxHdi+8CRToT2Xz7Da/46yxPW5BYLkjqmCTfnLxM5X+FEYWwgbEOd6MmlqlCJE1nuh3icb
NEJRcCY+kIVRgemiBn0C0/qPsUQF0SCG2ypjNb4/VYwwmAVORPvRSnlzkQpt0rxAoLx5xYJgM7Pq
MMuEg2vo3mypwVDZAKdwq1aX/s2VLEJrgBvNQfqGQo3raUnFVYyLfwC7+6aksXd9IP1vgimX9EfD
Jg/lOKaOMCYiUQhlWHVaUaQItL2Py2QR9n/Rj4c9Vyp5UKk/HRprCgqq9fjX2mMhvzM9Wa7FFO5V
mAbEcOIAV3IF2NBUp2qGC3jeSw8K4ao+fsnnWwFr8fhJ15kHz2u6z5Hj2QTuLGgCOnul7+jc8nFQ
JAC5Wp7Zw2yuNJgi47EfyFzG8agkl+rxiHk/mpMT7x2tMPDXenhAr+Eo0FSwPADVZXpKY8asdqda
eWKIzf382cKd1lKuXFqeuEkrqANj09Jf/r6pn6LB3MR3PUvsW4IhDiQaSgpMo8tb+wxOTfyoeh8a
3NhavueLY7rTcJEzkYOfJtN1+QIqT/LXVWjaC+KPKC96TFBCjh5PcEc7IUA5RBiH0sn2UkRzmAA9
bhuWKQlwnSL+v6IfemKziJDyl+ql5iiLRST3EKhSJahLSJrvGevqw7414nWUCO2nY/dj+NSzmHqf
XNRGlVZp2w1Kl/A1oDC3GDJFWw+R66NUBZZhHDbX/tklZi9kBRz1JCSAHMGywzl2VFWYvdtwkgKd
/Lxm6EDHi7sBCaCtDlrueWqn00QEp8Qq/ASX3ib/rEjGqJuFu10jqMmRZK5wcDg3IORgTU0+gegG
f9IPKq1QkVHFwPJOjZSVSPVS47L24UG8XRQjNDGCzskj+MVFU+Q9zArILmLnVaFw6AFhXUSTOQQz
PNJVJzYel2+oiNBNwwQ/ZVZoLyCzPC9grOXZofqxL4CxV1IACS3TdiYzh//DVOe1qYEIXEC+qmul
JHYi7hKXrFGzqfsrM9B5GAfxSWW2IC4M2o7ekliZ1kI0EF5qOJAv7nz8CwIpXWPTlLhvxYAfFtlb
cSYybfp1Fy5Dx0r5m/Hw7i9gnSGCQasKFc4xO3H8wX+3DHAWtVv+1Juo8oDvzmfL/V5yCiTtrU0z
1JKc7+vBkwTlPRUcEw3B7VqDOuS2n90svXYDLX/G1wsPxIlRJpLqep+9YlWqxNNKeJ6X93Ww/ZOY
yxeEM43B1XEQ8qozJny5TRFCw3etF7F38W0FHq7Ncpr6TFVAvrv6VRbIDSpTtEXEAJ/jnbgskUuc
OGTAvvfxaI5Oa5OrZTuWZ4zgxV1gWn5xQ/DVjeBWYJGlTCPQXQ3Yb7bETJzpysmzBJPIBGEyUOVl
fhYTaBWRzz8RWqQq19x4c9JTFEepcUeicjNOdj3/8DBL4QhbFOuG7R6GwFW83eUdc5G0b0/14y9H
5/l8CR5DvjN5t+WkItnw5kdkWYEj0WF4hkWvdas+j/akRbpB5B3tfOiv6f1XsOWcF6llGxRTPG9T
NjRmyhfT0jfDYVIUXaJZRPYLV5gKVIuqGcj8BbfwTmQbgDAR7x6d6GDOoJZIBpRYeKUsgY7bSQnZ
PW2AErOaRrURcAu55IMb2rRSUcKeI45gmJ1/Y0O3WaAAQWDy3zEbQS0b3qlx9doHRajjt9Riejqe
cwU84kQJD6+6odihPwetGbxNepGk4TYrB1MkVn6vBLO7GXL16v1iTbk7bBfrLyBQY1bxJlzY+6V0
IJHinTwBmtRAdUf4dKIudyOPJoDDZmL2NumPsZ5RhThFriscdIxuf8wdVGY4b47wUX9KUiH9ocV1
SvrZEiIXMZ/zJivganODeUQ06PZDI/7tI5ojS7XpkyG2XZB2mGZHOxD7qeDOxNpI1W2RMpE6tBF0
8M6W9YCV+kRsfle35nHl84wTh+G4a3sZO1WMyxaKS/R2oLRdP3lonDd5DUrIXoN0BeJuB80zTvph
1detvv5kbzPU3hFAdfpNU9Klmoebc84YIv6XEaKEtZqDg8qQ0iqemUwAY7Jv7zIJd2iMejEQXv8l
X8q4O/YdYVkCcbLqXJBc29R547GocsuvQ66TnmkAHrxaMGh+HUFfKj0PWnVoD6oX362cP9oDmaIp
1LILTr27AzE8bj5z7pvNTJldSpVndI3RMZFZyBBbMtm7vdJmGOc4aa95D0cu1OFhrxme8dofrPx4
zy74a2YZjQU2tCWj2w8rHPAo1scO0uGjlPl/eScnGYYMswSBPhMeFaGadtiYpo2QMUT4TXxzm19u
0QRIWvFrrzsL48pf/ON0cbW7uju7TuZr84LuARrNtMCZZB46vBVL7uDP3Rl1ZzKUymJn1RpyX9gX
LIdX4XtfdNGp9LWBZfaQiK169ezs3NrrQ07fesJq8ywSjrWqr3Ip5KKCl/3SuxAnvblqzWBquOGD
HGUkrXCyFWJuMgroaAkyGhZkrvjK/A+m2iS3T8EkkYLbr/N1IiC10blzr26r/z7/jfmRocN4bX5E
6zCnQlQ5poggvtgmAwiPErPSGKZWiKrwTmTt2AMnK+FTiY6PfveR79I3RAbWARvd+wanrXBcjdts
REbrzHRuysgygncE3D7vDBKq5JMMeTi6Fyc+8s9l6M4RDo6JLz5XTQXzfl6jQQZDYT0VMOq877fD
iFk5XvMBL+jAnkrYEbJPdLlVolaNbpbISlEorlNOrF8nHhQZEWVc63yVQuvPs0uJYFKUpdEfzcmM
hHcREwS/UTKVRRpvSgrssfJQthxf/TscyTpAMCPX/cBTgEM6F8zCKFLx1xJPODAOuSxuSmEljFQh
BaKh9zriGRJCtaFsz26S16pB/uz92QlTjmtziaXZzHko9R3doyLJEiQ29vm560FT6q4icR3qhkgN
EAWqawCNFLOwcBqSQsK62etf29H+7CKDfKVNrl+QgjBYLF8tOgFcx7NDRDGv36uFDwLmvjuwBnvk
ckp2PxxcphY9d52bmbFekV3f99sa8/lqu2yh8aQAb/yiSe1gzL6CR0sfLvBd7oy/RRsd60V8k74C
Ap2l6n371ho7Zqn9za+T01IhB85BEfmAOglw10mFYXLB0fNFPmxB1l+JeugVwyeVAfifNWX6Q7ku
kAYujNsmffCfbmYo0ry+ho41B4Sp/adci1DtC4LmkvahonyfNMgtlUmx8OyFtxlEY2p2pAfN0GvQ
2ljHnHEbgwdtfIVxdcRqPjaW/9EPpmWwblXVmMRWKUQLOkwScJjMUdjzZ4HsDJd4DAJxYH1927pA
bj9WMZMH7bANXT1jtbvYtbAYF0w5TOTmejdO1MVrIQ1RNhZmhqPmWLfu4jXG5ccfzuub5kJa3CvV
H7Dq5W1CGSyADsGMyhsgizyJGf437SpLZ2ZZpGWp9KP2xQS0x3SoUINYDZm09w7cu+t2q3/4aT7E
o+FUnlPBv3v7IWOI4JMNDtgMuDCD5UOamJ7bkECTKB/y28HgFXYum72mdiz2j5n+9o++E53IIKEg
uLpV7rK3eMFsHJksi8gkKF6J36mvoWJXB4C4M09ubMpypT/xaRcs6ObmYbiht/MGS/JsaVkOiEn3
CsWLKhewurEtZ7COihNfy0EBI45pCkW9fTHls3CGOW10xwJ6nZHLam6mNu0/LXmjR0wrBG7TYzUC
ggCMkwYGWNEhsTr55CaK8NNIuPtq/awnpuUttMIbCmdFc6fOZq9ppDtu8bH8m6A+asfqJJW3EGoe
62TrlZycoI5ljV/QwcZXoSb5UsbH0S1Sz6z7BH5rWhDnQ9smtGNm9slOrVvSXxV0k0GxU9Tj1/1L
bfx4ySyoYlQ2PltYNmmRDPZVZlLaPOqHJ/IANoAdqFpo4OBhEp7Ab6OJGhCAPN9g45ykSPXz06aG
7fzkVMireLaTjBz60tC37js8iXJ0Z2fbuODmnZLd8H4BhabpCQEJ1lRkcTnG2B68CE0ttSD3Ndf9
LKh2uB3SueE8u6/zAbQ1j3lywCB1VIBWBytf0ZqjmBt/TXARQGPcX1yzDvbsvV9PlzAj55IvXLtI
VsLQ8W3qAr7/V0gTvezjCOAryc2lAH33Xz0vOmdCUEVhKNhIo9NT0apaOOC87qirJE8fNNZv6Wh7
lxzV/Pf/sLvXtwX+5z8AC+d+Yuckbi86fX94m0wXn6GfXICHKmpuC6XwWszizpeJYYDvRtHNmVWH
1EeCoYlMznN1u3ZG8LzIu0a6ZaSi0K36nej8lMIqjPz7CNUu9nBlnpwTfAwfGn/VOwE0ar/1yhli
HXNaDAo63H/0+/2CSxsCT2j7DNAiHyHH1h35VqajLZ2tzYLHDzlWc6RUi4qC/LUO0BBFz8gMo6nT
myfVG3sAibnfqp6+XUvgiZ2dPcBpWTfKMAGQisb7lFC+qSNoZFPdMTHSp3/h9UXirA/KiIu8lytB
1m7Bqxx7Kj5wuk1vkuSpFaA98m0NMpsL866mYd3FEBY72pp66IEECqc8+A6FkZ2ENeSIbr9No1Dc
v6AdwTdR1bjbjWtOe1bIYTgfZsTjySTuT9Y+UdEOyyicAaiS0REAfgJmgq9vdB4C/f6/aQhlSA+q
1J9bNhntUwLcTkTsu+VwuqQrX8LBzIzV4M4Bt8g4aqNP9DjsiAIX9Nh88uWI1jBkdiiz29jLORJ0
Vq3lgFL7/MEgB4UMViw7QiiRHh+nq23Vzt2L9q+r8TMP16WhWj06AdtRVClAhJOWx2z0b+P2TPsN
6ebWXAOrtIuC9EwjcSjxiTKyLbh10ESygLW8fkOK3A2VBnP1HWppxezw6OEfZdDCimRs+a5HS6KM
3doeJjv8mTHsrauL14DJca7oAs54zjoEvQ0I+M78ptbvyc6bZLYpiQ1deWk5Br0GKJ0C/chyBRwY
/iyfvVhtFw4WnkxSC6VQXWfV8QY6/apotuSBbDWDH0N2KF/KthP3JIMGktcEyKDNJIUf43TozlT0
hncXoLgvo6iO49/EjC+oRaMol/oWTFdXi/I3An85vHCzeU0Rh3onyfwAVSUlO9Qu4tntEKw6Jv9H
SAsxSNdoY9vz7GnHmTIPEVyeR6edOw/cD044Zq+X5whrDXp1BjLyGG3nh46G6tdLLDzIn0Kp03fq
MD2dQqUHc9eJgN/MN0BqvzBrlqDGfEAFfdOSzlaP55XDcNvCsl+eXPJZRtgLPcvmI9B2YxH6Bo3W
zFimadJ779yRpECab2/WD/+Js9U3ngSvYd/lHjGXDSLvalf2wPt/gY9R7mBwS/pbeb/ZnESkPCgy
Arn4s05mIKbeYVCn6RBqjtxu7jFuM/q8LotoOblrCBsl/b+sEhEh3be8X9UTf/6tdb4bGuhnK6W8
Ejt8QcLM6oUs4mei3lrhLzz5ViAhVfE31H8yR1W2tltRpY+Hvee59E84DPZMBxU53p43ovgrt7mL
g9SRIFD680xAhOO7YTgGD0wbbwAMkmkHFhDLj3uiHQCM5GvdwdDHXWREci3xzHNOUR6qGe7+gXGs
FIv/wwCId+xLyZwRsvbxNV4lu7DZ9A/NF4+ArSYLZPoFyouvzdmdSAMEvq0XUD/HbDaInLS5Lcw4
bfQX7TDWemq4D80EQqZs7uK5VL7wwcOc/rs4SjJFNSMIxhAFuUG3IThdo/hqRCDug3HQqoqFr7Gy
IyGCHawyzbefADMtdGzh/dvT2khhdkKFhGdYPe6m7C0J0JCcQS7vcvDpkYDwBbMtkztQEBYBk18b
jCv80z5BWmUbYnVOghmJ597X82HT8GS+NqNqVnYQSm78PQefj4TuUb43qIEX8MJ3ODARofoDMSPq
as3OkK9+ad0FqxKNBvy+3BJ4Fh3CLZy84g87x/+GvBjtKR8eoLKzJGclcjg/mzxGqmFIpyvZyHNZ
8ECklwC1A4Dy4osyrJAiMjNpx6TRL2jBP2gS5OfXufl//wJDuP757f8Hp8kBCY73c5j/Yw61BLgl
oQJIzdCe72Ur/6Ys0Ik+th3OGsJcCF71qAy3TV19o6yea0CQ2Z4YDOZ+nNonpSFo3mDqAQzgyRq8
T4XFnj9sD7DMdllit0DFk8VHpypaG5ptVfkRiDH9JjnOU2ahaw0wgTMYbcRFPsObGK0edDL4r4sz
y4NFQxYybhI0PATXc7qmN8LaouT84VKR7bZcT4HrIzg5PgXl3Hs8ZWX7LY14zF+gX/YyU7kSwU0p
fLg7ZVMpoceTO7h94CCIlo/5BpDCEWa6gCUBV0Vbunxr9ijZjRvssT2QTFFpwuCpq/u9nIY/fSSq
aaC/KE0oIEYvJbhI85mcC0Zbg+fYC1nSH62fhy85/sWmGPsAEDo/NpH9il2InthOvmwzbLdR0xvJ
cKoaeHIRlG0O49tWzHHexLE9s5sPeU3+tnvjTP/+VOBlx4u7jy8fu3CzPsXmXVxkJedc16NhXPwN
7Zk+pbCJ6yzd+volP4UWdH31tD8+PJAm50Ke6E14axizRXEM8IfTsvIzUKXZ4y/1RR+lWV1yenr7
LW2Jhcql6ebWPPV2c4s3Ix7UrzTMAVYnbbRfJMOv2pfuNcvYPUa/w439AYEl3EbLXrsMrPF6PGKN
WAC0f2MsP0Q1WpT778wGqpCGmT9V847XfCj5Hn3UKLMSK051HMMrTdiJwOpsrLYzZr54a95DR5yw
/YZFZH1aZZ7D4LCGWipmGE9SJGVJSiaew4qAcp/zyBLAGPYhLBn3yb1Awm5utH+g5B3YQs+Z4RT6
Br2YdhoqsiLi+caDpCHPrAK2AOrBlMqmbjQ4P77HR/TrPVc7QlZkGQaHn8aklEIIsQtBEqFEVdSo
5Z40EECcEGmdFy0TFT8wR096qzIIOQ0jZswkJbTmQk/jB9FGE3/dNap2yeLN3nnekRZzLukQzAXx
NvWGWXlHTRNzKCuYVNS2GCXZRQRMpImf1DhbTXyyUWubIinABedZ6UYsNsg7IvvELUdgX5xntfTc
0J/emzYF2kxWW3lxxCX7AbhaoXltqPBTFGCaqCDchH7rjgMM5HJCrVR6PrgtYvuolJGLRIj6Ob4y
aAiU+GcvIuaCumPrEnKjbdJK21Umti2WtKxlmKMqdGKBulpRaYzFW4GHXs8AFdpB5JjzHC82KAks
fYuixm05yk5GOR+Sj+3gdptbU7CXV/jr8PJGI/vXIdqZznQFw1Dj6lDdcf4ugS2/WqOlybSfwyET
pRyGVjq+42m74pFApVYTxiHa2HMLB0VvJ1Q/+XKnYQtkEgFrN8114MP2LI2xKdUjj16eZNElMvWp
rEaueqbzswidj7Ma79wPzxbR/hTVO7xN6fHF8BMWE2jjIajr05kjs5J8VqyGmwAUJQDIHjbLaBsW
ucZJW9slVUALGTdUdzJJlUHIWLWjFH62OySYbEdOGePsYCZWcECJcMX+c6rF8mp+cbo1rgECM4C8
fVhmfjRFD7ZZsuanU1UVQKBm1t9rxoihNMN9djpR8q87bV8hkyFe5n4eGQxzrQLCPybO5BzIR9HF
aYK2ZbqVZMHDvFdetV6ofPVelLKXUafbrNKH2MfQP9PwnHl/V2kdY9ye5GyeFYxaER0zhBcjtWDn
i1u1vC2AokRIu6+WTjZAzJHXwe/m9a6ZoASWTj1kyU2H7X5eqWU5yUT+rj7JZWXMGQCvMs2WVYRY
Jaobenl+6yALgtRTJ/I5JTDFIPD1TcZXavmHRm9+2mc6znHtPbaLvXHOE1I4w2zQegg3irUWsokT
UALlxaPqRQ0JA2mMdO/YrCL5LhHZK7Xp/Gdy+JtKJ2cM+010+q2KhhmhQt4TjXcbXLuymGQ/wCWZ
0huzIZNZZarPSfm98pJbxZD61iv2GRc4+PYVF4qaXOkNvN+UpZ9tDbvGJjuSo9p0a43EDJmnbHDT
sczQqyM+wxlECajZB9d8unQh2zxWQrjsA692VDvnG+CB4D87a5BfvBxr3jLjP8rC6JjnfvpNfyDR
Jf6CqcZy3e8cb102eIQU9kL1Jt+t7TnuPye1Hq+qNzLe2NAbFQDDs6tCku2BCbmBd/Vu17h7ht0P
Gr4DiLl6Tl95DkFIWadYyX5l9rLivNok6rSLrXEtX3XBcArpQwlS6o8JWYUy+EmggMH4ez233h5R
ill6pTn1i/x/7b0OnEHmKEKQX8l2h8NrpXn2v1G0dtmKoiAZizMFi4fTkme3uNjWZHhZafCJeXQr
9OtQY9hcRl/Rlu3fUDosQAw+rYQ7+hYCKKz8VRZF9JHIJr2o7ZK7FECkcFAu4nZ+P1yJBs9fSgUU
Vm3Wz/8il6YvFzJTHeifW7NHSk8AedZMTfSKLDofyiFbqOvm2a+vLhIjV1XgnNSjyxmm4ZT7pzFF
5J2FzAjNIertcuLZjvYUODNaUITxBqbEq2TFZWEMZFFzQ8tFMDnTIVNB/C8T4BEGhc6M0vbRuz4h
9OmU/eqK831gNTS84h5oIqcMqy556Jp9HR96iXyjeeYJICE7yD+DBWajKqJZn7D02ZqUr8E7a3XF
DTU3JnQowSdjvlx9+65MVu53GjSjQTwdXSoUK9pElK0bPaqYYJsOIOZpuvjnjwbk3f1pnJFFt9uz
2AdA+WddrRMY+XigNgQ/+IEqHNiAOCtu1+qdhfneJKv8gMOF/2EsdsoALdjNzWZlTtlDEbYhuSpx
QuTA40avXN05Y8U2gb1bf/YxAmkz2wLICo0X2pBe9OI42VNBxIQfvy/FTS6oC7Ai36BTPxDi+3kT
ddz5UvEdJ6WAmwBOOZ+/d6m6lBUkb0bncKkm9Dk84NrrstBjNWsaX/XZJYNdzO5vLpuMUPxba06s
GNK+ibbj50I+QyMsiP1xk9DVTdEantVNSLUrhJZpQi8p3ArHfSNDqdQqoYceHeWtdlFzoeWDubxF
2Pvv7LBxj+XBAYKi7PW/2lFx+yhpeeM3vEpCIQpwoN1hk2VyI3vUw17TToXcsfLuoU5EuQqXRGKR
FZQHWYBNtx12Brizt7gtW99KEL2olvK8nO0Fa99N1PyI7XWcJONN0p9JKKAx8MMUnHda9iu8JlmC
yw0ue3WclpteEfnJ31d0R25jyR94TgCaFEpyv0zTVvadusmmWHpxcHBWA7fyagtZCIFSEvLnGriv
/70KuZkIzzbssf6/E0vymjmwgYMiNoAYjQsAx8VkDEHzyWo9skr67cqWi/35lGoVgSGP7IKabDI9
favuWnfvYtZWktcPEk64xDRVTW/VxO8lphUsyRy8ESAwEgv0KdeZ10Z6fDdl93V7vPvmHemlqfxw
jbX+ITzhmjKbu7jZTLnfrYlaYCdOaBAWycQ23b9zqtzX8jWAMQt2XA4AV3bCJdphaSZP4zikxHtu
kjEUURsr5/gR5O/yCRdsVbHN9XuPTiKEQUKvdSNpL3tDGVx5XR1LyJY/7dB/tO1klIAm7cUo5uQ1
bmJcTnSrAWKtP9M8AnWPtquzGxMlqchAH9h9TTqqUdFgc+UhYyNHsccCGFUV8ut5vv1v4KQMxv6h
VJZHjeAWxmh03ofJjyttPr0fiyMR7zhXcJAXMYBfXc5xAs0SAhUSRG/qZXj4tsFIveNx7Bu34whU
aPETjaP3sXWx0MTd3eQuDHqT7PsCtePsHNWXmOR76m95Ref9d/2j7kpRwjuRIhmA2XcXT4aQ6ri1
cvn4nBJpYj33BtkKwBQ1YrXESflAwbNmfQpLVIglWM4H81bHZSWRWaw9Lh7a/GvVgvTmzZ73HFk0
gpVEFv1sA+UCTCItVpgq8AaBJrtsiMlJhF/WY0jAt81JYfgrGfShl77XisoPFx7/mQ0bYaztj7iX
/PwOjnXOiNLsVX4h2Gi34S42U6zUeb/rSOEtn+m57+l8zt2QFLNYvcVb8FbEHAZO/cJfx3GWCfGu
OptY9mkTlQ6h12adSbJKfL6gMxQbdEv+5gTapKKzJMRPGwrX9PPFFoorFZa5lrfOYLFATfugIT/s
86N4vWOT91oU8qH0mIXPJ0Ysa8gbWHzPoSRO5LBmdM2e9hnOXbnKKQ1th5HtO6Gl4AJeDvu1yR7v
sK96zj50X+c7osQl/PXW6UMEUAzj2qreRv+J991mkL7WHlyaUJR2WZ4kIfGORlaePhOBFAI/4ddu
TAhaS9A7X8uF9jGATQ+Pp4bDsWrRqsUG5oQmzNpcnK9a0u30XZ7yYvElahlh1Rp1REXa4xU0ksDD
HpHsKFKIjZPvgjx9Omx17D3mDJ/QL6Mk4jL1ZsUJ2abs1qKHMVN2qImVHUlnClb9SE8WteVREVpj
JSIUPiOv37G5pIblFqVKHDvS8bXJV1ZSEqULpUj6TXqcyQvpSBS88PwNuSl43ea+lvQkRYP3J6s1
2dh5c4tFhzrZa4OVGxtjH57WxHzSrmgOaPXqhBC3eoghQhtb/xlG8t7pBaZHAK8rRHPJwzCm72mR
eQQv7J8BkyP8DSdkWTlGK9UR91KhKQw4YEH+gKcIUTqrC9sUuVSzuvB+7VmiEID19MmBcE5wOrc+
J29V4BU1+ybygUtp5UsqEZ2Evyo2dLBDTObnQ6J+CdJMouR7YGNNIGITbloLLKjI9gFauklNZXKC
taLJlPURRT/LkBYwynDvF1mijTfyxQMSHT+KCcEcLKk1UpaPCdljXR/JvQGZJdsiOKFHVGR4YGGM
1vN390qiB8ab+Hj73OGp3u/WET5AUCe6NN+2vcO/Ov5HlJn1RkJMKnVn3eSx2AgVSJcuBK6kawLg
PB0ep6jwtoz4Y1YMLsyInG4PJn8JXTAC6dwKcdy15Xv2Ub6tl3Iwyyh1xmgZ3APV6Vj9gf7AtM4H
t6EzRG/xs/1S/gNnY9slPbBctE1fcFfvY59DYp/SFpa5XhqC/4gwgx9uCPAbUlfYqSKXd0J871Xv
2kt9/VvPHU4C4w3kz6O7L823Eq9pNCoq0llsXhTGWIR6MjiJswyRRqckciHJYmhQY67xAMIPang9
QMVc3nfxeMnMKfJ51movxOCkAUOmhVYX4PdY2FgVhoPNx+RHHmf0NXwVS6diQpjKEk9ti+LQz5XI
UVqBis6x/bCRnCl8lv9BZp8JyegTcJvjjCFCdUvGQeZO55FxaPjIXif8megXiUJusB5uvkYze1/v
YJWmayBQBAmyso6FTwUhGNNT0Gcz41HF76glonml94ed7+WeRnCufpwUzrPdplQ5nsnHtz3wfONI
0ouh2vSWMVOqYPaihBB+UhSnbRuObiO2Mf17C+Rzt98ucHpJP3td3r0yd95Or0H/H4todlab9Won
BsaEqb1b9/UcZoDksN7l5oSchbVFoY4445defV3CuolAOma8e7ISB4uDs5flxKQWyH/dHEOklFAh
q05ylHIlAvXS1d3vP3/nIny2YssP31vM1XvHySe60yKwnjO50oVvqkKKqFBMiSOQj9U1nyTPzbnB
Szgb+SIrK6algIjlx9VbwJAHum98ZpPcMPPom1Y0TzdgtCYCEJytF1a+AISWYd+pz03eqpBGx1Ag
IafYG1HjTViVPpXLSPfk/iLUfzock8+R0AfysV7ZsOup7NldtqPchTxn6TMtpoKwwTuOR7V9fP/L
POb5hD1x2UVFiCURE0bEW+jNdIdgdLSSpqr/FXs6f85Gh6Wx1pDPRxmWFOpfeed7R3bPKoHsPcAj
bC2ggfjvRF3Y0Adh9JT005GdXPmuODc+uS0riekk/2j+TkZePeY83giZn3nPR5TThOFelzdhMKHY
6srvtgIwe1NK/6qo4zM4uAg/yQTia+I8OHcanCcJbNcO33Mor24M2/O0pGQwSnwhuWXyyMr2bRtv
tniJ71mMVt9CUN23vTCU1HHbv3j81UfO9OYJ5iVhKxj4VaLAyJGSTbx6qy4+oV/lpvmOR0tQCVZ8
wh1kaOJRzl6qREh773p7j7CoFKYhuEhLD5jQCsfemKfoFmzjPACbroPmIPsZ5VxXwTOGrU3ofTIP
q9nZur45MQXaTL+1nuT7MoTlEgQoryZg5irBhvfT/nLRIFEDsWDp2XBHLvViYiCpjPeyQyUqGORx
SgSNIpUAa0113Bmh+vSdViBVt46GKeaHeqGMMTiTptDXzUanLoZX30OAvKx/W1Ns9iNmCuOTdFn/
WgMQSgVsw9RiGEzNpd6d1kwcujRDBA4NXiTFW26gPidHMIJMlPh57HRbmBLEwfKZ7aNVpD/6E4Oe
pz9NB345IFBmS3rmAflGi9UZB0317v1y7r80y/naSoA2HsS1dieVG+hCefksOh4xYptS9IFUS0Ug
Plwoib12fWaiUBkI6ma1UYDndsiL4TI8MGcEaN5qNu2q11gqtr6YMDEqoPmMVlJ5puR0zW+lFzce
Fn6+NMtljE2gDBLmxr3CnQwwZoJmyn5vhmbCcgeWPvgrJkeH6sIgRIG6kDag1Ob6kmeLJEaR2h4h
gVSmtno00a2cIOL95h5Ee/X9LORSR0Y6dRtYMBMvc5SL0j61gtpXuwgvPoAhzyKLYG2SBQf0yMI/
1Ovl+WyKlcCyqsoWyfp0xPrWZHsv2NUTl8fQC20cT5OhlYeFtxGamgKvyoTYdqi13mFtVSrmg/R4
yCuwzphdWwqs5vtShHYVKRJ8010+/6a6a/hs+FUzGbMet4nf8ktN8WJfDFEEn5WPacb+F61eEzXY
UGxXvM7ASMTvJZfQ+0st2XrhZwX+QpvSmLK+I7D/ZnOFajfvzDwQdw5pq15O07aw09Y3pJ//NYaV
2gSQitXfHcE1c5lyYQYTAGbgf3bTglDPWhh41fqCojwbtitFzp+gVbtodRn7JvBPDok1yn1uLpJ/
9SAFhhdiO4jWrlxR0zJxPZgADP0GudqykUkc5LeViUFfmiROeaJvOcFlB+fjd0CUtieoFVzNlA5i
iEzx6B93xridbFgUllwN+woa21akmxwFNSm+tQqfZd2BNlAgySLkI0ajHNbEvy2ClxdV+d/juteV
HU5gK9U7fIeDvFB3qKfYzmL8wdKNNH0lY+VNou3HZWT7XwKxe15+yCvlhPpIuNP1I9GKGmBozhJS
/7+KDwfGhmzm3GPz6J5mMPvzA++NbSzcJIRu7UIr554zdX18JOcQuWseQyYrVNQVeW4DhDPykPMs
6MvBFBF63cUtN22pn/67ilmZDGGDXrzE9frSNOz1YjtCyGIrlvQ89tUiYp+ddNpGmB7A+Je+sdny
OIeWPCir5bm3vhzaGWxpUD7GZeSQzDJLu66OOeKQ8e7Uolcb+YR7xuUEhJSPLXRRZ4LnrAELz6IK
kPu9vqGC/nmQJUSF3i3TqD+IOF82jXu43tSRIY9Nvd+grZz85xCMBFWJpeyb8D01Pex/8gJFXZO+
fOMEFhNZQNB5hpTdkS+CY3lW7zSZI5+7fMhFs6LGCn7NDoFzmScMwAzbw8Z6j62ScAjjJM0sU+dM
FJdr4x51gCREFhumwiIAuFgkGT848dTzuzd4iFdLrHvFDezezfzr5wjvJFDX1K8PCaC42aATNn+o
EA8jCIPM4kUVKDF91D0tz2haBdlNahbCqEdcfbq3PiHJhANXHPJZiM9RlsrAAomMe4gUDWtRO5Hk
Gis8QeSEy+SnzK0hgfn5GDXg3k1twDPpBXvSPJy5ZH9KwDW3mc+QdyOrE8krCl1w5YDPjGfeFhos
G1ef5TXKr2T9cWtKk9s3TWVCQCrcLRBu+KwUrux6ALejQkmTAVbGuLvFw+9gFjCIjMTuv3+p7moT
JyopQDurGbXhffD39HawcTwcFhRhdGj1XoxgzhliIANYZYqSyK6IWGiymb+c1+7RyDD4G7gwtcAz
39UcE64ybGMysJjonIe+NiCJPNgYcaHjSwr56SE3xg/Ta+dlOZJ8b9nSITAyqr2RK1HBer09H+eQ
JyqAJ0FH5JB0kJBq//s9rHCqh8HapYgnitWx1cNRVk0uxx7U8j9C42XTuSbFaE23RoyEpc/6HjTf
5FrgDcXbjs5M4shzzbXip82IQoWNgmLpowDjaY9OiwkwT0eYA3L73sbnc7ZIrQlgpxQvyWNj0W/N
A80h7+6MLUgK2N/uH2rS5TG7B1R5CO7kgQu3iiBI4a5mS8QQqVvBp1sn3DEgB10jH+SIHH7NqyeP
X3wYdu0dcpADpAfNWpRj58yTzN9n6bcascM11qxcZUH8vwqu6qa+MixIEeYhPiZ0/Ee59rvonx89
C3mX3tI9lTioicxZDygvRcubK/Lh9D8zLjMyCLPv39W3dsVf2JZSj+UJHtwTy7oVcU0hKeL3vI6R
2SGKTqyb+9c7SZeU9FuUgYw7tG3QDk+h6vWsz7d84TP31MBRkWXv45UpgRHvqy3OxqMqlFONZOgs
j8DC4ey8pwSC03NGWwe43khEv6m6Qi1g7C+KKxqG9kdaon1G3xOzDLfc1d43g/qkCKimLK/wO1c2
p8tDlszbGXoG/Ga/haodE4vPF4QMIeZX62YtSxVM4vOsBpjdStKzQNYOg3f2N8FwPFPPLks5aKwu
M5CEGiK5QuEtb9E3LKLCyqQvHZKTXMEVO++m8rAL/un8525uNj4eLtPez0b2PiVO6OmLrfiE3S6x
vm11Z5VCnIR6n8b7+U7j8AlLprsKFbtVq879vwSCBDv91z4hMDp69jDKz8BpvG2NJlpu0/wCpn3R
6QAjuYpfWtL/boAspDhNmzDAQMoH2ssSA+9HcTcrbG/nZxeTKtHh26w4+Se3GKeIDa9hUT4gopwb
dvlkeYStBFkh1BbYahmjjfNBiWkNCy2i/sDsrgoZskeVJI2wyEZS2ZKE9hTo2r+OV4TXgHHgO44s
MiuzcYGa7fAcMBSAzGQZGjzGmmlHS3uSgOUcv0Lli2PZh4i0WH60G2s8WtjzfQO9vFIUk9Za6RkP
G6oHC4cGnGiS1puOQDkcFcPPOFds5ZKDrOgxTVvHChIXuJzS61MquFuhNFRVobVglOtU85qFbsVA
SPGL9/Tbe/SCsqjlAVT7Z6ht+zv0gs+vhC6nTUUJFK2keEFqjfhoFRT9zwEJJaLnjSqIfgei0bKp
10grGjnLscSChtr8TdI3FVLMKeAZ84++Rz0xXlHbYKN3dm9KxpR6Pu4KYN8IrR7W7H43yEvOTPmc
VSVI/vQUpBrmtNHRqBsamcm2JHzfrmhYxqQbSy3US3jMpBZxZpZMoI3muOhF2ucN7aFbPwVJQpdh
hX328/g/H5IODPfhyVT1TwZnar3l6A6mp/3L1ECFtmu1NU5wrQW5K80UcX4cLbRMvTd8hKvIkPxi
fEyIINj82VNZmv0oCdw2/08rcoEixoxu88EX6jGka1lD1DHfsYtaZ/k4GPwbv2P5vQyVew8zrPIS
YIXM8nJhm21gdd2/Pf3orbjuoSkmCBdzSWAk87qhB23QXTI0XwpJiYcgLoUaA2jU/srq5f5LUZAk
Ncyeaq7xuuNOB9+Fh4SwFbswtZAP6GzfAmGUmKVjEVkV3zwU8mUL6WLoFAUnlhZFsrLHbu9p85Sb
zmAXcVVeQoeQspH3leH5MhjUxD/KGjwVMhhjrLygVFLvEz8d8JpoQ6g/5lXxTULpdC1RRastThxx
pFsmyg+TtZLIIE/RyMEA3fYB/hohNJbSN1168op0zUex+a+xh77ig3VN6DWehvlE6NPUR9sDyz07
KA3yZqO8lx6G2UdozoL0Kug6CYS9XpteNVq9tZXTtgfGb7HPlp9byFTp96kiNmT4YVnnst5nq6Rn
EtKFz/st0vf2nnatoe+4KgF+Ko05nkfHI1nZQvoOiHepYRu21/nOP857r/jICP3TX/63Kh6TfZLr
n8cm1yJU/c0vLCY6oHcWmmuYetd4M7BzUQqIzmzBKdJb9FR0Os+NVaTY+br3B7wvqQE0HQCUFkg1
9f9afh/nVTgXFJnlSmlwni8my1UkNEk8vHqcpXdPwvwkL+mXcR2FCazeYVCITKq2A/pjioJ3d9ZL
PD3dAiPN5nguZ8t1+O7ovBHwXrTNWFNrpWY5kZSfXhC8IUA1ZjLkVHJlFwwId48nOsdhnnpbHUoT
k8Bktgvf1gb8ph5r+qiPSn8iDXDK+KmMO4b0n2HF+3Ui+X27LU2kDYcaU8dOVJmqedpb4w91nYy/
dCHg4dezuW+iYWPSMQMYU3YbHuW8u2pEc2gTuwRahEr4qxlV61WdHst3ugZm9kM7TU2AXiTC9vRb
NJKeRSOkELHA6txvW29KLvbd3EdqkQ7Ng0uanpHSnooKYj6GG+6g5Bkon7rCKttXasMd3HVCkQ+Q
v0bnOxFuxMSxw9uj8EmTnTum/gWfQr8c/UF9ZMgd1J/emych1/5zmTM1An1b+qxcLuHYpnsoupTp
MC6VN2/QYQ+qBxpmyfeXw1X+WRn48ngObSMsQz7QmB08bG6zmRqQ2611wA7Y0Xk29H5o19TyXLAQ
Ildxb0cw1GYU+HtgyOeBrtFJ+MUwBeya7BIdDAB3CD47tKb5BPSHEi4pNa2u8EQePw4/gF2cJ7zb
wtRXaR982KUcN4AupjTdkUEcfSYwPv51JJK6I8zSNHBtat1EZmT25Dl5ThTJyPmTnRRsejehmlBr
z1HUqU7C5mRh/a7jHQ0YMJA+Pv8w28l4XGcqeja8TJnSPQ+EkCCX/TYPhuG9MxwVKOMyALxEyjg2
HUY6eZ/a5g8qaD2dqmRZ771H5XkQq3Xk50TiNTNCwm44x2l2zuwcddXnBSuw6AUMy1aQIwZR2LMd
P/y/ACw7FwgTeMGwrUm8l93gkYrnTj25Bi8+9wsO4By8ZY+ihJ+znzVlMwrKsXU762vHcFIREx6Y
4HHuWbbLkgGOycpKuFCqjZ2ByvH9f/uvHghrt8JpvS0JTB7z6fvCQ64o+S6xH7vTnID0ANXYx0yy
yMDbBY2UTNrlXEwDfCI7TlUWUuY6IT92GY162ardgLZK1Uyt5Xs0nlnLnOyZnudC8TYPMpcKCPRt
oevwFNH9AiRQ4j+5W6RUlbR3V103oid11P8s+3z9fOkQ537M5INldBSSRunZkEFWKFOinZav+App
sS8cSLZrKd2kP7bewxEAZ4rG8tgZiQmNdFi28liaMDOqoAGXlV2oG1acIj1SwpzSlzRicQ1IgLHL
gmpODkMjo6q9AVgi86mMLuhgHf8/eq81+pV4CoqejQNHbXW2cF8tXM/25OIvjjSR0q+azw1LVPfq
iVs0fIYlttCKx9uc7h2QU/sA2VitbFNdF2ooLiiaiGHTIJYBllVeCa9Uvk9meNF8Y3ac4Dp3acUh
mBazbHfehdfqxdWC8wkBTMZjykXhn8Z8mj2inbvCJ9UASHCgbN4oulXAHu1dAuMHJZI/3b2Hv/F3
7XkE0/MLtF+ucXhmknodABBNZ9Xc1X+6X2TILAuurMnzIEoGbkU4w9p9b2tBwNaA1BLRa31sDe5Q
x0+JV08gWcpTG9MO6fDMJzfM8Gf00g+X4cH/AO+kr8srvwDsMXns/S6AChjKo4NECLfh6tExSRAt
senqBMy32tzstDKQRTBy5xjGmJ8OF7wiiUqpmZ6S+KJiAqDB8BtlNoWfHa7rBB3JBbHtDXGP4VIT
0Rf3juwZ/h7NrcfH9rdNNRKHezdtjMik/SyQ44nBdfIWn+bQHK1aoZo0nZFrjPAg4XMGWdwzhmJp
fVJ/+ck7sVeUtnzK4kXgi5n+dw+c4k9uEV2WneqxhTEbtsMAfaKZ3zobDrgiXgdfUy11nkzHDWUP
WywmDjQ5StInD6Rz+ULfPo5CCzDzqtaqbmSlPJL/VAKtUVEIzChsGkPX6q+44W25tGi4xzdwZNER
rCOLLatb651GO12uuGHrOpUU8RA8zcurPiCbtr7o3cOvMB14Wfsp/GjZQlvdB598TPV3TEtCaREZ
YDOZ2cVxrvQZ210ure4L4q6kbR78sEoKKy67ba6K8sfIHVfx4N9FGEa2HPUyccfJEcRCj9JQjwx2
k2ZXMcYoZOOeVmXuafWcOmkxq4Tg3Th2p2oxrj9RC/0MMueAdREBbc1nT75cfn3feSh+X6nVBcLB
lTZhfMhg2/Dr4BzXdX5VMCVwDb6FVR4hsY/SAD+fGY3IueYIC9HGEiJtsVJlRvqsDrKg5kOZnFOS
JNHlaTiS7Gxb6xTo7OD2iXdFB8M2ArQYt50oaim90LoxojWcy6Xd449gnoFAcOpZpXwT+ByTbSV0
IVGA9bHhpnPa/RSyJp4zfTJDhRW8e+weZM0Z2KkTw2iQbNEfIEYcvqyiKWkZkRtUlgyewNE2os9k
WjA/DxibHjtWU4lFOqA+67mig54ZvFjCpBW8RLu5NFRhxnHjNTguDnBI5hCbaFau0lqY0kiw0Mlb
Aw+eYszq+s6Fq2p1rpMETNFRZTw6WmmfloPdv9mVuZ/i/V1I2d+T8pR/RSnbs48Sk0286C1So+cP
6lNN18HIxqEGDrUF0F9JDWd/lWSzq//ZXTtooOW52bMut7VmGq9gkpD4/4SKEY9ekFS6UJYblWfI
hvuwmwjx4DTnUuE1HQw9ppkcR1OdQnXhqUR2aZbuittmxnElseyHlbcurYw2YaNKeWzcfN/8RvD2
1JZXsOV97UXEVHMk94mt/qL+fNg7vHQzpGCZ2dRb8/HuPEr2cB+yOgy9RLQ6Vc9eNrIgf3xuwSfm
8ticISoBVX4mwiU6AUM7Ds/p5D5dTXkeVcSEfNEJdub7Rgncy375RvZyQa6uJ2SnIcDVgDSZ5ZnG
hX2+3UaH1AOpaPUmumzmxMaln3ihzzIe8Znp1MOIFUmReKQwFirjRRm5GFNEVEC5mhfR1tpzoefu
+xuwPP/sh28ZPFu86LY4CTHNtNsqjBd4KQoGotZm/aCtSIrUwnWww6LIpz9XkmCBaMiRv+WdoS1D
LN4GUDLecpltkc0v0n3GykDXYWZUbvEkL9+LpLrzey3VJuLX250ubrMuaQpT1zOmgvtvuTTOcIu3
Mk/Asj36ph7D4f0YEUg/d47yPXdUydIqI94rmB63I2FafbLBHUpR53n+sL1IuEwMLBSJKI4dagtN
B+7YPSXbhp/VvvVFSL8fDrp+NdRq1H7PfRTk0Flyo2tms2uCPSIfx13QHigTxjUtTGoNKJsHq3JV
u+yHLbJ6dBH0LNo5SC1E9XjCQfDopMMn7fphObp+nQChGmtDKD94az8OHnJjyK+EXkQp/TgjxRPC
Z1HLZ3Q0cr7Uny1s+zR9S/sBCchqVGjIvmkVO4wRH9HlgF1p8T5Y+Fgp1Ln2OHsoY7VUkQN0JP4d
nwQs3DQP7fDOvq0w5sagVx2UVfffb7W/hlZNZ1/Sef3R0CNae6lHlVKjBXz0p7lT7vUfvBTHaXMg
5Wu3HrzDuOtdPyq4a19A/VqlbXs8ZN3q//QOec0zT9XkQneqQlWJTz+Xtj+wC8GAVJ06IVQGQa/3
rxYp8llUx2bPC/+dDuCCSiYidnL/nO9Z+HO+EHl8D2/l7uzl0kH2r/fTEwLsso5xdVOE+tyBXrDv
biiKzVdl3FVzAngi4GgAxHKfufvbt1pQfBdmk3ZGzRZ8Ak6QaJZNlm5VvwLHsKqD0caEW8xU6CQJ
kYgALc6nConolNhhid1ZBH5+fy2WUS4HUHIjX9ZqXZTvc3kttlgEBP7qCDLqRrD2ZpT1gdrdPNry
1921yAWL4Bf7/qJtF6rKvbhPJhuGVw8FgswpM2NefbYxhud4uUYgtfj2AmqgzvGDLoTFmQPRXg/+
xmjuQN5owDdiH3S4Ce4f4EeCkU0NQQBYdDPi0eP59I3/6y3g/o0IrJsGS67MsD6DTcTU7DRMTp8+
m4O8y6Kwh/u202+6zV1cOIVM+dQsJxPtnG9aKnbbMdL827HDYim2XH80Ymq/ym4bw2eq+vtxwFdx
AP/qii29P692R+jQeqfd1b6Sum9JlDbfF6eE/zl/vhxHfM0itZ/rjQu9l2Q6q+a+wflT+RNj6AgK
sWb3ALl2l+z5Xo8lRphbjstcDLFKZwHTUNSHsRW5JpONCWnd0szPF//b6qXd3Q+9ELtsRwKmrua4
TNS5I6cOOX7PtR6Lv/jV89aYJINnDecC9Uf7RcM3o7AhVGwiR+jxqm7cAKdoyf4imKD9/lhH5CcW
PZGhsiwbgX310jAUFXsbCNSYamJIY9U2+wgFT0qs/UXVlsREcL5KtVhMR2kR+4QkYV+9icVmIAdq
DxyPrPl9qhEydxL0Ds803GtzxkdetQWNEAk5t6H8/CwSFcF5iiF3AIZVKnmtMjcw2fzoB/Y25GNs
twlbOLUocRmZ6znQEzlAAp+AVC4OzyrR2reXi5ZT6wVuURF/46Mo/+Fe3pZGhgFJ1Cr/b17FV+w4
/EPOYKtm7mFHWjCRikQLVhjsdhpIkM0uctkBBwE+8MixclT94UAjprDVgwVY0GgdncDKXXYDyn+A
UnPSauXZAFdgdr5y1pIWOpthL8VpAadMeOsVKH8EEgyO51L3BW3TYWtGX+Xun17l9g9wgQN88tzC
3+Z8tgV0aQFnLNbYjwi8TwwkfZf9tZLh4hCTHIOtNKBRlqIVfneAR5VUl3GjkFkTCbjcVRzag5x/
Tp0wxGBuKASDJ/0yuKRhy+NA2YrLth359dzFQzms7M5FxJNyxWZEs/TP1xgVdF3XDNKB/ONorr9u
NmMWraaQPAL1Q4SH+D33FgmmQjKs5FzRGBk7XSxxUmMFZOAAzCdvp6aLNSCBkMGNMYCHxEOFfBSO
cJec3FkYb6XejdJ6aWzX50qWVnGK6USZElU9NBT3NF73HkJwXfG79Hj46fqsoA3OY+f3esqWmtFO
CT/+yExYa2d1/OAvADdTjlgmslkIQC3q8DI/qfZiJxp+v/bDE1YvZLrTpoyl41/GSwU9dz9hDITJ
fNlVXsdltokc/Q4U3U8EuaZSzDd9vXAYkZXOBROmQEu5ExrK6eOkGEejKCRPcLy4t7ENmSoRI612
93wGO0AsZPqXYaXJOBQ9ImPQqiDnj4+3ltcft85pD5bhmdHFPmx/QtBTkupz24sboe6VdITWHs/q
8AqDoGeMnJeVe6PwKzrBPVaLvBoj+46BKUO+3pIavY2PdrCDBy/og5cuov7YmQPLqYSFdWKQN/TA
6ALYUAIKVxR4diWunePTlIWjqnmbWq0hBD50wykNWkaXjolXrwDKmFmfhWu4JQoz/FWT7qht5zRc
YjswuBjWTpuABQqnU7XysM/ErWHNVT/CB/TteU/OlGF174S+xHrtsJGOI1kqxUbhxv9Le/PXSSOS
+WCP/n+atmy4tZmDQugBYPJ66B9R7POldgSshPS1h8KJPhLMCHFqXTzBB5IR2yG66eyuiU6viF3V
tSO2xhw9q7xyE+COYdQMbpFcJs8Zbi8usoPfuLX1toVYBHsiRo+ROtaWnLmK5KPW5Q6IFcabF6dK
5nB990fq40mmUZBoTf3byHnnqAeffBAyMD6Q1ila5KMQKBMMkysHNGvkeb0rTHY9o+j350a2pMEr
b+3nJeZImQBVIWM80IAkh7DFllLzzJtGExtbTRHTpYe/Teu9Uvxz/8Ks8wzcdPDahB/dUo3xa5WP
Ho9XFSD7JyBw8oI9p0rXNMqMYGIJI7VHeRkc/gIYRotUSzZ26yAHBzrWUIRvW0E09DUqSjXzO7jU
g2dH4XSMo4vuQJCge97g/wkP5p+Q4i5nPIKbvi/p1fH11i/Gd+dpuGgj4Wpg+Pau8uXepcZDYwMu
QZSyzgy4jxPyuTDUDMwkWN6ptVIzbybbIu7EgcRz2Nu3FGtzKrV67bstD7P0BTZ2GdEEhUdsgqzi
OltLCZlkSKa0fomizk/URzoODdfHLCHxxa8UiggT5+6kl1pzFDhQZM5plV9zTvsJFo3HWeNZk2rB
w4kP9PTx+VLS5+g2DUtiekKaidOssYKyyJ8RUK9hq0ynqJp5BMGaQSJhZsEVkNY4va5AQ+dXrSDa
SqGJ+JXPKU2iniPEBqFlkUc48DmeN4S8KposB1hqCKS4A1WNLEg4WIcFgbzZjt3/zw+tYqhA41er
0P3Z+p8mCH2p/unvjoEv1gfbhL+ingtSjJG5nFyxT1GRbUetYyeeE83XmadO44euVJLnzgjvvBdz
0+W1ZPIbAPdArFXoTUVoRxZAXmOYThCmssGaYQ4f/TC3R4bycwCCmQeqEk3XP1AYFS/PikrOTs9J
hw9h7Gi3RSoVXBOq3ekiJJPZw/+9PJs9TND90AvM7o+9nPcFtD77E5FuYj4hzgTRBcV4huilAQDT
E915EoI00W8p1It/UZXoBiUKsfZWzhHaP2woTmdJHI1r5svJXrUYhfYEveXinXr84JaCJEoktAnV
FGoUH8dR/8AG0qI/l2nwRzmPb1VBBv9MkeuDT19qyVb56HZ+JH9CPZEP5lJp6xFG9jg4hmAjJb8A
WrbnXJQa6B4l2Xjq+KrTV4sKcVj0FQl7egv6Dcf3VZPyxNspiKko3NnOwIm34NyLY77Jho88oom8
PSCVcHk5BMTUhnWCbQMPhQ7ZhmPzx1vXMQrFVE3KsBK/Nz5LkWWa6Ij1R4TyQNRlbaxI2cqgapc3
xI4/2VR9hMjeAVd2ya85E2EbU+WDP0e7JumZruIkO7+xoDaq0mRGLJ9B09B5SU5iU4tGd9wWhDMZ
3k78zyD+XVenY+2+N3h5W+nsPR+rQ5Haj/1woARj4b9aF3hrmkAulkn0gpQwiSIniwVUerPHPPYC
2usL4nZMJ0Fx88khFHDq8FKhUNbJlHBiB6MsWNyFqA5JQoWMKOXR117HHIgpWvTPv8hATAnVU1oZ
JW3G7arMOjX6Guxf47vQ3C+xCd7cpg7nM7UFbFIDqXdvbwde6w5xzJTORoLu0mx41STbAUS5n4pi
atb/TLUJQMlHwrLVT5g6KMGSmUuPCNutZ3g3/3PqExWRwp/P4xAQgYIyvZmBlw3uZc2VFKmSz2A8
U59gpI43gEkeqyh/MXkPyZ3xtliL0WqzV2JLD08t0vdn3rvwSc1XJhHaXGERAh+v6AmLxd8S/8uj
vO9CpwVvParRhSn2a8zHPmt1zAOilLCfpn1Bo3O2NA26dIm9Rn4WLQ22pNSFEIDJNMEXMzDb1Wwp
KBvRE2YXK/NCatvfaQQKGcdxxqBT77b+dC9TvcBlC9jag9JN/vYA++PLJOOKdMGx1D/lK2iMgdsg
kuv2wcMr4K7qFrCdKEJK6aFr7qsDqqk6YAWPLwfORkp4EKEmXh1y0cvqOxHqLPtCwveYFLoQ6J64
RoHvkXyLXWVDN9Ld4VF1Ks2l1XsUNfPkv71E3H6BCzKv4GakkH+18Pw9/qJ/cpEEt31yeHGURGcz
y6abmHwcSJs8KE+aKmWEbMHziCfxTbozXTPJkn7VK+VRkzO7dUaO5hdYD0YQPQAJAqKysnGo/EgW
NRYqW9ooI45Hvw9vitQ68/HY19n/7COWUqHRPugPiXCoqrcW7Prc6u7JhyXxUtn/sbjBDHDNl+FW
4iGYC8nD+eapJ4DR8dMWpgKmuv6F+HRz/QM862fjf4Xb7ajTJ9SfyEd5TtABO98RJCL6Pir8a+Cc
JDVr5lmCj7dxPgT4UtJXnsOyCOelR4IvAXy7rzkFsiOQsllmCNQp+As/3yliS6zGtRyJAMNKfen6
41tmuRW3AUZyAq3du84C5P1Q/BPc3UiZBhi1J8XiMFz/BRv713nr8GN9P4DkWyxQubxP8xhSXWZK
YcIGHEeoBV2A2bDbdqD97HEsnfoPv6rZYyvc8FYbeNu0VS36MZRp56cu/d0SEoHYcPTQJFl2WFMB
4Zd6UmHUvPhovIrkUAQA4r2bXjBccLE7GZYzVBYewyEst/RbYy/kyPvZSicFnLNHc+163oeHSrjJ
Rn05Tn51NSkhx1vXWbIPm/rYNc81bOFUMCbTyr3ThKF6JKSitPhXQBr0Rm3PV8wHBP+Q+5xmWMqe
vkNVVihAXklvXVInQO9c2przMbJbO/1BEN37scOwlZiRshbsXWpEkWBmjLlfBu6LJD1nYF4eSUWg
FX5xEgLpnto9+Z9fy2UMH1aciZ1PqrssidfL1O51TV2FH4nDYONZeQ+49ct7NnkWa/W0l/VfjJUQ
FzV4d44ZZeuhC7Sq9KTGMbpUY7JUZ+9bidpzbgoED3Y7+U5SxYFvlMvutIFIRibnKbbYFnqPXatF
1tC0Xa4OSjH21/Gi0iY2TR8fPcewTMqenpLgu5Sklk+tp7fdfiGFHfXYZj7WHsOQRQqf3PTNSHX5
h45Io36YlaLtfXC9VRljZFGsd6FDgGGp3bT8ePIWMYhkcm7w6tTBmIYDIyHNe24siqTPfRvZU7M6
adwojtkZXln/t03nJLZCFZ1whPJq27hItRmNlcc17N5enCYed//CfCxeImSSYiUK36uLJ9hTMdCw
OMujrvwAqnFwMP0hDWbso2oJ4Jy7ClMxngKWhrHebbIexUMcIwtUkn5uPM1sQ6GVnr4eEvKV8dS+
b9bw6xVasQWkQFrpUv4+xxClE3jagTSrXRVZwyjyeoa3fEA+zlNXBvCIJIqAAmT8fFhoUucD7+cF
HvcOs8MXgW3/Fh/t++bBFiOmPAbE+s+lrgWCRGGmawn4Yw7YkTilo2x8cvGLe6ZqxiayR94myvrX
tb38lk9mkCW6lLn6okhmDkoVQuBP7ySJnzfFbPxAH07CPHNph6u9AYFTsXYDwJqGg9dQhRiFjdhO
oJ1liFXqyl07C5fbceSIlL4cMLPZQ/ie+z2R9NNR4BdhO3JwxJjwxG1IUK4qxURNZyIxsfq0SGvC
37+Jm3qnoFGREHdWInI5LzPleL0BOXdJHXV8oZ6Jk6NlXPLlwym00E4+04KT1xPPxTE8i27F/dFH
QHJI1DV5TJWkUxK9W9vhP3oPayB+7Hv+DfjRs6qDCgQLtbOItl8rDGfP6fvRSOILkJ6HBevAr7Qq
fouLZXi9DBViLNR9Z63DWW7U6RifeeqPgd4vgpVCGC2H/PaIUcrWhC8QSu5rVyqu2N4fjnhVP4a6
Laml0YPCb2B7+VPPBtUl/ddenRqehunwDgUzAIP1MBw/nRtHlR2cUZUfLF7qd9vU83I15wXD/K3j
o4IzCo2CxoEV/bqgB1iJ1mBiIx4AsbvHDCm9Nn6sVL9PgSaViIRZph3NBlz0oOHmQTk/RtB0RnDY
IOTSlbtrjEDKk09f2Oefeu08E3d95vKdHOOdnz0Gu5bITJMjaWZdgCRT9U6Egtp2Q3XzBy/5jeha
d+QYptHHnvX1M+DaS1fqR0/o6KnmkcPQWBIsnTv0lLd6/0JJXhdg6I0XQnvPFzyAp9q9eN6eBKhR
ealSfT5cq4vE7Tia6iA0teSyiwOBHyVRQAgQJE4t0KPhvVhzDOtFAT6Yy7xpL7Em11Rtfo2mnbjR
RXfweTq3ZWpGIl9MCr6Xqb79VdOMj4XqwIP2dON/QzBUgsc/u8gSF7Js+R3UBJyQwPyvJHIyU/MF
aN0K7GdznVVrEclnVDczigofQflNzz7CXGwiQjwo3tqMcUtSkMykQ4kXaxcCKuLJG9evRyD6XTIg
bKYT9l3xaJPwFE10rm2ochqrLJrHRzHFQYce6YcnxGKzdgy4jWOwaTD/MhHBiWhZyl90jCGCutl/
ZvxIu/NrH1+wYhsVZ114zgfUoTKaLEwFpZPBbPGldRXNuN6PTAJx1aTb/R8FlWSXJyjX1P7zF6Ik
Y41uia8iEMc3n14hcjrjnGK8GEaUmE9tVAkcRxUwvM2c1+lxzHW9l6AvAmlCs4TWIiZSCZLufU56
WR9vN6iS5Ez9v7TKHbMKnM3RtZPIZtygw36IXGSrgHserc0d4S23JfxiUtkd9j+gfUU6VQ3xc01e
0T5x8ybqm4S2VLepuHmD+MlUQiqNfw5hLGHO0SjoW5BQVRSHNQadQZCPdt8R4SoeorNKl2IrXCOE
dq6WyP6zBSjQ+ubDzvqJGJ2y362Qb72RyWThVUY/WtnRztdnh0PIU0jsmx7k+rMVdX+2Avx6QZTF
ZcErKGvG7Nv+kTRqiMCOliz4CtpFOH85vYyUQIRRUlEsr2vwjy89K0vOcf60t8bEHsuKVZozfnFb
sOuxbQr/AIPnZvbJNT7OWxnD9ct/6RFtKSOuBLuuh1E7GvtRTFCgRBQkJNazn3dpa4rshKlgRoE3
lPXx/4tsBVIC0hldkuPlnFwLTDvohiG2ouySMRUQnS0vo2rK/K72yKczzvSIIcrRMbBsCzCzIghX
JL6m1Tc0j+jykkyyiIS/9GQepCazZonIHMrRT/V9HNVhmYebpi3OcA6q4p3GOUJG0+AdlueYhM9T
gvNkmTQdYINm2I7Shw7cZrsTnBBJYmEV2npnzkTgoUHesqAZuPPD1iHUxqnZzAhE/YSby7YUxCOS
53L8iiHHZS/YgybXCpYQX/+Wbt6JOr/zJOznwsHvIUWAyy6vsiGCkqI5l8xmseiMqronpzd5YGko
Gkre8y4sMZB0y27z+VMBPtZs2us4aVgaX2hL39gGb643IYoNVeY/xP4hqw8PEZLoHWhMnjvX8vtd
qPJaVa/o/b4BkzahWATciHAPdqNkdWnicDa/A7rpbjbOWePcsiBHFwi60WmNwnvjteXCAhEVCcz2
VrN/qMUQy4ZCke8Emyv89J2nLFmvEx26yCr/4cENmPykpEIBSG1ub1HEKbRtqKKvihBRqDbYOMPX
MVS37FlaKatDpzZeKrJwXZPuyJ2NM8JsvimWCypY/66uVgWcJk/KKQx79Oc8EbfVeOgskiDNufgg
cH62WrO8aCQoLYktKz7WOK2dcKgOZxqBgTq/PiY2edYUxlTmpAs8Wy6HTnpKSoIjfN2wDuWCIYnu
5EAHPbPuHCAZOZqTySVj4vrpbfZeu/OouY+BUTMU3PEFc2DSlxFIKlxytok2/Ofq22pLXC7FPoki
w9aI0YD7Hel4CULYDYzyRm98VVH/RATVmbkpYXrL8VaRuS1TKQp2u+l1CqUnfHszviQd+MV1VmQd
6rKgISjUIJpwOJrX0gb2Jb4DAHvcauPuMoUTlVREUspLQCr6EkjRe4xqYxIVZlCoBmMUEy0hqpZp
g0lZWOsK5HsxdAtsNADFBYMAi1MRNN7c47rCxv0OTd4xmLP0s1vjQzGnCykoc0wVG6NNaHtYijkP
V3keFdU1A7HVthZp03nHuYJjxl7MT5vSYCw3eYe7RrpSykSXvqax9uIQRsZTKcEIBZzKJBlIp7X1
KRey8BQVklPmUueh/LZWwhp4HsKUBytpmE76DfECDhYGlVg+Mh9fcBfmn28ED/4/80zgflF/+ip2
Tik5qOA0VFJTmGRTb5LRyuXBX8ArG0+6nzICXEt9Vi/tJ/kU8TDN6tPVY0v5+4nOr2FqhsLQAizZ
MVVugurkPrbYml9rszspLsqQ8BcSLRhlidkh2WtadV2DnFgx9YtC7DiwlIzC3OD55ilv5TIJp2oR
OTiLKwAChrNAV4FFVIPK38clpfI/PvgeES7XAHjIpOyQrWIz8xwtFNVG/uMKIAfHT+zgFLz3HLpe
mXwJcEn79eJ9OZHtx+S/dbEWmHTEVTYrrCTSNS/ovTnJMz4xv8qn9DIyWxUloj2VThSPU5nDFDTw
56CabSqrcZmlgjCvrETv8Ax26vtxKTE9DJxCCr58hgvDdGsSNR5Bi0MO6DTklkWkMlgiUWDT04bb
29BcvmEnti/dY8aS0ytKxARQEC3lUeCja4MkRmpx8igO2zzbmAYlDfxOtNc/Vp91N7/NHTtNaLkc
LUvXvmbUw4TbnjFSwhJQYoCuT/WY1zwLsxTwvHVVmXIv3faHeMo1q5qNh8jemOHJwkwiG/ME8ipE
pkYqmitpMZygUmPCyAcdANV0bQWtXgOJkSYeLuh8wT4ENjR4rTQ/8sfk35B9JfSeksOOJYLwFfQI
Hphv4t5Kyib+D2onM/7v8OHY8HhA+f2DnVTAO8XubegrcCmldZVKQ+fRSmh95hiXIRx24S0Eawpr
2y2LXORbiSC2fxB7EqjfZCV0D7V8DYKGxQ6lXKopQA8IWEgdh3EDkRo9xpxtA4tw0OWBWFV5VNlx
oOor3AkmDx/GMHdV2AUPr+ndwGPbbY+4eIlJdeJ0+25iej6Tzj/VvNX5anD6qBcv/rDthwSdaDVz
dOmBCPKxqxDvpj7VNI5G0NdxMpJvcZbLpAJXNo7Mbhdds10IaGShMBrjWMkzj1/gK/P+dhCN8Z4V
yOEa4IvqiFcutF6qe/76U2DqjFvpJTicImjaOwTgVozr/Rptukt12cNadstf5EZmLKUtWm25zi0A
VvO9GJXVc+Spc5kQ4F6MLhPJB6W0KKHzm09vm5TjDhtBuAwFC0UXsr2aK2hxeJgWLRAD0Gv0EF0D
27Xha+h077XyEYDdrvPnjmfD8Smj7rdDUcFfJgPsjyJXVzlxtTaaF5c4cyTIkafyAf8od8SNOfh1
nGWcZ7Ls+d6irz6+BoKMzSXLt0j9RPyjBoKHv9J8PMMHQEToa1KGq8xfmT1Bz1aPu59AghhXJcHr
hbgKUPZVlgXcMzCNx/GR30g7WtFPqqOMVV9vImaYj86n244QbFnp0xGKcq0w4kBFhKRy1fmZBjTW
rDeN8IR59/z2OW32UpRigu/I0j6SpylrAv1LME+atNHVMWv+TlixngOqN7FdCkXWgJWrC14x6FjV
u1C0eg89vhdCWcNomfWpuVEkRxhRNs4rlhHHZhGmbU7i8mfDF808/rtGbJUoUmo3dQnA3LnxfgOh
BN6SupelHpgWpxCdskx19CtDQjWRPOhP7UB8oFn5MOP+XaSflnaFFFqbmuhMAxJSW0yBO5hull/8
9F4Bee6nrbMHqxGNaKo0wU6Pg0Wb6v96FnsfsV9kAIOrAF/ytQBGIOqR7cqLgnD3Os2kHyWZn5CV
k3U0oD56k8hMH+ecHZx4KGr0IPmKQFrk/me9xVdVuC+S1P/4rrdqiqDvc8690PgL3Ol3lN28Q2Io
2ofUwwHIjaXyCdmS+U3A/6Mu1uVp5nW9P5uS8O87Ur2aIYJe5DS8cnq/5pamknf7by0LrUfdxVDJ
7IESfdqb7RD384dQuQvca6umKhdoBuSBkkvdFlA3yGVg+xHgBm0D5IDCHV7js6i5Vka52hcQ/Cfm
6tagQgDIvt1g2IgCH2q7qUMdxC7GqRY4d4z0rmpIqadrNYCW6T9MXi/Q4qRgKSwG2m/+Q26jkTZh
++JoPvg4voVUoH7Wucin0epirObk9+0O6PQKmz4x7zn3U/nP98cf91/zWBc5m6uqkT3GsevXw1kW
Vk+Dq0o2+Mv2De8iCxxo+Mqn3ED2j/ZJP7XUaGYnI29KnTlfokv/nrzBKco0nKwpJMiX17xM2J6p
+u6MgBY/crPOGUtbBIjjNA/3Mg6a4O4ZWekLD31iUP82D1QO/Xei7rXQ7jkRPCWce3S8Qc1SfTwt
MGHwWBUB5t7+0lBqVLHNZCpsjmOsENgumQEvRemeBMBoXEJjJPauxyqgkzCCS8hiUoc0QakYhd8D
q/2Byo86DxtfxBA150vxkLd16cPdWP8mOdaLj7hzyawt4oFMTs72R3L/lpIT19AgM1VnDk4AfHEG
/x8lkm3fZTRk8PhZKQgvU4KcMzJltld/uTA3VLxmpkZTG6UYfAzSycqPiNDQI7H1vVjR7waK7864
5rKsTO1hwXhAaRABksVel82BsAKiBtY0PQqch+pFc2YrRE6472u4F7I4jOKLu7ELWEGAzRf0ZbEX
2m5IVj991MgT51IE6IjWwB+4ONzDkWNEyKLMIN6p7br7vqdJKr19eRwGt+rsbHBlSLnseNZ7WST+
VvuDOy91zXZwRsJC0aQr1EBxQJQrgttc+t8UwlL4zM29IQa0zGv0yl/T72RSSreAN6nQR0T+IYLp
Oo2LNl/4hZ928CDvUZyrnCTWVXg8KNL++pL1qR8UCpPYvJ7OwU8qCvLdfVjcYzfumNnH9tYsmiwL
XYnBG9lgsTtu6RMzgNI+06KsKmcuNYpDr+axRVJmyeg5NKPg25nstS1U9kuimOJ41ZJKNNuLYm2y
emCCawS6E5BwUcvW8R46q0CPkRsxrcjZvk5sv92trK2UptzGgkwzuVzdwXeiFm34Y4BigvQfaKZB
QjEJD6+lc/fA4T+Vt2PtZ0VKPqu5ywfxO1voPNsE9l8fygEwxN/WYuJVDn74+Ke4WnEmthrGrQI/
xnXsBkfdjk/crl8S8IKWKwov0oMDCFr+lmQFYJhyniqf0VVYLQQROJEo06OG41coi6+2piaQIv8z
4EU7+d3nEZV59s1rAkyVjd+7v/iaxBdIhYlz9sJlyp7aGejT1XrZ/Ri1W5Gcnube6qs+G95buaRu
eMHxDDkS5J2+o1dSEkJ7jRpxwrh0heYltZjUwIHLGMHPkDKO3dYqxTQe2oxSt95xb20f4Q4XIz00
szLj8eUjT6K7ymFLOE/Gov27caBg6eYuAgYYq2cNDdYh6dloAgV2KQnhg7loJiD12rlxN7dPpM+z
odoJ3re2xCgjEqzwsSGwrUSuyOTVr9fpnUFwb8F6MdGmZHIUvzuhXJ5Y7vN5ANIPgOjRXDSojgNN
SZUwVGMWbnhEFLSSZMrgpIk6po/9DvP48jRmBRp/WYVoSw9VlaFyOwgyF+7ctFn6O2pCBrDIdGYn
6ZLNJXjKNmh/K9yFTB/sPZheRGzAmpB32n6SqRf88E/m0BiDXuf74N1o/9Mo3yKbL5O1opYRPHZj
lpLTPQLl9vmkGn+N48rnpar/cbFxk/fgVIul2P6MXJvIRnFVeMvvph+epL6ZG4StNq0VPbYbncFp
A2UU9ST3VT4ARu+rDfpCu9cIxM7TJP+rdvfAJ64RfWgynAyq++NEAzD93oZH/FWKaNMeMHwcoTpb
OsTggUFA1w7JezNsNl/PRuJ2JSuk0vJsxdnKH/+7QotSLj11Y+gni0/Aef0hWGVvhgeT481FgEqd
VK6LJYgVMn4CziJ9DyYTE80K+or6PjRUgHufKX7+KdlsW8MfPZFcLasaikn/z+EzlGbNXivW/9/h
vcvS8/Jxt6LccTSZrvpBPvEOOzCfDPEuIlu1DI6WYO2vpQpfVXNKgBpHngeVgheac33DCwfFmlmF
nhsT37ab2zXuvfqqPVnbV1MxyVj2WECYaPGSvTxo28FLwOSyIUDyyS1Rb+b2N6C4V+KJAUaS5Z4j
HahUbBgMFD8IJE9kW4Ueg/VhJABjYzpdysR/OBdEWC5CMllVCU6foFZd9NYy5yutpsMUVGbSfgA2
30nOw0bMfxvIYVlBXkuOs6oKed/SeEUZ17eYj6c1ONnRnSglCxVDBN24zCgqJnMu3kVA0w9CvkhQ
nugtKytb0kshQugF8adqK3XC1I/o3pT28G5XGVXZAdMachjVPkUrBHlIUxvwhYnDkDNrLfYJIGe3
HQNgN5E3eWk80dUrKvFC9gKWd1W5WC/tvwNucCa1QYh32a6nkkcmEBqiJ7jEp2WfBRf755hcxwC2
F5sI1WhN7PdG/9YmWKkoUMM3XeqE7Eq8Y0qYuuntnTU5yvKTpWx4grgUWSHeC7131IgayIxwVWZu
vptLhld/WDTXU86w2PSEXt9nqVmD+f9QYqD86OEJ/KhWH8xXq6MwmrReGLHFBYqEPv3b/Cxrkp9y
ScPWtiNDRiltAOmyZVgKMhtBKrXSLXs9ZfOfyrcnvlsfGbIUbSXh75sCqs8ZhzznZpwHX7RP1IOC
ciz393D5fhCl9XyngPvPC8JGv57uOKGPRrFj5rTqAgC2QLjaJ7cVNa445I1NeRmOZrdDriNU1xEg
j7cNsSYv1fHq5kbi54usVzwOTmJWubcYZwC3Agszn3IXMdoch1RPf60j90Li8M2lSAOSzUsI6LoN
L+yt7WkbhbV3X5s7lAoOrgRJPQqdtG6gunLZ1g64Yelc7eS8BfksJ2CCU6Ka7VBT5l4FYVyICl5m
ZUNBYxwd74KtF6iUATs2BeeNBVFsKLsV9KVlMUb04fDhSval3G5F/3QvMyoYRrllcVioiecyxkvr
a2M0RByK7alKVYWjQvJIz4isw8EYPsF8LeeYiBiopzmAorvXVY0yoXhRkQ10eHlAcwrk02lHE8A1
dzdkeUUJxxptFSmncoHMOFpk+Dp0c6vd/9MqRWrvP5TFnRpvk2Ch8Y5XUnmKx7gliSfzE3H0uObJ
1lSGB996MnqckF12Bve7H1qumhlq8bqF2zu/BrvsMcFCT9Eg7rgmX7r5jMMQ9MGAE12NTXc5cVIt
8eVZVu61rLNn7sUnJ6+M88JIaTkcXUeHvxykrcDYwgB8JTjyTK7phVy4s9R7TL18R6MHr5WajBxW
zHRXuHKww8iUx/CZoEivnUOXk2Gcw8dn/9D/1/6UUpnmzxOToGw0HS6cj4QTxYwEyTsNH8jtWFof
SHu4Wbo/8M/IIgBoFi+xzC1G4DHoJ07/ahlO9+zUokaEjyqUb6U/J8Wa9GbxPpOlHjtFwdWolgQO
7FUfd05CnzJmVsseY+osx0LkzEh0ldNJFAUesrqIgfS5oz3pK+TSqNwuGzzJwttDL2wyvizAAwAI
XlLlWKk9T5PNqYMj/XW3Vqz5ZthNMVt/f5oV95A+X9lCpUOVJGl41OjBDW/Wvmj2aqkxHaktcKjk
oXF4ZtRoz9m0m5rhcRpe46KCofSZSlHjyi90ZrwIuaUPdYBIfvpQxSjvrPGXLDfrdUo4Gk/FrI0i
P4yWTEZbtNycPiuCyriW7Proy8vkG8iZ8eaKsk8sSBEmeRj+lk4xj3aV9yDkxtNNtjmgrQ4ECO3j
ZswFjvMu+lZ+60clnUbkKLWsgvfqYTWLCAQVVntbIu7z9jEPa/0TK3EJye9FH9OWy8B9sodn+wDp
J9TRrcJ0yLfhzkaXJiKzEUze5osBPYsWL6vLBJO0/7ohUe+KYAuz3rTPhh0y3YAq6bKGLZEuKlcf
cKI+Q3MrFge0D5CjAlAmDkHbpxL7Y8INn2CU/wUQwAuIqZWvXoUlr1wVhv83/aVXpSp0dCD0Ebhj
VOmbMgtcSNU2x7yLzdGWDfujs6AL3oql4Nf7f6j/QgVMj09sEQCPmfQ57zrCTkLSBWFQ71An78Ys
oqpOBv0nvDuIs64qCkHHEUa+yoFowVw3Te8Hf37V7t3CU7rjEQ45RG71tuvC63TTJW012UQhzCPw
srFCIIZWXIGv1e+sJ51QWwxzNQhzP2RNG9IKPHlS/KEe1L4TltTacCtA1RLeBNZM2VRXh8fPb3uF
AUCR6sfMTj4fbg5qcDNQirrtDhayUeMxNPR0+KYtHoSGPXqKYExHlOqXughSOdDXqoThjiPf6Yfz
jUnLlyt3zf5IfbIMy29zk4lFmk5T+n5UMkmRwWaXPzcuVro/PtVkCxXSuJQtyPlSCXxNyE6fhZq0
JpMNMXwmN2uc1+PDEtiPu0EdeCSqJ14YT8TmUNNB3+M3peW9UVP5LUAouBZZBaArtT09FdN8Fa9h
BhrmGkw+czgGxzrKOQroDOhyoSz99uaPYjFMSAoRBd5T0VlJq+i3qRYcsaEjubg2enhT13wjPin+
BZOD0snBs8lmDd3AgO8tY9LYrdxOsmR0XG8iiMT/uc9kMSuP7Q6D+nbb829oSrbWIM5cztlPfk7x
X/TBYOl/4fVzZSlolDTXd5z+Zx1QxtYSZSJcGz33JpMZlmk+SXtEp1WIDWj96VWvYtsYJ9NhNBLJ
mWN/EFiOhy8qM+krzYZ6RIyqUs50myZmiddaYeGcBzfTcbDRyS0fzjNdJwYVNYxmJ8M7j/B/EkBz
3AHc0iVDB+D8Xx4CwDAypiOr9uoChA97l4KrzIs4r3fFmG1xQZvUNHQZavgSaO8VrCTeDH6YjEr9
GnZfOBlQupM53oeLtZ0FZCgqLFH6NWGBQWSXTxLAHBKydzCeljE6ZXASYJQQH8dCkOJrF9BAHrzk
5AM9MJqOYLETkL4bDY6RzCg1t9XGmsRi/f1G9AjJjkjAqfFbq6rNl0UiTk5bDMJw1hHvkx/+8waZ
aEiZDDxvC1+NfqNaH2+32YweRTa/70lCVk6N++ZknpfA0y1LcwOowycp3Xpakgad2KDUuLAm7wzK
M5NFTBzvhQYDhLW2HsG3ijGiXwvm7CmnYZ3R02VJmWWgxvcNSUJp+q+PSQTmtEHMiMiTt0x4ZTIF
wlPeEiCIt0NhFLuvYDWfbMzotyta2yFHYRyNzNqjXprU/jrqJVKPUh7WylCP6dF/wVeZ17MNXwPh
Ze4zep40Kd0Inls8dUhcTNRItWVcDf8pXHVzwP0rhmXB39ftdoOOjjzXIBNv2QxjseCGrm1wQ8d5
x3C3EwHjW6PG2cZpP4iH2noDVzIO01k1Ta8ThIJoydFZxEr4fiBcxoZJGgqFLaTC0RskecYIE0GW
DBcu1NGhu+T1Wn4NrTMVa4LF5jqIiBRAZttGVd5G4na9Qkk2s38007eHP5ERyMQSWuka6DWxMLsl
M1LdHXUO6Kyg+MsGeO14HTaMZ8Li6YKZmT3df7BqwifcVTkc+lBDJmk6XT09Lne/ePVslQFgGokD
lpgNUESC9PmIBrexscyXx1VySn4KNLbdSDR1zohNbYCgGSedUebJ94JScGUDyXBe1AJKtQvsmGlx
gfn7+0CetqJtvHC2ep2upt1gOP8P2rlRjm7cixA4NzmIGCB/RjaTu+tFNX2sM7LJzR/BmfcLt2h+
GJwFbCcBXi5LMx/RwUTGo1DzZm3OoJo7ICWbVDHbfPm8NUNNcftQqu+2TBOTqiZ8g4xKD6kOVYG/
yZduYnF/gM8k4gmhgXqPWJQ1kPQAi3Gcw0MB4eODbpGHoBdmvJVBHx7x46oR7fVxMRX121ve9EYn
tCGu6vqpEo/WjLwRZrm54bhztUVvkzrFA1Oq9EyNSCC8uDQZdjhr6+pbcUCkh9rgWqDlX7utuunN
LcefqvLYt/LXAOj8aS8fQy9oM4ABwtqK0Gp/RugMO4YT0sb2YikLOajydozhdmzFpIFoxUCt1uyK
yVu4BnigX4W9Fpu4qtcsUvG7+x57+RagcVYfoXMUDNcYg549PIrmNgPfG8vdvSkIpK73UyCK2/Mu
azRp+Bj0xfZqOMWkKfxk/ZCt6m4q153GowHNSWh59VWBTaO/qobmgxdr7UJA9sDKwI825Ud7YnHg
HPW7DqUJXQw9M7pEdKEqO0iKKNBsRWaNPGRNm6fFS8qdVlEiO1BhiEBiIxTGL1yBZrhAhmTiKFrK
tj9pht+M90TrWasG90a2ZvJD8IHIwIGz661E6t/MFh4cr38P01GdYvxDH2v64LRWBf9kOLRMN1ku
csBRTo+pHC/QbWVkk+r/BRCt59cBBnnDcgtbyLefaHjEbdRr8mlHeUiBMmxgQ6hkvwfKA6hnxdUe
3ctJWMSbYcrxv1L9ppZXMP0ZAO6vgRzjMiL+nlu8ES/efHxxjJgus1cS86HsrHTWSnnIWwjv1zXO
bZEUrJ3/r4G0KNzvbvV8J3tlKwcSplqMnU1zzxR1RTSbJtCf4CSrbWs6EpsFET1TNGGe8k+GCBml
5PGBmNTnGBG5TyoTjvbHhsZsUJuoshU+2tzkIvx531EkJzD40nFdcxi5++VqbNUIAJPF0lxvXz5y
cD4hzo8RKlcmxU8UZFTt/a9d5wmYqSY6kb7r0CVffeWocWIt6xRipYnDFUlVs3G9mK71KS5eOq7w
Xr+KvbJ60iu8mphODMWMCxTWpwGvEGoMkrOgx37/SpFRzQeNizwepEapxHk196Fbgtfsvm1VgVQ1
2pfneonnO+3Ca1XjgkZHpO5mSATjhUlPnBTijiyWbBKSFxLGc0wup9N+zjSHk1X0wYDOBCQAQswS
I7xLQTlsYjCRFm9jW3QveqIj1CK2eKaPiPaPfQ8WevgKoNgIe9DyR9y9/81MvwFB/eUr377AxW8J
W4aT8W8fOpH+WHkecu0YdMiaCZXN6/QsRdNyhA9oeaAK1MvTLuC2NjdBA9TX2Qef9Tcj/RvYdAn7
bEoIAJkF0kAGMmoGxQxISNIlaO+XmjVu0A/3Tl72/yRmFyoODFbXcf8kafx3FhyoowGW5lODewaN
a/2TRmxKIoEwW5vpvAxpzYQhLmXo7R/a6lzqhqzRxDVzDkoufRygXjib3LuVvj8yKfAlvjNJikx0
VHt9qQ0nnoGUal7DT9TYCdnkYBij+hOQH0P1v7+JNMneKm+GsqPv69zJccl+5q5Cq3tpBuAfCf/a
Cq9eay9GxXZrz/6uER1Q50rlcIxqNrkakms0t7N4m6gMtsGN2B/6E2Q46vaOPu16mdo6yI8chxdl
wWLTMebk7XqJFKBnbfVkAvPQEbZ3bf+tEkHLDkMszOHfZv9EjbU/ZPTaHOO38NGvkPLvUd7cJ/ZX
dU+o88VXgAScKqi8PkUZyRUS6AyxQWDTfnSFbJQ7Sg9CuA99URLLmu5QOU1R1ZvAi7Zf4Z49jrZV
i8UF8dYTvB6DkmcTdTQIJYdcOZ8ZblX5cbPbtqBDRZ9msaNGPNxqPn9s4512yiUfDlKftvJFVXHz
mJWPjGvpIFz4WsYX4wUZJG5IwhsPci67XPEg5PEJg8G1S2ID52CmQQ6/ncSPTtPygNBg2mthMpge
nn+KxVi+/tYx6L3PmXtgVKcXkVm7YOCm2JuU98SvQZaUytpQkfu/9w8o1qSbxKC8Jcr18FVsp9Pv
1NY0jgcUxPiMfRgURcgeDsOcYYJpytCBgPvebN7XUdNLww0pjre/qpEDCMCiwanA5ASVG2FfiA14
7ZmcfwCHYOAgGQpri8UJly0CVobJkw1v8r0bRdhDQMqGBhD5oLOgQYOoJUvNbdsnoTdBnmJ63qt3
+n5vVowD5dOAtFzMdNyBzntnjq+j4knwwFkDLeilbeREojnfUu3XXhULMLpn6rvsG4Mad9nHkFfw
ApRPuZOnoDuP2kxmvUOt1SI0YK9sJ+6b4xUDXTvXFMS+vjBnNvCtRLyXhZaC9p5KRmr2adqGNsfa
EG7H3NrcYjcEca3x/pHjm5+lX0sEO9z2/a1DMhN+tO2DXBRX+w7nIexWRunOBtMPxcWJN93O7lKJ
fbwWVjsM3m5lS2mWXlSCdhHDKj5QxdjjDQgvBvQcWBKe8Snnl6cEl0TgGyP1xNASKdU/NOOYKi7o
RCWdU+0r3bYuAEHujUVIbkv5li9d9q+vgbZRLRiK2Gy3eDpKudYscrgtnbe8RAfHECO5xOpC6qQ4
fjqFQf/B4847rrXnpuUSfk6n0CxSEP71ZRhKaFu1KMCW6F1U55kcbL3fCkgGvVWcR2q7VTxgPWJU
/VRisXVBhVebOdGSA3O0JXpNqfag5yYDBb30B0yGUodH7F2tfPRgP2eISfKsoYx1hIIY/G4lhbBS
jbUYtfPNl1GsbV1b1jqClyDFSUUPm+ve8bs6WgKqlVVmFKrDy52aj/XOLgKATf2gywBf3cQSMnwP
LcctyZCWK9C8qiw1i0t55w6wRahKF/6W4A0fNhHEo3Raq8jgzYUoK8rnJ2p3g/hpJ3emjYW8/srP
p+et/9m+Ajuq9+iPbeT3Z2a9BEbnpNLekJPsE7EtcZjuvfl+QlPIsNyd5fLlv7EhENog9xeY4CUC
bIT7UhikyqyDbBRggxy5dekcc27/HlKTcmwPcU3P7zf7Gp+uN8XlwMo5aV+efAUhqMRpdENij9vB
rWyFVKVrkjC6si5SYqP72TGApHqO6XX6246Pc4HhlI2Fpjbw7MAkDMnuQp5Zntgr/lWwJbeJfXsR
t8xOh+n6Qw+5uatrlpUO+NPs1GI8KGxnlR8D0qYROFzk5PdYiRrs/9kC4Mzk4FVenC4Xqe7nIhnH
U0nYe+VIljEuu+8fZljHHwqKn1V22CAPmEybF0f4gPr5Pl42H566db6U3KOhwwGFqGLstrvrn4x2
aBf+83vWjJYEU3s70cdHCP4/zXbdnCY4QceyZxJcrMk/x7JtRhPn4vrwkGaEq06Lwcyz8eb+P+TF
OuIHrY3FDdaOEQW5G1MEsD16yu2pzp22K+oP/gkMRd56eAgL0KAVkoy1dZXDc8IEEKzAr4B7j8Dm
EuEUh4BuyEc+Ds1sVMeuYsBJewEVowcvm+BbWFi1+bluOi5IUiSzR4vQ4nQ37jy6aPjnKkMdL4Am
d4h8lrMZ/QU7lEfa9kNvI0431PJ5wwj1PRhM1vbnGMzt2+BvI7T4h10zrnhZbi2pYXAGmoDHuNvi
d0Od8JeOvRgbHqMe3ds4lZNz4rKzcv16sKid6I8UHMT6auSyvom88TV28GsPQCT0Xu+JlPgJ5Xu/
wmd8BLfMyPILEfeuH1YryMK7FuG6MWDs4t10x70UDSq5ubdwlQSsDzHGdwtVnHB7TxrOdMFVupMP
rFnlSIIsMwak+7SfdtexIsgHVBEvzQ4tBHZODHydXHzobqsXaKNQLyP+ZYfuPmHohmldMSB9z6O1
00erSXZSKja4h0iR9bY1yyv1SNff+asl34U9OeMi2hlZb6v9AhgOY699bWroJfZvM3iPV4bM+EQ0
In9JCammWMvTdGo3pCMOD0RmGczWHE/IkG1vCvZ/b4Vi6oCmKgEyDtM61NIlnlLBP0icpC99Ak5+
ujmC+bvo5ygCYeNjyJxxJoI2gWSfwQnpxQapkblGltziIYjhEDZYsqT1pdtSV6gDR7WwLZNBIrcH
b63pfS7kn2l/tYXzWN7Vqm9BZVp0hMlvawfpP4K+mPV75hJBG5rhYegra24ips9HZH9kJqjpMIFH
zdDjbg53n3iHrrjLcqXFPxTwlEE36RWhKYQfXzXDnvPgB0kVP2GZNPpzV5WJei1fLuKR6N2z9QDQ
5rn7Acui5OVSvCBhb3nHh3RF/aKCimV43KFQ8jx5QkIEV1rwfDhksAsSF0iLoBXGPfEOOt94hG2G
wnSLhCqxDiFjGKE7PlUS6wxUnw+zJwjP6X7wKw7iOZzLQixAt6uGKYiYz4VXN7XGa6sXH0tHD3LL
CCUzE6gLAcnMRvszzYoCNNkyfpGM8YsK5hyn0gqlNn0aVTttTykqULRz11dz1XOwsOpKV27ANJFk
T0HYP90apPAaJf3ZchWA0hOvUi6N46876g4kch0m5T/DI/mrgx8orzeu0qOWnARxNEOeb7xxBbaC
Chd52Tt9Jo/dnmdLcyotOHcHYFz9LQcgiPexDe4RUv/XfMhDhK+IyVFGWP4N0ElJWq0YqPnLUgCo
CkRm3z4EkEFBJifs7ZEzg+WwQ/N6Gied0n4oymLb7sw/4Z/odqHRso5fOIKaVhNILacmvdSLiZci
dn8IutE/v1RQSiKB6uFzbsp4Iowua/irm0WCTCjUHi3entZQN6wCFrPKxmcYfXWiMsSWeaAAnaid
A1x72TxYk2FDV/jUf2vwbzI21YdOictT48MbxB0rylRE8tPtJAhabRVrarb+HLaX3/sfXgaKSiSq
uEf/tinPwt/uJvDm74+gZUKZVvO6iniRatXr5T2+NLxO2XZOfSu2itCFtVTMcdtHvgd7pLAZPxbj
kaG7LOO339wN3lT8j4/qRJ5EDkDHZbsK2nq5yLPEb49uMVbGvDGVS+EIVTznFSTDRLpKXCyjfquY
DQRdbB80T13EU3Sev7lCqJUXYjebmHBWXI195KLdVwhZxcuqItoS9+dL5FpEuyOJ/d8kh57VNnNX
RzBlWi/9nis4bq6MCZ7Vm87OyDNqNYWsEYy3AETpmZM7rQq7NbOyMlX7OwlbyqjHDsZBPAokVpu/
dhSJ64BTrFijKL1TIb2lkMyoo4QF2hEccjb1VEhr1bIvGtX/QfL50dxdSgRGij8DCDKuExG3lq24
q2cq4jpFyuJ2XNXUilcBk14EtmrF0FUH7UxzMt3j9rNe87PhxSeNT0hkyxoemuAC79BkZVvatE1B
ONL7vFyqvMiO7JkkMCbJiLDe286s0Cg8gk/785M6gnukd+6RW4e0cEAm9xmu2FSFfjC2lagXFq0/
ok0ra5FPTdHWriB7oaElIntNseCPaJXgKwskv80OAXFYym4sD4LF8NgQYoyC/Vhcx7xQ/fG1gfn8
6ptKHBdq+5fbKBAGmNPdTSWzHwVTuj9xQwcensPcOkC19YjMMBV6yCvjESFGeoNqgfdLlSmfEFQc
U1uk6A8Y4h+IdmoyB56oqNra3xL222Z4wCwQKcxVvZkzVhgqNHYSdVUXtmpuSpBBurLedKY8IVG3
O9NG4hdGvgv0OHMx60xer0qSCaiwHTyM022P88Ohg0Ql5CSP8GgOi5qvOYVqyNUvJOMtP9CGI2GY
/FclfbfS//9MNGHZKqS8rgYrXPi1LrHuhYcUKzE5LZEznwyozL364h5BIP4rOOYPmB2xX64Qx5OC
M3+OkCVoGRCzoutNY07h2aI2ZEIi/tXrPkimAyCQH4mzrz7/+dRSigdBnGabKw0a4Fhp+EqFAFzI
GCmyb7ZdGpl9ShkrSE6PkgzPtUNW+YayRdchxn/DIIjva7xujFwEFWhyvkryOj5VyyMmQxj6hLRZ
rvxY2B4AwGkaBFmKIAjaWMqTX6ygkScc1IvBXSXVtmlz87Ltha5HzBq1I6GFLdEv4yl8cWONRPAS
hRGO/b7D4DFUyeMuMaLLK/SAMMP3cFf4ufV+zTC8JyxsURvJmX5gd12VrPXawifVpMfVU6bjMYiH
9FsLHh3qH/ME12zVDb5JkinEi3lnpg2IM55nOmC6cu5D0VHF52qycBPr3xIDf9Jh9cp4P0+uADMe
F2SVKh3yNrXO+k9wxT7M5JXdRZV66WeRGO/FqsNF+BxKKa7ptzYg4M1wCmKHnS4cKiXH9YHjeBUb
qxy/jMLuej+OwMJnOB9KhrGEWJbP6FzC07gWdB6Lz/j5s4Toi5x00nZjp7GpJTvcjNNLvIsxZsJY
CHq0caJxFs1Tq9piCXHaiwsdZC+/mFYco/FKGCESVLKKD+UzeLYgiZCJUUlfigRbmTN4bb24EHHI
UmpaeX27VM7cDbz4w2U3J4MR7KeFCXRi+a/Ajy88XZ+ty2+IylhVAugjF/WD7JdwF1oRsAHc6KML
OFCJyPJcxmH6Yj76p+Km5uUWyALPmxIae2LvuR68UQR8TRN4+1L5Lm/LxtRvnZ3+fr8bx+9Ea2qF
BaSuhMH3uZpCeMEr5MJ9tmhZVDNJ9yUzbKuc9rSWiXsngKMRnJBM/l0F59IhWSvOwwgX8a5/xY6Y
lIuCocbkJ5FtB0mBV1neHYVlUUMxQ4R2p/TYAhW5Gwpmt5QOyTZfswqWX915PQNLlNTVyIAe+XoJ
SsxkzNnBSb4f+VZIjL9EcTnR816SKDiF384mu9FlDtf2LqOb9swkfarr+WfuXWnH6/lOFMZefo1T
zDVfcg9WcSpdHK57+XCLs50mLZqQIk7vbYIIRsC99dH8R3rNUbrW7N9n56sBwZGaCFF3ihpfpP0G
MfGfyspJl6QRtAJ3aItg4iU66/R6FrXkC0ewzAXYuW+wvHfrxh1hncu+1XL+Df307mIAOc67m4ZG
j9TbiIQnENtkFxZRyub2pLnuS6GwzPHKhG2Oy7F4w5L7lzVjlmsG12qh4TcVaRHanchHf2c/2PHs
7DqQHglB0Sgin5rqWSzf2CrVBPHiD/gQ4I/TpCjzgXzMM9lOD5DxmVLhrNPY3QoE+VVT5WcFJorZ
+2UjcDEIib1sNLuiIw0MGU2uplJVRdIj6EEGVJgLRR4uTpd8ThXl+yLC3coguLVbdoBtlOwtJpsp
di4vDneov+5jUHJWGtyL75ZldmHo9yD4d68G4jVkqPlGNrBoFNTEme8fS8xo+Qblzqaoc6CrqysZ
z395FYgk7QhIaLJQvv3qdkVPQGw/bl4l5aYAKNN1JSh5/Pl2GS34swTDFJTJ0BmA1H4af9OHHaSd
Fz83/rtqZ+rHzVd8PdzpUpCcBwlwtucjkOCCdURdHT4pa3ERwMJySbG0DtC2kFiduZGis9O5kMCU
yMxUfpjZmzxlWEn0YOMGBjJX8O4UZodohMhHE6hGxVSs3hX74pi9aTTVjb6zI5KEFqXQaRWdDYTp
5AdFziwV++7P39WZAg8DSoLK84tzGvN2wtTQs+7ObsifXYBkyq7PJIm39F7Qy9JGFuIsYyA71yHZ
vLRZ5QZSaCubgWx5FD2iOAmkdjn1mQ5wxJua29cHqq1zd3vElMVfT59b3OPSpvwltaprS7YVHgAz
sT6RXI0ZhsA0ZE1/xGK9buuTsjdADZ34UM+JExXQcLpIdtzjdgmdgVGu787RyYZXPH/oqB7hujZ+
Y+cd96/74XjedXKfnY9SB5HbNLMIb9Zw0gGxVOfz07NJl+o4ogxJV8GKMgNejMd414mheGFo7oda
dn+FSfGaP4E8CX0ZW8gzLTZJ16MxhmQ4Oxzc26+kgyDrar+BSyvOzQusWqOf/oE0eDOWbjbQoH7b
o9E/OdGKUwO45GJZCHgzLi0wtznF2xJRD2Ep0iquHkMpq0+jKkU1e+RzW4USOsyT3AWuykvHqawv
zgnPCc7L9D41aJJsMW8zVLt5wAVyVJHfEV1hM8fz6yR1HSwnGRDKphFX40rqtHCBMpPsLRYgFgIx
7i8P9IvYqLKg5WtbgcioIGYWBxHMfBjB19Q/WUGOb7RoAVaB31da1Rzk1JS/ygJLB2Yj/q6Vfwb/
zYE97FuKkkpuuvMEgyxpUOXUy4HsirDq51Qe0CoHefAIzl67ObToR1SeHhm9LhUqHUg9+3oia2ud
NNiOYHC9RKGOG3VR2Q/VX9jyXpPfe0R0mryHrS0T049/0uAvwUEhN+0KIzlbFdUpRDSNQqHMJq+c
y0YLw5C/SfyyeHWlmDJ5kw0kGqCy66cnU8VJEa31VpgrMnI/3SDSUCH6jIy5h48Z01TEX+Vjx1CU
RSfeGSpu6iP7mGjhovlR5SP++7149Bbnfyey2oK3WrQO4wdmdOV7DMdHBzDqWBJ3oNecZHmcH875
M9mksousgN6myGSnovUOklTk/WwlnlE+zikZ3CetJEbRE81A+qRjnTLATVrJJ0cTqcBe4q47QdVP
gRBd1goinwGLe1aH5AFMCa0mz3mf7kVj2erTeFabrBEQtZESyL5FdB/FZI/FCIEeSecOM34jnzZK
Szpx7WFWBCk+kM3/nWPVqpI6FRtZtCpQC6oGkNs39pYFpVZF3I3a5A4n9Elubhzc4bJ3ymL+SAqj
OtfAhttDUjWtJTZ8cHMTin0QpJzWGdSvvX+BNMgfNoHaL5e+XzRLXqHLWfpiaTjBDjITr2yzPBBj
4h03u3GsUVTfFChi8LSqX3YUIAGck8zjWCUhHLX/9tvPLLnBSXY3gQpvB4zD4ATwsYr0rLaJsPcU
rFAMtJ1XHzFzHWbs47yuXvMrrinLLvRU9pxn1W/xKvLrPM/lMAj0ujBE9ASdPkkpSH8B7SNhc6Bg
W8gPiRwZk7Jx7OSMu8CjrQq2FoJ++YTE7b7+M/0kdB6vCLJowhFyJw/QBPH21SiuTmo/+ZYeu1vy
DTtX2dk6X2Om/oJQUKSnJNRAlXEmgvXIyFB3QrKPP1JeZBUy+im6CDZqk5JapZ12Fuq5jyqcKv6K
yiq6cxC8U9/D2lIMC9UOrdEgfnW9aRICZ/ggVzMY2bT78XveQwfwyXJ/bX80VzwJV2/wQAhbsHFD
+NwqVgdfnXPcBhnQ6VEIVTJxdP5uz211siXIzCOGJNhXkmejYXXcydz8Ef3VrlwMlewGg7QiFUd3
Vq5AQWJP/krCF9d002zkTtBKyFK3BGpygfcI80a1GX3GRnyX3fI9YHeQexpLcBxEMEpxX8g15mjd
NsF6T0OvxzdQnb6TAHTQe/xpy+kULpxxO32FXuypomS9cuaIAEz1xpoE5VLjYtVyMc2VBhWDTkxb
j8QeHVcAGh1JgBftMMrfFSbCXnv6NuEMmHJHfZ+u+6JVr7VKggGfjGKER7GdPbCgfJYpvJiLvtVl
yz6mV4t26NVWiwP5bPpLe0FpgR3xRvXiCobSLNbt0tup5mj6qfEPC9gh8pr3GQsUnGC4pG0OjSSO
3dgE5Kst1D28FaotIinchGOBOszg0DvULBjgjQ4pgTosTVMxYRK3C7dOELv7Nw7HDnTPhlqD+iBq
My61iZsRb/C9vx0b7r6MJkB8A8+XJ2KrspN6Y6q9oCu+pUbQpfU0cpuA6YdaDjmNKuGjunQCFsae
6kSF6fbYI1QTZwCxGCIT31LCEciCDNeN4o8Z0/hncOOSodPbEEizV5oslx4C/UyEdQIbFRL7EXnC
hdwToBWsXh05LdCbAlaOuET7cTv6z4J4wieh+2zNQaHvKVEgN9HVOl+MSrF98TuzC+NnZKgbJlNe
gVNgv9iZdrWLeF1QyvuRK+w4qdaanDII2R3TfTklZwjIzVd+51DQFT77FP6c3KFsLlBqQnYie5nw
bFrlA45tJldGqmtLwHxrtPL9q0RVCpIFxJ9YTunLvMKOyuI8HDKwpMdbR4GU//cvAGI+kyHu4I4T
iu4YfHw1z3vZEjXA6n+p835tTqzPYDZEiA/fhW+FCKawMXafRiG0cMnbzcyGikPFeWcldaepxEtD
GsXsTWpHtKydp3e4Qr7CLzVdtQNgiYNFRrHKeljv2NpJyyl0P+S7nHwsaY3NjyYPUfSWvSDtCjin
wGNU7By+cT4Npf8Z/XY2+dhTRACt0eKjSNGlzy3WiYOIh+9d8yeRwU65Y1TSSouzt3uRo3MEg3bq
yEl8Zz8RNQhoUB1vs7ck9QIbVwvmha4rThIDJwKX+1/n444WsX7cnWvwdjofX9w9vIjK8Ym1KDsi
cvw8AxQf6JqnNRZoFhyjM6eGya2/xdBXhLSWmlYC6JFDKKUxB8XJZh/mDN8CNF8yHOw8QV72Znkl
TmKMq2KcJHMAlqUiAMMgaD6hbqsuASHGpSF0mWcnbEB24mD8Cv2NdFjbm1cnLBHRuNCK9/3PBWFs
XWFARosAqvAX/GwZWokD2PS1NU3DHL6QTkpbLI34nmMFPyVg8kc2J1Rm3cREKG/7rGYV7e5eImzE
u+rJordhDOAT6UauSmD/bUlDTIlGVDSDnltbI1AvCExTPcRsRP4upIZ8Mm3YiFBb3wCo3kduF21A
dTPsf4zKwUjPn2xmwddJqwz8wWrmULRA3zha77OjRosPL5wBEaAMrxVlxSfSuQgBw7tcYGJmMd8Q
n8RTnBNCWoTWah0GwXdv2RiYNbdJe4qPXC3hFk2FaolpDyRutQxTaYV47DJzIwkZ6pv9/bXAQoYs
wIc48biS/gvcdMOHNXTpdovprSAJEB+NXaFTjCBFLSv5lMtuozYI8whXwjJcK59TIvBkJEk/oujS
+Jq2sqH6Qa8rEIY5FwzyZblrw/s2qERIlui/ulO1Ha1BmVxo1GbJDgZ4fujyJBUH1lQrxAln2Hbt
Ablqpgwawp8MOwDsLOh9lVL27VNgvuSFjcnSLPvb0Wa1+c0tgSEiMiCN/Y9BOMqDqgsB3o2z87dK
JDkFoIse3jA82LXUJn8/WUhs+V22XqooRbCCQcz9SH6w2a7c4CvZt0P3Gm15yDBKWWTa6w3Q7lha
vwFp6i/JPP9tuYTv9iVi6M4k1rVCUw93lpAit3E1DGoPaf4xOAC78Q9a2eIbAqSZqz3IaegLhKPo
vVAOs5pnwSuL/HkZuflI+sEDe+UKUSCJAiNcV9EJtcPQ1Zmi5aNVSRjARitewk544jLTeJDmJ8dT
FK95KmQbs5ldO0yvozPeKU0HCNcFZZ6LaBZDzfEQBrjbzyT060GFr9N+Yr6L11+OFJGwR5rKbKt3
MdxTTyBbepwmS+Ew1O/JYxaxRKUH+gz3kXBvyK0vePkkRsBLnlQKooAWPuFrLzNJGOk1047bQjE9
Zj47D1olZyP4F+nI7k3R8GcmobwJ7sWS9uwdtyhlwBh2v7docGFFbll1SlCe0AGMGftYClOFkWla
qYcfN5yiTAbtWtgfwV3S6AiJQhbedv2h3yZeSFjky85nIBdbaPwZQAcB6ZbIScKJmKJAobmNxKQj
qg1c94Qgns8nsT1n/YK+raFuJiO1Q29IoVOWnnnnWOXGxbv+XOFV3FinxySISFu9qPGLp68PWENp
+6XUVAojLGyndMsVb12M0dWvviMcHjFgp0ck5uvTT1d9OrJMG8dAaBKiyVdD4kWvExb/Y4ZvSaSU
nwFor9j4JM/x1tvppiW5ThvM/hsUk+JUrUIDYmS4O+k0arYQLE/Yz6PGybe0h8UqKo57BX/fxdCG
+0j9A3Rcg8tNFf+6p037muNQNTsZoZ7v7sqQ2qnS+fO/GPQtTdanckKxeAztYsnYBUOqwBHBTfUb
iAjNETw/X/xyft7eOCk2YSxA3Urk7ZyFxS9cANBOX0eV0JKSCRDSrbALgeOZPWeI2dUO2Tayd/ec
R8ihn4f1wXjb1bQYsdTkb5RDcTzAQt5UkLjixteye+EFyyb1PVOtasV9UA7gpm+Ou57AhOJS1o08
k9Kt0asWkSho7aotjK1E9QdvUekUt9Z0ZSYtp+zvbFUnvHjuTZIF5Qb9+lHzdyDfGeY0mwC/A7cM
gCiDIq6vhM3FBWlUwyFMKb7JUJg7RJYXyDOcztH3EeRS7R+dSga6xb90ERd0h7VJXH/AEC1A2S6o
1zQuQlxPLjhdEZ7Rg9Fk/EluTFjezlgmz3BaplMZwxoR3ozvhZRqSdI3Hn6HUa94uRNCTLsX4YuF
BMMjVKdBFxaJhH8zMeT6+AXBZJZFKB5Jf1GWY4eK8cF4S/e6oXMCnBQdD2dwiQA3vWEN7HR4bEHm
vaspLVhwpfUSsRthGW5Js4KxcQqP0wUj22+H26WY23RD+v0wx/Diw2DdZ+PCzWlPvBGtSu0BB9r3
VO9hTjo1w5IgkBgGsSkwpYeKT8gR5FOByTujzEbEOABqWcVLBiCGxvXfPiysjFzridoUBRg+bGxy
fbr7Y05/lBWqS6tVBvlbcHQqhiaFSQnifT8uzfWg+zqzorZ7CrEwvlZk2dvkDM4yr4Gk3sox/nI0
WlboS+wgXuchbHXosBk2NU0TbBIYyABbbPWsBubKOZwI2r4ojlneDIAj2ilCBvTAnCy3JQQbvkHq
5M6leNw37Y94iTEL3RveJCivokrXZ0b0+bCEdebuJ381wTesumde2WzdQuzF0Bbk7OmpASYKNgx7
ogX5BFoGDCX6YVx42WjKldDby0p1VB1HsA9wzy4VknMri02i9Wk8UCBn/MxRKgqrJbWGMWSk2Wk2
kpxiunmlJ+xaTqU+mzKfj+hpVxcDvnqrx8J4hQZtaS4LSg9xzmchDCXss4FA+THk3JUyHVNtUydE
QS03ul+p1CdDrw+Rf6vgd2RiUoEmYs6GYJFyb+ZadOZ/pDF7J35eOec6+jYFC2dtak8kxZQrO8yT
79KD+KDg057h1PSwY1NtDpx8qY5XkRvGZ+Rou7TL1LRzuRj/puHey269bkm56uJiHH7sdDH07YB7
dFtq3xvb3jn0pJma14Lyo/zRZtiqBEml+3qh5glXEqYfpyFNDUx/sUvEY4RC+4y3jVC9Ic+O5UsL
xafkyioUxX4lad+fmpiFSI9x1TPRTjgArQdYcaoq5i1BdAW84iCq65lfhFLNeIwUUGNcZd3ZZZ5t
uqaEx2QRHQNXjw7QDG7cYCpbQhmuwPlg9KvNFmozhv6iUZNguOURbAn09llTU2dWoREqpxlg0bHa
yujDWvrFD94j9mYhHoh6pLFgWST0JqR7phy910tKmjhGI7YHGke+sHNUgHmyqITmoZXn2JvLX4wr
UtbyLM5f4B4YgWKcih99gynPXOr4LdwFpyr74SR8KB9FmILeOKqrKnq8W0R+YbPl0Yjuu+0DdGI8
2k5YZ9hjYfqTDC5/hJ4XAnQIgd2ScaC2zpoap3NWJuu3bg4hvGaT8PXqRLe17g0tFUaS1oUaoasL
JvRqS7zqz02iWFxkxf3KuP0MPeojewdWBK08rMRSDXHSFEOy2qWyvUhjeBTq9B3BtAsyRIQSvUvC
+J6dGCHGykzKbaHpEFBON7ia/rBAPgh0ZUSGuQYraOILiXc7joN2c3PKiig5/NOfRoCJ1vq/+OYF
mULdP0m++4xScpDGbCohqSJPAGPjEVUdj6Cpmy8Xflju6HgZ+gYMu23EO5OsEGrOovAc6aLf//bJ
Nv+W5ucR9SYMNLxZdNZ+KLLr+uneo1BCeHVWaEERLWiqNT7WYt+xM+v+UrfRx0w0t4GdHhQf30SI
0eLWzB4AVLRtvXzTJs8EwWH7mqFRHuQTyw6CmC3SupkJf371mLhRQnRq7sK9jit91HmjMEu0agn7
rgAO1wbMyR5LcVcSbZweDc2cxYE+dBNmtAHMUFXCYEiMfJTmsSaae+R5lkVA1XKdr7OFbn+usBev
lnV4bURQOltECNFFxP/0K7GC2QgiZGwEdRnJIt5REJtzEkaW+1hryxjidQWfxdV+YRzKzSMLEXqB
uLf2krOpdi058ADNWqphBl4O8sRd0Cf9c1xQErO5EJmivVO7owUaKf+ZiLpHJmoZBjYdANbmFj0t
6f2jqKvkEu1r/GmNDi4hh3DxyhGrJY8KQQDv7ulNYRnuznfHMQ1ZbuS3sz8jhj4D0K1/mzvEnvWi
QL3nE+nCBBLE1yQGpWoI9dX/CX56KDvRF/VEM+ZRi6y+F2CwH0YRPIsbE/jO+iQ5yzK2Uiuesx54
svA8oQpE4Ez8cAbSskIO8wXwhcKM941RmcwOy9PjmctX9nhwhcLVtg44Frw8L3kzuyBfZ/MbGYBR
YW36BmiveVpwXS5hfcyu0OVUYFa2F+v+JKayLyGfWbNuqbJPCA5ldQVVIzf97B5axZhrPnT4DJtn
IMx6CiO1Mgt998xI0FvXWKNn2S+ytfQAZMKhVxTXe8fw6VO/LK/kqz8thymgiJcJbxATS+81uimt
5itmBoaGfVeNkrxgOf37Yucph7HKQPEAxdW/yoOH6lRDsEtrw0jc1H1KawCphtuOpFacQ5wBZx/n
/0SpfUdc/Rk0HeMqNW9REp9Saa2fUCUNCzZe6fxOkp5Q+38djiSifl3CRPjVd2hizjVgdP2lJGv/
Yoedw0BBvDk4N4CRXSGN2ptdsG/y2TG5+/3xEDE4pkmmTYM4PLBn53b7T4cKty0le5fYbsdDrZml
ekkqKzjcw1TVxokUtNZsfRMgFa93zvz+X6Un6pITWyXPF52rtkPdfLYQqLioFYNYemm22BXUOFww
U/RgH0SfcUHT6oKZpBGsB3MraI6joZHv52zwOPS/EaevJmgcUADInFJKqVgjkKtxl4tnjvEqVQUx
0RbIvXWocAVL45O6+o1pyNm/t3cwfMtze+sTADKZSVFFss6dziNTA544nfGa88sxr8R9i/mCgkhb
FHOJM94UeNU93WBhLHC17NlrJVJ7uGjHnX/XXWgPZ/EyaFMjbwjscF5a54r1pHlSQkSV3ZPSVRQi
EAbpcrfdRXDNYik0SithXz9Oa8WrLbG9pu/Of4VRWSF2YBNEUF8/Ah5snr5hfvXQ6NYJMiFIzyaN
/co2RJpvUBsZNxxLhFckVHlWRmzimWMgg6JSEFV1ZbqTyUwrPgMt+r6zVTNVuCfAVtynWoTJIaFL
nhJMsPalQkWdhn+qUWm+Mb7aMmJDOEvno+Q0ps2xwsUEgZfcKPk7x9KMJF04GwRJ+sXvTczGRS30
G+XXB4SPSyHV3vqmLHULem/PdXJ4kEaYdWlc7UpkziyJEbdOzko/Jg3ysVu1rnPYy5k1GWt3Gj4L
ADW6h65zqP/OUG8p5zV9Iylh1cDdpwp8ZhL4YCx08RRN0JAPNRh4pgdMaf4/5k8sXnrTHLLnkePR
9uQiC4QgXPlMKvKYtgXnhm7p6XM7Etxnwfx9SBAIWNVTkU03B0tfp6ZN5H/fVQPV3DyylqB2yM/e
CyuHiiIMubww0gy++nT5Fbu1hRb+lKIfIYBh63XG5OOqrHjiuWSfmLGUpNa8EzQ9jAvLBMqm1TMp
Alqtup6tFP3OEaCn69k41tsukEbmj6eYvCk8sJQG+e0chgsgA6j1DBM/yey1A2H1NqjGm2c8FXLv
FpAjRlxr3+YYjw2E0SBgz+yoWCIuh4BfmymjlYI4LJ127kgTzdo97FUxMnHa5Nb/XusTtiOQaNzv
Y2H8sJbwnXltlhndB/Aq2KUArSKTVcqMt7u0HzpZGBRxmISAMGaISx6DmHy1lOzAVmH4tc++pgaa
N+e5bTtj9CGZkXjfHLrAISKPcUCrcwiZhvjJMgcq3z2fEA9t3752VoKq2BR8/NauVasVwdhQwoQT
ISWA+gpfmdykKT74Ixe+S8MjFSa0pXGG2BcUwMtujJ3k7ESl0DC4eiwVYycuNuQQ56cWOgVKtZZ9
d4xy8Yx8xIRYAr/Vi2ar3INs4x9VJIFBe6WiXbBo//rJspYq3eSnHwPulUhTvAl6Dn0PqvphUrTJ
1wZo4zKZT68YN/KVhYObJjJgjD5fWlU+GP36uWrezwl9L8XMikzwAIV5+GmbL0L+UcRVGT2pEIs1
Nzc8RZgOlU7aS+S/n4Nj7dI5vikMbb9CE1QzCY60o0ywSwwFZdY40d0x/rRp2XT8QccpCso6FcSf
2xqGXQFFLGBl638UfC6oUfFgysGLlPCFcSrqDemubAjtNZ1I4J95a4W7omdK9fMPebsdC5YQxwL0
8ZCdVCfhFqmyLhhEPBQIlZbC+k2ROAAyvVlEw3eHWdEzOyVOURJ0dDOMk/8cPwpKAax+eAaKLiHN
w25OuSBp13QU1xYS8OhXpnG+fonKecU5FCUmvbJv6P0mutZXFAfVHQmle3YPWgxJbvxS0v34ICnS
9JlRfy6OL935BtNShLiybb91yXU7aXwwzewNuHWYLYu8wi8m34CZDnVR48hLgH15ly/CDUAayb/E
VdlYgqaQc+bpzA/TssIMl6P7B5PXqCDgTfMtplq7gqjI/GPmjXpPUExieFdEF08yCI6/LjAHc886
2s/RX1ftGbICQKhTcEQOGEOqpmA3heceN+iuFVrXS2n7yJGsjyYySVLnTL9yeePhb9pLjQqrE1+V
m8YC8E32s7Ygjec/Ygc8TzHMm872gSJfLeKQ3H+miqLaW+MdQ14BVt/5GaSuSoSeP2n/cKwgeVRc
9B4sXxP5fLyvmEaCet6gdEYFL9e3pIX3qlDW0WoGTTrSE3qZF0qh9gdaBfrj9hj/FGFaL0SoTO+w
rP7nto+3x4d8Y7CYs01lAIWVGlI70jKVjX7JImutpL1DS7xDXGQs40OlK4GmN4g43h7KkelBsYKB
skI9W2+NFnsfSG0f/VDWupF5aW+CAT+cUN9Lv8CxtM5NFFlC+fhB0wHHux2FRnZGC0baWCeNw3iw
RjggfEW9LeXe5T8UzfVqKFlJyUY2jsixNxwF4getiNvpemfaMCB/Y4jDQxnCbqcWUPBqodUNt3tM
QyKJcGvwvbOQBY6K1lTZddGZKnmWf+JL9SDI6TpInFy5P/XqeFu2sN9D1h6haTKk1TiVyCGHvq8H
5Ey41jlbX7OmEO5p2yMF1JJlRurexM71z2reNSgG8a7cHOUAAVr0fRtGXhFbZZaBMZ4I9Svu44Wm
Vcn+TzsoQ72kaWP9EHjPFOt5YEa/AH1sw0pYalMLUGmaDrCMSeY9ZmYcB66oeQqbskbqijcsaxoR
SU675SxVdl1u0s+K9EhCr8uQB3TEaORNFiA+9oRJAHEMg7PX887W12S0uOFw8ZR5h1rVyKop7OCh
zxiTnxwKVdkB25JlYwY2zxNwvmNFb0YtwDFUJ8EM64XbUDTN97GU9bIYlWc95hUREFz0iFaw+MDQ
Al3jF/NFPPtasfxwh6WYNB6WrHRte1zV+enannTDLxPsZarl8UhIl+3QuvhyXveMs5t7RE9qTGvs
YYWkyLKw4QIUbL9VmZNwmIJV1AkDq6mUOnvO5dUnSFtGJpLGwKB9m4HuYaoUDSo+IO0rHStGs7BJ
3mEpKqw4EwnPMXLjy+Vleb2DkOblXONKLd7Jf4c50p99rAnfMQIFX4o2puBu7kBMHEg9mgj3KCg7
PnrcBS6PpSnlWJCX/E/YDkPxT5CvsWpzXLNXE/+G28reVLTPKqxs7sfHuWOXrIItGTYICvNr+nHI
j8/H9BgvPJCT7RewFcMmpFMbJEWPtZ3EdAISemEPCjsJR+FlhG5WHuw//7gZZS3DzVFZyhP3bqur
NF8DpT4s7R3YGWLK0jmaoR/DNH+MerOpuvq6nNtJRGvFaZzDWQnZi7q5gptWJwVSSJ2A0ynBcziv
WoyWR5cGrWtkRip5Hu0IWfz+SaMDnehgdEc9D9eR6NudDnn8mS48vnLlDVmKm28OrAX1sKK96BLq
Og3x53ABQ3ssPVMvKUMPC6UNCQ7leVexqq7cuTIsx5sLotORDBOHSb238q3U0yDfGq2zwZsB/Mz/
qbCiqdonO4Qok2tNnbZGFzB6NibNsoayqJve+vCtNaCfUEjYGhmHjdNEudSXmJebkKXrNwmIcLV1
32waLUpVus8OrHFPb2J4T+/J6dOF0ojGU+VJEMuFQHQzpa1MvuhUM0mUEGFMTwsOiAJuPR1UaP02
y/oBrFy02JGfXVm5UbJpYm/AqqGjZviDycPclXyAV7VxrNS5YcBgtMucPwBv0pWBIUThaJH7FyNA
fvvwQ+kxJYka5t9YnYzJ16HiZAYIU3vYqNgLgZAU8pPVp1/f2SDZrWQBiDCtdbDVLGC923lXZf53
LEmJQjviHGDhU6RL0tDnSeLASva6D3dsrQAuLpwpZUgOvMvyUNh5qxkb6ejDuvzdovt2VTALqQdT
baCcdPPrFB/32gADi1MPYSfPTI3bFogHkT2bNTVtAcO70mGSbA7QzZLApubgcfgxskF0pxxMXzhL
iT5doUNn4+mEuugrZsnQxHDEe8J8J1SswrAZyjg7LiRwO/AI7ESoR+02ssYNEw2uyTacHmgGbKMq
EKnlusjKEfH2Gg/IdmX7yACVnJzwZ/exZOek44u6MKWdEPvN9jKk21tzUIlxGc0tksyWJdl539fN
KzFEBy9R7G03cBYnn0VAzmcjbgvDU3nxkdMMhKouWgaxJ4ZX02BaNIMJbqs2306KwhAq5SPdfkuY
2Iwsfc0rsJ+YhH7QNMLVRbxnQcscxGrucNlVNuXGVU5pJJG/skumk9rmDGkFUFlLEx/tGc3tocWl
iB3swwZ1gTRssGcsKPi+hzXG/hXAo4JTdSDb9Mmjt3NhwKj5eqMpp4gETsAuTklBSL1nSBd+z5HO
sMNxpDmn8OavQVeHsiENEnnU85JUPGfrCwIb7q711oh59g5TsoDEwGeHeV6dlxWB4Wg8uvb1ZyML
pawEj+1N8lKSOq6cuI7iIr35Rtyw8QD1XtqbSwoec9EAWH9CDf9vaxXLnhy6z4vs0qOQsoBCFU4i
ZGEMUX8SKoy1M/9MiCuNaJZkvdPEMogIcNDjorgdFGzsYjQ5MFl4skdTL1qoaziLTPCQ13LOqx4n
VW4wzH2wAXFwfbkgTY08+ZuP/9HVQ+sn2oINsDdXukmFGZUSaUZNqVrNr+lh4dH2oS+G4fiTYQgm
a3dFdHxdoRAX0vi4ReDiDB0CfQUQcZ75ySBUcaYyUrBSr+GYKMaCHK21rTZIXNQBw2L2hQ43CgDK
OWbRJYsTI7NQKOho13ttddFCWPcyKgCq+LOf3Bn2ZrhsmpNanXpAop12DDmtG2uu239Glxi+vQtQ
Hk+xbNXz4IcEVSSRKU7y0clMXZ8glCdNfSJUwKrlUpW8SbX/CWel4eW4cVFLwMvUV5DmzviBVdsg
/nODHMhIEWQoX1mYG6LVCIVXTO+PJ8bkruCwsUaxFcHenCqbxjIX7kpN0wTOpRsqj8VMct1CG2Un
j2AsE9i6nTIKXfuTrztkNABJc0a0wq/uplLqH1lcnMLHStmRLHjp1jBJwGcpqkp7wNZ+fxa1aaz1
JPTBzKePoZgg6mHGcRZpl3UllEb7eFQ25ekphGAQAuEgIZ617lhP/31QRWZv+3foOs56CIov3FBj
d7btLf/cffr2ANe8ipw3MpjrPRS3tPh2Wbp90KN5pXaZ2HE6dxDmDJbOl2zIa7HblqIUbNEY23do
6UNY0GvsydCYRGFYDB40OepRkCe5oHk6kCwrBrFJZo6SZerKOD30yIxBpbF3tkYi0n5mzEXEEzFG
BlIdiX4naU/W0Bjf/S16lhmxg4PMo/hFPGQVjzO09fnNTX5PeE8OElAxUgGi+eR2N4f1kipaz/uW
V6++dTTber7wO7zh+vhgmB5l5YP6W/QUHcfgQ5o/gzc3mGvDPMhiNq/Sh6mZck+C4kyemEeDFMy9
6z0raR7bEL21BuiCeXuRLhg0faWYGhRWVwQuss08EiRf09i0nXE6BCpDdptw1dakJ90hLRSgFYxU
GjLIgsu3nLKq7QTbE9WMb+wv5mm2EUaPWNKA1m4IgLXcEh4OeIt5MTxbDyLIMMlka6QTl1W0oOpR
ofEXiAtBv2KTr5D1y39VyuwuzAHnD1HPwkTHhNPAZiPfq4hUwIdcBaLBpmucDaEpDRkN4qkrE01v
kMA7QX/ZIltrvTrTs3KPWSZ8S5nu3xQt45zfKRaNJHcZbye8hkRhqkw9U6SQExo03VDjseKa9rVJ
wPZZYtlAHFSLzjSLWpUprmwiu6GJrH1CywkuwvtT8u+jwofwRWwBdthAWiEkMtUTvo08EtJp/OGO
q0wByXp4bTtED4tWLJc4gqBklvC55HMkNZmP3GELnf79Qw9WdFSkGJe/+he4Gy9HSbBr/5c3Tblp
B7L//I+pQStfNtGqesbhCGh4gxYQu9PAbY7/hY3Yk4jkYprPrdT/53Ve/Xb0EbIdNY3yLnuPkwjI
OufPqplVPSdzNgpfmF7Rx3xJ6JGkrTQ5+RhT25FQ5YBxe2uvDAs9P1E0jpgxwsh958KQJ4RWlmKU
+rmoQHguoYTCycnhhL/Ohtt//C3l4TfO6nA1g9aUB2csvViwTbyWU8hJsul0QUUDKcXRVybum5vG
8TrBZZxI//c9KzXJZLKZ6X6do3VdkJifJiVPdNktqTlAw+gLJJ8zb/c1ObHH3KbngwClxCb+6j6T
1A4mXNyD953ckT3nhBuynT+FGxDKfZiMxwollmpFYNqoTA68U1Ixp5huIhStwfWNxQ2FeSShq+rC
dzmMppstJQrKbFvXP98Yw0Wy4+7jR6FnvuyaXpY1Wy+sU0PLAlj4z1gP2jsRI0u6jkhYchsPE/aV
wF/TNbdmp1gmESRvRoEj4VUSZ++yN29TtjcXJnGMe+WOx7zZNlXq4Ek8kls3EMUlCO3TCfdT5z7P
iQ/A8NQnq2cRgm6S7ywMfyS0KVR5rHpVDGGZBI0hSVKpLEYxUxAUdlgP6ZLkhoPEN7+0hh03zdbF
lCAWiZ41KaTLTLvk8kw5ahB+7DbOI9gljP5b7G8UiQnsyW5u84gedbBYgjcpSY+UV0wWzaqWyrr3
Uaog78zwFY5h/fyJnWeU6JCiAn2hqlwVVQfB8bZGYDS0gWiPOXAyv9Pdsv9ptyeK4NuEDHsTdZ33
hg80EkL7RyDnI+qxmJnL94x6nWYfv7cK/oLXTenz8JqDAKJG21ZcPCSohR0+cY68F3f4IhM78p9x
oQpFMQlenH0gU55S9pxadbAbzKz0O4Br0F/faABV8+PhwbRE5Oozqre3V4JX6uSO/IQHU8hKqwig
oJZMgB3f99PIoZAroSGu2O1Cn8sQp6cmBEeFfqke9JDxEK91x3h9C3j/hu+alaMEDV0awHKKMqUG
ZHfn5g6jtJ9i4u9nwS0I58fpbOnhB/Ds+cLWprCGphq6BUMYU1HHDd3he89dNPJii2UF/6XAeGig
TQcl0tNIGe1Iqk8IepgmV/ynOHbbyfeumk/DmcOSHjyXdvPbO5lspoXS1R0Kkq9mOTGqp9O2XYP3
v6PqLXl3bZnPHzmyYKOytsyWqHIWHZ+XBcm8DWvGalfd02E0K0V+EFzvt3KFpgviOuqUjSdrxmDK
3n/4Ewt0OV3uqUgpHzei7vWBIeni4LtP1duajxxmbKmIxVA3upBk4Zpf908dCF37ZB4xRJ1jVSfB
yRIzIEIgjJSP0JcWYh/o7dojFys/nWywngPozTE7PvxEjodE9CApDrhtwoHql3Zdezm00+bjfBUv
5c46xWcew77Pwcc0ptmJraKQqYddZr7MwrygAf7jXo3bF8Bo0jrm8gEYkNg2R6EQslDNmEHK9uGs
3efV0pDb1QYQn5FIXQMWuWAkS5h22DD/+J07hN+yhawqnyM2ZaaqeiHUMz9jUeNeJqP1hx6itfwJ
RWtTfKMvGCCQgNFmbo7e2ogvZ7fjzZvI9hnd3S8oJp4IFZ/d2uZizMPBNbv4w0c8L2AQ3m3A8Bft
ewQ6pbJdThzaDoMxPJ5+zJpqyyzZPR/WmfQXd9wtUOPnXcxtLuiJ8bxwznfYyw5lAycDnzLzyRbj
kCesgZ1rrO5hbSBXBtzwnR/2TOXzNhu6iff3BufpJuYG77reKI0KY2XMXV3hbum+w/2M6aZeWgCS
DMKFQbWWCDTDFR80Kwxqka7U2oPzBj5Mw120UGzYY8fusmlp9Fb3sGFK/aWOGbwoh1N/GbFiCD0e
0Fj/ms+Ic6/BEq+k+ljo5HSnJ7RW7LYGwgoU6IWX4vhgqvTnb59jXAVu/YsUqCnYurfOE5G3pR8C
vsRYw659qL6wleHhuqQQH9UqOTt9/slhLRQ0L+/PnKS3RNfjahdmeGARaYR65ujmg/X8ORfS+gP6
wvOlIbR12fHY1tujGHgUHo01/Pdyt6tEMVhr4n+LeMqjOtYj9LG6pAtvcmMJzDLJ5TtSJyELKcjm
tqEoKHpPMTSbLL00U7jj2tPOXI3XkWjJXmLhLrfozXAbLBbvoHZkQmot+o6a6ipkSUYF9zCvQMXQ
q2IVc8CACVlyFTi/i2YixUjwGO8iZMzb6buKn8cmLxlQ79VQBxAVDsioMsJ85kETMiIkCOqSYSTC
+2jOFVcaZdqHizaROIa9o6H+euzUSXPTq+85Z+D1xZyQzw6OStyBKaxLgJHhdUgtfvS0DFcIHVkx
+QappQZl38t/1uiFkpZjhsemrg7mBN7CGT3SKwJdx6mjxZsl91tIzDxAcWa1TdmudqdTru2fqVUI
BKlZ4UVl1NSeY/UZbUsdpy3Yvsu/5Tb1LjdCbg0XFuDhsgfy4VDpnn64mMCRMHdnD11TB7TOpLZS
2jLc6Xuf1wL58kOfKqbA4CTtaGhfI0nEu/V4y+7HZLxvz6THxf/m86v1cUBgMN7WTNC52k5CkbXN
g2Oomo7fwl69JMXTOT9bvOu6e20PRRB7ziAoZT9YKxo0IOHHB5/i1zblvc6a92u5HzwvIjaDtCnW
TcSr+jADHbNaOnMc6L4ckPbIX+/nwq08RGa4wxE/bKsFC1ewEk99hYA3ooKt/YOc5fQPrO+xnsS9
MPvY1Fl4oD4S43l+Sv/UL0naxGNbKkGEdkfRN6ZM03/yYEwiCbDSc9B+fXXxHHQjAkn0jMaeT8vI
J5JJWT/BMxmOYQvPjX8+8JYYIP9EyqW/vNjO//ThhYWpaJQ3fBqWugsR69CM/3S7da75ZnUE6XnW
q0I+ID1F7atOHu+mIbIe7leG9+O9QlsOWvN+W7GQpICSjM51s20ovIofaRMc5k6N4NFKDIAPVWYb
FlVZUqRNtWLkmOfU5Lu7fLvcaL66Ol9y+NBj+BaZEfTBo8+rS618dCj7fDPVw4DLF7RT6/eDK6Y2
ueDA3WuO+lqSTN2XYjqhnNSERUcu6ngSOdPUDipqdCLXC8ga17ULYHAxh7UYwBLOx7qYWRyCaHsu
GgwDkcECqU8dFBbSN8jn0bvObf35ZGP8VictISzI2oJvEC/rSKtqcpTq1iG3Y17VKjjIsBvmbbhI
8wBh4+XgDYEusiYqqxrpj3zilqEOTAiV0q2vzl5EpUcZiAVbOKQi/BjD+fCK1XqD2JHb7OEs+Iyr
58Ra6hxncYhLZ/6HKdtdHC3bOgstWhvaFhlCOZP44vaUW0QGUpWvB2FeYujXV/kYjnMfJbXJcUgR
Fv2entxFZrvoYukN8Ng/ejIeCtdOndyhbIToL/IoF8znlkAq6IsZZMYkuIAEY9NHYjiK3lV87cYB
ESCnJzci2Uyxjag/0KGRBboKbtqHAYM3zXGLPg6pDgM7FPns7ksjxYoG7wIi6IFS8lT/x7hR56rT
hWTzVi6zln1jw6S1b/J0xDX/QCMgqP8bPw6IKYy40kL2b86xTrM4BcTQtPYqZOAHd/mgaViLH1Y/
h2GJz6/1DOSiA9tD2BBS5ferugRQG5u6iLglgV/rqTgMP6KMQZMsUandH48KPlQ+3u2tHIw6Jwtk
FErRx45Okvpxok/TIGLGkXN+FBM/pFK1LSn4cYqDisc4cFy2dJbHlpyWkmkhFoDM9PoPnnc+sAmR
839DoTDBzeFTTvVPSPcSAcdcEFvLvmnjAQH8ticdSnHqzde/FmzTD81REeozXx1LZkrkO8yivzKB
V5lH76lgI77D1ZHTkmi32NQhiYYTphxKo8YFTaUFeYUc0zDxlp/3kX0xX8sEfrSstas0J/OJe9KU
SkPdI5LlBKfhEcQgGSdfEHUZskS/JZ7QzQ3GvJLmysn28hDDx5/Ja0iPint/x/dYzDiyAuKURTuN
9OSXgPP6rT0jszqrTbgzD7vvysje+Ar8mPqcE4cXqh2ueESnY9xRmO2lTozVze06JVsrM4YujV51
kA2IQ6qeQr/QXE+fs8FZtNzmFaj882CgTgYPIpdwgl87owmbm9dbIURY6bi+tp6DDGtYcii9JAZf
qGnAKomJpJ0kau+c7EPwn0h6CMT6AociTIKt1Y5eJ/FDMb8ykuI38OB9wUlziePBNuYwg5GdyFai
dyqlv0WR35YfWr/wu5OgKDSbuOoSQa5hU9t/MPYXiDXGmL3Lr9gf1kY63RnK5Ym0SSwqP8YK6Yor
gNdZ494BpQqqHU75u1rqWd68S6htU/vU/H+T//Hi4pVrEouUfPtRI2GtkMWdDVT5bpt9ju2zsF5I
92zJs5BP3Snl88hLRD6UEkuNA7bPLzikzn805jWiweG6fDXFisUj34gWqczvN/RtFjOo6ShuiQwe
tylP6RSf78Z5R2ggPFVmLamukfMPdxrUdTgjeuagZPcHJihKMZdpXplF7lxHWI7V5Z5r9xhzDFUb
mh4MMcbQfCt9qy9i32FDN6UUyp3WwTqMzBEn2SPd3eefzkxTaobpbU93ZgXaGGammHA+R0cnTIMK
xgCKcxQZhsAqlYZU1r5PNhpWhy6BuFr9AURLjKJQBP2DzbgkUIo9VOpmeZLJkEnyGGsK0F41rXtM
VOqk58XwEoAxv+Z6Gq+secopifweCgaFvcEiSfQQwPv0RrAXoSckv46RfUF4gBsageYd0MftrJbJ
7/lgCVoVLcUPH4r+SqIMHCtXed+z1UHkjGmlp6l/8riij3nBj/v/3hLTwBnajueFbvCA7hegq+JF
2cPHqQNCzXiLni3oH+lPYFqMy6+OmSjS9iM6WnPu78R8sAw4vpRj3KarUT+rjgea3Syv/u8Cfkq8
SPcL6fMZ3mtKwTj2aj2NLy1ZNLORyzLMD8RIHGmFTvTjaRUxKh8i31CrAot1fiGPn9pZyK8nTpZ2
eGquw8+BUIJeGCdhYlmP4oVYso6zXMMTc4/Qmsyk9oRkn3xpjVG5QGGNjjFAglmzPc3xoGIp9wCz
R9kc8xgx3lt6j3PxqcntFEVGDaIFFd8Zm3bdl9vkKqVuCsfR50cH7taiLuVf+gdnjSN/gQKdL2nQ
mO+RDOP8t1O6NzELSCLM4SRPCeySYB9cCXXYHi4ykjf1ej2LdlhEB1W1mRGzhedKGYGUKMtVZSb1
Ct6tIhLN/wLUHvHGGkcv0npRzocmhVwjfm7iPYmQKIZvSE8w++5aL3gUX0OMq36yCj9dLhVIZbx7
Xjwgv6HsEcMadeoPkDc7A+axu0D7NUrP5hrQMn3xI6LM9uxk9JDoUjLxK4Cbq0WmAg6KBk40p71W
6PBToZuz7CZc544fRFjZMQdOtvZMteizlalIFUkmkYE9jyNxW9SkHWNSwTsfIaDYU9E2bsMOkjFk
jtj0Tmc+2eg5nuUABIE30mMMoTXYJi2f7+OmS8aWyVczzVSMMUZsjBeNhIW30R0x3PO7f/CjspBa
GOUFdhYDtaYUdhJAimmvVZO8DAVApz/He7YGWpK4bvvHapF4IpjTsxrxUdNqrSB+bKPDkPGWySg0
CuUKqFUxeKAVQyzriKM/4mBYvvLhAc4Q7zPDQWrIaW5TwKNIEr/QSF2+uaClnmyusjw1BOiDqUbZ
aSyTrqHYnvQ4JkDgo0AQ1wEf96Cq+fiszyVcrBXBCnN3tew6QOq1ioFAFDYkIGK1U73j0JRuOJfC
mTZdgBvuFHAuQsxo/1mUH0igqT4h63uowBlYauW+uIz84RoRCEvW4gQwQsZxWD6U+m+v510/ghjP
ar6eVUnXA2N33vRiGOgf693xGpn2qdT9iaC73GyP3q4S9t+aWIowaOfoNPidmwfnbbsOwLv8RzOT
3YO98E2mFqvURi/yALOQ73lfDns89ES98cTLeVeEheTQoTUIPjF3ufmULKicwCpqdX7IsewgBeGg
7mvLd3Ri4O2pyIBjKnCxRNKzBDldYoyhtTHA/NKHpr8+AGxEgwormmLgq4WVr/RueEYfLe6qnX8S
LpoTvQZe22BbTOxC1ztusATQpnn7oPnqKjLF13pAy9aKf5iGXmFIwwWXzx2Q4m9J36nB780FF8zd
vaFqoMqlGQkimMDJaexsv05lBg7P0pNkQ+fNra94mysOG0c0d5E3saj5YK82GRThe9ldhMHgbygz
M+gUZbgBNXZYxXX9m22UK1LeWy6Ok8LnDmGzfbL+w3d0MRxJGxBA1dGgh8epP0w4NiTD1IdhDhAM
W9FG5lC/B9eqaS8uDC1Cqcqaa/uiyYE6adzNBZWz62RWBx4xxlS5LsHCjNT46GFDlr2+FtK+zVyT
ENLHL7ls1SsBJdRMf67wQetNQlJm760bYpxSagkKuEq0+xCg2gHpyMHMpds9N7QX43GiN88fQQcU
r66aOOKIjjkelYAtbhlUOICIPiR3NaFVu/ABj0zMNsCFCuN4WVB3OLxCkQCwmlP4nNdA2DGB8PJ6
TIzrmYrcX0WtY7PVdVDfd8mYx6EIbCquWJFkLx50kRxpN9qVxQ2v6grsOUsAJ2XMYtTPdbMVFdt3
tUxT0xUvcHM25sWASVc1NJWycO8GWIqnSYOQyrAQB7zyvKMCdgLoc5iZIg8yaqf1H3hyAYDWEeN6
s/NS9jmD00rUW/o1ISlh8Jp428Qsy90QIREHiJXbaErwIDmvcKB9vDlYNOzN5m0aqKdPAofEmUQj
CV5AhlJJwJxOA++eZOA1UYaWGNTO9LRXuSGVa49d3LLEaERR2cyjXsu3pDzlSuPrrVGmQHy04O1K
zUGkdtt5F8leZjx/C+wDM+hQFTScb98Bze6X55Yy2H0/WKl0q5Cc/ClAns5o5UAVJMa5gptFYMoT
JM2rM7azxmbxX5/q0KCr3q6GEvtqThJPO+2pg7C9SScx/pdIklZV72vikwM8GD6A+xhg9vT4UoCs
/x5flYgfMnEC1Z81l9axj+DzhHa+7OWxxVxHwsG8lZQwbe8+Bqa6CCMccfGVfiaBx/YDCzLxWq6R
GZGzN4dq1XiXfqsxEyI5Egll30kLeDENooQ8qUKuzpZR3VJCmAS/H0JUC2lMyIYDhQEyRBFUGM+c
mv+6r4IMGl0f1eYqBdBgzyWNeeyTa9o1VFCc+IEnP4vPdJO+LuQn4zrZqKMjI+9eDGPee8ayvkhO
HM6kzWjaDM4cpSz+W3emZLLWmqZrbeKTjIBWFhWqgV0XLlKtjoXLPE5ZUPOTuR8egOIRo3HgqlME
rALaxaw4dYwHXiKzeWTJuzCSHpHG/Ucuq6Vw6yov8OYCZk8JeZuaAdL0LrRRPz2lPxu2TkssKXH7
AgJ5sxnjA96aGbdFHWbEIsrhV+cfRFzX+b/3DJHS3FcY/v8kgLPVn0TZYBqzlUL9qkxTZUpBHJdE
Gj7xhYlmA++P2tfaPgHNPJZMl/+HilmMLqzef8cE7uZWOClKmLAMu/Yu7b4Ix5oe1SqK2+jOdVtC
QIgW/kimErvsLzSIvn3X9QnBpZEgw1BOiZFaku+/irXVV2d7EFXXA/xLbvbmPNxdl5S1AdKecbci
svS2jYI+/DzO3WUQBeSwyalSGi5PTn+SCmdaAs5G6FSatMFFftu1Gqg7iRFFxtl5UnrqxXmycYRO
A5Y+PxYJMYLA2X0wOJY1436xpLUU79vt2fQ5Z9gmZUAjZFgnciA0cK8X2AdX1Xg9G336N/DdSG6V
Nbwe7Oj4LtmlkVHOklRh/wsBqZ72Ux0QLLxngRzy5+mVRkzLmldhawU3lgm5W/wnd07OGRgp1LlR
fwk6MiXPZ0LpXZhoj/syMktxCHxlPFmbYBof5fQZOGjXKnp0AJF6eTm1crpVLbns/LYq+5djHHQg
LOc4onQA3kYiNbh3Q+V1qWftogKxzvJxkuXk/Q/EAta66tO8v7T2/l9RvNWKLYTo1WJzLePK0lAI
vRWya8Vi8Sg3oR3QtNFxY4VN100GFpGAedNIanu9Xc34Ly98B+aVz+AFLsIFEFYtz/BFbUni2rbG
GeV8f4gT6xfEA4gA6uNG61pB7h1C1RV6KSMJENd4iKoRJ8uc26Lupi+DWsZaSUFzKz2vA4ZGb/ga
1wqqjktta5SlK2/ziE9zJ4LvQ9k0VWn+uoeYMLoeNR1lGZbbYugx0H6IA8c1lzvEhQmsLni7sMvZ
taAtEpwxhKbBvERw5LSQiaEbK5+0S9t/8EpNfVk1g7vHBEDJdpkxjy/116gOnUU3KNVyQnXPisib
osP8xSWwl3vuFYZR1EapEiC25MgIQhQUgG0zgmGElii9r/Z277FfUKV/ECZQr20U8if7ENv/0FXp
70vGV/7trIjlLBi2nwrzvWTJjiO/PpPur5g9dzshOE9vWKWNfwtge5bWi0kY4WNgmZhdxX+NrMrn
rX6hH/wptOWfr26pSz8GGLmc+EI3gmlI3mZHZ2hTm4JuTfPvzEq91OH5a6UnM/0OAADwsW55WfuI
pk49Xjnn1cxivNlwMuAlf7wOhELv2ctcak5A3RVWqmBAHjp56Svs+Knz+q4BqWtb8xY0wHUCz7GW
91dBh7Osq9vd/odXyqXPbpC3GOKrqlM4kjfM7Tl78bVU9+1DSnanrUWiuZxD2/NHhRV+o7PnseYR
pUTRAuuBdogRHOaCN7AnfdfEu48c7qWGdUcLgZRi48w+GGpUesjeSXERpxsbZZQGBOcS2aPxMyOL
/t0GaW9uSwYitQkzZxFaF60g9zYe0drcI7wRW9DvJe0mg7kLrbGFphuvQ0UjPczot/XFstPmqtSf
ysQZZhKg5hf56WGej2+8ZF1Zs/vgSGaX6fABYmVwlQPbDWx7pMVdu4zHjn5MRK7evdHLOpTMEuxJ
0Uf4KcXkkYZ2DPHEP0Esv6n2ZJup+vd7Rhz8nmS9s6gffYrNJVYr6DUQ/Kba3otlq1fJqmcGKzt1
oVE0U4f/ElD7bOwS0GyZ83WUjuBjpaYIVSrh3iGObnT9xpHzwbnhobOPWPVbmPWwHtfpGDWmY1n+
doLbtCjH+7u3dtxzd/s4YbpQIJXCogoU/wq6NUU/zADwIf2tflqpUMh+VA/yl1w3I4ti2jNN7Art
C/RbN2kGcJD+XDoeksP6lE73j6oZPJ4GcnTEUCHVSr/KciDXRjoRRlaKkZcAXmTpFQwAPR73iOyb
mripvbKRSmC+wo7rIEnvIJK89dQANv1cFjw8IWm3fbxXNcd2ePs+nlD9eJbapDDloQBd7gdJwZ6G
aqRhn7tjfPRWLohe67ckQ2n7z9EPaNRVh1HIp2Y2JaNhbOdkNT+jHvSXb5AKJE9DuLz2T+P4jbH4
fgCPIufBs+Ngztp6x4ZA2pvC13n6yjGw8PLQERWeOQrHTKyKtSPhnT7pBfXFgeQ+aGH0Bj7NdXKj
e+9051rGdwD52WJSqokn9hrkw5tOS6rRBXRgbdzGMRPPNI2RiVEpR6gQTpkLiCp+ENXN0yZgo/Y3
yizv6XGgGzvGQjh4JDMsBODRfB+hp4k8EX+Hif+c6jAt/AU4I5Gbir/Z+fmyWoQSLixtC2JVQaZL
ABh0DNyvIG4QZwYpoUM+VsGQSbr9LLaWf+un2RVsckVXUhGj/qYEvAf4QHMXSgZddfpS7CQ7uQmj
KO8mH1HiDLEK3t/rp29TC98G23QKl0FJzbWjwGt/jqyHy3gBfMwTEAM47ukc6A23iMMgyBObKyyh
Ue2Qf1AQSdCToQOdizE/ZUf1+h3t4/JT0xbP4Keo3KQZtQytRaSAbutQPpTJLZ6FwUO/qxk+2bw1
/p6/hu/4vdEGzxFP+oQiLzYjr/TjmRB+H7ZDwlCjReUhOe0mpy8R19842ZNmH/TyymVxD2iF1SBP
xBmFoDcG6zVhgy5psfH7T1EgEUV/Tm7+CRXwcCNVbvDCVcB3tL9xqajXGWEuwHox43AWEK5oyvCk
IYkWFQbbiIJwdZle0cq5AGKrcZy7ZXntOnk4dzB5ENfr/YmvOHZR7QsEvjTEzSF+Y0HbNU3jeNSG
qYKb17KVp1APzCGkRW366qyjecLQkJMveKKJLiwi56zZ1EE9A0HRI4T4NmQu/Ygk4grduP6kG4Jg
2EyMplnUnF8ZAD0yyciOdHdJC5nErCbWa0n/Ay6MvuHrAutwaaLUyop69ENUctqLj6cOSZryLiHi
n2q6dXu5IUooNhhMCDCsb1RxL/4GDhGU6jhLToPn6q/XxfO2nVRgRl2sE0H+HyA71xYWZuxU15xf
XaN1SaDUuTcvGarUEjZz64zk8ayPO/IGjZ+jJylpqWo7R26hn/+1aglhKNtfBURCUX0hXPZSVFi2
9ASf90Tg+08CNn+PnzCeN0owgXruqDAiirZ3vYaMo3zDzSe2uAyI9wThTbYGKwV5Ytv99YWqsHKJ
JJ5Y2JnS/oYsGIn+sGYBODSK5xVAj0XPRU8ML3QBzqB5wURhFFkMOfFaOTOMrqtzZ9W4n94e7bJ1
NQLld/2XiBTrgzcsyFKTC6vf9hWbxbBn+yDjlM0vfQ3Ks1F94Iu7BvlpsmXcNWXNyyerMy7EJre7
Um7gBny1cgyzY7aXU/x+1YzCJ958oBMc8aLHhHHnmdBot2PlmbOWsTCPq+H6AbfFM1wDlbDu4th6
fO4csoS5jPBivxCwBqOstW2J9xaffwKd9cCi8SijmuN+7+ovMKnkarriEW+XcTM3C3TuxA3T7wrr
lZISmLpOr9oqoWj+NkW7d1DDaUANwUA5jpZ3pQ2tn2y58FXmw9U0zLrJPnz70nJoRmxbB1Ock9Zh
MF+ZFMGLNaOmp/16Zfw2DacdKUBHZs3Z1c0XAPJjLm9kFZUNmXSF1vCKRPdeqTaxivGTYDDWNdcJ
UOX+Lc/uTGxNl+nDHakEBNzPys40a+mA0cVq5rnMm1ichihtU4Dd7LkVgXvUIda24hU8iRReIcdE
gSnVdeC9soj8PeEcivXeVMjpvdvEUFequE1z0wPuDOWn59asWxJmbEBqCKkVDqd0P4Sy20MAqRL6
AAa/IXovl2qDr+dJYg9SHg0MamHJsB22e9WuthzGYlZw2GTbskMO1uHdRf/HivpVFjS1ImOMeO0T
ZOaB91GkwaOxjVmBa0KhEXjOUQ11KT63/AlzimL6nllQCT8rm5WB/jZdc9H9drjDarQAxKGofYBY
s6eGqEsKa5sGRkYm0xCpl5i43hdHIcUv/Ex0eZook5lsUSXXkFVEcPZXjmLKD5cXoLGz0a6yDjTy
+If/I/4YTjuiOHvBWqJqJkWtDGrOqtipc+7amZVmUU4QStukxVniorusFKEQSBlChhrOOK7D+MIu
80HzJDK/7wrjyP0Ea2WjrLaJ24gBUPLS5K+oijG0lyF+2a8eDkmMZ38PvIgSIX5nrBkhUKGtdrT4
3isDKS7aN4FJmGwp50dNA00q7OgmsdSooEcfbxXPnHdTLQkziCLruFMyn3p7DazwO0rmUqk8rIw0
qIxSOLiXSPtMMEDaSUhJTZPy2X8VW0HFZOFrgLz1rCCqD7j5pY2mFEmDbEOR5uMDyfdEm+NPOoMy
SQyLvf0UjM7JpmX49GK/R62dWZLvFZ2a07Blc4ajgjq+1xMIdRC2T6b7yXU9JToq4BDH8kPHp9Wm
SWeD1WRPQIKueeTMGsg2FWOsaOCSqdLbLdn/qISeTaAwvTEMXBM71NvNyFpz1/hvY8iQtaBRYf1y
qX9KpPrpGw2IdeAYqPsFA6hSmk5CZWcnfd7IJSqNsoyAllEhG4LHMl8wD/rIEIV7GyZSejGo09lo
NPQAE/VhJUKITRsUlK6AWm3sXU0O9PSjbgynCBJLfiHzK8g6Z3e273hNSyW2DohL5FSoBczKUJ5L
Q67yUDImIPnGKZ8IWMQs6jHOemMU/Nf6ha/18XCkili1+bhYbjdNpcWAy/1U8FylZKthGhKkcT44
yOa7hm+viW1gzI5q/zzpOa1vP+tweW3eMlAx0pmOT4ZDTC0IwAba0Zn5j1+Be8cRLH9Iye58NUMb
MxWYjcNQV+glG3OKU2tesPTOW4WYTsvpiCRXry1ofcTPdE9/idH0PYdtEUGrpHSsOMnkmrw/0PCn
6idlYaEQ/wmr+yGWz/HjpXWbrvcPggpdKkypVTo82dX2ChjoX8iqblSXvO2yrV8pPGkA92BGxwka
Mi7vWnumB5TMjR5Nqn5h5vgY4ObO3jqTrp84E6O19OsPFCtmOe0nJnSUO4vIXIe2Wo9JC0GCfYiF
gC1tjodGePLRsdneBrOxX6BEZmP9/ZGqguHcER7Rm86DAyO6X9RCddccGq46iITt6ExbQxXQrhzp
3fyt2CBs61g17BpuBgHJZZYOcBChnZ5XoxCMxUmQe6YMMN/iZnyY6aUAA035vC8qlnl7N21iAFWu
TTIY6W0+WwKgfbPq7PR6VlVJ3/bHAYjZJ1Z6frf5g2QNZ1RluPKDGUrdYifV2IDGbX07bT3/MFHc
MqsxeMpVN8/NpGVlavZpE4NRHmSr0YA6KfMejao/Bak7dvAtvQD0frwhSKzQaJ6JlpKQFctXzp2m
xQDvnfjjh8hGou09xaVmmKw/p9nbJmQ0K1iV5JJRk2j94DFuPEAZu+7dyzmJDCkKPp8TIKZPZvDZ
UQ7DNExGPKVTseCIochRO+Vc3E7Uho7nIC42ObzC5S12GYzANN+llnfVYqLTs4X+F+rZ95WQJDG/
OuH+34X6Kgiw6Sp/49I7+zdw+ENLbKW27DnqrL6pA6YJlTfp4Ru0BEfLTetLKnnqx5PAkXGvKQAS
idjWLrsdqnB+wy3iPsEYyWTbmPubwrweC9iC1tdP6X7Q7v3BBqLGr2azZcHU2NnsTyKCw2i6OqXc
pHQ2XRPJRCnmmMS2O8Wq2Gyr9kB+lUNGiqwE8zFD1X27iTq2WJG24P3bdci1GoO6SBC19jRkiBxc
MjZzdlaEvjoKU2x54ARMO/VcPlkg1UZDpDzSZ3NIuEIp7Ik0O82KO/a02PDGHEQZFDwvMqmHhFdf
J8QlBvzF/8hwf2eWu5p9rjr1jWF5w0/LQy+LuwGpL+ghznFZ0bXN7nG34e9Tez04FIqPY+pDajIw
qXEI3RVxEXlcrh53RWEzQ/9uzw8U9u8EWipy4CofJ2YQdg3U++UHuA3wvX6LuEbcvUBCghFi0EN5
3iMbFKfR6is2I5/Bq/stj8Ns9QVu1xhD2aNIqwFEeMr9VjHvhX7czMzuwncUxWQ3x1c+OvfH2G0a
nnLPu9EVzV4nReH9kfE2KzZaj8GR6J9hhWYW5w+5EtcZGNpLi3Wjv3sigVKXtDzUfROaMl3XyLY1
TQrZZj1x9NwGd9TBjBoEa9hlNg5pjqVx63/oKHgWqRmaJqu9bhA/55km5IjEWQot3z4Ml8QnhhJD
wwcIdt4ih3aKk5LyNhsQbrh9j5pT9YOfAILhkGS4JnctIici05T7DTw3eEHdxa1TyFs2cHXxo8Fv
m0zRzPe7s4ucDgju126ln+l1U2/ZdXCsX1ciq5WH2mnUtfH7Thz4YYpXpr/S3ObKVoJHyUhx+PKO
tf1T7M5u0j3RTh1oj5aYlbLdZMBbS4XgN2M6yy5yMzTRQLwfNeDH8BOssiqJtwFJXKBHDBnC5Deu
OTL41G7pLOIbBy6GRObxn0c/kHMDtfqI1aaJ5fgKmD5CZ63mY3R6lvTVjOrD6ixdvR0jfn9e3Qfw
xdSDhBh2n15M4LmJXldE6CK0FKX8Fn8+yXYDdgJVq7n2Yk9tt8LhEpX01ERwyhqU2DDFcJh3sEU9
6lQ/sGQ3W0gfPzuCbWBniXUVrL8UkoGzRcsEzKn8dp6rNt+UuBWlRT2yCgopCw784Eair8bVgH/S
UDKImWX9DJ50qlSvprZQZ3TDqOrCW507U0AC95kOndrWgv3o+NYRAq4i4CTKky75NuuoxG1lCxN1
JWxe2Gh8Halcz583yg3Nkxzz7xTM1lSrTuhVNPp4BzLnydzUKjCTojmlyxAoXkcbu3rlvLFZ0cVo
3HCgUS52hZ+E3CIGflcOS+836FOdPyQYph53Tn8iIRAsHVXmM8uVd3wo4jnK/dawW664NID/AybJ
xvXxwG3gXU8c9ga/LpNQCTTcakVdTVvdEJSSWthqukQNNIW6737VRcnQVWPsse4ivcPrNg3T9lQr
98JuzOCTK/VaGvO9xvl7mwVwtF1hRVbIZtHXcjofJDVQC0CgrWl3f/MjfFC3wTOkIme9tXkeXzYE
4ZCYnM+6AVCJX0u3wjdN23fkHjaIZlfgeJrghewWkb/WvFnJc/a3JqEwknevBH8sfxkGKLw3M0Mq
XItgGVKZc0xLI+HnTogEk8cN/1weDCXWMBNjLtwLLeaJkaxof5Nxxfyl+LnBtEflXHqvNmqp2IiS
XnSyY03sUAhIeo2hJ+7FdruC71ru8/3mVapimVsUXXoPnGl0NQJTgvGVw3dl2WjMd/2muxIB1pb1
qCqp9UUwq/IWzCG3LT852xfa3FPHTno112vXP+Pn7js83A6R6JAJvoHEuOYUdtkfi0gvt+bwDuzn
7bpEPbVtnLOZ/bgm8RYSHU7H7KhhwPKo7xpc/9Qrwfge9SsB1lqrA8ZigvM0BfMmZ8k5+t/GRtDO
uhsW3TOEQSZbOd9eST6kwhZGt1Mcq1zMYnxA4p+OpHkrAg7tp/jRE8Ee4LoCC78uQ/+3WbHma9X4
oZjB3oFIQEZjUEF9xADNHzE7FQmuUm8TTCAAo5oRh61U0US9iJsqFrTAC0RM/rciTt1x1xA2QpAu
F9vd8OH/dDWSpMU/Ipy3V+DTNb3TFvmOwsfVwlcwqiywVy9Pv5o3+M7NjtQcGBSCJPkCK4UyT7Fv
UX3VYBsiy0x7WDzEAw6nOxZUKRZ15OYtqEGJeq0IvlOThrfu5KtdiOdPAmByEY+JodCM366Fh8EC
FKabYA/S0cIVq5JpydQDe9Loh/N4wBHWx1kM22FZOlJgGYe3wD2RKYRjlJFd0BEQ2A9CGD3FbK6T
pFp4CpPTK5vhcfFgcyXCmxciri4oanQdBGRAldg1NSGa/1T7Dd4Ce2rnzRwCUPUb2M3rbjPbBIGa
NLFCG1RnWhrgs8Uctd5PaUVsq71F60I5yXw8hgLC3K7HUOjp/PQujfknqD0xE2cEXNnlMCtS6l03
EPKGtM60l72mnwF4EsR4Jy08J5x9IbuWrshnU6svKHIUVNNkk53+jQBqHs5KmTwJD4mgQlI0MmIo
BGYqiFWk6PXAEeRJZfvvVTdNPsZZtpm0JqWOgq+2cTRsNnBaZ5FAbdLDVMP6Q9Z18BuIG1Dfir7v
sq7O1m5Y+QJraZyEWj1/tQaBO3hgGaoPTQ1XJstRkRwf+RJ+xlAG47aItTYFbii3D4xNQY4lEDil
aPAIkFDSj3ZupLHnTeFQxh6HdR1d6iy6n8+vyh3DCXhYkjqp0tzxS7BIQnw/9Q5ZiCPbaphCSXF9
BQUc4JPn9N0zBB2EztvG4EXTYg2NluzlSewDaHX++Sj6+/w2/0N84eEEAiZOFLU4K9KjDKFz4M/E
PcV1THRK7h4wV0JznWQKx9fbvL0XzQmnNU6GulTLG7kSGSnApVqjrTtwmdXfJIXmSSYbMsArKE14
EvRoRMHlVvehAhEeEJ4/+vzzz+eDRqZ4yDigGZoId/L94ZznBxVvcLi4tQkrKLyX2FQehAEioWB+
gSIdLKsC/5Wq2TQw8+Hm2I4LgPOIxMsdwozcWBYJ5LxgY/+mprKon5K9wPzpO+564PXLW31iwItU
I3D6HcewhheIapqBlc7VRjNErjKfvY3QOmeFyBklPp9GkzNRxAmO3Of80N9JGE7NB5AyVlbuje+r
VhaHKpIQgCP15RAghO7uzRCG2hfESKIf+ieNkeOMKYxdcOln4KFsP4nnh1kSxzv1B3IxjA1SWHT+
1/E8QERmQL5W/CjJ19GsZFcawV291mhNdkIhdYUDXeQAyou+i14LhrVekw0KdYzoPLKBZ41pY4jd
P+YSDV/aSWAdpeHMtBVYoxiMBMvtveEgoz3UkS+z1n0KU5GBrzkKgRR88PnWJb52G5ZvFFT7/BpC
DKGH7kXMa6zrHJ0k7aXqzlybE/PaZdkw8HvNqnEuQqANHe++51jijav8wbpPk/NSNh6hqKwTU2IG
IZeaxQ7KUEZ7+aKnooUTWZT10umHRKDDR2tiyxMkNckPdOpdqHb9Vz1DgiBGF92x6VFyik7YC07a
dIvCDe8/H8AayJgQrHOMV8sUlUU0NZ140aWYTejuNZl8+Hp3gAzU9/3VBAJgRHQ9oWIU4D2C5ZGJ
mQ75Rrg5gcp6WGo+GwWR2sE1QbY76k2nYsL7c+XHbpzjzb6xnbcmCsWiMAxD7Y1iDxpWO4Vdyz1M
r9oDdxfo9cJNo3Z0OzqlmS9zjyd0Mg64QuupcmS4WSkr8mDQ2Pg+oXpuS59pKBzB7hFKWHEvQLOx
OL7BbaS3W6hao3hB8PJ8hkct3P4xcHIb8ZGO0RIsiTHRSCSk0yfi8iILx9wqXuki5gftnAIVoxyG
M9GkuwUXfEkcHlHU7K+4NwyUw8ptdKZ8kE9/ALPHlFs2a2xrKulWlqoY9JUe3M9wSHRO/K4gJYlH
PeeYN/M9B1khRFZaPFxfylvwCX4qTN9AixcBhasiDjEaWbUB9RF2Uv3/Xy98Vxrp6wreQSbiPv5r
zlchSmeXqQ92b7nt/0i0+u9twOrSlCrRUC7e6RFyr8twleu7AMJffHGAyY3O5IhhNp8PokNiXkXr
aPSxVANnLIzDCpLfA6K9OekIQ4vfUY/WIcD93DXRo2/uPlBS2ZKN+4+mJQzXrUQLUXCpRRd5rQft
6R/Uidkp/CX0L5CtUSq+afqVIONG8s07oBHu7Wl55EY/FToI5rPrRlHjH4EN2sdTOnV3gMhfQTsy
tEYuOwkSNER83ot27SH/G+I8eXuLBoctjWWowxOlhxSbyypU/+r4B9t5mq+grGiaMvfNBQIICkCk
VcQXgEg+O8OXrsUGUbkTP/eIz6+GVt+KaJ2Ys5Orgfx5bGLsOMC2jz24UOriAf5R0/jJXK5217Rf
XZT7b1gZzCHb2PdBT5iusgV2B3teOI9Cyu2QBCIhHmJrUv/sZ83G6MnDcAmbrncEXdGr2Z0G76qw
IHmVlqdxuwYsQJsEzmb1xtBrwLEPCK0OI1CT5kFmFyBKQUUZBDq+dydimeajCAolMYMucMcDvGA1
btRO8Xc5+hr7LUyp1VFTwCM+UKPFoxx8xsGDjaPQdIC9J+N6zPbh3/HSeXevrldUXS7FXTP8yefS
LRXKIeXplLuNFLEydN6KEztsNPByacHt023pHjcGlC8yuvpNPSa9a+ttoowlVcmZGXdAWPYkaBT1
Ty8DOJQQx6qD7ZERN0gHK4+vcHFN+mXhgIqdMhCgRC2hh2Fk5ngRdH0NKkc7y/tzBEWeh0slKa7G
emjqVFgfsGXIs09IQJ1AFRLufzYYA4xoJyDOChP0R2FNvWtQM+D8Y+AIxiT2TH9xVFZofuvE3hxc
YZe1kCEZXwbqmYM9E+3jbRsoPc17gZ9vX7Qj5f3xj7QuRdlOYFJHZGaMr/3w9XwJnoq+wSwA0TGJ
iMI1P2PPgvTeW+5KF4yEAlFQGDwL2Ax1uN4merclaRt0NC8WeFAD71kCMBESHFEahl2mRQ1wdRCW
r0EefO8IyVX6+CfVjZQd5ROiCWOy35f0teKXp285M5f+XItKWuY1P5JESc3gtETmCy/vxJlmlahY
XspQ3fYJALO4h5SbM59T8Hd+rKQ/zAiQzObiGAbxhG93jdY1xJts96OAdoodxxOnqYzEdnPi1UaI
dfjEcwQflRAfGuO8FUvZFJ1JcK8I/wsp9vrYjz1YMgk3rrT6v8HFy4dE3Wpr0FJfHEESjf51kdBP
Z4u7p/tVkvSRTOA8imR2Cy42bwNLZ+H8F48lNtaJyVwKOWEaXrsP2yrQPfarYJT5OR/gkmW2iX/N
DKjxwdV0ZN5/AzPA+387/57PUemWqg7TdF0Iv2PfSEP9Chk7etK4N4/+ZLIpJRvKtghohNxYKB+x
UeNcJdvMi2+qfFQkyWUq4Jpz4hbl2r2QKQahM5SgriYMDhn91wPjnveNJE+SUBr0WZjgVP0gHaoY
SX7NDdBknOF2A2EPYMgGbELplFAyfu+yHyLMqvh7T5U3goPBKmZ5WnlLD2vTQsyeEEjQQ0zP+B7j
3T7afRT/uQQhq+CqqCEN3j5viDORFIMRGveOKM2GUqtaBCgqIc0yYrnLmlbhxXAVXs5PUnS4f3mn
saezUSxF6s+kDPN4uRwyvo5oBblmOXadK2KZj2/C01jNyXNi+YK4zdKbYSH2KWovDg8YXZFM4Cb5
rP4EWtp5VtlDMznbOSETPgC1fiJ3lZkt0kZgSWufMTm08BRfNvJtKkHOuJsPLYATK25FAdQ72T/8
egn1Pc4efAm1RtKaXiPRhXyl49qOckNm/svBQLziNDZ1wpgjMoSRtvCY/kt0ZqwVLV1t3PZPeyuT
rgkOv3Hq4Fxl0QUUryBNGtBjcb1LWf9iw/tsOpRb3bHoQb1RkR/DKHDOOHdZiZmDHeR7KZP4tQmR
2npNtQvQyIg5wvy39EWXKPuN6rQcNds4p1zeYclnHwpZpCjdKEM6OAlNVB+QB/d0mGQrMLsCjNxx
TTMxsIHk10UTznwSg1eNcanyokIRqSZ8RGr5nUlRwcr38etqhE6aa2XfCfSunUlROzS9+SR6t1G5
tE/Mi1BfKeNDzLy5jK1+7zuPANCphLHUA9VCWwxLbm+CV8b+TIPRJnY2/QZN84SQErvCfrVGSVhg
SaA8FgJZr5ReOYISjPlX2dLBL43Q4CHNqqUTOQG9ME2kUTF45Z/ovtbVHGbKwSAIzPaH65+0CJk0
sa+/AqDHoMLBo8N8e3xAJFluXXNlPp2lCiTn33Amd8oo3XzmLchruIRThES2Le09c5SEabV5H8Hc
2ady243QAI52fff/W3skDI6U3rdR6MMy4HKT7WZntgJEFj3YWyWgdGXMa25MjEzMws2iy3oFT/JA
gIqtocYAzdbWpGrt57gOC0w7qxL21fskdjZNXlVugPVNHDTKaASKJZHDkVdw8RoLwXEtWHJAbc86
ogpF/5eJ0Ao9YG70i6oBUSA16XmNqoYyLatlmm7d09Hi/fKJJYCQUapwwNAkD9ayochFTLakCOGW
vf4Xgjpzb0eNUkt9NCCi+ZE/ZzKIRo9tzf/G0wXJ7jPlKqKPyPAePHtqprHfFxfVolA4SbX1f3/l
UEyWgh6mIBMJGmHjx9T6hd74vJsKWfEmtK57jbLIYhXkCiiawbHbqTpS63pVRhTFmCOTY6H7x6gc
neKG1QOafMlliNWd4o11POTAQWKnfnEeVPElcJHz4XHDQEcMAsmvsvD8fIqhPpFFuWxfE92Eh26r
tNHBXrJDcrSZ9TK20g+YkNBXbCZyKVgWvaK2kepRcJy/J3xsaQieag8g1v0POqzPkradA5SsJ7Og
2Wym+XfVHH9jCKriiVygEJvqXNjd/g0wzo4Z6cSd+Kp6fGGfcMCAA27fPcRm50aUhvv4rGPP+Q80
soqhLS3Kl/WLVvtFzxP/HxaEGLgo2rCkbfxeOjddT99SvHEjnT/YSqzOnlgDX+zQQfMefRUsZHDd
6tESae9m4AJRwVU95zZAecM3LvSpdplUkAfShs+C3y4Lr9eOtNE9R3WVJ3waVTB7PlbeKRk4G58M
o79mhEV0y7ofD9UVs3PE0M5G5NjRbe7SNagrqbOm6Ow/lO0DGy4CtnjWOTZaz1WZL+DDHtdOM4CF
alfqfgpGyIUnfq8Z04sVpnw+t/NVBOQwbPQhN0k5qkkCU7s4c04vC6wdSDtrod9S3RFBWZJfQj+T
lOd0/pG62Q4UT+XEcMWAXR5rb/s9sXGGEdtbF3tO4df7er9mG6alLfNvQk3N8aNDj0o3TB1UhWoW
qXkeNISMpO3cRwz1EkGqMrp5kpw+o/N6Mc3vcHOaYT830tSv1VEHxrpq6+hxAHnXCBtE9kCNVht3
gtnpNLS5bbSPqhNRQYvENzr+qlW8H2V9gkDoiZkf8LhBNEAX5Zb+zBD3p2pa3ULSF/34RkjBytax
U4eW5jkIpZ3SCKgJISLV7EU73hk9ggKOpdv2fZ/ScdQu5I2d7OY9I7HZ8MqKsRN3z6TdO9Dnno9/
wKRnYwwVbM8Z45WtIXr6D9o1tvWCiYHl4E5tRGv4R/nSBy7Z4BpTUYz/ciWcQSdrB55ioqrRGFmS
gC5RiBXmGbIvFIRtf0AcoOJGESed26Vj2D2yyL9HCT2oPDdIq+bmkL0PrJL97+wlcLZTR7tiw3Wn
2EZxlYcFbre1BrlmRZTlvDBqvtCVg3Y43CEHFLYL0idBpr2ZV4WPW8dj0jXDrAYq4wXuP0ofYkif
FBvOIF2VYl3gcPSadnLImltqYE6YUJACGHpkW+CXPrG/0n+Bk+ydpDg2+JqgTojgyK1PKpjHsZlg
Leq1n++xLBSdLYk8l80TGnTr1lVHalgieBaDV2P9W55Lyo+l5qWqlfq8t8NePnm2WnbQePZYavkl
xOLmZZqEvcmvfeSEwWi2caotLC5rb8u+XTEIj3GVJ2Ay/sIDo67/k29rwgjyna4nkD3f0YsVpaid
e3HRvGwHo5g9NC+8Kh+vAawJiy3XN4rC7uCEMoxXltsPIASzT0oaQW4qPP3SHvrltYnNJZyZQmET
LPysesfttY3nYfWvKa75BmJWegfiIy86/sgBN+4rF4sU0NAVM0BBB+oHzOPFLYRICPhHuJj2sO8y
Q01MngMuGvXPlqcZRtJiQ5V/4FggWXfq7XKcYjS6MxedJI/WZHLi+W/t1RpUORpRqkalKDcF53v8
QbS+Db4xBhZ+dJHjE0MWrCvyIzMudzKG2Gfc1KE5ikit+KcB1RhOu3O1q3a5zW5Tqzu5polUQoqS
kW8JmW4kJrWwPZqA3QwvmwRDnkaF80knDpJ67wDXf9RUZHf6tXYt/Ah0iIdlPGRmeXaoa1rjeAC4
wLZBkmW7TgWXC+tq9bpAZ9eRkB1uuQeqTGMkz+ztG6+r7rZjy27uyiSy8Vsi1aVR7b/iVCQxwLjS
PuRVJLWmfGcP1SIlxtkcszgs72h1kywd0Zv+F4JqdLngReRcxA1t2AOXoZRPDVeg273Glsf+Bxmr
nX1gxzeySrZEHRTQ1Jvpip7eucJY+d4b1uPclyQxlV6WBRTtwSDLRBO5tkJpRxmnxV6Q2x0Y5eAq
J+z0gsrJ84Y5n7vsdKPt8ZfydFMMNWBskUWFqCLjobIqOZdAzw2BoQXUH5kHa2ay/j4jRQI7i+qP
pGl1sLcqRZuPd8++X/FLzlHrUjPxmjcxEyqizVrs8QfQflB2Q6Ha6Wo10tScBrBpxSNyzPQzgYx+
Dd45b/R+8Rz3NWVw7ZOYydR1HfYnvT1TkYhRtuOP5o8q/Lt5LTCZ6XZpE6aSnmm1OFRXopqHHHkF
VN9X4u9XTHTkkBESTGHDDe27gKnc8aeXZ+QMJhXfilHzbeebNjna8p/W3hBPuH+Hl5gEnU/Wh//i
Y1JsCctgrZBZA7/4yzE0tiAT/IZEEKqvuEyFjvOkhgOl58oj7nT6KNvfRnOpT6noogwIozsMU9yu
BG5kLa5zcpNC4iiSXFYxI3SSkF5FPPehvTVkf4AevBl399tzH2FwpPkcinX4R7bi/BmXGmQPihzU
Yifn2ZbpD6gFR5Nhc2w0P36dji0r0DW+X1mRboKHvbbo5ig3rIylr+UF0nc1n9pq93qtj3mfAhBM
T0bRCf6yeyyx0Swm74/SDG17eDOnxBZf46iYp8wKw2J1kvHUiruzbgB62fJryLBqAWsAC+LtCUtU
gCIYuyxqihU6JxYzV5kBbpPCswc2wsUVb6Y2Qz2eCGAFdv4wUOzACiVa4f1Vl3fdHfqS8g8H6gNr
t3q6XnuxvXKs3m4qmLuyn2C4FvuH3ki1PL9lEFnUloJY6EhJD1s0bj667KUYPAvQoXTHwppkRFnx
daFVeJQHUDQETfvpjjC5MG1cjQPvdZq8xMXyv3ygS6ETD7azQofC8kClmCpbRklRLLfeTRzWMYzA
qfeUS1tFyPouSs5FU02SnGSHnhJ/R/1frM30xhEn8VpSPsiZQNhN+0wSkPsAoPrGJsvXgGBhpS9t
tjzpCUs3As6g062vxIHjunC3vvHlUyfZQ92UviclYXOgAN5jc0txRp1Z5xYsxEAZxNTDhLHEMbm7
Rjmi6xR0lj81LLsRR50pzjQ554bFkJqBQg0nV+DUtlu+O+JL2I9kz+kxiutYag1WWxGNC+KF5O/F
bLt/ZO40kOY4kk10tntnIYRCf4e7Tj5pTiFIh8TNSW/f3IZQJf3yhJfOFPJuqNeiEmF8bOGM2mJ2
MSzM+PzYOgOHzq3dsaWDLDEk6zco2iQFQzQQtytF3S1jwzVAZ2bTu9iPEzQWdMX1iR0sHiPKPSZC
whWoE9IMrEcLyDqBzaMRvzsM85jYRtCoE+CukV5FDTmPjWxgThOPLghOeNBYuzJIiWaSjXHcz+0L
x/INZBfuf4e40U+wIKAWWO54H1I4YhJufqhYmsFhlB+SHHmRDcT5BoVGaXzfzdhPZCUM5i8We2Dp
yQn5SoPUQ4piP26D+3PGjfb4e6zoMos9cLhll4jSitaZjVJUb+kPk6sBezXn1fEJxyQA/5zh6NKD
g9R9FGMoGLBjt5k7WWhIXcQ5kVfQllirLvQW4NQN7Jr3uu2cMcPkuzIPC3yXCIfT4W6BzCQd8pZ7
5uYrdKh9PSCiYP57DmpBYNEgPY6HmpdatODZBdyfzbbsOJRUePlEz9uaW3fV2iMFGWpOH8PQonSh
TSZxuSiK1Uh2QxE1cTlqreRMKviWVxLCddd+GK4e5b/vYwBBrdnbYSfcPTF3+eOV/eVokxfY9I+O
dx4rcudgWz/Ssnkctia/ZOpTr1bM5ZFVHcjxD0O0DIgZ3KCEgJ1ar2CCXX1m6x8IOLxc4Kc6RV45
68lp7+WautN5trOlw1q4ltf1/ozV3KBM0ZPtkd/pv6/v61Ntbx9NqKCWZdSIcTJ0RlOiJM29oT9w
7wXqHe9goIX+5H/I+1QsCEcoC0VnDkWIa/rOUi7X10Z0/eNi5HvGu+FOXy+XDTA2bwv6MIooRcYl
E80PbjhYP9r5aKwveT3zTUmljHT3Nj0WuHBocTUYpRCCCEVyvlynK7jbg0mdIV51bhMGU3Cm1tAH
K+V71O78eq03hfLIBqZgyBjR7jOudUY1i1MJ+EtMF02n+jFkxhOB8zZpwIOkJVf2quQ0MayKT3VN
oXQY3q+MZiVUZsxLNOtMPSH3Y/dd+hQSPqTI1F+82BER2CC0mV44QGwlwWQnUOi7bSJiu35qWeCQ
9K87s7a4rOO86DKZ7jsuX2e7Dskrh1nFdTZiWAMmC3TCe13XIZ/wGwRh6zsg02WUMDIQ63TaoSvK
4ZsuU1/jdEc3G50bVnWOrtplp3xcgZJY7H47oPfhb6skyvKYEbXxlYnH0XwMyxRpRPfA0IZaVJdI
rDe2PELG5eXGUPetQD42AtvSVsXItqhd9avEJy2v8kz/E9HZOhJHwNIhqYpzM7YcLmzKzh0e4Z9+
+2TKDa62O05g4RN1UvOy3ZQBgHslq6ak589CSeL+LfK4WjImWiMDRdDLdwyhNTwDsX4gJaZaybfa
+lG+nYWnjIOa90EcVZMAf5oNE3Yb8WEaiAN362GiM0+4u4vIKTByFZRRcbDpXtKyu3QmoxcR8ehN
0c1wmd+T62mNfHjeKhNtHVWhBN1WEXjlSKXerw5QcCIyTQ2fAKhtYSq9EhSOvsNjs9XmO9qu1B/n
FxLWBzHE32us8lmTDfSUfkLoItLQYRU1h3P8tmwMbhR+34l6Kas2km2Ft9j43HjT9WVdUgjYePte
keQ3K5HIbQNHK4i9tp7vaNXW15Xd9izFBBRXD/pk4rSZNgJh2lkafu5uxFiJEBET3CxFgg+7KbUo
TbDzkJcSZQkbhoo5gocusblcOjRa9PJMYe15635aPnAQqJYYKbOYn9zo1OsTIv2FNmDMFxlVVfCU
/mmDrprBPK7/BroX3MS7DWv8RF+cH+TxjfXh86Is8V3unB0IZciHviNhLtEjw9p8nxS0kjfd0Kuv
crETpw1PeEf7FCHhvibO+QSHI2l3RzmWRUEejdEHmTVcGXozbP56Ua/DVV0FenEhcwKgOcsHa7iu
+GGvwA2a6SPZIpbPLHmdn9/0EkdQiavgMDwLBXEJCAXQgpu90XZC7U6xf9HZQiD/YV3ab7g0E7wa
LJFfSVL8ZI82V7N29a04Mys8qaG2mf7zISWdNNOxpflP2Xuf96+t2CqrRVqrnY4oAZVEQDXEGe6a
PJs2DNEutqmTnEhXPNKR1o+lK7m/BO09x8nEhaQ0czBZUFL/UFQ75wXnsjL+7MUmj0uY986Vpp6T
e5I6cwZ3aWCDvl9JfQrYWIRPJdHuaBalhbFPHeI7LqhZ2Rpxo/99qYI7PT5kokt7e9tqVOXF5r1a
9Ltf4R+S0UAD6FSNpJC1OG4xKMPaNf3qTUEf445reOwBlgXE/9HhdtYcd5Tl+oSr95uKMV0EfpPH
qbEkQl8riJbfuHn/h0MPFnmQKZkfNVRasU+jH7KYszuHjSB+6d6P3prQlMa1Z5IETdzox/bELavW
xYmLhJnxI1fp6B7mJn3XsDNwabGKchGKt5OhFz1+Bu66y37/H/mccPqrvIatFsV6UMvpbI0kkNb9
qN79sHXRnF+ib0RV+ozN3yFwXTgzDdQVsKUUJb99Tiuun5KQXaNC38aAWCEyLchvtUG2IaVGR4kj
bRUjazwz91Qi2HoDUtvB+vyMpSD4chkdE8SemfFaDf4SF+8QSIChvFIvXti6xNb0YDgtIrVGQj9n
CSSauuUz/B8ah1uO9GBdIx+6ScXfRuUAE24FQGwmLLUW+p2kt45b32bZc4UZvTg6Ar4GRyErufIB
7KRL8QY/PLoS2xkBAGMicpqg8DeHo0MKx+ht1YkiVi61l2s7nBMTuROCe0vzEuDmdsGtIduCAnAx
jfZF6iL0xtVVTwEvhLfNQuBAUGLhflhNcsfRNVvbpnChWfBr7Di+BLx3E76b1Bank4bPtMceyZ00
kyDtq0/DN/xCARB136kYGFP4LvFAr2VuyVk68Rcr28MCPZx17i0p9DevIr7wbk+V9dx3MRy1/6nn
KinYCWLAFXxZWz0VQJ8UPLB/+fi427svr9IM56vYphuTNBsOFtb3Pm6EPGRK/ZTIHbr3nWl5jAe7
o4gb3onRgcPM4yR3thi93oJXLyEAAeqoJdkCQOPhuEWoVO2iqt9NX4aIa3CAVTbOvrIT82SdEmI2
Y4GB2yJulrelk334xuT118J7IGSQiU6BADI17ngM1DwKUojpjF366mzC3u//cg3y2x+omFjv+m9e
nA2kjJFCxd2TMfkobCU2qICFvjpzOFOTuOCKC4psKLCc7E3BWdg6IrRoHH+NOwnxFXKhp4oC+xiH
1u+iICoSJa/iBLmyRJEO7f8negK1R7U0wje2jFktqewREugSsXxNjPvUGThHA7/uOZ09ErmdOft/
6KdLsKxzSxP2Ezj8tGzJ8d8/BUabk6ewUXMkFbzF4rKehtNSfMeUjXCfFKzbTrhMFK6uzPoUvjZ7
OSe+lVVrvTjDTJnUnyeZPG75US8TlKxlqJP7JpXkyMyGyQIHaLfkZWhgtYRBkQKvg8cUXsMsmT1/
WZEaKq7v2DgTHncikDoNYmyYWc3oU5y0FtwS+6biLhay58h00jGlFT/v7hvrsv6EKm2AACxVHLJt
pWifMB8OzJFb88spFuYOBDmYHCbEFkmfgSZWQ5QHp1QFnzwIh5MhDCbNBM9kyO5AfIKQDD4XvREX
lBZAJ4iby3Nacsq07Qb5sofBlTetA5gN6wUCO4hhAdJiOPrngW1U2N5NrahTVlaSmIiujE7ad2m+
R6JBLqKy6PuVYaVqn0D8jq5SAZfiAKlTLYH32AioY4eV/YRTxNWkXrrInjFYfNFLLE60G6ZV+wNH
6l44PfU6YIOHbzxpAUL88yr6udJX6uqYwRc7UCxLi0SM7PBGRj25I10UJKs66g15ksFocSZhaPv7
R2ZCaYAHIyBGYc/x1X5xQ7K7AMeygppbBeZ0ZjgRaAYPFgpX680fJUgMXZCW6xIlcuBU8ECbp48/
g4b+kb7pS2K72lXQU1/E7H/5fsZZ8/YwFH8qF7sCHwV/yGNFsPArYlEVaQJdeR/DATP+w/hRRBt/
44ZFjabG8jyJXCCHKSIFb/QqWzDZmqvsXGrArA5z1vTURx8BrtX7P5IAvQ35K0AcICaKlF0L3W5W
Gym5rWh+aw1Tew1kBWOMl6uQAybh0GNcg95ByhA/SUYRVWshrgnn/Kk2FnzBiyFSLduYLmkcBthN
z44RsF6zdSacUQuMNgwYrqr7xsDRLget2Xw1H0QJoSg2DtIokV4axXeolPH+soUkddVmZlH/P3xW
DH9YLO287Tzq//7fazYn8NiYIpBuf01rOxhWquqg935PfuNJ/Eoxe0KvqyyWo519e7wA8G/5Z6IC
d+oACH8BMYC1U2ffOWz9gTuvFnOw27HtiXQ9zmd7i3GpZ0uenQSMeulsC9gpg3HX261sD6wW8bCi
+ggMfOQ+TWE1MWwvEe2obqjb2jXdror94HbiNrFdzL8QSKiakMe/9HQc/Zg6syEbzNHwKJ8dc3Yd
vm4rNXhz6Rwj7aqC55S+kKvPZcqJt9P2FC9dNL7cau3h0yVx/mZRGZ2xQoA+EwyXpj54Y831jeQ9
NAWabWHlX+Q6HtBmNYcmiGSRBU1q4BkUPqO3eLwrlhZFCqYZMrMIIDViPL48h37L5VvuCkTciFXV
0Zwu4YTPh6PE+sTL51y2MsVLEhUOUmYGaeYrkUdeEFqk0awwNx/IDERmM4G5eGD5XlosgNnpbSgF
tAREaYYVYyyDQbQBpFa8aQiJOyqtpcX6e7pBPNMAPuYxPwxPuYR1dWPbTo7+HBs0QqWZg77zYi8l
ep/BVCdRE+rTZwyBaBCPF9ugOI1wPA06izJFwoAh1T3avbXjqsuVsztTuxxf0IwT1UXH2VUTIj6G
DlF70WKXxVuwvP/1B95GmQFTr9YZ2atcLsOmDTr0s1T1r6zjEGDe5fRiJUPVbUTpURfjnD6LvARx
Rzwfae9MMtkc6l25YXVmQSvr958GIOrnmOKZjtf/75LDbDTZ6lWmqGH5B2ps+EGEGsoPqVz/R3t+
gCL57tNFEZkDCRjOJ7v/MtwVXWA1/ypowqqOpmfYIqT/CwrRvRYfu9Nm+wRf3g3fQSNBg+ERjePA
5AVyuvFmtm9n9e0YBB7ewN5cHkS/RbIAp6IXwS2H92H+5n9V2CQvYR7OiCJ/Wwt/g935IjAYwIpo
LM2mDxy5lnvlgBYuze8f6zxutbDcYw4SMT+6UpgWQxCaNNNbHNIzBd2HU/4LyLLlUsmYCirFiOt8
P74El7ayQXK+Ev8RveE0R/tTbczRTxZLFOnIREh13/hBDda7QM3i0+PBSJJ/YrzmkpyPsypUgriK
+aJrL5C4whT5c1EZ+kIUjtRo3DcK3ZUuqnCbrkvMUE2TvctExosnLS5z66ZGuxFeMXXxuSRL4ijq
yCbfO4IEiO9+OaeOh1VpnBxFKJHkhcMgmjICtnLCXrh5DT6YME1AKDaNl1zLhdif8LQuqS05evY7
Lfy4UQrLENyEkGF3MuL7+l0Zx+bR5mvpazH/SrvgsGcKLOCIaOj+OtVIEDhBwlETK0cXz2Dhjo5j
JgoH3X6WHMjFUNERlRyDXXJxa8vpmKibRcA3a0dbrAi7e7CfKKYTWtp4V/es3qUbLH6wzgBrb2U9
RW6Pw43qrQgbofS0HGzWWhugr18uvyT/iO0WQiloNvuEV0B7jjRFFR70uhmk5k8v/Cd1aJwTBTRM
B9ZGW/FkEahwgKv5HR/Q5a5gsaC0kHdYWxHM98tt5bHxPMfzcjvFyqCd+w7V6gqh6RUE+DVNSavP
tzwY+jlXWtnKMH0DxfGEd9Hrx9mpq+0TXvQrJDtDg634vUtH803D80WVFkwZGa05ZCCFMnopTSw8
en/I7Xw06xsHOioH16/S7ccPIkmrl9MWEMNj+hyO45svZpbO1+oCoBPPwZ4IUMVU9zf/tYqxGfjQ
SyA93oAD5oDxvI1Yjl+3glo9SzNKM1f3zAlKyno1cXrAzKGDV38ZvxUkVKZ9HNvKcMrhmGQAA3Th
1Wo4Sv/MsGeUenPAC5XUUMKL78dkLzL3O8YGj4WL7bI8qx+e+/HFuFzviuoV96LBg/MVuyoe11R6
2PA9jb7CkCrjWfOte6X3eb3+xxP3jlW2+nXUhTfRKs7cK0yCw+lxgnI4Bk+vFeojKEez7+caqCEp
UcQJhY7JNGpzx4LRF9qedeR5nVRC7G42gqUuOhHmUk9nOiK+u6VsRMOd+nvWLYvyVr4iFZUF1c69
SRPayPKmF0P+pqHstIdHFKx3gsYcdkhiHQzqhq8mqyWbqQS0WxUFYCZHBiawcuPdwwM9Db+44+Kp
j0n0hUrXVjYVjibt+RRhRRCqjz0336mJUlaSm491QHP+bgbN2E6ZvpI4a705w3cFx0G2EA1OoA62
doJRn+0tyaPOcrcW5zfZn7B4P+prsmduH4JxDZnvcE9xaIrTTitCQm6nngsUuWSVzzqG2QJx/HJW
u3nq5CgqUFHhdSMf+2t9nqDDizaHpf92c0rsOkesAK0HL3+MFKQh1frVyap/d0Au6UVxeCM6GqDd
COXPITxiT0UKp4SEzs36712CzSl/qk0szSc/dL0cEZf7w7pUyGlwNBVpjmcV8+FyBoUezmCftuim
vvXFvNY/wKau2D6kIj3D3SALUJL89GgkAilB+DS08H3ovjSPq3hRqOCNZtSMfQGw9zOFkUFKSBoP
Ybc/y/038b6pBz8FDgm2Mcy5pLCl4rPu0hQq4jeob2NBNmRXlyZfQ+ounBEbQ+m04HPTdUrq9lsC
szldF5KJA3jdRP510RbtwaZ9R/F0CN7WAlhkn9bRzEVy15aKKbKuVGe7WdLLc12yKnQHX6xhluZ0
nBcl+WBCaF5+ygs1kBDG5UPtwjC7/UvdUyRhMhm0FM3Tau4iqmeTzplpoyL6ikjzwgDyvfZHPam4
Xsh8UYCWT6AifXUCsDTB4H816vThWcnyhDFTmcAjgTAXUzA5vCPZJ8AmjmPIhd2HxbKOT0Iwt0ZR
tOpNQ3EFbHcww9pPVyridedDY4OIJUaVubHNKv9MyuSW/kNuar40CJtiX1BFiFVg/pw83WGYZBtd
Dd4SUNpY6lAIdes+gxQZWoCI3WvVrovYnvkfrbesyhnfo3A3ORAy9WNGh05h3ydAlDn8Oix7o6Qn
yVAQeg+ryMZmry2gKFOFPldhN9c8DIf+j+Z8j/gpSMws/S22yLMB9ezc5g5536uCubRCGVs1i/o/
iu5MX2pHdf8Upu6Up+niZ9Ys4EVuoDxt6V8mrdY8lV+A7gp4xrUndZTfuia/8RWhxnOFHG8fKwJg
nc3mCxLZbwuJnxdlez8KYy6p7lcLyJ1knajUhAfaiTdPe6LibIfhbGWLq+52JXaIUTGILfLLjIxB
TB1oKrj4X+6cwozqaV93acKGl9QpXws4zIyEWPwFV2kXs4qcDK1mT7vgFrwaN1JqD3WkkJL5Er8c
H9b+IluxUEZLs3UHEoz9NBIaipadqF+Xk1jnaAGax0uctThIzThC8ksTVFRlKVbLBkff9DHc7oO5
jOcEkmAOeY7cbUetNaRlzjFQ4XgYop2L35C4WycoEwBzQlyVCnzIUFTcHwe7+pBzyGYhCc4zaqnZ
t//cLR11LSfL2vkUZw3XPBzn/fcPWRHEUShm+v3UsLfaYuwpxWBkMshMBEbfCwsZTT20RD8bcPsg
5FO3aWfrn2mxE3UQNk4s8Y8EkqfrUzjqYZrTwSHJZcFjW31fOqEn75ejvfzymj+wolhzSleFaLRQ
8+Ndv6A/QNB3jCngNvwP79rX/iqqcysvLx28f6MByTS6I5BAqo+QYgwzQXKiEdXYDXuS/rF13LsB
UEgYXWOMYvUL6p+BABngwudH3v/3oMtyywdFoxTxz479w96Z74r5KYlxaYkGTuBQmc8kLohz+7Nm
Gq1bNjnTOeKCRKkD9I1z5LvjvVgPHfG6Lgc36REh2zBqIMMiqQFEfHCJJXKRyINjVMU8HfudS8Wh
VoKtUdB+XAIf2Pd9fEPoRW9pTJwUK+UYevewx6ZZRa4ha97AOm/TExHwQOU3mTXSIwW4jJX/Tz4Y
7E0QkfN2BBRSvTS3Q1wCto+Zq1bxntNpPSA8DlXLTCXC3ElDYSb4hxpfrQw1xG5LqNE7dPQPdu1Q
R9HTWkMtbL53HPni4UY7rg5xefXoQ50d7Dyq7DUx1GGkOa6ot6VqdfxRzmoENBsjEuhZ9Dsuex5w
cqLU+dQh5rjJTz3n9v4z2AQqiwQv2sDgyetoXz4kh/rWy3equMv8GR5e/Ji5RNLtBTjWVWIphtKV
xpwU5tcGXYfbCoHhitNUP8LhRE+Qk4QdOHIVvxfccvhhmurueuK2o/WvX1KWILHq1y1QAMlmUjhM
G9YfCWPiRMGx8WDKNCN9OCLKAH2kkBg3iw6BQQJmy95scVc7grp/olgDGO39CfGz7Dk4Uih53NXJ
1LJxi8Cq5+W2TjyHTMcQtK3Yc0X+Acb3eC6iBPhSkiPcJ7hrnXs8cbmzKYCQHk+fLqEfT2cnaRrf
kUUaiJDfjPTx8oVpGZSwOS/SrXXByczAvxm/c0mI2phsb8KTmDpOFYC81i6fopfW2roy8COhai7C
LAJUrWknl9pHJq0RSQ/QGibjWcIW9o0Xo9/KBWicHAIeC50dOcYnlrcHiBwaLZjFe4ZewGeBk3g4
JbOi461Fw/Lj4754ZIOMNFcQdy1Jl2xbYYTgKtFHWm79rDKKp0u50ukAbF76zINMM2Hm+oUHd7d0
sQ1CgKL6hS5CMVyt5C55BBvG/tNKhb5PwAt1ZzbCC1kjZtLgFqRz/sOOohsbgluQdEhHBA0F87dL
sXcbrctUaXcxtLu6WgReIqrDTzl8chFrVqwFAwK+P/Dv2JO2JwmuCVe9y8XRNky4uUfJNvqKvOJV
RIHdWBU/09AuIH6bUWFCi5zayU35aq7uv9zKiwXEg8KGM65mtAQdW1ypZ+13F2GWiAFy6oqtW1Gc
MQurwk80UT/7Y0UI/KhxcOXGUwagccVZQWDGnCu+V5tSNWo5PSE3kLxNJ5WjqnFxEmfPOnKZXs2k
TOCbNa7F2Zus9GxNh2NEay18HOTeOE0X2uW15o6bpAQ88CT/xPWq2NrTyU7R3WQ+cvAT9Fct0gtn
pd9tBUtsXFiXV1l4JcWCi6E/KmT21MXRrvPxOzjqtwFlj54LeuCd7HU36pRU57ce8MxKy/9RllwL
z/ic4SplXEhDnrV+5H2u2B4sJGrl5rEa9KpuUg88xutKF9Rc3998ZZrrjVSXXzDz+3G8LZhFNfOL
SUIx/HpXDxtZ2Upig5lA1CNtHed0hrAAYH7Jz+BAy9SvWKmjvLMuG7A7p1O3RTQgt77QIVpyVYVz
8kJU8Xbx455QRGBxUDW525lyf8hgrqGYpmfGaTrzboREAH03Gkh0qrUmpUxC2mr2D6ZmQCXJTNmr
+ThykYZSMH7VX0utXM/6+DjOv3b+ajC7ohNx3iGdS9i98C39iIRwLN+QiPpBho1EGGMhUSPKWY21
8xr4yqsTS38qwImhBc/X9QGKFzMFPTIfRRuJqTED0p1KUE81ErCrttF5z2sed3TbRcnRlyA9Dqt+
xhaCbonggiRTG/3WqDs7xrB3ZE4KkVDvl+SxnnNP0rzAyr7hD64bY/J4HIJjxrnJCH+nLpBQ/LfM
HzFAVSlsFD7lnzS0lB+EtiReNOx4ui3rYO0Mpzg4gEticoFp68uZWG8MF/y3z1nGHptmmoEdJxrr
zEd1+JjDOvtdcO3Shsdui8h0g6yr63KxPGv2DwgtC17ZrQbq9NNdQOLn6WesBTIV//2rT8Z/2oCi
aK7DIPx5GKa2Tubhz26CfqzpciIhEDiHIY7DsDaMZJLE9owRA2NI3bo4dNw9cpix/EqTG7VW4Zz8
gdAFuBID5t+k/AgQSvuXlLo7aevqcCJBFPM1CyBsWHPw/xhiaFgIuLUnsmclqVVf9QTNzg3V6mjx
iuasafnLM9GD9whgSRXK3GzWY1PYtfXFZs4ALNkSOyiQtesCQ46RYTQKHGQcC7aqvavl3lsz0cr3
Gl13zI44O3GCkrTxzrwH4WScEDNUSzzNOeBAKXlQumzY/SyGVSV+Xo/GPOJmtto9oLfeuP93Xpdd
mlAqsXKSbj4JlHGIccmQqQapG3DSzLNkJxl6epqsPzxZgJu8C2NFktUjQCAER3yZsQlFJGBRCrRD
Ntr6a7PdOCvhxR6DjRDASeSyVIQME3nNq496hzDnOhihA6NmWnuu4qDlpgD97CNvhz7Ro6bDI54M
jlCSfOWaC+Yq/JpMZ3xAaT/LG8OwM4eThvoHFOei+Nb15/8mXGh01R7rC1Ls1kxBeTBHhJDIII9z
W98iLJy8p0DQkhOULpb3s8ffdlTT9Iox/Vxm+JvACnM+KWgzPqmRbe3JOJwreQdHsuiUYxPzk/Aq
ti47n3g6sUaKW/V+PxIL305wU6NqFPQceUtWrfRQV7Wo30RGnSLKsnyeMryBCLqCpL5M2CZQQQb+
3QJ95yd+frFF5vW5qKS4GXJH96iT9CpJcjZTbJiwoXCLokp/cJG7WfCq/k/5i3velv4NUtWegV4e
85qD20Jp/cE3vGrA6HDlPGfQfpOJGaHllmlorWO5gC2P6CM39utJjj6YIzy2o3JG4QNyQRPhPhwk
cwlCwF6X2EweqTL9NNDM52mWp4GMYgrYlynALhxcCDKqvWhVQ/kjWNZbSGfl1dx8pAGkJrdvOgax
YYBqWoC3YSb7l5ZT0mu5LqYpNDZtJTWZ9ZTwPxVB8uwAA524KSrRcVsCaciw8SCqBu2yJTskFcWi
k80Peq1P7i8TXTZ+yFpNzbOsK6OwUq7ueigun+vrFKXsIh+Zh06a+hTPnkD0RYH8r8TT/42+6era
y8DFdPwdhRNTA3Effjydezztb005Xeso2C+gjUbCcvoa1e7uSYbFHJm1nCD91xAY+oo6FGRA16cg
DlVNO12rnm/l01/zLHizEWBNVT8lL+H4USuRu1roolYdB9/PGw6AsW9Ueopdlbrj6v4jpoS/P40f
CG+0LtqwcQUedQ06IDk3zxXGzozfgJenJ1Rl4uwqxGWaEui6Hy92NUbqgAB7256LBANrhE2cl5my
NGTZbSy1CQ0Zqj6tB3Cv9E5NIbNikuCbFNqjBFnKddyuvRJN178XnTo49fNunOqQm04UbMJBQEro
laF9dPPaeVB3ptIxzEXnXVSjyoDI66DIMapcP3PS3ALdpVQwb8Yhw7naF5ropBQpq4lmLGokgOGy
2yCl2rB9jQtdCV4o38GKTWVk5Sy4x3gqQS6D2+UHOKC6baUI53yyp8AcDwVDc2aa1TTDUtjNS5j2
XAu98VJ5Tt9KKglkhds6Ov4AcnHDqjuun0HC9uJ364sSwUCBEddGiZNxnRhu7iEoSLDSkwV3KVm+
76xXV4JoV07gBBo8r8aqAlXS9VLYtPlk9Fiqf2MeYX8F3Epob3j7tN1tBBAEp7b1P0PgfCCdJumB
GswUpD+gU4pze/BOrqO8ZOSAiuIPf3dnJj90tG++ZIFkTX4ZGB3JwTd+NjJ1uDTgxea37TsNFWE/
feaU76Ip4y6B3qYaY2T2Lo30OBfKlqzcVrau+eFOh6jtJTClXY1LbuBC0xZjSY+nI+nngFMwz2d4
zP8/tTjvdl6OGHvE3ygYQaZQspKWEkPPs6kcqMcwm3Me+Du46upG4hAojmtWLNgNF2pzvvlgTA1a
Mgv/TyVZ5tbbzzpOP/RnsXQqzyhfjmqrQZpx/mc53TEHu3FbGx8mCN8DtqK91pbKxypMETZp55hw
KR5w1+QTDQHcKYxiRDjFC/JaNaMffv793iC0G5F9gHBG/1Tb/9KBhQP1b24ytIXzsR97PZ2JL3vF
9Vfay9eAUpiwfgVrC/XDbn6hdPCoDODZI363q/GHcJ1YhnG8vieHGJGdHov86IZawCgC9Yq1NaRr
BpL6XFvzpV2KrEREgZprUuGXxUl9UG/NChFzBsdooMtDU9xok3qAbHZzJrjRqBpIr2thscboTmqR
N/53fQpBC57qQ9r0tfu/ouTgWR+2Sbu9rqc5fWv82UMWOOd3sdrRibgUuKVMEQNCnmjcev7/MG/e
iWuVo4C18u4zU+WxrazMePGAXY3ZUE4xc2KFqAAIWx0kbHQOgBMS542bCu+NsYfPQis5Bnak7Uyv
Slf9o3o8YwvRF1gvI+fCbvOjMa+lXsJUF5eCABsFGfISVojkDZxy558QPbh7FI2NMyI2Iozow2hc
7zZnpB7I4RcrJ7xBtqgKYU0/LQ85zCD6+DUNOlwHdgF7N3RKPXhr1EEP20WOJ7VDGGi4edm38HI3
Wqfzo/dfREe5z46LJOXvW7RvmpbDl5BUzAdfl66NAiF2AmNFJZcpnu7Q00KcdntPzcdIi0baNoO8
PNGm6IymO43ATXtnwJy/+IewX51ACXc0jR4Cl4ojGPnTFFCkR9s8+k50hDMTaS89suypTOBjEl8z
rSdgFj9vU6Gg5h8EtUJK7prFU2q1mQT19oFITFbYJhs+omESF74rEP3wXnjyAkaFlvCgVip2SdnJ
BeOK6EpgG5oNdlJifxWnmPkZ4IsFhCB9BwfTtim1yL9+Df4Mrzjv7ItnOiB3O/vbMtoz2VtReamT
sbWNK9Q14mnY1P2xv7RmZMdEHkKz7G8LrGjuPH3FJ05XoDbiAdS4bVgbQKKYVv35cUU7QWNOrYgm
4WYd4H/dPti/EjcMHhNWk0Rm0saMdePQmiUBvXdLQJpKN8ajMB05BygpwD8Gqn5BoOskBSDBrq76
qRMI2laMvs7LGnmHlfLW+G/oXdKbQEaUCPjOA/mAUUJwZCx1ldUKzbXDyDT4F7rb5TjAzBg+kjw/
2DcRL32S1QR5nQHdvR7khHtnNGangxTl5VYGC1VRCHHESJOxsTDyokDvmiQL2bCZCv8zVOsLFgC0
wE4pgHpa6M1SMSVOPwC85thhIvHP4W4Mi1Xok+rOIYakZbAjid4A8KAZTLqGCRGP8G6ptgYev0h8
c4lltewxm0qDQeNp1oS/gFN3gnN2lmJz1KkeR6a4T16Z7OR1ZA/0bRTpOv6z+iy56ZRloYlS94mV
ye68JF8yuJx9lQ+IGF1a+p5ZFCXmzs7rYoivXMl64zSrAQ1W4bNzq6YeMejWA2u94V4nkpVXcsEl
O2YoohrINZLOaaMB6pUTfFVTqmCLLQJ4B+mdcjiPMHfLQq5vpvSvmAxi9yCe77AzW1/1MffgSieS
gl5zHFRQHUyXRPuF9jd43Ka+WreiIj4yZDGRjXVTCJyG9yfZ4AhxvcAvPS7LKSLjkaF0S+NI1hyK
qbkZWY8F3IKplrti1fEhpB3WK1hv/DQBKWuh0daYeRwmYIBalNvf75nly4ZldTlp86GiRXy9sJbV
6Kk9QaI26d/U6NHQK0H34+XiTRaEygGJ8HGSJh/Cp5JtEEmLUxKovImuwgBaBPktBCShCNBZWJuk
puFXPh9J5wUtPYDVbk2UYhvXFdtm22o8W6zVJTluUMw/c/oBxb2mfy5FLK7LjkNW+6RHj8kv/vP8
ecLmTPWNE0yHbOkrRjyyM7+4ORn539ce07Idi6tKy6aOqP5sZqQovVEfc679YcRpWwPMvez4VGI7
6Dbyvb+zoUJ+sG3LzLaj2Lj28hHmfekbPMabKx+o/JleAv6G0mNqG3ljZt3rHKaruMnwekwli6Vl
pVUaDy2vLfjbveV147105kULliihg1EPPPHlwSO9pB8TwCBQ9ujaWDEiXGogRFKzKDFoHlq7NlRG
t+gbdeJFN2ifbv8quO/oO4HwNHr85e95lyqdk2AlIAayaXlWK7JbFQECldq+VUmYFhLhGMXzAEqS
P8Qp13UJcC1ZigR47OhmR2mKU+bMo0QTr7tnIByExbq5X8+aT4e2bv3A5odWKn+eOxkZiQZ3OpS8
8XuHCYGMq1GW/wp/ETjmyrPMwRbltfr2TNKaY1gwQRGb10efSiQeC3dpmVodY8/e9Vt5VNLNzQmS
ciLyzjg1tRKprDt3v4X0DlvKWBoUORFfrJ1cueAVUZl35Fc0piT2uVCdbE4kdEgtq7Z4QEFL+usQ
huQgsKZKJhM2HgPkuJWcnIFUtq13eR6njVQxVHXfVFoy5H1zdTE5A9vh49NwplkfPqHNDq16esiZ
WP23t4IO8PyH5oaJnDYZBmlJCKfn7576dpzHO2TEsBUSbyRHxjbrBrtsp2Qpj0fNUuVHuDGYue7I
Vo9Z7MVv2WQwjAhw5cf2pE3rymu3J9Y0OE8q6sDnqVXUfWliHAIM4PdQuURVQmvtWWuVVdJtr0IQ
aGYuZYf81JjCgcx1Vp3E1CSK/xT7X2v/UXR1PJtm5+fIU/uz+UPozVZn1IbB71JUA3mraH+RNkz4
3uNjrsAdLpIRgCUg06E4ZoGD7MGCcT1e90ZKroyNg9x0SdpLt4LVe/FjONaJca7lWx1aubCXyXps
3gjbCd1E0JF5rZQ+gIpKEpPUvRM+49CJsCXMg+gTJPQ0UVLJapizMsAILP9m+aIm0t1ve65pKpEB
Rkk0beha3E+bkcvUQkLD2nn02SXn4IUGD10NqgEGoGTyap5Ow+khL97CXxCCjUMdIRY7flejMYIx
OwCcIYxFxa4YdDGhmTuwPQmWYxtjF88sf9CTkk/Ho9lV4XkauTaRY2hiwvovdqEe5xMTEH3wXYjg
r3zzLipb6eXXabXj8dhWrQZVmTPSTdWh+W1gzBjgqTPaLADZG246MvRv8QPqTwiE4YmRNfiyLGYV
mW5gi1U7p9CR5LR6LbFw6xGNaQ/xkRYJ+PU1ucGA3qDu+aBSf0PPsXFG9KmnCk+FnLoE56k3mIiY
cz3PdclIIaCL80VimWM7Nnsrqe5Ff9yY7jYTJx99au+1KIuZKVD0rB3Y0whrDuy1exbwVkyCu+j+
vn+DoJ6nABuzAm8/0yuebYl9Gn53oteYDk3Fe0Z9fqK3ruA3+2wWd+wqANqfphcD3HXf/Rs6R3Au
9AvmlP/Ipy+z1qYPBWqwnS1MqeHbHamxLsQKRw/eUdAy8sd6egs5Ei7PpOIkAE0lopW5QdcoZFK9
k+3Cups5syucZSzhOPZu+QJsF9i3JAbTUsKDa/glCdYxSKBJ56vtnoACQAU99Bbvu7gphDtqtbpE
ZS1Bf5ZpZQHTKw5bAjn0OxzLcui2bB8TvAn2+55y2rUW9zXwn8YStOsvx8tEQ3Nllb606zBuRnN9
rKQ54mEKuOY7QsA6kZn4rBufiWHTA6DpIuK30GHAGKfBI+18q5yct+uMKOnTeLeug4Ny5KDehbvl
Fno6bPasHBGzaWVHff4bYCGTWMe+EPxVzmedsOmeHByTzFpJcmqxG47YaOv2Ig8BmOxQrX4LhuLy
lGmslNcmhPZqMvfSNWuxXezI3PSR97OULDGYiJqcMe5xnaigOVij0cli9b8G//AY6KqBT3Qlx9Px
HzHWKNh+DQDdpEaAUe+8owHL4Nak+Pou4BF2wFwnfJLJHj/Ea4O1Z6h/rvegWeWXBVb4KlX3iuAk
ejr9IPoasRBa4wv7GQ4BwmjFksQbBJ5fY9vPfX5KeyRgmM7IeAfRd64nVrFBGJW6BahYcjqZepkS
yTpH/1zNfft/62sW+OHprgFb683tIP80fMcU+MjjK3Ksejlgkzyrf/CmVN4IoyLiOFaEF6Y1VVLR
Wp1qkvaXz1rpDadCUKLoDAjd/fdrP+tgHH2h1XJkv6TVLPyxtRsLg00GssKTVzJYR2nVbSA9fTv5
IeSwHTRA453MJHu9hTR59PVNN6+NM2y/K81ugrJMTfvcW3Gml5unaat2cXQ2yzuMp008DWSQQvXV
tMHs8kq/DLkQcWaS0w+OGqMbph8OsYsv7b28vWoIKaC9egRGfA0MYdU8UA+IJ+jFRdBlGE6MNVcW
PzOt0grXbmh5wqk8pi1BLTrzatRI3g1n8EVUEANR9+6xZFnIs+p82XW16iXJTTpFxVvDPElpIK4E
eZ9HtS9f6jTEJ2TRDcUxemq0JWUIn7/jSWKC2IxmeLCy9PRy1tl48STe2XSLIPf4hp811siue62m
bQCFLnbAB/o2ANC6YVU/Oq+AeHDPTS5YI7+ZOhltMrSvFdAl5nZYg6eQdyN3wmT8nMnbFuEXPtie
ijppxTLTMxBHN6u97Di1yilWbJXngTZ+eXdCqMp3pikfBSv0uu2ntmaIBn1toKfzSTkIzcRq+39A
FsZAF+yDgJvoaEWIAztLVcC+BcEqHack9+/cVHZiGyP/5WWouDzF2WQ0I2YbE0x/Bdh1IEIuB/FK
BymMMHJEkEpkMCzCJTq/fBrxY6JR+WwjOEhPyh2vmKQprfYcseHiNnhiArGkZIdgYtw9FG169MSM
9IoUJ0LzezB5TIJ06uHN7yyt6Hvdnjgfh3qvmuuKItTBuKrODvtAes0lzNnSn1wJ55oNFPsvneF6
/T4licRsDsWq7lCxCQZAaRGrdqPWKq/qKu+n4CqEHSl+tBbwhhPvutdxLuW62eeyljG1upEdzOT+
iBVOvOLqEEV40fYkD5oi40ejumirfLB2HPyQ7wXSvmpggYVN1iHsniJ94ZGY0Vw8gx8ue7V+/lBE
orrLv50TxxIkgF3KgOsNISVgEgbBdWgglbeOGtYMNDaZzi5GsGVhjRUsDcMf0myl0HPtcA/w3ol+
8orLpnej0cJc3Y7qbNBDALiEwdqtoFORRfJTMd+3zesZZqCThTGasYlzt199PCwYXB2emaqdvCc1
nZGWLQB8sdeOPEYXeQ6yQQAwVJwdwkZkJsNgintjHXmg1ToX+S1cCvZgtxJdjujFHn3vNoK7kg3J
sTpd8z4UgR/4AhDmFCC1UpvOaLnP3j+T0qG4TwfOhsa8fVjCw3Jm1ObKbGffVUo1WHnSY9PIriTF
FkucuGwK3j8KPf633ErlixL1bbBQNFQcfnl6nsrPLydsWZWQhFtPILDkhIFd/d3u6qZuu2oSZPP0
Prx9EafxI67Sw+PyUY44d0FQ28rSOCoEf53NgH07lvXJwJqrj3/+EbHG+YFiTGHkmwb7Yg9at6/y
y1XDl9ZNEmz3s7eSxqygfCxFtQkzo575/FySsfwS0UpiZCgM6MsS+CAx1/JJOLSlYeOPjgB6+k5a
1WC/oBwzoFyokLKaQIkMVMudhFwoMbOu4yt9ldt18oVcNDalw1du9cyVC+/E3X/jLR1YzbZdaGjB
bCeEV/bqmIRtblR5chuUXhDjf/A6Vn+UeTwUtxuOzRraZT9N8E4u8zxHbSuM+m7P3pyZIQI6yDKG
1H0uZfb2gL1IUwxdNbVVh1dKqOw7PBK8WLYs9uLcstORdYTrVI2/RyzJISAunh0RquSjhIE7Lfud
gAYstcV8pN0DGQUdCqwwn01ujwwzBl9aC9+Xhs+fWj6zGl62HPQggRmck8OoYnkstCm3crZJ2vxd
6FlrZ0X3xPdDnTGuurPjwmpk1XRbIb0/nq4L27kixrG1RJOLyzEshHSYu6BYsDAv8yu8Gbdvc48a
z1rMT8YHC/wkkSUl36JcpZgnmV29LQHhE3iZrqUZdLZmzZJlGOlf4wTTTdsb0qUbLveylxitGpCS
pKmw0NacrZG+T0tjH9JFQ3rrO8UNdXAej+zsdz4wYx+dCNukZfkT1nJEd+iaxJhISITuYTtHgqIZ
e5MV/FcPuLcDJ1Rm/HXMJ11Iu61ONkGKcoc/Gw4eI23ZcwORD14x1DzOUmL68Ok9NVwdHHtx3rpL
VxOUAjaiIfXLhV9rS4cpZckgxBIAFtHCJZb0tHae4WAbQYB+DtDYASkJrBBcNvNSvb3vDnXV5io9
ziTb9+bGgrN32v9sUOg71yVeRpUkP3owaqmIAb9Uj76fzO7/WFajmhaA3TOfmO40U6ICAlz6i4fz
V7ylnLnU02p4QZpXvToTXpIBMev85/BjXYMo/qgCKbULCF+VxQLu2d1MVU7g2MBkNYXfif9cz1hG
nGlHe6mosuWUc0+tmk4NUvuhmYkETI34pu0bFmEVHUwGYxA4st+SFdXz0wzHdwjXAfwVQ+Cumc4A
c59e2hlbba/+4vtGvWfE1v+4SlrGtOcXQFsniBWnXLu6eTLMqYnwc6Ps/gn+M4WgEMQmH+7kbiZT
gplp0o9PuRzGqZ/9JrLaztNCxd3UnMqymUv5INi6l4TM7UCyrLIXyqvwih9Y9DeHGlL/Pvx2sbU5
4ndp0iU4MqQg6NUYZ86flS4aE+CYNs0XaZj9D58mybu44sNiHvI5fWWlyTrV/psLuNQT14KB/XpU
h85+AhE0Cjr0as0p20fcDgA5O47HHRA9mUkQuMmTemhkUd7xdCJ5T6ZjItm7sky23+P5NPm9TIfz
TVM9OEywKQq0yZYt0v/Z/XOzTGUNVXs4mHMuBYPbZ4Uvwd24CU0UlDnyTKLDWba1S+frr9To1bm3
MiEC0w0ZcXc/i0FLoGDUZIf6/s9fkOCT1ntn80Xoep0QlZkaJn+a/8QNPJtnNEQznFPvA0EEbDJN
Lz5ESva/d/wT5kpnxOw9Q6peuk71xyloVt/T+z8hl31NgscBvRnO3lZfvOuxIf9axd0MKadmkuJK
BebNohzxWcF898cLfhu/VlRcW0nxPqK/kBZtpejm56uNpUd08DNJuXwvYuJy7YQ1cn2rKyhFncFK
IHk3fXvvGRvWxwWw7s5nPo0ZwxZ6pOnaF6qgUxg6eAo7VoNQcRCmunMXv8lhgDXm+FUUkNLHigs7
AdASNX+vbIMRRdnc/DbKoGlJl22k079XTPQwTxAEL+/kCcb/6fQGezgrgDLnsD/v4guRRDLZaQhW
FYfs1B/JObkedKhj9bqJTbxpu/WU1m81JQaI0N/kcB/3t11mUnqGpKooE8FfvG5aDlfxK+UIu/5B
9WMHBO4nRWC7o5m6Ip1g6o2wD4TUu56Rw6+sVw1f6eDyIyOueoZvF3qbTa1Q6Ocf/ekH88hS/Wvv
S1rlSUNYvgePQrGlaEdgyD71YzL6DfkkzC4Sux4FqqDWZ0WeawYiZ8JISkyojztTbZFytsbtkmn/
olyh2VRhmJs9SH0ag91aYs5KApnuJWduWQH0FlvPvkEaosWEvU1yX5DIDX2KbFeTLVg0vSRNk16i
mYEaMQJlcm2X3yUckiOELMu67oziatKEBQQNjuH/xu6fy2/Xx+d90H/GTLVIV/b736R8rdVZ3nBG
nhsr7gp1PW2X48V2wYY5dAbILkVt5btUlnPfL/B4C6CGNgvD+uA0wOK0S35fIoXYBLItcl7tEsWW
nhkfVLHBr5QnfiIYgvIMYkOkFtdycVYxP8G+utmVUNkaDdCxCJGjYQqH4psQFTXLaYQhVpzWOenl
gBI/Jd/R7oqNsH5zN99/VOOZydpFUIg8c5JxCKMEi+oJT9RTIn6S2diWLQMX8DfKOWEw1ogz2Ob5
A8eGhO9kVJDsGe+v4/xUBt2YSL+EaODHZVVtvGb53W2UMAUHwkeeDxJPSpzQRbS9ZDdmNMV6T7e6
D37GFDrkGYjb4hrCviWlRkEgtsfma43pewrIxfaXRvDQLnYAWiYbnlDANPF+cs2Nzvu90QlkHgHM
pkuSyIkElwXb9BiYx2Fy+vuejBrxApOL+/NDuIU/nWLuIlXvdc2qTkhP0pwyMPzhLzzW1sIpbjMx
tb5u7tlkJ2aluXjm3PT8UIyFb9srRGgf1GVBblLNUFJimfpaiPIeltSKfjt7Rwr+UBWjn7wBCtXb
QlLbMODTeRXBRQivZ8PTW4a8i0LyF1ivD4LSnVYRYmejMjhjJ9lL8Y6cZKQQFnKK7dT9kEqcC0XT
a8wKsBoGE8yEot4eecrJuqLYP5sbBDVFoweSGSxTFjM4kxTsun7IPxw+BravdRiALyGEWG95c5GO
8yF/VLoi4VKAJrlpRzuD/kXnn5OreRQn9GC5do+PldRbCwc71+VsMYficZACBOXdDfiIemD06PqH
JH+G/Gn22nc9oz9j54FAZJAWNRIhvuyNpVrB9COWv9TDjUeQFMLgTpgIYx0BXkybudQiTDIrdMwr
JN5IZz8pE1B58ns3iyOAg8OjC+Y1G9kyjrIpDlmdlop+cZkrPxs6BXGbK4gdWsoEVdeoKMcXEh8m
+mihVa5r0a56/k3uBhfRQIsCs0qTh17Q4wd5Q7p4VdokeHE+dtxivpMCZk3yoxJAUtW7tOHys3zV
52nnRI5xch6SpfCNAvXpOXQiPqmIdyuMDSWL1CtHKa//Yd7lfrG/Rv9zi6yKb8H8Dm78+XNu/iiN
tFiuKBZmw6bHREbAL/r+XYbhAfkMrv4UVX7GSTop/TeWP31NfwtUnI88nQ9+b6N0hBmr9yrW0oz8
mzN9kj/a0tHoxMVdXW2cYImB7is3pZHFgBAjRuosdiVsmooblyE3NFL0Ua00OQlVAtHtO4EHvSLx
UPkot//qIbsg08IMe2QEGhexMpkCDj7fG+hDpw1IjRUtfpXhJGXTWYDbSLczxuJEIyR95njt74Dn
F8OtPJwgccA2gHfZd7XxLuk8amsA1DRTNnsiOJ2tL53fMjFxdyiNp55ZFDS0vwY+jf+E2cUmzhhX
R3TD4wEsRJyfiTUyJmIB6nU4xD2ZXDX/e1GPF6jtbIz2NjDyY0jlIqDb/IYVeGn2V4J2pTg5mroH
pgZhW41kP4dqgKOcfqRmrXbdFtqOiIPA/tD7d5u2RR6oOY6HQ/HELKgALOyFTyRMBS5hjR9r+jkF
Q1SisJZeiJIlYTp4dkXqia/5J3Yu7Hj+mVtUZErbs8czVTlpt5Ia6UBvYiryVV5VoOvyAY0r7QoC
2T5gholvm/FTxJvT8r5RIPddNhnBGV4PdZAGMbu6i+kHp0jDtydNCS1gUMmIzA3w04legn/2NpZJ
NmaBIhin50sUis73rUYie5ZQxSIXHMRegJYs/9a4KL3cHteNWUDZD1v+P1NPBbyK3R5N7ldBgkWc
27StaUn4ZgSBpv54BzymIpUilECtQRoWgG69ra0PBjZlAEj44lwx3j4Ltx+NcNHmcFeiKKTJHTf7
LfjxRsesGFB5+BGO4og5DGHSgct99nnMCS52IeKdQQu0ZlfJcLfGzNhpVCWxq3V+w3OThe9YAQ2x
Fq2QGMTNgd0DNRzuKObPzVWCuY9CW/0x2mgTHu50Pq3QBrRTS5AKIu5bzfLMjHwjQOMDDqUKqS8F
VVolALvmQvMWhRgeHNpNwb/wkTs7MvSsa13Glb1KJAxew5YIcAC9MFrHyvNX09A1ReD61cH5czZO
672rzHZIB8zPCk0q9K6+LRfFWo9xF8bzLYRHCIcXLaPS1nlsLiDKxZAI/7nLRVL405phtgSRehCr
1RV+Xd6iN+XoBLahfOG0qFUwjgNFuIusnwxFa3WnC+yMwyCKR0fkLoq1LR5Qfi2eUU8iJFOF78l+
zPS28RWL/Av470QooxliujYJrDyJ6vc+WcQ3ZX0/ZuraoppOl5WYmA1L5CjHwRqoRpImFMl0LNGg
LiyGHdZrNkJp2hMp8iboMCbXaA1+0Ft4PWOeBvV9pnuxQd2L7pQ9S9VUtYhsDvxNKdstjmZr9W/3
l5zw5Ub+ls+sV/W9w3iie38Jb+j60rLPfx7z2Oe/n9dRp+nY/FxInk2l65hBZeEZh5ztPM3i8TOM
khtG1MhhEkDGC6drp2/qPb+VEaC334SiAoiwNT0lRE4PYL0GgkJtEWu5qY1XMqokIFP3xp0gCMy8
saFH/Rh9WacJD87TCfZw434UruDIuMHYJZwbep47eu4bWBduLSfElzE0whTKpmya67DvTrG4s+oy
qZZTDpXfZHLpwLV4wjsVZZKm51snDjXBzI7wRd/Rp+Q6irbHmre2XP3XbLHfsEoRVwiKETeEb5w4
DS6DZ9HLXrLgjU9qIVkIeT59p5gR4toSeIeAUVFZE2q1Xnr9V/D4HwmzT0Uum+/vOjeKg7hIs8GZ
AOZJiuxExYWOCmNSaWXSFrimHRDqrZ/yrQlq4zy8UpoAMdqooyQFYaH7nstAd65AnlazsVK8u0wD
dxjEyQr0vl0UKtQhE+gtGVLmugA2IIRXr1gEEVzigWjUI6BC8wsZEyV/kK66jOQ2wCOsem6LK3i0
FXckTDtA8g84oe0wuqVm1nOX5DWm50NiO1ltDr4gpc6vHX0CfcxqiMGN3WZcjGjakR41FK02WzdA
VjhWRpkVm2t/t/jFacc8YHz1XTzLwDaQOl1YGkqmL7hp4WFa9Ttg+QQsilmqeVZ8hyjKTvghuVYg
Xs0oLy2aRvlahzcoiYRJY8MuYoSJa+1AD/UM6VhHXJfosHfYWlSBmkdsoZbEJmz2uMTvU1PSTffe
KDG4UCQ+l+bQi8ZdUR+xl5+iEzoFiC1Rgou5A8ntxsRx97vkKDy5/98aLdYCyfpprlA5CHvjg7fZ
jM4hv9WyAx1KJLzQUfclzaA0yvy+SuEKBLxwQFCpaX908VSMmV7CPoo5EE1ofuDHnHk5aVIHIH4P
C+R2eHfa8uROdV8EPf5y6LPaxBu+xqytwdufE1JrPL6sVR29ZQibPqbA577zFNsDR5CK05vPztLS
Z4b8Ba8AIfWRZ3q5AzaY5Ey0UY7l3TYUsQnQnhBowq5MZjECTZwN1E+I5LDKEgzexIlOv+zbprk8
Sg2XzGQEbVnxd4iLKWzjSTzucB2N2x4P22+NEmU+OlpakC3b/nJmk5kIzv9LMeJYQbIQ/M56wcU5
Lz3jVmlvSJ1D6Sciv7HYyVUNac7ibsxXjaUbubzSQQmEfs8LYM7xV3dleqbROEhBZU0HU3K5rxLK
93Xurz57s0V/SVotktX7CPLp5K29xMC6bB96S4buslT5YHOsX2iI78616cNZZ1Urf/EbxbCwpOMK
S8ynQRZ6ql7CAYAAzEhqGBaUIWehbshW1JEeZFmnTSj+4ANizEtwMx2yliHEy94LlRPwNDoqtzwP
MWRrrJJ6YMP5brcoW9L/+AlNElz/8LJj5Os7Sm9oaN0Zn8A7UFCaK49mIa8U4qnU199jkxRWxeh1
5R6qo49Iv0y3Mtc9IT8nAx9YWg6w1/aOxb9eGw6Q35OntwQ5muRvx86RKFIV3QoKiozn+YI5BtAV
oeqVSFUDWN/Q8OgWoQaBV2vb9qFtnddOQ4UeU0qw7Z0FnWRUmkzKkZBIHXXsk+Gnq7qLPAFSPkcP
k9MXOPK0Mmbfb9QIviSltVitNtQoYPoHh7QGjg6aVIpYYD2DV5uOlg2urN6yn4aXHDircBDClAoL
JVqgEuRFX8YIZVS7zWHHbx6fJCZ40ebNI6D322uqjEQEXJrYLFblcKf40GuNAzie3S9+Wrag24PM
nJGYhQC6iV3vvQe98aSlORcdszDtDLftVJrqCY82VGqWIqRrWTTSSyUQ8vstetnfzhl0LjwQTHco
XEWKTMk130Q+L93YOC8VaZqnjzLYZrLNhEhP11H2GnmYEroTnCeQ5/yDEtAQJkoelBoTMZHXKe6O
cPnLNMaVrCeYaLT1TXTaX7NeSBlxvAaOGz3lsMqinZdD5yPk2BVbVINM+OeSI3C7wN4JkXBMtcD/
8vEbM1/qO5x+QTCr3uhB8NmMC6qzje/qeWu7CjJtdlUcSy33dJQSSOBDjgG63Y0LK/szuJKG/Xv4
E2eDlbjrdN4fgWERKL6uZKep8GKhUBlbv/fQNokLn5wle+mgwNH+Bi6OxzGDNCdh9T+exJqIoLBR
xcWPeHoLtF8odhcyXEWt78jxseswub6EDaS2oWII8HxxxUp4pf8CCGcVHqVlppKQGiN1K+hn/Q6K
x8VQ3ROiCTkACF/xebgE2840nKEGhEckkIYwlRMs8ZC45iGdaM/3ZhpsA35NwT8vUBA3AQMdqhYT
9yTDHCyRTihHatRPl9RvMPAaCbQG+2ApXxfQltyZtXiv6tfM0d4bXyWKV+O8m5h3duW7hKmYBbqN
72Wu77i5RdEKX/zAKahwE/M0nTRgl9m8hhlq/qgL0QO5fuHNGc0s8oFNi/8BQPng4WwKtQICXkCg
DUHj7aK18BzBX3lRfdW+zIeJRq4ybkTxMNWk5ZE/l40nnzC5X33HIu6wHR8w/XoCQQuiKLEZv2Sx
JBwlm12K6PlyASlVrsNYqVAwqTEtVdtVCr2qIAjF8mg2t/XqCrsYPbbl267x5E83ig8Z7Q0PkL1X
DqJfwih56WCnTt0jOJ5hABjci6PdUFJrmDFKl73+CCpu5hoIjbEiVHcGVVDaXxJmd3UTN0gGAobo
rjwJvLd+b3H8jue6VQW1zhM4+gkm1oSu274Ej2uiWh2sYfVzn69yn/VNoy3Pl6xf8PCjVGPyXyCw
8DlCxjL7l2vIWYJulMxmmWQ++ZylIE1KdDVSVgTr0X+WWW/j2RqztXq+bWIjDKFCfLVhQIRPOaHI
++zOwS0kUQgt3knCOE7QSEmkvYhE6m9NotJtbxcX/vT8q+redHwVNf2WzM5JqAaS1lk3BiVQNfJ6
jSWNL8rjk5HAr+vsuArbFW0JhAyt8Qc2j4x4DyHIAjfmgNDLfnxLerb+8J0t7HZ+t4JYmMEwW0q+
V+fNCjhP0uxxeVRnALOJCk7l6ePdTA8mfY9fjKWTRAB/hJ+63UZbbf1OvbaS6Nr0V6Iz93mWckOK
jCMR5XDrur4pri9yya8nbWbJTkk2tl62b2HQ2gHm6PnV4yrok2p0U0aPICWF9xGICQ5NqqCssBiF
19uP8MtzLGCvvf9R8Wn8y87uJOTm136I39z//TztCL9VPF9v7eEww6cqJ24Wi+iFiFDNi1R2dwWf
7Xrd10qyahGBEw7bimvQQRV5k/QCrXJJm/GlRs1fgoek0z34E+adv6Ke+SK3MSdZiax78fE2OWc9
yxmMOE78FhWZFQaUVUkrUm7cKRf10S1Ltkv08lM6oTcdVesfBH3QH889CLBJzWVkzf8Jmj/kdBru
qTc7csuKmoSyrLyRureUsKAZBRf4jL5HiO1pR9FscCK2BKkgDOoZqN2Ong9BnmhZ3ozrVB7tiJCj
rDKjxUAXjkLeiILHXsG7swowcJb3QcXqe5x5y4aPNk9zLCb7g9w6QRN+U3iRWCEBw1EME1ccsNcb
RDRQlaMkh+ZMFaOYdwqTgp2lu2LH1Owookp6+dpRa1I/wQ/PQrtlLB4jmzJU649bKtpEyxe95Ms/
v/VGBBErIMQbdrMOQ4iqbq8oZ9k6mILBi2/ewGXznjWL9D7GhoizXbTAVwjcNQy3P8bGE1rAjUe/
+bpVwpa8hRGpMsqh22kl72IjeDtEC3zHRMq4pX3QCsm/FTV2x+KgzulUp6Ju89XwdmghO7VGj99D
YNDrJFaqU8BUeAAXEACsIHC9VYYYre6DHiZrn0pq6hWrV0zPHDtiAVWa/alNgjSJyrN0QIBkeuSp
GZxTkvBrpwUWYgAuYvlKCIxU2Jo82PH6zuOYp4uCzUz69aRs7LabPV1FiTNY1Vzf83v681Q2CFk8
PjDAliFCJEOB35Eci9+ucbcTrT9umKU4ZsiGWUEgws1Uhh0QvJB5Y47WCUlrSHsOzpvrgrKkaWE+
AYUriDQoKje/5yM2TSX4+/A7ZZ2KbCXHT15k2x0HMThA96zuToHDNBpCs0pAXL9P+ahnWJmtrLIc
rY920wrf9bS8LpGmbh4Wz49p5ru+vSIcktcpeoXF3ts/akYO+2I/NCgiw2W4TMbPN2OkFGpYZLcE
XavTghs3827Asz0dYOGMEfC4I18SGm0sa5FPAKYz+S/jY1UT6AmCblG63amalYc9Ed9mbg3ikYDq
wv+vfjB63w8l6KL9CdEW5z2MjWUF2DijNAQi5VtB6iXwRoNC6AL5vUj3BPdYY4dE45NJPB03jfDb
wUo7rDuZW1zc3POp7QXC5Xw0X4ryYLoM4lwYcrAF5HKexQumOD56S7CXMvQ16jqS5P5czELKAQfv
rBsHvU5e0kk9+Bz49nJlR20Xfb/tQfzp/krBBV5cGO5X5iFGWw22/HUAMVHzosc+cVENq1V3cmpD
yLLyBpqzF/upfVvETnUl8S2LeXveMDXTdEFfoBic36tXMY+X64DN9SstDhwLDr8gIw9GAX+StVbE
j1R1oOIElJSnnHgb1074mUce34R16KZcqN6jM0NFNtVD0bgkqYtnZdbGqsYJNLOdsJAE5itGXUPF
xOshmIH/LgdYu77JvvIAtGBuIog+xyXb2eg6QCEBfpHWiE9ukJMagCnKXcLb/NhaAX6bOXoy4qqk
zk+CyIu+lbSoSObfcoOeJVg80fqq1WMpoCh/4e6SIExCo0U8J7hTZEAFwNky2R4kSpqtMDDVkbOJ
Pkdvy3r0r6lPODsvKlXWA4KJdXu4Zx6oooB104ydeKbltXaZEj/fl+G2esapg/Dxf68Li/4d5jJT
jazSaijGHEiEvZzgcClY5E/UcD1ZiEf1/uFUEdzpp3dLy4JcO69MvvsXWbc2DDbA+jl5LZm9fCcH
3++68SLLI7KJeBJyHZYARFMjr68OYXWHu3KE3EwlgKcKLArUxfwqHoGKDez4Mqo/rwr0z56bO3y0
NhKrGYIEdgjw4y7SLqaK2VcyiStRDOH2IvKCZP7AQoWRMgwkCsW6hj5WSEYpnV69OQsqlw4WHfhI
2NtOSKadyPFQYv+PWEhMrCXdAJOhW1hdzs0u+7L2X3kKKh+ECB1cryZgIn12G3M6kBy3CH+QfsZk
7EYdVfZEy4hFH2nbom6ESPp4qHcDexW92LqZFgwsTgZv2iawov9OqGzVcBP9uYIOpaTnbAswSPL7
LtTc9qxsGHDr8FfSoOOtDtKSUSJp4EaNeea9InZ+wHkYAOgr4UoXBEELhkbDkGo0MZdYErH7Xf4r
K8hcjjXakLO6bZgql2mBj+lCLOvrAsonVaDV1Gj37TKXaQ9oy2bVbpJWTxOAGeJXG4eZrzy11B7W
1Zo8C0+8/36RvQCcpcUTtsNGZWTLkAZbatLM+9VJhsoiw8Ls0CGzj/Yb++6iddU3CZxkzWYzZqFl
XfHqmO1RLWMQueoQcmSbI1wAB473+TodH9EufFsU8NX34aGwbv0Ukoq0LiEvCtU10+HlbOWYQam3
JkZ2o+f5WtWtwAmmKaG/yRhs/cUuRboeYsaW32+amT18/o3arLEIIdUyfxcgFbHUXCr/yY+Fwn6k
v/WZFCChYAaJ+DSpdxxQOSwScnZqadPl8IPnV+qxDg4AEOlTZWzn9jXgHNmTuFqT9ma8Q6av86EI
K8og+3YHJogoGonuG8cqRNtZYgfkjZMS2PTPfy/kGn1LaC7uiizOm4Lgdp+gOkc+dPIM7qEXump9
UaH7o6HXg65OnPZXrtLmCA9T+oFDAySuqkI9YK2QmDEld4iKJdHdQQOWB15AhPPpjzIGj4HGVrfu
p+WvdwdWmnQxb+RYnV1vtGoTUt68ma+ik+rRO+Rk2FjzvedPQQbu+jhw9f+hdvfyFEmfl5t1/Ivq
VpqPIMdTtyhF+w15OdU/x1XPz03Wiechg2DSP7MiK1HyiPX8d3pCN3toDOgSxoW9OwW+DLvaDu6L
2PpeHjpmlj6jP7G7JxHYQK02C7QfE8Ka2OiU3X8QRVoXJOMcbAZ/vR2FTPSG6B0vxKruic/Goj9c
6MZMqLhZSLerUxuKFgCZXZh8rPr3xaD+CXU9XCazxPO459YBsoMIpALog7cILCrk/A0Drb56AGuS
ae9uBI8v+su1uXm8alPdmGVLWbSCAPufnEuELs92E6iWyPFGUE+l4RA9Ou1G0YIAzBPZOrAuuqD/
v7X6tgRJLHL7LHOWyW6bqFbkh2CkZG4gGrTynF2Y+DDBHAJMzJh98bDTMng3BTOZuy9pi7ysbWu2
Gn0ZPYXPdh7i7SXyc0PG5KPH1jEqKXLi3gk3RQRioNsgPevC3gCIMfrsALo1PKCdwGzMsD023dAH
tm+Xb/R3r/KINZlLYMpCW6zQaWzUJDjhYc1IbFgl7CiG2C8HscyTYxxnXkRaWGPuwcqHFu4UH5Ui
k5hoES5XqGaRIu/qhY4+Z3Xpx0pZbjmpKeNeN18/tUbr2v2zeEYq1n0IqR3bmRpwOkAmga1HL65p
y+LvqadNnVd3IrBfZX4K19vPRqiL3Ud8jGF3y4w9UIn5fkXf+iSacWRCynOny7fIr9FPUMtiFqAG
OVEI50wmAsKR5AVIHiqlNvbFqSqlX4CNQbw5uwgfOKB+Oq0gU46eCeAnLj05kNiKl/Mda25QSFiN
yeDDtBUv8Cn58nEDSNsyy/AHSQ+WQ/GVPICuZOCUTNKo0uLWhXgSyt0XVWCCKG0l80cBcbw9+zGe
Nxz7eMZ6p1o45EBoAzKckj4snkJ/7TUAh3nZBaO8M8LxUqdEnw07/YVpGz7qjMCCuFyhdhRFou7Q
NY53Gn6zu4zAyCulhbfhnfxwgGC/w8TT4xyGKwf1KX0c8O8vC1dXshLTMdiZD9LGIFy50AwdbWW0
N4mzaSgA5WRYpEfl2b1o0R0PKuLK6SHOG3Dc1E25tNfsrHtG1eY7rAsnDlcy8bK2UqwUAacjiML8
WCGCsjfAAoKqj49918rtGOKCldCu8u5LlObDFK9gogbVVvsLuJ5adkZO2Ea9gmZGjK0P8jVvhW7o
yZBUy9Tm9pyrxluPRD/IWsEAf8z+r7dwUgbWXKorXX6VIIHetBia/zwwT8ez+3jzL+lOqZWK3dv4
PUFCmxWV5NVyC7pFDSrDz8lQl92F+19N2K4Bw0ojW5H9nHoPQ+cku1hR/K8pOIuBrDCfush14pyq
JEaFgJ8pHfeNRFL+BBsbksNRH+0PbxgXHPB2ACvlSIcbQk9KyWcMmFRvcj83mAgnfq3rijr5YATh
KiIXUFnEpFWJQGf84XWtxituWOxHYodLlFgvCioDjxw/ijDev0cc86HgbnHZgUZsJzoOfWVWjhwz
SBZj1UoJwLr9WBB4ENMvWy1NCBd71Y7gm4TQ4fPl0/nwH7Wwim4D6ZB9VkQPcTrDcrQ9IsQBnn4H
32UXrBODNAGcWuRDyz9RFVOhTfhmxTlegR1Z+s8eAc11nUdMLJiez+2sPECQvM2uD73f4NOgv79R
v1dmKCygW1XqRQdAbyCe7MmiqhyJ7l5VQAymu3GrhVte8ufVR1sQ+lBgXxl01pbi0qIW+yGIpRsR
t+0hLpQ6jv+ipQelukguUl5xWqds8O0DotqDcq0stucIWuhIfG5ZMCEpyzW//BUvrA46dU0Su6VL
Mh+qGxMMX8CWwnEFuOixedk7EMxnl19bBB18pFotyI0wGIgnJ/UP3Hv7crPhAqdJH5TZy6i/rsW7
oYigJ04lx5NdoB6ddjwwUZ+hZ1s66SF4d+f9ZSQIs6IBztlmYJLLYQxduKHnms+gjxGdreWmGNqS
gxnLRAUb+N8zlBaZXKzhzwkBoYkzls8j0r2QEJQfyc/zbDFDHLHD0rdKGAB1UJtVfiB3Uah2aNEK
xQUHjwcnYADkod9QZPFoMynom248X80etAmUEJfTWaPpwpmc9NfEea07hK7ySWmlY6gVRfht4su2
nW8uUNwNODKnIsbafWDI/LFUv99DTFzB0zJY55Z6SseXoLYkVWEWRsih92WP9CRxM2fe46Dq+tuW
8cj7sBbFJjDxOohxuQc5fyK0XVTR+CnqKs9SOiZ0lZAKWnmHYKYAEF7Un1c8ov9xWagS3PAdD8J4
68BkELLrJtcPWHPyscR+8/RIQfZIHh1G/4kKtbZtfuVT3gOLL6W9bDhsHnT5BK8e7/+b/E5PpAET
KLlyekIKfPAJi1y4Wql/u/pNCcXBiI5tSyF7CD83m5oWCOX+fgCmcjjKcD7qiHYvlek66go81vWv
iYgJTA/2nGf+JrHvnIfNzF6u5WAbmDj321VLBLZ/nq+rJ/xRTSp40obqm796pyZ5eeAPHHv22Vtd
4n/OMjifnHr7XYulON3BS28QqQaXv0FrwhJU0CQNMbRiWX55l8w2syz6fyIXp39v+jM1aRC26DvD
jxDs0PheKCii7xJB3T15mXJ+VdxMtUfyJeJ700/Sqt19AIyMgiBkSfH+wd2c9wIULunG9CGK1mCV
CJamdz8kerpnsUllu5tVl5zW4qILng73KEwbLkMmnTAmFQNYzr3/Yj3X2/IuPHYi7nXr0K9Y4zFl
Uue0nbIpdnyWttA5PcpJhEb/xRU8OJhX5wucMBkLM6DX4vQSyPcJiws0iVJiRb+4q7syLAMI1q3I
pZ9F8xyolqedW+YxLI1IABtEvyS44GcMc5etTh/W/VgGmlFRya/o8VdkiH8XFWyqNduO1nl9xH0V
hR+vJ7R6L+mKDnVxxDZ4ys33IzTgK0LQlVjlUY20Rj7zKlJ4ZCQnDYfXhGBX+/hoqfIrZx1ko9Ku
WdZszmrO0oqzp+/YiMfjgyyHF45SzprRXyYNYnQ5KDP87rAaIIUlvPvJQCIubw6VYEnM/1IFNlBp
ZaHJULRywEt/mXsMYF0YcX0SmOxR2jobjic5bZcV8zxdFTcCM+vC+uClcGLAdaoUatiAhdLs+HXd
8YDc9PfJlqywEJdYj7U/lZ0/XtkxK86dXd8ix7iKUvSVMEdvfK+VE9/KeJe21RPjic+pCl68QlKz
qPZngos7QScuf8YZ57lY5DaanvM7mGFQRU93oDLaqnq4AZJxSQtKgS/DFLQBlntFMdqLzoImwVgx
j+28c4Y+nqXvnUoyaBPDgyq+D7lD2+FvFmzGCOKNxhzVYRO1qW/l9/UJLhHEvZEn80G95yrfpxwA
dgUASHEYxEhdyNyh6VXxLEEXFvCR4xsxiOJbnfXRdkjckNq3W9MiFzjyYT68gmH7v36ZbmOg3UIp
XGLGoarC6NM2YV2VJ6kd2ZMon8wojFrgF3baCzZFwXfFPRwSRgfVu5MpDxrgo+zKSYKZ0s+LQiuo
SOaC7e6C/3tHbWCVBMJxWSY9XHDcVHr5JTZmwiWl9M2j6maK2oY+XA6oX8Ggl+5YVUb29b2rcEyX
ayVlbDGOH+fQj4Fyn9YGBJKwze3lb+fcvIUlx1o7c2ho20wDRrQ92HkuJ3LuULBk99wFlkop+XYi
2nHSl5A08x3gvM/vtjuB0WX7g1/T6IekHDP4yniuY9U6VlF8ETlXNKBYvc5APFCui1T0vyO420lk
SstnLFB8EGFZv0AgHoQ93EGPbiucj0tdvatb6KwuzrZQxBXkLpMdhRnLlbbd/DMfpnvYMfcEqxcx
izN1vahEF8TRCJ3m4i0xms/pXOq4/4jBPkhgKgzsmiQJ68c6tf20A54ZQ+7PdAN0i4zkaesBX8QA
QNY2z2tYPLFWQ7ThOGrG0G5N/wdCH53LNjKc0fFIDAYR4qpidzaJyd25L15W8cY0DBeZbiRPc0bB
L0BauY/Ej+IXefLF2h10OMa2JclvpfYRgiGFYgDLPwh9ZLkvBnId0UvgLnj4tJwC2oMwagq1coWP
LAyiOq6ncrHATwiQTjlCmtxnx4BddSskES7wSq6uM6mTS7YXkDohFu7fmpFkyydE8+svNdZ/1w7m
Abiy2vl3ZpKDRaXF5u/b97HLQxgLwVqJ6e2tJof+RtN/q406mPDO+ZxV1Mqcls72DkJB7oTOv4eG
WUAExtDIOWKBJLe7gJ/VTIOqnBnh711UTAq7NfEu/BeMsdyUAetCmkes6m9rm1VXKG0yqzQf/aUQ
UrfwDgMOJBnCEHgK8s0UA45aEgIHlrdjucUT6Z8R7C7pxoGn6WdFafbdQ9UiQFtzN/f4/m+iM/W0
f/p/rIGikBKlFvoRK+qlOAUiqF9/JJETd+atOL+dWPFp5GaUs1vG6mAKd00yBiIfU1BCqmRwqC0e
rDM/YNxN0QfuXy5xl1jk4VC5iUgmqM4/UkTso+TsmzpgZMwf+pMPiPEha9RaoXeWTTnwRSMGTidI
yCFW9ElfJoB+Xhj76qbh47D9DWdKp6f+NpCguAAq1tuRu5UxkE9RLSxFWUDmJD6L3VjSwdxRlDWH
eeZzEJHRrKAA7k88tfuZJFqjOIZ00fyW2eq4k9ObcWe8lE3TzGCeHoHFeRqw1mmakeZUdN7fqfsD
JsQNCqRpZa0ZxUOWRlb/xNW1kdntCRHZX+lEenVL/tOuuzYWqmIl9bqE1rcTes92QURW71t8Aq2v
SkpEHLYII0y9Rb0mYptDRNcIpvRVmlHhgtav24INC5xohfc7yNtZ8UxZPvgBTPMM+oZw8XNhzyQO
ejaltS8Jh4FWiMZJn/6IWwNYnyV/aXPxBryqz4/J0vJQwblebt/+LQ4DTpNPKsdbiWodaXpEP6Q9
3Z5z3bfQi/KUCoYx96qvPWA/84b3pVshEfFPdu+J9FW+iPFYMZo8Ptj+BjdB6g3i5SNxo1qsmRG4
SjgZpWBD4TR4qILBuZvmy5rKZMiBBlfqgxZNaLoJkqVG+eOhzujLYiYv5wQ/plpEUQWqoqN/YN9T
6vqZNwXMJNqRTKaIpCVNq/VO3928Ci4kqndsmss4P4B+aSHxIsnewjTXb9R6bP6O5+IrlsNQUp8e
hYMipet9OaCXDXIq1o4yYIQePMWlT7393IWtZBmMvdAyJT9rTy5ehEWwiCZKqplkezGpi5aioRkm
T+NTN16T9focn4XQjQRzJHVTHIsaepFMgx+9dzch7eW1+VybVCstmcS8mMoEvGUMRDVxkF2xcYtQ
VJlAALTBkdkoECm8WbDW3RuuF6qbh67KDLTewySKsyNj4sIUf5yCBUtYwTEZ3FHF3FP/EbmGcJ+N
2OthW8WxIm5yFn3SAGcqVyzGGvstEohKSWumfy1l3XKAur5ENNfxYU42TNfiboygkn1VA7tJZ1c7
Yq42xsavSYqsfPsRS6FzeOk6gZRK+G5LLKkdkQsQgOGKKt32YIfYSIqxY4XjW97GjkeDcZfzphKp
uKWsBSt8MIC4okNfqj2y60dFzoSeXzdyn+FP8Xs2qFquLQU3aqMSXJ7jTvBH7kdbXQUYsKFprxn3
NdNzama9xGXMob8iVl2Sr9GY8aS0cx2x0XcOMWc5HW2LMikp8JPSrMn7bhtYmhb5PnNWsq+TCs4X
bX55jZoZj9BlcGHTdCYskb6Tgc3nT7XUa3EGO5IyX1EUpp4CpdBuvc3nnM19vwrRIYJk1ntFI/++
f5WK9V+o2vAgIXGP5eGZgs4R3pEVPpJMwTspx/++cQ7rZK8Sh86f/J/eTNU3gHD0HZSZR006Uc5x
3/JulGYlsjTy1cyEeHmFKmyAl3Ar3+mM9tc36+5h8bIBFIKBWAKPSE6qE0Lh2VfnmWjtdyTpL+Dw
LJKBr99xFqdoREaw9Q0a28XYu/NjpYzA16S9IXRIgLoWwcn30/EDsykN+tH7K2xjr5eFCWgWoxDM
I0EHAAUaKt3xWNCCS9Ow7KS2yXKZbyC4gD9DLW23pTvmJEuDg4ydD/K3e6sHRaM5aaVXwE4wAHXf
96VQzmQhN/HFO9mFyVZiGABfzJRmMMbp52jGs5rVX/MHqt9nVeS0UxSxsmaPnoPfh8Q166DTfr+M
B7lDcdrZqrMZvP92Tx5R9ClP4tlPNMMPgnyiGkvulMvHDf6D+jW4AdQPzwlOuum9LwlQBI0vUFsn
bmavudeyPvyd+T0YMhh6bzjSE5M2B9v1fX5+o4kQHncpEy0ng/xQZR7j7EL/Yi3nHfF7wOpBGpp+
oO3466Okr5+Jq1Gzqf4yt/xRxYIVetPO7aQXM91gIWCHZi/jYKUAuzLSbXH39VcLNcxxDnCsMlp5
AQvJVBqr5gq1ENE5nzMbSi3PZeOhPRzpbWWIpYYj9/O5hp2eLTkY/VnR48mdx5+7OH0peXA1/J5t
p50FxBVP1pSWak9aV65e3Qml3sEHGD+ehIRd0B6wxDEuSBS5d/8oqiZFIexzxToF7VhyjwDDToqR
JRF+Kr3DF9+V24SghUb7kMJuM1TIAfReZPfu2+NVJ4gFYBocbffPC8PU2C4/a9kWKUKhZ2MFHIxq
7sqwB1mXun81SJpDPrSbgNGZlsPYq5F59wzZdym2VTCnNHvjPaekddgMGTFKmtABxQYSX+sbDMJ8
Pk2tH9qboXDxPKalcHU3BYMmKqlo7nRfEHkVAqS3xKRQj4gAZJyb6ilDPmEoLAAjTrMqa7oaAMRe
zNqM8lZr6hQtXa+6Jmoqvs9BUM4gW6HyrtLpVL4Cmz3Q2wVyZ6Wj0a9pM1IRDQtiZtZz+GgVm6S9
z1OHYtph2uz0CM+HdZ2QLX0+NpMgst1SEGfxEChFqScrGEArR3znIX69L328wtwjTyY9UpdqcHMy
9ef+sV/+QIgDwxoY+HAcKWWe0F6Msvil8PVp0+/QM6uE1V0wdU4k7AN1sCB73byv0G7r1H6HWqXT
wUHQi8u3oRNf6xgkbnDlfnTf7iXBvvtBWD+9XVfXLOfXcBBJBIQLo3WisIfwPNvQ+JPFCYzIMWSd
CkKktQgdu+CvTFMPHgiLsS1XzP33vHzNqfi/WzduZ9przMOfTPqbTyyQKAT9S9l0QfFaNd0ppMaa
t3nyxzruvLfuqwL68AflxQ8FJUfOfs9QXWaBULH3EFRIN8axRypyPRui3ld4mTirRc6TW8teigjd
rW0XPhNrzl4SNrskAqUgTvr9z45DzyywKs4T27Ip87atNB17Fj5hR0XPDM+nvnJRinXmUL0uQhrK
Md6qB+GuEuz7Wt3p+7p7HPp+emXcGuLJBfk+JFvKUUePcv1ztHHBCT3V93CZuQD3BNx7LzAx9V/6
q1GLAClFLKigC7A4HIxz7WY0/xsi2wXyuaNKPPF4eC3gddYxFSrMKk/AuFZE0lowyytoEdkg9TAt
LhoLwmGgMbtB6/p2mzR+5dHxWAFGJ9ZypX4TaDuztr553DP5S512Uk0ctjt1Mi2OgoLgZ/DUEYg1
HiNy6czNjniBJx8NbvtBb2lFjOCMUXZa1jzxDXK/ywmfn6g1JizbKIBwVKP6/ut88gCRUGz9+tUK
i7iiGbrDAU53vFsYuum9Ze2mDLtTYA/gZ51aKAVh1VLdmgNjRDa4rw8QRKyPDRyb+ic8PGrsRnd3
AOlDAJAJtoff2CzzFeZzz/cMDIinPXuI8eG5yR+EtAI8T1kE8lstSip8zJRVRLxOolqISnodu85D
1vsdwOarOBcng7M/WdSzfjJLDolqr0mU7WnmVDE504UrosugYUUczQhMYx+0GmhWTuOF2mDBVme7
rFVbJN2xDzisqYf0Wh02VQw+ajnn3Uwa2/l0dRc3z+qf6zTmqvGb5hVHEiWcsN7XDZI4SkeimAQ9
eEt7FBsYhw5YkJ4kcGHwHFA8MG+IlVUwbUcadSl9hhk/6702ZjUFH8Iplhv/9K7FIC2LkITAhYz3
0lI6X/ml1iRIGwgkYCLibtagoFl8Wjhjrl6+tjYwIL93ldw6D+wzFoTWPBZDglMoVWviBOCn24Ne
EOHrSg2zbHyjW0pJJVDVc69x/IaHmzd2+yBejAGSTVRoYNRVvsuweVZLZodxZWYcNRADCYhdhQdd
JWl3IgH+EFLMOz8a68h4hrUKhsTkDj+c0E7JskcVD5k96r/xMRHSBsNRG4omXaPXrnZlmwOQK/R6
RzDNonEEnsLMpyTGpeH4TprX/Q+9+8Z60jZPBQx0Qp3BcYiIM/uRkuvmnsye2SW1DJgOraMfSs6f
dsgIASz7wPegDxb8imKsPV1vT+yW1gFvSfnmu0fk42ZXwqjbmShJ5Q/KuYLW/gI0FtseGMYk5q2K
EWYw7jc1gWv+0NkJl0/cEjiYSJnmnXPBNrQX0XWIN4Kou5X4x3OibaMm4Npkusmon4FCdM5lqG8e
HsPY+VlOdLdDyWl+GIWM4glxTMjeuOx7wWOtK/xYf+OO5DN9Ue1pRsQSq1xl8MfBAuTvmI3c5zLc
YGZwYkuyryE8FlMcH+LnvUxqPuHX3YPGo8NqdHYi+bQvWJKICZ0NEdIK2tPxUdzxh+1BxPJ8Ff84
5TDcfQEmPX01dXd9TWnVidt2U2YlKc2PRIXYQIwaEQ/lIGX+xBatHMdwfZLu3+9n+tEWi2h0LRNF
e1AmtxCDiKaU+oCbYIlIM/rZ2Z+AP7st71uCSiZ/3xxWmNiKOb0W/sbrG1K3L/lOfR0DSvlZCitx
odMIixtfVFkpi6RrJDNIz/D/q0ggx2J+E74vfc9ygQKe+erlHosmLei/TMvjBNenPwUl1y3Ka4cG
5og6KkM190w6nk62Z3ih45apUky1ekuTF4LBi0hrMJZ9tNjY+1truCc9dc1JuUhpovkn98Z3ncVc
sP7G5J+nFaqo7XKNKIDZhqClZ/9OfDDJMgmJP1jJjfufew1ZOPtDYH/ttnz7dKHXMU2WyWNBcocM
dApnd8NfixpAW0vpy/AxB2OTw+2BmY/kta4EXM0B+AFjVUmLiyQCcDa73SowBiDmcwGs5OzwhRQM
qvSQQYlLurITdh19gM4WJgRQktv+SUA95je5pdMe0FlsbxV9XBrYzlOhRjM0tM3gp5j9bAc+0CDl
0hLAKbJjb2js1TfjJTXyHwiKpVu+x3iTEIAD6JWVUodGenwYFBwRLTmQ91ybdrv6lMLN6MGHAJCe
9VnDLzwrKh14VQZBfp7vL4g7oRsq3QoG33rpLAwXGGKwsgdT1VWfErf8fGRzvbRu//qW38ZoFJHM
cAajIW2p0utg3y/CuCuP/BN2ueMR21sm6M3WlehWl2hLAvA1kb2GL2crV72yHVXTAmJ0nNBJ4qbV
DZZbUrkCTQGNgugNvi9wMX9FQp+a1JvwB1cdAzHYjrClHcQchLS3tsGdbg/Q+EYhFi/oxobOlKuR
l/bAA8txVOa/w9zx2uRNseY/0A4/5O/azw3n+G1B2RUXSzcBEXrMU34cA7P4kJEtYsP5UJfqS42V
/bDQ8ATSMWgADGzUNHDugU/3AuuypmLtzQLBwmUmln6ecX7YCkZ3NFCZXJsin9VI5ifCtc9TGx7Q
8kQNaMmS5mdXMpeCCxetcqTyDZ2Q34awF2VfF3ZYausqWZLbPGHTcBIFGARhiwpLAZzExcRn7JQT
8qbAwfsMr9oGogU/VX2gZ34qUQyGQWe6Yyec5yCF6dqNz+Oxq97x7WkMzmgD8/4j842GA8gm/Enn
CHUbFl0ZEusfoMiKkqRMbQcInH2l01NgXSKo64D9gTovUyiCiui1mhRgNQ/yEp576vdTgJhHs48W
oFGA9qhNmfWmgK6xe/LMwpHM88uybiNmFx4n0Wo3Euk0O2N90xhqg3dfO1kT1nv/XRrvgDb6pQLo
oEFnEQ6Okrwst4q3xRomxIah5NE7qv70jPG71gCcW6QavWUehtiIhNdMSESHik/vGR4kj7/X5Dun
qVtuldtWkd/evSNLBof+WKAkaQCXXsjphqRXvj1RzQhe/10JBUbwWeuDp1qeFvTjLkqlNCOYBJBs
QNOlOPb6UEj5Ygh/I5EtH+sRlzMZKiG78JBTd64jp5T/RZ0qJ5uaBoDPggwey83SHDu1ZuwT+L6z
W2oxYqNzseAWbaHgnHZ0XLhOifd8Tr7zBhD5SxfjRmwdwDIxOvxqZo33glkzGAefDC+azcrPiT62
M31XPC20k9tfOB7oAIgxCocEof4lqyCyFdJSqoeOpEreb9OIVOpiQ8o+sDffHEn3ur9qI+JVbrkO
6z99C4kHihcErvmPAstw3CQ2Gyan/LRl/2vD0BbBv82kE1vNvVz3G60GZ4Kc7jWf92qNUPhgcxAM
2HiObxLwPgwUpyM5pZRAw3bOENbgOh042lP5BPwgORbp6OaGjpEMgNVg/3E6poi3ViXG3Aq7Ex+3
hM1nQfMC7X8iRoTkU2LKdqX7TfYuK6D5WUe5zpbFheOCcy91n06IaNU14YFw1otSL+pIdbIRa5eR
SXsE3MQCTqB/1mYkNHNxX5MEgSWrEx//f++hRY2EFAzYPdTCrE48+gunKt4lramdcfao9lHHOfxI
/pOI0swIy9GdnZg+luY5UXNoq7WipVN7edni5a+HtvX9tKpAeIFGQfgmEBBKAOzCCp7s7z7sSHW1
GmQmlIkGPCcnlQUoC0T0y3fdS5sFyo2npf+oEgD07hOnDf5XYXrRFG5E8ll6U0TcEV+VEY4rvXrO
tqso7yJ5tZ34xaPWlm1JA3mTPEd1Oa6TLq9OsgklEoD11MTcNtRcYkOajtvuwktsPFJRyEJqBOYW
+ZfE5TWgp+iZsvDUiGfA1xusx46h8pFxlI2+1S5hySLYSbBe/8GiwlC4hhyoUJqzH0FrxZaBg4YT
j2dJFFyxgbVs9jDBH7vN9bk2SCBWlVH4PVwpyvID1fBimV+rOf1XfadkehiJh9/lSzaap6ljZd+3
teHBGoxPruqAWzyy8vb1xj30ozVH/WGNKwE0SMa2CH8lw4Xgjyxsvygjt/owRpv3djxtwWnG+b7u
X7WZca/BTu1xVcqwWxSxmh4FNBk2ukB6QEyvXwKiD8FYS0241X8Hjv6Qf72xXQ7fnOQyP9DxtN+M
E0fko+GqyokK5cEoUoHh01TQMS5x7Ip//cAQNdbaGbPCkEojsuLvtlnxBn4y/ZmE9vbQpV8lO7yX
ZT1Y1V8HK4PBcpcHNPq89H79NpOIOe16xj9QmQPuQoua5xKYYidi6/r56DxigHaCwGxuJmtzDpkx
m1XhhFPbe2TDnVAiPqkAk2Jin0luSXVR4zgIq5o+eR9abqvflIgRoxEu8/GxX1VCPe8dA/mSbooC
KMuskqD9aJ6rMM6wbe9R8ATTp0hDYL67u7xxOczOYuBWNzh+cXDjkVYBv4oxybnTkFp7k+Yyld1j
cwM27XN8tyHWDjEYucy8B1BcPSuJs5bWm2+iaa5HMCoz3Zku7+QlhvCphllTny9Kux2FO1RjNTrI
piq6p6To+8k2k3qh98bKPkKHy43egAaURt/QZtiu6ypkyiHpTDdQIw9owpGo6iPa28lX1OpxsjJ7
Gm6MoKiPkBo2U2qdye5UPk3esWU8AXg8x2sRGCAVivHnN9IEKz8QuxpyUt2rBxJ9pbEo8b7YjByo
vU7nvEDznpw2cfylf3MwCRCt06DMNn9c3Kid2DSbxCNjtgjgVIJI3DsT0Oa0lJv5Pxn8Jd/kVqwA
Cy+U4qwmbWxxaM43xWaPKXztj2dOL4+tZHqOLvvbBqEBc23DjfiKj8R4p7M3IJtS3B0Lbt5kYQEm
++uiolIX2Fw21h0yz06WCwzbdcHA9ZjSCwgDDtQpSRYoY6HJNAWcLwVLoWN2bJtpGk7jfW1eQidL
KqZvtJcxlBL/fzE5HJ+6pqJvSeb+/ok1Ckcn13VttsigENt1avekpvQ5+gCyJnWKOa8r1RXDBzQ7
TX3wvZJgDCh94UJbbr/IZMwWOxGc/Vhg6dRp6MlmwIYuGWaonMg1IFlckpVqRVHIYwsi2TJF8s71
Gzz2FL+Nt1sfAJsHBGSmWycjgFRr6G2AGPaQwbIKbxE5Se/7qd2YQtnWmib8QFHh8XQQSIIvR6Qv
YBBp+e9oFohaUpp+073Qg1xE0TkT9+ojFMJaQQJBUFz+qxTl9s+Bo2cH5frdjvFd50kOGpGP6i4V
h8BSXCKz3B+PDnOC3JEEx4r53DzexDUZV2z2Ly0aeLtNhf42I/12CpsdqQ9itRw6ie4uuWwFUHsy
Fo6BVoY4DPSkj+viZGPsldinoG5QpRbzSCt7f1oOxbrtCsIqOcHokrAg0J+qFTnQKuG0mNDOJOnw
KpWJJZIZudCp5/75ORF6pFekmYiiFQ+ruKsoZcTniZQJngtn2+k0WHoP+ewVUCefNvdtEmD+YGcy
fvZkvXp2OWS103357LWMAXfBYliumJp2WlRdY1Oqy7e7a1flBHxSYcTjB7MEXNBzf+yH6gC1Pwyj
ETOrfQ3HimZHPAQ0rHbBjl6LWw2HkCbsJnnsIiXzdiICJeTn7Kq9xu+fnRWFfoYQimZbE0AidR+4
nkHbsXatpQD0C4xXmP9M3DOmWQAcWDl85dKuE9OoU28vs/AfK4E6GGd+wmwWpRd/6wglXp4ZCaz8
GNEU9eP0WFK41vhEy8Eub4MoS3ZxArlHobx95HhPzoO7/O48F01xl7GwHo0YB1Wknh6Ho5YE5Rbo
VH+8bxeQDnxTQoEktb49lCFUwn/hjex42Z9c0M7HemrMnD45RGSgYIREcJ3QfC1W/yjqvumbDAa2
UnRY8PPHyNqLija9OqMSsajcpF8+d5p16Kueumn0Z9Sfr4yfXRUSKdjy9aB4Hbwb2iHVApXpthmu
BlJuUV/QmRc9nqmaG2/AlNx48GKCWe2+P/YCLQSsGI4QARk1hlj8NQEl9f1sSa7+eiKFd85/kw+F
LqLtRv74M36yRtKtraBC5mY9bqyTZy7cDG/LKp95Tm1/6cOYtMVZ9iAlKXsR/vkpZhA8k6bJfbsJ
VSn965weFHaiGIfOEEv5MlxmM6NFoFf4TFqQv1VA60TIE7YLlF38yhuFAxj09QReK/4JqYYhu4kq
8L+rTsTG+rV/btyp11NTsQpuLhIPugF9ewsmQoNYZZ2aZ2w4y19Hq7rZvIxPFam4odEN0MUAZDZc
FavwWTKVKhJD1pyRBHAO1WIwcFnBwwiDhqgt75eRJnY2aHJ6zJZhB4YKtq2Zcv1/Yd7Mj96MrM8B
FFY4UX9jnXyJNobaVyYnJxVMGw/mmAI/vOwN1Nx9OeQG2LiRMqttz/u85/ObQyt7NgyZwS9QMSej
CJoBrJXtKaMi+tIb9k25K4CvBn+MHKuW8bssQTneKm1umiSZnmOrWkaq/DAmT5Q0SugILAR/W6K3
sMc8kMqDfQ5190a96fKAdGfmmpMFytYQcBhgKThLmW6R+fShjhz9rX131tzSD+90/I+skVXykTjd
Xs/mLMO3CsH2JMvdizIFnQng0QGZ7bOMtwRQ9iezwY7+MB6WkPpqnE77RGhO7F5fQwaI+u3W4jYy
zAR2aC1p1ChmPL7dLFfTLQD25VOriRYz1afeTsnvB+LpGz/FDJg+WNrJF3Wsx9l5NxSXpScUDXcE
NRJZFQpBsBoLmMbHM14zSE/1ZJKn1y2yFquqtHW6G+50q7UTXR1+pkHJwI0Xz16geVvER3H2GPHy
ZGX1Qdya4pd/eVxevu0WTDv1fcDOWjenKTRnvRiLge1hROE7iBLxPTD7SKbh8cc79EkTwLI+H/4v
PStDd5b2tQq6Sm27Thv6ooBtoFzupy369o+/bZZZdDTP5sAfDnR8QoGqid2VBbraUp0iXw7nBnWO
h8cYTjednOVZFb/xksNpTS0lPqiwRkT7wLiiFJfGA+C9gVjXLvYGTdPnUe+nleS3CtOmvydgrkGl
7aaTikpMvThrhT+cwk5fhDseTnD5tNp0y6/74B00l1ahKvVjsv7jd5R4GcgVDjThBezZqTx8GYmF
RlU6ODPq4VcX9dDhzaa/YG55V29cOcowPHlXsZKU+0tGbuck2uG1LfkVqjgA19xUSPFzJrNZ9XyL
erm9CExc4p99q2ZgH1VVhRHQ0ZzKP59/Cq5G63Ev3+EhBOfiItallzWlJJOSFwA8Opp6P5LvoMR7
7k4jiB6aOavpSd6ue5YCaHCa3RZTB5F9B8vs2ByIORcyVfZmanVVCbZwhmjPmTw28OkANVKKscpR
M4c13scMWbmcToRnPVxFFuBwhxhMv7QJQnMox0VBcBynUglonLM2kH2mFp79xGh4Wc7mX4P5dDw9
gWlNe4aHvzuhr7SRLbUV6ZD0v3c6sMzqtqAwADv1CK9BCrASaxCon829KGXs108i9GMZhc+S4p9i
8+xWwbV57Fv3xTi8HJCCDRSC5Gyyopl3huXGyR5MUl7tHF3aDzvXJ5s42fdeG5KBongrL4uck2O0
/DqR4hFtgN/lvG38jYV4BYuP1MzwY6XXud0VFVbxQ7bKwDs0PkrtARwb/dKaJ8VtPNvLwt9V9AGe
h/MgvQ9xv77ukGl7TNQ3MmmO8NXXRKdLFcp3oZsSXQCSqJf69LHpDjnZkxRD85G7M9AF4w6NQfp3
zA+58DX7lcZG71vwWJwRZKG57Nri7WsKyWSbOSVkG1XFJd4IZ4tMnXyvyzQqLcLj2tRDyKIstUrr
AbGyvg1AUGRBvuwIZ8hXzDLsis2QLRrtLVgoaqHIYKvX7AstTdYT6nF9F/QigPqNsF9SuXtAQA6S
ufOnrMbIHpUMfpfTtPrBhu+qbd1JosGhejMomI4Gg7s9idu2z7DksCZ6wB4agmlt2RiMsa+98084
yCKgQ+PE+zsNL0z/W3QQImCDkNZkS44ntRbHxyXHzyI0ctIoOnsFQgrg0XZs7XD3bUc5nmQotgHv
SB6yRWyQ7H7gyZaMUQYTFLQ+FjANZeZqZ2/CCozLEKpbBGfm9+XhIPIh1jbT9/gMChP1ibbD3xZ/
aG9c5W3oa341k4ve6sDc5ncD29peX/x7dXPN5qiKEXasSttq34nUGIvTkWjTTbAIdiOM/8ThXz2E
IP4ld7ZQQmCZO6bt7tZGPxZfvlstphxg/q1I627DGn+5wU0kYqJbQWXFvN3rfI9Ea3J+LWdv3iqq
V9QHziRraQdBJ5xRFU8D6eLPg6+kxbQgY2TAlMX+FypxMnBWy45izjN+65Cdl22mqfuUh6qXoAds
u6WCDpbJ4Al9SdHxzm+yzUiktNlNXukP3wjiG1QuhQ0e2V1RPUbiQFGMjurl/CMUCBpmB4S9X8iI
ZfcWyWsu15hzbfBqindyaiappYjKHDCo1ExRmijc4mnpIQqBJ/QWGWxLBxZBM8eG6uNSe0pwvwrG
pxbdzFBJWKdDHlBEcwzPkZYBzIU8klp79V6ZKDV9A9ziYuLTQwb8CEJIrhPQBVZHTn65trGuSkqG
Ur1Hx7I4dfjNel0knmZ8N1hnLMIdoZW3YGKeu4BZqadPZlNLBhhiLf0P2u02Rr5zFRZCHbR+BNnj
cDobTYno4y7EoMHHcso8A/32oqbe++2LDU+1xhE5R/Z1rritRoFVWP2V00dkhvYPdVeKqBh81nGS
Yag7hPJAh8SdGUpY1XrH4a9zQoF+8jKBBB/FPAdgtx+W2RUDqNcTrvHk0LGsEUOOX2sgqjs7v6q0
fmNVlHscJl4dq3RWZ6LisaDpHQjOvVeQbIxPexkft82BExuKpkVNBcHOK5p+av3N1oSevRJgXS8C
x2iOaRTWCbXietjw1j0dswNJY1JSPuS2O8m3EuxidIHkLfmHs4UEtaoZdGauk6Tif/3BwLld7hkb
OAnjYM84V2zUr5QC04BLET/lxYK6TljgkZagH2cQEtPmf9BHTACh7YBFoMKMxlr0ghrTTbTD+fn9
5qExXEADdf3HqYdtw9s9f7YwX2WLLGLEHl/3K393MGJ/t87cAPTLKuUoWGikWyfpt+kg3lorAypl
1J18OAmsimdDHGVoYNf19x41x2K2/c2MA09uQOgTHGSYT2mBM4gmtPMqSugAAtNFu7iotBIAvuzH
9edgnAEJDWp9EgdO9KkQ71WdZ58lVr/VnDLJYA8I0eI9kJ6Vktx89URcS/eWje4u2eHIuR+QQOE4
3i1BBtqBse+YBZuyqKjlHi2EPJMnT/l6TRmgSe7tBzIPqcE83U5GZDJtwSxhQ5t1oE2H9DYlN8am
ga7kaMCbwjSH816rZLD83JI51XjTwQzJDAxmsxKHN/IFZI3dBLIWJ6QXHL8eolNWc8bKS8n73Wb7
oM8DPPuQ+/L13tcCZph7LuTYqa2S0foD8L/RmlYZK1PpOMUjF3lWJ2UjAqk3MYfI3yF8KwtI/mCO
2uRWS5ABzZAV1zUFCPQhUI/zcB1bBDy1wLZx9xPYC/0lwGDnR0RMj0cbIaSSDY6z5KXRoTaBAKqW
PjavIzIudhnrey/oIo1yANFxe3u1w74mBL14bBpl86xvMleonbyWJ6AsGRd3J3o+1EU0m/rGgtoj
j/B84Ssg2TIDPxC0X6KNPaXgR5voMN5DKy24/RT46BkWpxQgbEZNkOsH6mN3/5gvb8K0Ya8DVc3Q
pQfIK/vltqXGaw/YeQBHwD7EYuaLlFCIIT22+GgUhbiapKTa+LsqVwDionAQLsKofSNn/OyVdxR5
tUH8CgWbkoMq7PasTU/6z7p4NDEWipqn9xApHw2adCLtyZSiZS42HIr8dESP5gbbp6fq2b9YC3V8
u3NoELCYwq47h/hmJJAa6JLlXsy9f0a5jGAGenE5iEWcVJda4a+oxeUDLVK2cP3R07a1cMyqv3KT
IwBpEkIuygkr7/iB99qHQx4BWfIs/X5GNGCHBuMmD/XgLM8MAn8c/CxZgDN0GwzCWJ4Ud4vo1R4J
eukQrCv+hhN3DxZI60vbtvBt5UU1Oy7GAlZr5UW7CUnRNwhUC0nSqY7yGkGXcYLlGGUOemFdmJ8b
BaJNVatC326RhaoGcqGmDAlfeXXjeQfj5wzBBPVan9VJmaaZRT3qsXmbG0In2PYRxDydVkJFvZGa
SqaVt1ISwbD52xix/NJeljlylBUqOpArvsYCEJlOPoLjWfwvL5+AMRcJ/10Quk6PofF6RLUngXEl
xBY7jXtPtvNyYgtkX4dIJq7USSovEZyuZm8TF78ymjTK46en778Uj2zRH99NTlr/sn10+TJpcCBX
bv1iwoh0xX3gRnX9Eu0nqrLjfNPz6YWPTpyv7PGb8DoZFFO3txLssFrKwaTBIY3OiropfqvIras/
UQ0scSvXGDVXLLwe54npEijTIvZgJ0YsHBBh5hxi6lMcMdHrrEVx6hxIXr88U3hAVmECZqW/4d4/
lTjNd37LgF03V00svRBlm4XEwY+tRWegMyp+FXkJ+iRnoCWoVVRdt8M91SOefRZXz9xm7nJMj4uk
pEKaRil/PiZje3UV6FR1wiRNp3wMyrsrcM31FFVAb4QtpX3KADeg5GlO2YUP/3RcsGYuHmx4Voh5
k/Nnc0ctjuWB74M1U5UtTw7TeDp01PtWjx/iPIodiLlNVmvs4zmUtNc2vBvglrYt1kEP5UPL0PwV
Jgi4/4FUMWzwXQ1hYKwyJNaXOaU/W9ru9slacmYyL+fRbULG2sMWh1ANKs/uuWKp5dBp8AJWLGC0
zxjTGhQa2PSObXasCIau9ZJJF4ny/o6FEkqxYpDXeCEJDOtnZORx+llVIqKmoYd3LsPL+IurxxEG
e1ttIxBYNLAG0nZfrGtmEIAlVtS2A2huuNeVKQpVTOktwglHtEdHjPIrhMcDOC8WMDvKVLqAurL3
K/UML21GSUJhRhIWej/eWkwWmcvfKGfZRf8j57uIeuzaxayBoeWkrEenN7SSd0CixBp7BWlaTw1w
SFbj2hgupfNcUru8+JCI+jq53+80awp8tXpI+MpbKSixikaaKbjWFT5P8fvgl+VWCgSmHlQNR0SC
RUP6MTv4m15tqH2x9Jb3+3q2siVarzIqWqvI1iMAVN6kILSRCRbNjnqsnq9AlyF12JVFd4XnFdA3
QBVEQw+1abqUZiA8jRHeVthFtCud2dBzdOr616mwPPI6jPErmiifL4E3KOlHlSZlKvEghhJL6NNg
54lv4AR8BCndLF7XKjEbupnkvJINqgAA1gHfgc9zEFjNj/L921ZlfwDXUlHhF2Ro33lGr+RK+nw7
2dIye0L/+cHbpmHwmS96DFknJztiWgcCjk/7OM5inPhWisxYbYhNNL4a+Uqmjwd71u/w7dT39kZl
sISuhbvjRXZXaoiKjNiWLe32c7l0H16HT1YlqWg0OuO7L7bGMu60XhQsBiBOaGxYEIfugiMH94j8
Q5Kj+bZnoOLJnJGIFMhpi8H/i00JxsahASBiuBH1lNDR69FDnrfb3w7Iqfcf+uzQhOl0V3DcBPke
i+zxXsgetIvDJbvGpEpgNoo1xN2INwmcSS9jmX09Jk8fOzV05qWaOrFAwCVl9tBruYuwIr0AHgdf
yOjm/EYcRNSpRAlBiTaMwPAg/YSiEXdMUCZSZgrTDPL9rFZBfG3t/BnNv6EqjnqSGdj/j4AXYUtq
qmkAIoSA7N6g3ySHZw4ZaSJX+APnmEElKcm0XSnYGRVlnTMFmB2MupPfGVbnzKzr8t/5XPHQlmXD
helNLV0vPV4texmjIQuojqOFxH8xK67ILbl25fcBFkPxDwiCQvlhwghFCacUMoyLwgNTHONrSdjF
3Cz8FoBP2Kvd1RDO6x+0QMZzXFHQw5dbc2eq3jVMLUU4aULJ8V2lUnFslOuaL6v/AgvjPUJP0rlA
STb81SuTdKsG7Yjke3Ld9VaTJjjNYURiKmxYvQNjzWvI6QwPtOgUVaY/KiKxVE49oAlNphftrsQ2
PEnfFYW3ciqNbAd9Wu8QHEdZfVWC7xerp0EhwIbp/COVhIC1rdOjF8kHCFXzNqLnY2H+13acquk+
dF7bJkXolfqFbBcv3wd+6Axd0RnTUTnnHcN3zusCICzDQAFKaAXY23DP93rylOd9JnUffinwoMYV
1RR/potQWg8XbDWc6/FcRdFBQdezwsfpBtRHI0Cd+F2XKizVuZWbsrgY7W0EEAmhlHy/igROjZ2V
5aOqQYdFsnEzGsRMCcpFNV6uyZaBUmxg3mVqicCxRmAaBPlk7KGxlmAdrpjUax3RXcelKSZWOP3f
9lfpIfy1IFpGyvIirm69dV2Ivx9vXLYe4RDHVLy9hv73302DxZ8FnB0UhqRelD3LFiTNqU6UTVzX
W87tO/T1Z40jtgzOsK1VpIjVojNuNMdUJI0YcfCP22VLtuAhsGnjMH6IcKVT849JU2RRHpegGimF
8oLcEk3sEOF9tIGjWrjNIXTtlS8YWRPU5qcf21Wh/iTGtl4X8nw9ktnK1H2/DBbRDOhDMfQi4xE+
JmlWMV+d9QpNN84vtQM1MDph2QvM/p1SYxtrRdPQagwwD96FDlGMrqJQqzgniHUkm3S9pfTIRoLL
pFfayKt8FvW1hGC+zFcPywe+oTFSHAh2jXbaJAX8WUBYCmtgVU6+O59EMK1gnZnD2s/oji/fKQSj
xQ/lMy8FoetczvoqUYqpYtSLofXuXdYDbgE6gvRgdBKWQz1syhsRIXcJDMcpzydXOCqFb9Gc/pea
/iVgMKvaSGw49W8eyYdtdE+2uMVgGX9AhAaSGmp9FNjlA+VmfvzygKV9axStp52IE//4Gh1tuVn8
rwFu0/JkmOZsSTWxFeMXXLni3IZtiBydDeFLhUKst96i038WQePrZ52EslVKlG6ozwoNM13h/X47
fusRKXjOXWykOcVhQVOxgYHb1gkFFADQdOeatMs+vkcmNguEOgKgSt8lhcFOAc53gYoXNfH6rbSy
xCKYHois6wcJtr4iACTleWPjcHOvxrwbvzPee58Gi6Hew8VmQbhl4J8hNSa/ldeBugi/dV9Erp8A
3oVwEkG1ia3E1izoJLMsWJu0X0BhxI2kV3SFl7ds2G/t8DHRKc0xBCT7Q0vGT4PeVWpXAOxEe6d9
aAZRShv+InKfwf1F3KHmzB2MGicAGWMUlmRr/ktywI3tBiPRfB/OeCD/4V16YtNXFPcQdVVA2fdK
KydGmTjb+BY2HmXy+YXrMpfKiD1vi0KSNjAOYRliA4HHu3rJR2nVljW9nqiRVZOQ4ueOQyt8I0lM
r+fnTTVXd2trV/ii2CD57Mv33i6kVZJFDeHoUogWnZmEMo5wSJ03lXxN+/6vuWzZLicngoHX5zyt
sNOeuRp0BLFmAPO77/vmea6aBcCj+Zd7o08IhoXt1NpS/3zDuKAm4ZbhX8/zqTh9rGHvQwcQjf//
y8qj9c+WQhwFFyvFh1gg6Xg/zcRHFY998OYLpJTq/SO+MJK7V0NuIAwxN+vsrI459Jvb5shOx3Pz
bPkmqYC8lzrfKMIiHPPiwhc3/1cIzzO9UyZQu5Uk/UZe+STsgjN7g3BRah3PxQL5haTE9KgDyHtH
iZKnAjSL9IopbbIfxkRvZFoI+tbmCu2EMpLw6e32ycYfWlVl4mLT19ommcqZhqPf7sF/e2HAX7af
IRs47T73N5Yq+ZGfccKwEvXrjoygphL3eR3JDN+eSqIIXuatsp8pX20VOm0R1IN9+ybu4aZo5KEk
0Ex4GCRiffW3F6MuooJ0E6Jn6jirOw40xijsuyayAfv3cmQzl+XdFCI0dJYJ79LL8pl3p3lYErGc
NwkA6PiOWy0W5sulqIaEeKnpsvOkRlSMDzZ/KexQlPUECnOqeRDLOlXqXIn21187BBo1/hBAuUz9
R3SDIRbF9rxPf+5edUXUUYWRMLym/YaR1ojsHnc96DYwZ4FtTiarLOm5fNfwsVK/pxjDp27tzwMy
PnWefLNOiQU+qanaFfdT/Q/QW2kkRyp7594IAjVjSQp05XfJAFSmUnkxoT6R2k0/Rk0pDzmQlmmQ
m9YoLoGM5KCMjtICA7zjaZqVj2nxaaP1VN0QmPRhJbhNvNsRrWwnzibQFa5G8TggO58GgArPzl9G
annMLcJ9gC8a0Yf6TT2UAg1eZowTOvTvWSbGIQAxcKeQRxIzDh7/rUBUQmKC/GF/Se/zcT2LE4bJ
ordA/dWsBgJoRcL+GiNYymw7vjT988K/qKYukPkTFfWmbdfr+EUhMG2zENcx8FeZBTCuPq5pib7+
gC+Ymjkpg/i+ioTK89ZyCLIOryc9pF1NhMCq2F1LZbH+xxJW7M632cYPYKITuKrd0xfdsiTeSIM6
s61zMr1FSwYN6d/h9S5011UDQjxlM+qeyhS5G3sbkelgIXYA2eXTQES0qPSy2wXfQn9TSt+PL3Mb
E0qUym5SIgI7LdZCZAUewSv2SZ5/xDLKzMM1pl6aEIsI96f8rKjukNIaXPDrL23FblgMpLIHeQ3Y
T/0esYoFEFd5YNIXy/QZQWhFm87HUbblLo9mnNnA91SDRz+HrELZWDve2ZIdo/OMS42A/xfTx7cX
sU4kvEHJfwj1xv36nH97AuMJRa8p/cThfABhrqerEu9L+oWpPFhyg8b/6Tw5saV9hRjjgmsYq9e/
RGD5waaA9Qp42e8ua0YHZuergRsFLX4VXvtwgBNFkl3l8I9KPEf5+aqmz4v18ig29ycjwDT0tzF+
/PWz+yK9c9u6A6Lb8QtJ4/sza8H4ooAJhqJdhObJmfiPoSNRmIQBYXzZrg9k8v1KarxnGOzCiKiV
RnkBrGVZbP0tuGjxTocIWDduLodaEkROAEYNTa/uSE/YyVd3cST3HFdMkt2GRt6ojDPzozCsU11q
eyJ+9043FK7YYpnOMDgdBuMKDkbc3Bxr6hm3XTn91Kc4V9/AOpB/nbMYphvQbOMC6EUsYLNa6y0D
StQozq2AJdjgOHeYgxXS0YXUUNNVDn3jTDv1cn1ckxrH/L/LoYC9rSH/9NkBm9zzIR+WG21tdX9W
LR6u3RwAGCH/JZxRV7axvKateOBrwXl3SiPdC6SNjJrv7UDxcG0l/QzHVhSZdQo0TMZ5pJWcpXPc
DB5amUbAf0dzoLDPTjyCkcg6RC5DWq4oFJAxGSIoPb4BiU+yo32CMOD6AbDcIN4w2ThZjh8ko/OI
/HpBChV+zYPE+h+nNrWwe31UGI7SN6DbSEjjtFQ+R/dQWH25QcIgBgLnv6KMDwu6fjy5ZRczx159
kUgrmoLSUeNQDPnXf7oSuhXnHjG+UvD4ulqxjomz9dr8NU+uACHNbxy4WG4gYDULHyVgvsrQ5CJ0
cotCdJ9l1S+cNHRuh0C5j++YydDhOJ1ld1hriZOdAZaohoge8FVef+g6UyttpRQUtDbvdpVv6Ye8
m/FLX+PwlKfXkHGH0DTtQ+Pb316wpRhZeEaS36Ca9nDamblzWiupBAUY4PVzy778vWeLhEiBJRx3
3PRv+C/OzpK3HFKCXJzyEnUG0krEIWnnZ0SvHOy3sad1w7lvpnGCQC7vyxb9AjXbzo3jl+2+umJi
4BsGvR9sRqHwZIMq5arnLEo3xE9x6T7D5nLMB697T0+qTFeqwXIz3Y40Tk8v1kQOLz0T6SIq6B4U
OEy9tUfmkzd9w/SSWtQhn/Oqv3wwRIxgkBvirUIZJQXIW4xp9XlMOBXN/EXxkNFg+8VFE1XbUilB
2ij1K+ebKOqKdVhK0peNHKUziksC0t94MWvtqCqEGrcd0MrV1+05Gge6bFH75+5XtEtPwkZ31aiK
TXIP8UeVBtY8kpg3qc2HK1AS8dsXCIOJNyVMnbnj0PzKT+qk2qSIEmY1iq7+pqUQOWwixcwdGfZS
zvWHF5wLHMQWKO+RlPBYGHwdAn23BSZ6w9Bi/yRRkukaP5UmMIOfYauZboeShiY1gKtiQCXCAlcM
xDURal3FU8cN6BMPclrHesrtGGpGPNBApUUHTQVKCxwL11WqFhTANTnPVJ/LCSp0l0gbYrULKQyg
qkTTsNwmQwpNQ0WcsjbC9LdKHyiG/vUd3m9jOGMbeFgYxI+1kf7ulgaHMNdNrnjEy9H5JNxHBRI6
7S7H85Fm4n8B407n2+HAXmYMzyrjpGdEUX7G2lDnuyJpMBNkl7C94LjVcSSaOevuCF5Njz4d1jWx
AWc1TimoY6gMEwwCBAknVbLh6+xwxY3kG+vcf0GJ/+dB3GqvUh4wnNQxkh5odHpucGomQkoB8zgv
DGh3+ZAmL7FahzareqsjruAemPNH/vI6cXFITqCYNgj933qYDHZoZiyZIKQoGI/z9E+KbMNPj1aX
2xhkk6GKiPC0jMlGRkk16VovntP84wlPNGrfhTQoXpQeAAiqPRISEpblKdiPdNyMV34br/5TaDyI
T/Bim30kImqcT5ctZA9m+hXHqTY7A7Qf4jp2xCwbFJ2gYXR1yEDLVfVw7fYYQLxfkhm9jymmeTQY
qq54UE5yIgdWtSaTIXdEy6CFoyBY3fHASeviH3+tf5ayHcFj2wMRjF4SGDG2Qzn4ypntS4uJjRe1
m1hbKMCIUoW6IiGjna6my4+2OSCjeoSrrLbQuUCUW/WvDeQ/hXSIKTd0q8tA1C8AuawDf6tNAJK/
oWYtuxC6Vr6ZLzuCUfQEn41z2kvZSyLAoENoisXFgeyxmMMfRJU1Pq2mpMDgNrnVCz9tkjY6sIHX
6eXXmxcU9lHtJtA6g66awaEH0rzjskPfsWa5AMC1+iaWw+OTSawJxpIuLWKsA25BuRxWj29CHY78
RqmphSjyYhXZol/Wd8OKjM08Vn6gRdddmvgXcpME3r64IxKy7tfFekIK1Ame2P3nheTm4DZosCYK
G+qozt+yRCcXRiBEjCFAhUlIzMtWbWCm6ATBw+jj429Lv5TVAsBdrPsyB6Hvg89oSVQJ4GdFyMX6
YNIc1p99Uux9DnzcWm9MvZ2Mtcx1gj/32K63idMVH1SctXB+VRZHu2T9FrevpUEQT8r8sbIrdRfJ
mWriSgqXO22iOJygTLag9lcYowMY3g/TkQz7NcBjLIoITvAs85i2dUsqybGTGCcz2LW3pwG4Cx7U
32p+Duob7LjDfFI3bGuUOT/fO/y/m9S936TAaQSK7ReJE5ur2Dcws9BVRQUVyr0JQLRy5FJjN7/X
InkwGf9clMb9Yz/HvoSmO7QPNmlTIk2GSSyw537wDIsyBIliT661mPV5Ki++znThlmsOAeYyynZd
rNvqgl0tm6IsSgorIK5RKIwnzFXT3kUPYv0x+ErmmE4Q7pAupuwAs96OgYA4Up8UvHHU27Rgmc6I
My3f2myqUE49C90hLVYQkRakAfegZfUC4ga4txOoecqQ3+ZtCrnu2Efe+zA0x9TuyFC+H8+V5YG0
yD/lhnxnxw1xFwcRn3MSezeYKgij0KEUTyV3KoIttd4eas2aOWg86cOWshyxFY46EAfczFHManO1
h11JlWVZhqqEBQXPgC5W9SAgQtxASFpouHawlPP9SqBCloXpiHYNGLiIVu+k9oMCoe82xfDlGvqC
dU3yt5525NZZ7BfCK0F6BsBdb/rN3ihsDumW9jGwIyuli71jMwvXc2FhY2FSnftAr/vq+6WzCEb+
N6PpkynOlIVcpke2e6QMmHhQA3pCzt2nn+uA+WPK7Ut5emcotfDrSxTuy1/JBk2j+dLtrMPwwYwF
DSv/blb70jYVO0n1CiR2rb6gvW847/6pBAZqX6R33UzwSpAFaUYJ3VVJ2leUQc8iLAEss2hVAc5y
ZpWbwFraRbhm3eBBGd8EJ5qk4JrGdG1+X6ExDc006phRm9AKRZRZy7HSJ7339UoQdmnPLm/tFsOc
PzaCQXAq34I3FbHmeYx0wow6SwEwzNhfTJ6u2hjYuvJwOVvEHf7u3ddoeTZAMRaxkMQFMcM9pSei
exHFv+zZ88weAFPgOSoa9ogGqDZC3D4zotdE0nv+NYIF65wlv47ZR5JkyWUJBQmG1vt9XTVwSYZu
LhEzwO04qnP0uwHA1+UXCIiW8RdaiPCVa9lIprdpRnW5/7JzpJx2AV7a3an4d75HzkN8IpckiJCt
UskYegCXGT0O3NHZnSzDetJBlpTemt4BW/bCXmFb+42wRulNCibi+t4l8ulJ9v9Y23pNGl8Hon8a
RQb/L8fUn7Uffq536Xml4nNsLFKGImAHuoOm22570L+8H0bHslZX6tzY67RmcrH/qglfotI3uh48
E6wqdfyWWKp7iTS9RMklmJDOUxgnSR0Mga8SXI/Au9/N5zs9WYaHRdSUiwIMS3JwFw78+fVpLyBe
LLOWADnRGMMW7jWpiCP/r+z+PcYBAznABIgXIcVj6CbWLSKdeJnE2dzlBDgFPQAP1hJjCL/QK/xk
OrrWdMGRNvSBV7712ULchvHj/OF1a8HZLN7+XfU/Jeeil0N9NA5rkzT3R0WwMV6p2jMnfa6/cubS
aDm62jqIxSAQqWs0tKqav0UKnoe1oLubB2wJMTxo6eZpdvIZ8u3KNPJ38uDapcgBdSFARkcscLCM
Gq4J/ET0HuFlo0GVSAGcY/MzIvhDzQ3DQXjU4JIT02udExa/8sua2/FzxVdpt7rGD5dF6Ov4TWwp
aMYsOcVVJZOuH8bk1u+mSEzA6l9hoWBVpn7ExlqiF+CTKN2qLIA55gqDkiSLEmrAoZTX5uirMZQN
kPQ/hB4L5yyUpfycY0R+YzgFSGMdpg/KTH/CSqsqDdr5YB5rCcUteXy2bvKcjRK9bJZskNTzi4dz
cK7GBpEeKKMrEuzKZObjSzj79dbEVqteJdhQSzXsA55XvfI0rdGbIek3sWqlelCD2P/05zq/5QgQ
BJsw1zoZ5fwupyUjqTMMPA+ixUietalqSQUkwgQ4TdmKQn90w7DORrJ8o/reYqsTLJQJNRrc+Shx
Xt4fH5G7eXfijrz/ne3kyertA/76WqNAh/FM8yUAxt+ZtkqGwoQhruA7vS21fOo4v6C+qzDYRT4J
Th/WjWIRh+NNRkD4IopWsXogOLUZipH5DIuQVqmaY6B0afOoDUG7z8+heLfgGt1SPnf9Fe2hKlmB
M3LeTV/Fz4a9mRUD51LgX6SE8+Yqmsn4wWXdqL/kJjNUtPdZGPCc6DoBpu/bSd/ZB+bWdPypVBWX
RHMQactKptsiIi+RMcmLOwAvdr2t24bGeopz87RgCFh55rzEfJ2IjUBD6q/Xf797FA98h1CwldZz
evrklDVM72o7v+0YcgH5wySvn/dYwYARJLrkMAasMBhF3nooYR/xHFbZhViImNN7WddKuIs7lvww
VmnZCZPEL8BE0xp6gFugmdIjhrRgOLoI8EbhZ3Hcze/1Aa2kK9gFNOB8gE9HgAA2i1CrGDHKTLMR
NDF9zKcB+LSz+KLlZdne64zB4EdbIW3YRqQuziIPNgpOcLSqbv2/AYJpMzWMaQOKCwVXQSrJSY4D
3H5OwxwwANC44W4JyHgMSdzE9xxVeA786wMnZGPlX28xA/nQxrPv9MpO8Z63ZQqex1rI3ZH7bYue
Pyg7fr0rjA+ItDzhx0/k5n6K/RAL++oa+NpkrHMB/TQZqG8+Py6zdQabs+jGmIajFwJJpQ1/VHVU
yBdgDZU/HXJ03UZB0pLGEH2tzIgYsWSuPJlcuNc7d+hJPnYBhYC3HmTOmC/zQ1jK2IXn7RuULhEX
B7whLM5TDJv9zMU+PM36x3GCpSBunhZd7SF9Fke4bz2pfF8MPaxIt8ZVg/WE2Yd+vF5bswl6JIB2
mUzH43cZk0JaAVWnLn15ZG96ymt3bPDLg5lrXrALwObogD+rIWv2iH+NXRB/judkHJ4JP0bGdnJW
PVvOs+CtAsL6F0UYBQukOk+xseKEm+YYkxcNSbTaHhRfNuk7ch/hW0jtN3dzDtBhqTREUBwCNQCm
Agg46D06BkE3DHuN5RojNaU+BxPv1CuhSUZUCROowX2deQNguYWsahfV/xxpATFhn9BQCtb1viVt
MF8m4jZ0k4W7bBWIkn+6RXPwSC93tiAVie5UeGDy87obsZduq//2V4IAv9trQAgUCEBWgCNY3w1e
Io2FBSO+Xgh92J4ug5pIuLasNqh9mM5DLKIvmTgnK64ErSoYzUdbZF3MPt3d51NKnQVsh8NJGCOA
lqXaiEqwL1L4GtY41XAuTFvRgvS9yryeWKNGnoGpQBgL7d8P/Enza1jLzNU8GAeR1u3YN/WpH9x9
Qxm1vSdfFBxPKQqakZ9eyxi3OxChYkdbjpS7D3mTzTXd6u/uNqYrRErlNnmpUfUh37B0g0Rf3Kf3
SG0mNW1UerS92sZDvZ1jY9KBNkjiQlM2cFcjPSGMr0Qa4e0GSHkg2sJCSLMADw3YlVPnToYwnt2+
eu6tyvEPLZhtkhQE4buwiXv15/I7VPoKmo/IHBY3lOy/6njqlbN8oJP4c8b42xx8otWL1E+DYRgq
ioPSWT9gCutsiZ/otUQX5Bpx5blGS698fgcLaJWigFBNQVHc85znDqZSocjvpzVFvry3vetVD4r7
BuoaGQaHv4VNj4tirOnpxa2y1hzrHCmv845fyPBVnWCXpNaSYKBf7pZY6zr4i9UUQr3QyhO3qZwB
OJB83JBLlk/LyhCOCfaKC6dMjJPoeH/WkKB9raRsxYtcIVesmw1NCvA5yQ/KP96DfVHTH72RsiHp
KtEFF2gwlM3j9cQ6Ib+5mM3LSL+WkNRBVJfdl0embfDdvneXYnpwTsH3R5rcmPRXr4L5Snx6V3ti
MjYK6BQxClNQdtvaZ459gX3Ndl7+uz3w7Mzw/4xrV5C1/y7qGU26sxy8HXaYxzI5G5szcKJwaJ53
7VClnu6AUDLjns5YXow7gqnakjtIR799St6tuJfs3vqwJ25TO7yj262mW4zoaUV1WpzTFO4mC8Hy
Vv1Y8ICI9urke57uYWFoMPS5T4xlUnhkbOKhiHGYBuhvQ78iNxTo0/6ARV4tBjdeonlPepxoaO6/
1izTKVTGGs6dCanY0Jds9+dJTrsCGTT8D0w9mQfqj/gR7+PI7A0jFzfdUrzsX6lPk7hA/lreVFxM
H+QjSJS0e9T83Dt9Hg44+fkSO5ne9ZPqVvL9fu1ylapSz75MOq3WYgp4jQpA9KrQWHlWdHYwS4wq
Jo3uvbr+HWb88Q95IU+PkHohRm789iHNQRNuKxa1GoI22Ia6iRcVRl6mL7urgtnIHq3LSYC2gm6x
2dBUvnfIlvsanZdRDdo0nZzBFZtGMdpU0pABELB7iPOefC3bH4w2/YcnXEv9qbMrw60H2LD/MI94
sxYse8Our+UeWwf6H7pfcAT1cKqH6LudY/ZLlZSeFLJjhfhGo64l4VEaYAnGSHxerv+r/+bH7u0o
fL9g5Pl0D1spKVR9bwhBraBHY5/fLnMlsG4Mr3bhVUqhouIiadtVi424GtWybWhAqKfkUfqmzznp
pawTbM7KQlf2gwPUmB9PD/8XNRo0ILoICcSe67bvgNSq+bWyDx0VCxbIfoj6fWiHWigtFCs2W9P6
Wpmmj3Sq2XzqJ5EVu+yvpIpiB76bvOgkKjDrcH1E3zJSndDZaPx+vFh49FxaKWdqKhCW0lNiKlSQ
RZQITXu6NZB1IH7OBwsGtVqxthOIvF+um/Z5rTA6ztcJj5zAle2HZyeh1kGu6gqMPQFAkkOBYagc
ocOpnz37rRioylEIcrqvh77u63eH4jk+ZI9XwBgKQj5RWBYtL/6FafKvq0YaPqi1p3pvHWPeriQ0
qh98bhSgE/JTtXMnixP618fwT8UrlZx/n7h3MHHSSU5Eyv/5I+ViMeneny/6PLkrzYuqudY97MYc
vX/HK9sBbTp9CBQ92BeNyR5TFDx3Ehlw1KGi5UotCTPMXD6dth3PLvUb6B7d/Xed0b0vkR/po3So
vldzdSlTkdbpIP+bB0pEibdldIWIJfXEozFisVOOr1ojsp6hv+wyGXezXbx1uXHKHB9Pyc/u2wej
BTYvaHa6EnCeEpDnR5d92YvJ23BXZCF3xiHZqNkhjELeB6PNEDmDWlBw1yshsX8ZoUnvRBkJpvfM
1+SfRhpPSKmiwlnJjUZH9dPm5uLOtARygCwNXaFQlwQJMyO3qgUpTLuzY07KtHBVJt39M8VtS8EQ
XnHAGMPOEo32sgWxJeCvftLIa6hIBlxWkGr9i8rXkpe42hfLx0WIm7OPkjR5zvommsSnUZ1BAPnx
JHvtfVzEyaKuHEZYyRKjC0zbl04gs284VF80gH1MuxU9E6+yDncBDHLhLIjmgMs5J+zKYLJZQkgE
4NZvbWLgxkUsPh5vwjValPCLi5D5Rv6pBFi66d9w9vMY+cPGhYNoW75R8274LNW5OBqH8/7FF1cY
kMCDwZVeCVIxnIGtmP+oTE4c0GRtlo2Nxl5BBQ1KCf931O8S7s1SfldbeuGG133FT09rjT4FozJe
Hdm3A2c/5Uh3jDfXKCVnaSUisuISXEbIRbeXLbv2HekGbkOf/383bU9cHEt5vJIIjA5yq4Q1Jhjj
JwnhJepSusAIY5cezw8J/qA1YOZr346Pe6As5nVrGXgYEuE/Bc+n8zb8iyaw8TPMU1tnU8aY6BpX
4/vwAT7fC3/y1Hf8ihdNiy2/CX5rUo4h4c7JKsAkVjTQMbWjGih4EOtuEuokZPNNwc4Y35tDKxiK
BYqv8XU/eNpdJKqPneOSwnqgSotb4/k0ia4QfqTNpExmz905xGMblpk1InSPhKmwBQt3NNhwx11j
2eEj62MFy2vHDOQKSv4Mesyj8t+czwlrp93tTllOL19zqbsgru8v3ppm0uACCJBn1TUVzDVajyvc
Icyiv4b0gzAXU7RsQ5qy/9v+YQG+ig76WHvhrIUEvnkQ0PAeWYNqwGaqkgLx/T8mH3JbCWQDL7T1
N0DcJYxQE00bvHRAT8ay9Mkw5FPnkd3V7pQK5DAvMM1WHJawqAG1WahyPPQzm58gYJibx8u7enCX
tApt2miNyrDrJox7DBSfwZMXXe2iEfhLnnyNAATYj/spxv4v+71E/E2p3UE/xNo//1DVrI9ZC8rb
lYDNjmS2XPENOqTBOmYj09s7zYIotMDWXjn78PG4OYCSwVGdde5cSZwd2FnRTz/b8FXVe+3A3d6U
oksiBIlxmFjpxi/FwLXrr1UBfu79laM4jnGxilSHzZEdazrjxUMCXL6n/mrS/dwCVPu0co6cFWfi
56xPN6M76l147Y1uVxoSd4OcxeoE6mQfoPQgfGBymgF+l+xevaHa9YCUfDdFoTIdIVqOoXF552A9
KUiMBGb8oRrExuFaVjmj70MsY90U/BX4FEy0ccPQ/Mz02xktPWT+YPzxWfiawIRBCQJdYCxP0X3r
ikzxYeHCg6aZznX8vUbtqUxJXPp+O4yzFajow6AwNr9FoDudytCeWvHihNFaFIOcqybIyTCA01r6
wlSnXUSUEaFnwIkXT9OWcd3N9VxEWQYY0yqV3jpPv0QLOPOzeGDFHhnf/TGmA0nmU+Mp/wIJR+We
tt5NH/LccYcL3yklBjVYTkRly7+lI7By4x2TBjLsI56cn9HdRQPge9lk8j2k3J67D6jZsoHHzMxm
7o/b4ag7GQeMIwV7muk0S/kzbPiGF59rrr19F+XEN1HDYtRgDbMyiZpAFhmESApHyGP6cxyp7PrS
+H+XkVU/8fYKLCmQk1fN8alVMOcWhIBfEyVEgtHbxt/g0lViVADaBpqqBRy3dG4dfdgDL1CnRwhv
lKUR2bDiHQvH3A04++So81lk3ICsEH6xzFaWBScu/vvFlgFs0g/phiNVXu+9HHcGpP1dOLCpnPff
KTBn1yrZMXUxlwO6x23uMwm2gvJpDsB+3boiQ0dpJf55TJr/aga1nXtf3hY0SPf7wbuSjyNLEBlM
z7VF7On4EIc5dmejF3yhad5k9DoXhKsAY03rYmZntxG9BfSp+FEGriRhjGugT7IT7Ob7JA6DE4pF
iFJOZdEF+LjuapqmDMBm9fmWPpebwFcnjCDtM600D/aU6NylJPdGFUgH197ULfK/0EM36Gv4+GsT
DzB1xt62nviu79UzKshhGUD47faBJfXzzMWGtQ64QMKKNWNz7s/arDTMCejxFu+8rKsWQWRciDmO
DJ8ic6BzhEvh00Moqdlcz97Tk9OCL3iq0EOcyeBXRKUlHj6aU3NVnWhGepBhK6XR0r2yQv8WvIgY
Fkb0UF6Z4D+94uL/ZScEC5LaafHrOJUewChVTA66Sp8p63ktY1hIplPAEQwj0N46/Y6biule1urz
o0TFq7pXJMbC2WOClYTBUAw7tAJWn613iCe3DSyFVBWuKP5CBuxTgaMkJ91inHsEVV6/6qqN/YPA
+nxzZ/ATOPjiQ2XBptvaZiBNT5zdubjKFSiqjmN+AXpyNTH1xo7s8SpFVElQSFp9sCcxjmu/fN1W
AyvVxBWVJJD+kOkmAgfo7sYKed5j/vlHqezM0ElsHInTJTsK4hY/kV6xg8Mnajfjih8UQjzSeOJm
DLR9zRCDioKed93x8FywA7w43tVDQGLh8XEfMyOAi34f6SSo5VdOh8zaiMAlAdOG81S/6iE8Pvxg
ev+ByCLPn2OzvwlUshhwuUQoPHPHEzwSYKSHZDANA9vInEssnNpCpgXqgjt3jqoV5sUSNlBN994h
+4A+ikW8P7jui52Dv44YcuQs3FsUK+8MzMC6U3JqaGBaC4Z2ipHGQY+VXcJhKatHUDjWdxON4kCk
z+IThe94CRufFab5LUktr11u/eivmsvSv5FshQXj6sOMtntmJ/ALokaoUCKUbA2hMfbpup5ntl3l
30uqfNqqbj0/EJmYM9Q+Y4+vD/rth5xqc6cbD4Q52FwHYVWcd5PspFK/kxTCvCJXiYySbRUjLtiX
U7VvCxd1/MTOBsCfv6h4iFkLAzoCMkF8OYmzP6DZGbCto+h/HXwC8V3zL6laYnDnhzvHizV0PCf+
/FK4g0alCEClcZI/FlqZfnAyW8c9sAkpvKGwMv5yD9G29dOhQXFh73hAA7Nwm5qpxgNlni7WfuLH
veb7POzRi0UxrikiD3NTW70VH8/p8HCpJdbYdpGcYGbREU3baD+HZVzBpbTv4UCpuEfZoKNLfxyM
QB56jzvKxhp5ilKIJwmP09aC2idz3e8t9EVwDZlul8KxX/LeIfRzLHhqDp9jY7V+47+cmyhEntM7
MUKzzu6DrpttOAB4vhn6yJ63MxqSYzYJ6SrxZXiz7xqcaLoKuM0ZL0JYMurp7IpxqEopQSvWPbfG
d3rXUWIsTMg6dU2zNLw/ppiKnH69Z05oI2emqv2FyYZ3jBs2+gcEntUMOB/Y5RtNaOQUK+8q8aa+
XDkdKHjHfM9w1fHM1k/xa/BVeFi0a+K38sKYJAfC2dNPuzg1v+oZfExxL5qhFwmKlHi1W0kWxuWV
4w5GaiG9pCSFfrKQNTCb/1+EwEi4JspyUf5sWsjHbbwNmfZwe0Af88nFHRvHDS95FHIGv/Wthkxl
f1w/VZBaxxhtwSfQKO1Qo2/xAPF62PcN8TFomTY/rzt3nbnXrKnHMYAndM5lXGjUHCvwyB0ygn7x
sJM5p52/EZUfDwVu9LvHZWbaRYLVeehYzJVrx4EhnK13aj87zTZeEldT6RJBuDNMi6VYTNDAeiBQ
ZncoehE0BwkLBbLsVURyp0909QRkKhwY4wewjNzDLS51KePvRoRpR4LWK+OcTWEQFZ6Ln2eGggRV
ij0UqfN21p1jPyUWW5flCni4Lahq07nL6GxuvpmuAWcyXaIWyY57a4euihSCuJXFwmMRVBPTFuus
MPEQD3waIrHR0fEs4GFBrMtqtdMzRJedT9wNq6+Tm/6AELYNXGkpWmyzrUfmBZspMycP0NajcvSG
uz6uD0r+5BP6yq0N3iKLrn5AZQx0FgaYqMzXb4lQu8XJMWs4xdKIZwE5jsh6YBsFqaf+5SbRbYNm
1+IywnwwKCQxm9AOP6RaGOvgXWZf1CyUt/BlD4O3dmUw0EsKQlwCROgi2Dt9jVOzzzDrq36eKNmA
/CK3PfiPKhI4EQ9myg13JC95rS8ShpuhihOWc4ziv3p1wBKb3pea5dNOuTHfMsVeEjVZKx8m/tU8
31LrVcc5lXfOjibZDIiFm4/5xrjI/lbpjpjXNU3rPqKxPo0pFIlXUI1UR9Gz7uCxuL9K1tL+uRPZ
C2VcEGUF0XuLKMoNYeULXVzPnXRPWUwbxctxMLaW5t7ITcIU0vC2e/C4vL7Wb94m4wmhVZ82k8a1
lqqRyISFbNw3tNmXY1IftZ0QlcKbVbS7ZcR4SkvUIYRNONkGqr6cIlTUV+zMzRJo9b2ZdVh1hETG
z6xy1ItF/ozmojGTZIwaFbCKqjsetScT9a43yyvIx5WkAWyvBjbDvDYkPua3p3vqL+bvLLGKAPQe
1Pmwh/J7ZcTs18LvdLfIdIor9nEj1Y8c9mltUJqmlapSAhyuZoj3A8wkYczSQTvQLk8sa3+4tX7z
TqBIX/aywp2gToWYa3XtrXmBq8/fZM8AtwFljn1pgtXxkAk9ihINDpQY+AqQvnSU/JvJ13gKHh5B
qr/SAOVI8glo1rCp5qZSEh0kaCysdeXPoeGE+IK0FnnRBSCtKSABI2RQjAVBBgomBvZJ73o8AYwa
IKvvPqNvHzwq6DNTCXv3vA5vSSAM4AsCcJip3v0fCawBdgvc7BX70IUH58RoUyIa8HhUA0wU+aTv
toIyLA/19Rhb8e++XqvWiOmpJ/Tn6wtN6PVfGFDjxmq0bT2D89GbIGqlC9zDvwconzDCHHu/QUAT
mz/bQbs45+35vcYKiK7fcEneYKD7q5W5Tm1W8HdMmiWsjV4XIzTc2VrpFJhxPySv+QpxH/FDarJZ
XBCuVqSyNFD93ylTdBAI/7fT2fr8AAgB5fA0gYr1F3l3Xo25jumoCVFbqrYJs1F8892zAnYk2iCx
KPD1Xyz3WX7EGDwqC0UAy5v60by4dlVnl8IxY4oqXJ3vtTGVZ5NWyxLa6mckLDmv+nESrWReZzyX
qxmfc/CcNPCKpW0pLRmKbHkdTujIV94JFDDPz5MBkODN0R2XiBv8U+RV7F2Jdg5JeKGoDmaEY4p0
BWvH5NcFHHY+ENqY8z+mXUzT1RImg6faQM73ar8VnF4Ap5j20B5JzzGIlH9/q/C8mp+SBS0pDPOh
xXDWbzxixgyerkjuGdCL0opkTMxoFkS6dd79DfKoqvgcMN/s+FiK0iISYXgkBdy0dK2KLKF08L1y
i+rzLHcbwSiib0JvPdPZB+RdQYpVjqfMGLMkfBdHhQ/YcB2KpCjZqusiCkkPtc47UK+s9YAE8YxC
U94doZwPdrDFTp7atFsFPC0MOpDosepUNwi9qRXCY9w+sQQ8a+pJhuBCuzs+yWrury28mi6IMjTL
Orc438b34MFbwpRA5oGIDVEIFDKTXA+Gul7gb0t11XY4yeq2PXeDk01T3bRFzMGytmQ9VOeBbh/5
GLSQjKS15H6O/B2SIgTrzA0yOgUn2ATtjJM3Iiy5s2YeP4sDZk171jcigw06sCNaJxYQYgyKlBzC
RMTEJilVZZnIg4csTVaS7B9nMWCQlR5UnZfII4OLfS8KYHiOGTvFd00P4VXQcFvCxaEjVhEHPD/W
WXjgrbt01pLmZ5rCnKtrldWmGIvKhQeLI6DMO83U5w7TsWYBQP0hu16WnzjAAo3DE229rYfruDyk
Tf3/AEokHxBcn59YBMPLk+UOeuoXGR4EgKockMUFRDshalYW9E1evqC8ctx/vy/acRKrBqvqOl2j
gAKK0vzGgwz1p9gnbI719dlGGN9pd6G1K+A57Xm75JajeuODvyWCBC5us70vzpGahoONyKmSBf1L
OsCsfPvfvuoDsUneyCRT9po+sFam8n5pLHcibgi87pcTNN3W36sRiB1dpFeTAN1F8z3LD606B7Ob
m04tjPbXdoi/Oup9iZsqUpBAAbrCvheCV7+5yw8E9DKYUWcVzJyJH0xUi+siFZvY5TsH3JPvsbi3
kAbbnTSu1S0HjzAQw5J8c+a+/BJ0YhsCSJEbuBXgteQ91q42KfxhhakoY/ng75UdSpUtWDGEk8Kq
qVE/NGgOVxJsnvWGceT1osT8Z6o7LfQe3Pyqe217CiKOiDadPz30IHTG6/gSFwLRYHyJmARd6nPo
+tG2wSkKwFWm2n7tGdPnyOrhcKSRgh6UGIrW5GFIBywJlv97BdLRfL9ZXsQkG+MQzxneedRGJ252
D/ezzZtffKLF7HVYqD30l+YmK1oo+9TtVpvACX1nf5mlZy92yo5O2lriSiihGgASi9YHBHd0m78q
p5gqgSMkUOtPtQi1srCzYEslf1/RIIDjhfUGvalaR6r62MEFlsj9DcFdqU8Iszh1dgAfXPTXeKF2
0B7xydWxKo8ayKXtl3au6mfu99JWQurRxlBSybW5Agaek2nXpQfhnsSGZUjEyTiQUJ4CdsexYQK3
iX5F/xtpk9VFTqmlQ6Z/NKKotZIAetWf9wcfKHM+7rL4tVh65nBoFr6YeQWSZ/P7GY1w4i9Ds2Tc
FrbfVj6O3YL0eUMMA1vXdE/GvUBv2k8HuDSS/BpuKJxq3YkIImoSEBR8tNFMpJTc29vt5MCJY2K4
PNhHXiycDlgPLTms99Z0RmJaLyg2VaYemIG7CPW/ydoGgBPXr2EicShKarNYhj4K8dpthYJbM3cm
LkoTik4tgxHErrspR7dfp2EjHHmXN7RcvM7MDTbFTyugb9eozMy7cNduA7+VGodYcLufs8UfJkoI
CpkIDTku7oHJGDYkI9dZwy1rs7InuDuvdm/FTLMWijbwiazZHmY36rIpRDYLWcfAEYA7hm64IpMt
u35oFAOwuWW1OaEgH4BlDH+YM5JOJkMJml6X1lwnMcWmW5CUQDx/sFor8qmgRPoApvjQAfHz108n
KHXxJHPhLaoVqxO1+FpAhDelZ0SHkOwkosOEp//fZktOhrum+DGFeHUjr0dqWZY6XOeGqOfvXHLQ
DO2VAGT0vFUPc+nkL3wm+lXf4qzWp/cX5LgTPwxwfLhwc15/NuJEhZseQlhgx8JMwjYrtrMVcMmV
T7RizS9Ox8028h/1QNc5LIeHtTDvK2H1aOK6tMvv4i+Qxm/f/7PCYsvG7tTGlsC0uGFLLSLenz/h
LOar/u9KeXR6ZPc6v6YevlDP9ptWSGE1Ep1/04NUjh0Uzo8WiFmLvlau3bOIaNXazo9A65EP692L
uG1mLHwnrg85lpgS6OaKs6zB3xy3B5Xi5UEpmSoPRVvxJr1fYVM+ZBl5QujL5w1gMW57W1OkkCCg
bWq/LlFDGTO9sfmf4WWAd7M+pHlIleY7fyYljFiLY9Cvj0FYA8Ef+UwkDzcwxdw3/yM2E2MzeQgf
gQnVqLaHCIqhQCr22DPnvl7ph2RqkTU4+euKqulwe5NqCcuAAO4kUvK+7m0zB9JVRywLSxQ7ZyPq
6P95/g/NitESpA6BJ3D/OoyfLuPKnTzmQpP2eJA0LWrTGs9hCecIa4NPEQs9j4+fo1pZB3xSTALZ
H+pMlwxcbSVjn4fUIz6F3VJ+f42J+sZyv1SH881WIJrsCzjEtZZxQkT0ZlI38zQlZeRlFHKEDx65
0KXRKjcpVjSA+46lpIZBiQOszvgB6RX0+JM8Tb6vhEyMLlHHtGKyLVDqPgGl0Uensv6DY3ULCJ7P
T+4LRhSbQnZ8pPNTu57bt/Jo2EPpnJ5jGJCOi9YIK4zLkvcujkH6MNoXbC8zM5bdJjtjMFJDjSko
mDY2M/fZbjYkd5G9u52KVU5dmkCV/eropppFOlBEUWTIa26RVuDPA888lJm/n0qIQftXA+XdAEXy
0GL9uzfQyJV/KMKtnDh3yTLG3w/At+IhDshrOSR7NYQ9fDG81NA7l0Oturi/ql3Z+Grb9XSI0KmE
DyvKyvejkNln6UVOZMrGBhHKryxdckdlDsqL4KmJ2xxBWtRBnrbbJZinbZ0/DqK1nkun7hTlrA65
dRDXfgyFM2vGsBPYlJCmBUhepyo/aqQbQl4u5satMwgtmiVvvJ/ZlW+Vrhn4YhmEbUpJuYsS/04+
0qH0J+/M/ESjE5L6s8mUFa0Q1fSGF0Nn33gKtFiL0nQP5SdJkO+HZcNfiZkXIrqRAWbE3BzAHamS
GhK/lhrcNVArR4UvrMwNS10xMqfVNmn1Zhz8be1j0R9StrVSFpizSey8EBkFgQHDPlvXlYtegHet
0krAL+kxGNuyRiRq320cD2WxxYPkn6LqUYGcvadlFk+WHHl0J2/upcWPnV1EIMAyMMtym+VFZdkx
VDKQ6nNYf/zFhpOoFoOtqyaihZEO4QNvicPXtFhmSpq9L/JZVVVN8e6vfLLD44Zoe0De4FGgElGe
SZggt1NbXUzMqK5DQ3Uevlt5kfiV3IKvOdzkBpwMa3W0VVt5lx/FRidA+TyfgXI2hU4Ai+lKP01L
8BGlDGRWuRk9VAPwqna2fiEyb5ZnyD3Wwwc8EqkSOTiaYdMWZzFWJteMUFBES+UX+HAWtA997MYJ
1HMlOGENgn/lryvlqcXhFIta2drZxMpV6IjvinpJinVQMnGPPcAR9/CZltrXNrkgmimk5aiXl9kI
Y7FmTjM+L94ZQcOecioqKh3VcFO1RZth1L423/VPcvYz6s1lx6qbUIJFN7akXjMR1aeKLX3uXheD
ogOmmoj7cv6WAryRYhEHwYIWGILRzstA56/kBtUe81JVP99FrI1Bv6Y8Gn09j+fbPGfbJ3zhLz7p
ii69TZVnvoBVV5a9n9ziJVXzd/3rbNI8O1AGcBVEjoKa6Vqmpg26ofmFffgZ8LTIiHGXNQwYydtb
fQZVJdiplDgPay3W8C65UKNnYmA2ueHHWz9kkFZLDmeLHW61aVYTFRht9DV7TLBKE9diCfS0axYT
vUzaaXJGbTpu3KzFTkobrqvOfjGG/u1RvIffwAuvbAEyfsIZt08cvDq1AXefA3QqKqlFBKtB3Jw9
UPkZM5Ut08QR1Ej+wovQtsU1qRPtLFxPhacWnEqX/yK7oxTPoxmbtlR7NblM4XX8shdzfIlhoCjS
pppbN1u6ZtdM40MY+3yYCt29AQgnYJlnNs7egJbL2gslF/yLu5CvIP6g56pAQTwcM63e8X9yjEDB
2OX0kxeL3RPlVnbhYbHlfXFAwy12rbdDjYxgQ5QwGKMCKLVXsOLJaN8hhkBpi8rOBcP63HrDewIA
1ym4Z5ioveJxiq9rfr9zP0WzeclI/xjCn7yFDTqOT5h5skMzOIIs5SlaDAMA5RmkIHEu7aBhx5rM
e8T1UJdfKeAZDvRxm2QhqP5X34OpEoIZWfsgyaAuBrbbwoKiGS30SAqpCB+ayFg2SgpuA65lj/t7
RpwVPFO5raSBY5StkwefstECgyxk+4gEnicdRPBpujLA9xQFLSYAF04whmfdjNySu+P/fyyNLA3f
uUptIFu2jDSghxH7vEeLzt0QFsu22lguum2EGlmufi8J6JMmItpYmMx8D7g01JnOks9IL7uYVNYg
erj1+rcDbswjNDbXKlVnKFf2Ks9b/fvBXSQFQ0jH5G23G6ZP25t+8KJ3DPJZDXV10yCcGC+ApoTS
HFGL1Pgi0BN8pQRSiLR3qgigVWZQQGxi0Vk13ccZbPatOiq17zg9QC8rlvu+uPl6qqr2TMXVHm85
KJR82IK7cJj8NtZP4SQdZuYVaxHnPeibrxnbLTvE02r9m3SlA+9AKoHXASe/6X3DyKge6t9hax/n
bX4BRLaB3xYZKVMCGQSR9m2vsEMrx+bOdRM/FFREvXRZvLmDXSLfSwS4+ZWWY7XzoMLk70+K/4DZ
xkMjmo1bR1F7nvQWR0FXKpXeREvEKqGJPyJXAhhLUbk5TQ2QUmXJ0N4nZBotL1bjLdQaNK7tCC0z
RRca/xdfFHWW83zAGxdNatit+VzCwOxiKTjDIYeKmePcxo+keRxjnT6j1VB5GwE8+a/jilx9SRWi
5S4srcyHYrBt6Q5F/YhaMHxopHovGeKKfWfYbqmuHfLJ2uUciijNekY5LZjHmvecpg/cb0BFWDUH
hAr6uJladWIkLj3Z137G76mdfiSYoCj2ZoipH1NvFQLlsp+G/A0mtlTbQokvUUGXmvXZK9NY9MGu
g3COrtrHhdveW0n6R9IRlcJGDyg7cqGnL6uJKBBh7S/8asRqZ/ZWNcW8N7RsbuxhdX+iVCOlLAYD
pP66klL88du2MBQE8zrz7xINW4zJ0K2RVNPkoZy7fk2zSus4WVZXYLYCle5QlrbWEFgUifPtNo9k
1+hK6kxmQ0JTVc+poncjmrymTdsrxD4l4imsg2Y7biy+TTw1MSpTCiv1uaH3j+nO4M8nAnIZDIqg
8hjslHjFiedE7WSI9kckV1S0QtDEYWsd2Ev9xLYpzJy4+5sn8XNaxaKuPVeOHdEu9DZagnE+TRPu
mDu4+kg1kcZlEgd7ZD/YzKykdQQNLy+mTqGyEj3bwfkT85rMNmJIC/fKnnzXaK6DP0OU9HL0Hek1
0tQvu6cWnsft1utrK6AZ1sjjNkH5bu4rfr4d6tzi2feWkK5vzDMD83bdBoX8212alqPFx0q1LHVb
JvzkjLKfntcz6JxCJdj/sF2ttsqc9fGeQCMWYxSPX7CUC/YikHuBzyjrX0+hRvKZoF3t6B+phjyH
Mv34rg7ayJTJdvqsv//xF+suWbjhQQl0zg+wOAw08HBgHplK9no+TtbOfSLIs88GVToJyU1re5Rk
b+hgCbfH4gF/NNYdCzmmxksJgs4+4CxP0FzxLWPM9vvqMFJoiaYovuXKPByvmFcDsGL+1G2EelIi
zzOp2aKTgfZ7yayDeaoGXJLSfnrvjqw/YxVilal0rByShgvb6NjER5VXTO6qrmonYYvpREk++6xk
41lvm1sWpBSfiS4hlJjxNADtu82nw4OJ/5/dMGYA9EQ9qwW/H3MExKJx12x8wHAYev8u7Xcbwwo/
imVP8V/N1ygFVQ3lXrqBvfLBI0FdKbypUmWhaJBesmX8RGK7eOmcRy+mx5T8AUQeMYkGw0twZ/LB
NCAqDbBhsCznOzEKNJ2BvQXV6zmZK+wxMgLwNae9LLTobR+z9LjDcwip/RLEXfeebmqyKzGnk7lL
YkiPo2dH00c/51AdrwlmB2ZDEXtdELdW6WOI4kercz43DzUiXCp5xnJ38bHIwLXVHJwvbWL9lHTL
L7CkVc75quogwMHd89rXt2Y578odKIbhEyzJtsE1kwOhBUcRKX8duFW6Lei3a18k2FHoUfblPpQ5
rNQ1DeufMzc0LbWcwm3FmaUzMoJ/ajtuWZPJ9yvU4es0003nlcnCAnOO6VxRAi8WCrcgY2sdSF1q
cULqLdCcLnbUI0plJxi9ttUY4u+iyjgwwPEobkwHvsH6Rk+/wIyjMZmiud4DbtaaBnECuPdZeJUj
qJ4f6I8/S0CQOUf0T01XYYUap2iUEEqjtFrbZoFAPEBjAzl0MLufoDYb3ARC/eJH2L0ATPPv0ZKx
iy8E81yUlIAaKsGwCFD9aVdPGh+VH9vhEUJl7hozMOXAt6QLUXovk5+wtbNCNBAXYlPVaM7fAiSi
g0tRvRLJsPs/VqvsuapcKJwCf3djl257Qbk+XCYyM8yvF6VcZanCgMHy7fsZJ52i9WeuR7HWoN9M
6StjHvnJdI1ddQwwq062/2R9ooJiuXtJ4TxIaZFpuG/R/6taJvXLZbZBy0XDykBxLo73GKc0NKfu
+GVQuS8Yvx/LJaor1YWE5hPz0VRhirhhevQd57oG01PIklZZTke5QYRL4+mOGGimI7QG+98DKk0i
zpkVBu4MtG2gQfglQEodbjWqZVDa3nVz9dP1hhBL7vGzWk7EZvvAUqkrRKNgV3XJ92ag65Y0gxGA
uhLVt/Z54kwrBGPPaT96BKSgLuMEG1CSFyIW7imZOu46k0bwFGw/7EYckR/0Va7aAJ9PxH4Vy/y+
BwzbCl8M9kLFh4Ya7vYR/y1xUviQ2Vq7MtimR9xuYFLFmFA1PJVoJexSf357yoChqjJB7wRc6CP4
4bSpcdQbB1WyWZWOWGI2ChpmUl8duD8yaRK/46u1/VE3ePli6McEsxna594uitQT0V3Tk7Hqlypn
6ZkDZoAnfqxGB6yvwt1IGb4CmMXmgC7ZX4VKn5TRJ4D8P+w6c2am3454vJ73hyirTK8e+RjLP/Ob
tuW6VOSd792sw0bXYNnI8+hu2x+vjIiOhmcM72QtjC96Oauzz/c0Qn7K0LCNtKGUnx5X50e1qk36
dW7IEeflCHrlh29WJ1b2z4vpHEqBKxl7hM7FzZyKswty+Hjyqczn58btn3/WFBHZrq8DF1jB5kRV
9MAEyytMX0ubyIQMYu3OvDoWHzXKhang+OafSrqTMshOGGxcE4PYO1XLAQ+bwuCvjDNMIs1yP43L
XkmoZSU+8aGCEHv4wJs0U7tqV3Qm8F/s9rC2DDeMwpSFBE41HM/h7Qv7nd7vZyd/+2WJkvP+2o3d
VhbCXlV562PR/9YPzYvwf74WhM585iMQabHy7m+CqzQ6Tr42JyCpmfOAVzGs/tjtrqadnFJXiNzA
9z7IuWvHoAk7as/KvIuTgczMktcXP2Xn74LUBnK+v0PGOl1I41bZxBCwBgFL6P6w4YOlQFdpq0od
lhICnuKRc4T0hbnvLpdy2zmD5b5u14EcN3I2uH/SfyvXrZ7FaImI8HrZ/M/NaCecEdo6XrfnYJNg
tF8vSzwEfY9eZKuBJVpbjepEfKNj7peX58k7d+bf5894TjqKAzsFxHvy/vwSeoDN2xj5s0qLarAW
qSA1msAZnAab0fkOi3h/A+l3C0yymbL3WLMMoO9lhBK3wVUJhoC80sz1u9sjkPkxiocn0E9XMm+u
NlW9tdBfcMRqGB06PAa1aCt6Ix4lkL45YE3nI3qpxJkjt5oYu01rhRHCRzne+zRP2TW3bkoWmKf6
XLo4qkuoajfFE+/3GgwZVTrYYUsFTlaZEr9mzH/M6ClsNcTN9x9Jl5xiSSgs3h88pEolzX6+24vC
o7ALyevvZ0JaFVpU3toVrbbjD0rzRRBRI4ghdiEznnAGiTFBa44jdLz0xNA2wx9ZPK5lyr0XcGwi
pTu+LsmCOw9Qe+A1HZerSIVt6yozORBSAXoZmwdGNdfll4pkkgtzcwhFmuTVuYbK+SWuYoSg/hIY
WCYdTshcdpofL6n3cvxYrFykcDQwDDWZ7ZDyRICGcBZTaGMT+MtbVYkQ7zgXVMcldRs0cawfPR8h
G5HttyL1/YD2zxj8u8spup4UdiARynejXGjY5gHiKml2oqD79xk3eHBB8tpNsVwflaoL6yTkdFqe
y8dqt8ZNc/3873IU4ey4yfyDHWAy1EFDZDduJgd8qtyZFROa0M5owapDD9XpvDAxMaX4+i3nlM3V
JASFFDtMBLqBCH4TACp+LLmfv6WGBozWRTBDfMYPg54idBeowj88QSNsmqFGx/7k2dYj/lAuMNMI
JrR1GB0mjd2UqHpn22l045UCMRQ2J0oeFfOEKpUqdUblDI0/R4ti5cL+DEDq6dUSXzF51NVr6Nq4
Ke0NSC3mHLXyrhFq5rQD3jp6VapngRIUhQPuru35YXhdwEdcac+fwXnb4obM2oKEWVUr/W1cUpr6
8Xea5CCeSIC3F1X8JZQw0Qprs8z/BFzs2Mk9TqrLXLQXJJ9LMqKly2qty5k7dJKPSxjZ2fRTIPe7
p1vhkA84cbtPD21zcWWsTtaKKtFPp9FhGvyQ9vZ15W+SSFb0wpMr0LoB9CXpRv57nT/Qp7qjpMBr
A6Dw4zV72xJpzfF6l3XlhhgZk8Yj8GVF0is3DobzUmIJauKI5bAby3bJlKBHsb+Eg8x3dH8sNOhl
TeZ856xVEiOL3lLVZ+AJ3C33SeUkffzDPucH9jzydrGEchl5yqJ2apr5qcnePR2A86+ZH3Sw6GXz
PY0GK+9ydE6UW9KUw1sYjmd66QYDc3KWGrbzH7rBuDdL7zb9S00aT2c1CPxv08PX6D4tspfVhKRD
1al7hNPf7S4Cm024JU2HlpvtYgxEypxIuIIonLMFmf2PSdslSMgr/dgUjppkHiiRvt2CC2Rl1tM1
jCYjuzhemcYM08bG2+5Ti3/g3sTDTXdjzKhem2WdeRhTY98AApIzDPveQbYG6alMbcuBMRLZ0yR0
vfvDaRUnbkHqLOZ9wzLcmrhrf1QsLQwXL0iDCoK3scJWpYvbXrISv38euuMgaOxoHyI+RHrmkWnO
17/jS+0ZaHobOWlAiPbD4qt/lBV+sm5wyZAetykoJy5Lg/JRncErXbRgirihGRNYQOB8SlibTwwf
RiBnUm/HYDF5CHzQ7ruq8hK3QUHjFDDwBiSpJmaUcktGfub2giaYsSFO3KLc+UmLmJyn6b6EUKio
6Sr5ELNi+ny/+T+BgyWYQbsTsXpm99rwhIJUwvCb4lOuQmrprSxUmRhJq1xo9sGGjR2CnPn6kmW1
ZYpeor8ajRszouL0Si2AMICfl9AU1XfMWg9pn7F+VOMVX+yXY2Z6WvwLmhgeXuf33VamC2Kcv6/N
sf25L2TGRavSHEVCBD/vml33aTfA9aVKgXLr7yIH5TQi3nK71OGAVO0eWMGbKpRtZt/+LazMAbcW
8PouroJuatoOojLu7devVFnGthpEDaKCuL1Mwb141Hgs302NRY0z8kNqdKXreYZcX3ZQ7JufoM9t
+Popx0yLVicLYsQdTXB1CJZ3FfANxl8WTNZ00+Y98tQqkzx7Wgtv+C/DxpLFXkE6Hx0OAbcpQStH
OBEMLlGm4rYky54iNgAqAk4xK3n/rm8nafHa5NXPJTzfGPJlKssfx6l1AFhZu709w+/iqhOlPC8p
0cEFboZA9bX37+fOkTgPcyUYWh5RAr7HWwdMA/5mTvD4LwU2GRfFqQLtIZGUZkOdQnV6N2xNn9sc
f1CWL6MNHAABCtyaI8ECjXmVx5uBjyrMFrwlqVASeDfUPelIYrc6oMzjJzC8Cu9nNnJeUi3O1Qgm
lVdA5utAbUKE2kCNozoSStAiYFZklAep3TaO+S02AQRoKMEZLwX4o44raBhBClKmy9UCw4rAsUH8
9hrMqUOU81ub/VdY36ZDWItQIWwDK0TxJ+0kwio0xFK05qPAzI53RqKqAXKE5wZMTWOA6asdvuet
DEjJmu6/IG2dpYfeHH9AAYYbpl1cf2zX2stiG77+9MIqYNl+z42n3y0kvQEzMvANgUhjZ8SSIthq
uvN8erN8t9T2w9IfitUAVKiw2CUI5vsdRUqw9WuTdaPC3jH1LqLpfJcmK/ZMYuk/HQ8HtFP6HkGi
iys5ULwZmtLXqfqYks3/WWazKaTmSISXE5JBtaNEcp8NooZW+00IYabKC09LYc/LZcXm9QHNzlIw
WvTsgDMCXordt4BvG8Ykp+ypPSck7toMtk9TMCbMgrMSAD3r99jFXmkx2ZwjqgKI0+avvafADWlw
UiOsqH7jJPpH8sISVpg+hTOXu0j/8Qui/6L2oOu00F521tYlULqYkuviqZ9eUnwgGEn0Tjzz3LjS
ue/+ngv4lyKt6J1/QNlsjdtj9Zue77U6nF/+pNQ8eMkFfsPSme0S/hanKOe6FBIfUCDm7eM2aKo/
sQGnkJaMJpC0v2mV9rem3L+xa3GbCDXv2QxuLuA8O9ywkCNnPmgBmswMEmA05iy+FX8VrDWzJRpM
W/Y2ASGirY23y0E+DYEgrHLRdPoqmKK2oaU+BUpzxYBwGPNvgf3BQOdRDnjXrCgmIAME7VOEgfT3
2Pr1PWycxJdzg4oL5fBFBE5J79d660/bnl/oSOfs+8FvbKBis5F+/id3pFjsSrCnH1w6J9Xe+UmZ
iqo9UgLJRPLELhVZNHe2k/SEf7o3DmRPWdIb5YIu8TnRk7Yi7ZIenR8ilc+9muJzv8go2q12GR+c
opr7p4w/q3fVodJoSlqlaZpxknmxuJbx/N0WHkw7Zwq6dxLHKgC7VFs7lsSVClyc2mPYYwKyXL36
R43Vc7QtcGbCoKnlVn3MdMz+coowG8/I51GFc/DR1vFpoXMplrataSnsON3LuPzBm93duzrp3RqM
hCs9R73BW0YNvLgm9359y8zx3ZEo2gycThSLQnFFt5pbwH2huGQ+Jo0TYVflLyfEQwaDTog+u1zM
54i2+WO/FY7GWSY03sZcADBtX7jNYXQ9SGsr3oBKG0kSQgsIR8XGkzuwz+JGI3p71SGoAwHzVNeP
qS5eWwkg2EryBi5NQIP3Hj3EiLgKEv9OCJhHXPOA7VVIpKGtr6TlbkHxJT3N2D2w+pT4bBU65y2m
64qSM9IyQ4yUklEkMpzwLWvquOUjK/cpbExss1PeXK0Bc8ejeE2GuxGmUWhYTbKxqj4J2Sn9w/4W
xlIAnMc23rwlpxt0CNdpUn9BMJY49o7rRiplm2oFzafdSWwEepre6GZtmjA3Cfl/6MkslygcZS2j
hJyesJ0vhZMujuXg1n1KJH9VdfdgPu6AD0XXwoqiHAPEe9HPJtM0392aljzUyKiBTe8IbjQakRwS
OoE3lINEvH73yhdz2zR4VUgDE20IjT0t2FEpbbxmFUWTqeELnvSlk1V+gzbnhU6HXynoRnQrZVSX
npEbEurXnky7dquzSliWl0sBGEIq87IHvhEduixjiRKRr7ndtFOromdqmq+k1pJOslMFJE56ZoGK
sBtM+WhGJjLP/fHMUhGnn7T0nc4UB53lu6hHAsbstUnoFggBzclVYH8WjOfKHKZyuHOSEWuWgiN5
FDh51s2Vl3kILjpflS6r1l/KeDaLt4etE9y+B+dL9K7ueVb1gp1N9ODUZuWnjm2CBs0VcL926fs/
8BxoFEKV2eZk72zj3xN2tXHsVI3yCTMl5VM7smDLLG83QxLwQsE6TjR5GnAXoI01T0413LW4WYRh
V56xhD4utkfT5vUG91pUp7HyPHIDwLLeQdijZ1ZSn1+/MhzuAFPpjLoQjY9sR+0m1Gwkj8Jg4Ua4
e0IgOIyjVrk1oJhRsLP/HwF7RS/BZscVJ5Su7M3kJ06u4FnTb+5lGFD8jagjVYHHJKmfy6UCIcV0
A2/fwvwgmFXkJLqxTx5bBWrXrxOMq16CMrpxA5gcc8uzvDyHAETcNc6TNGXkfR1udn6+MW+xXTTa
tRmoU4FkzZhOIpLuHTY0kYP5hmkS92q8dnbkzcIIPEQmGVvYxuWooFyMmdLCWFR21UwELqPcjKKP
sLRuhHH4JJnkH9muPpqw+lejxVb1KbqUrNNbjStqLllrwvaBO6NW3wWJV+T8rp2A6up0kejpmieM
aIxXaCrHxl/9U1yRAqpKi27urLnSVe/0mGuzlfQscHQd6+Q4VLiNp9DEY2ZSSJAr3Sha9Krx0vZ8
xH6FW6Fp31HIPfsOQ5OZMIvVHGO1WLFsymH3GTuOhT61I6MSIz7XXfsjfsWcxSBfFdBs4gkXZlIV
vETpC5EuDVkwdCAsSofBY8T/1yUJ9pGeiwMkXa8XoHgEMUAGWyBEEiR3pCnsydbOGobKK/LNY23z
Ffcb8PKQ2btNsWIUx7LunXUs1245hHB0Pvozj3SJSovohBEZA8UsQ1TS+0RgrGm91ORZE1cNH0qL
GXW37TQoF4D/O6rTFITz2JygFFrgn9IY/3eQf287ikw0Tk1uialW6hhl2RJgaZPgMD76Y6fA/9w/
FSapshM2Ohqk+/90YWZfmZ18Icy1rjN38KjFNmZkkh9mJ9O1K96uMLpqxSrCqwOb6GMf/SEWl8J+
6+oHqUvaPsIXu+kmYdBZHwWaD4G4eFeKnYElE3lyHePqMOjOh22OikJnxp3AXOjdL7iN7klNC85K
cb2AEw54h/5XG/hmnOu/POlaQSs7ocGYsp8X864Q6Nox8QjpcJPpXpApKODbtEMM0k32E4rU77UB
sQtMGOM0XN6qJr0K2Z8NA+6K7TsY90YFxgDYXydFMLG+zSFEHYVoMVy3Mjsrt9E5umpUo7//6X6o
wmQF3qmnj9cA+TZDh2sqbDVNfX4J15xtDIPXnZjKplWqXSc7yblLZ25nwjtGE6Bi2qmm0nbQN3Bu
EBiBXQiXgsj5g/lwf1FhT3SKCVTTP4lrThXqO0FIg8Kth3c4TaI7sCwRyquBNyVjBkka19pfooPb
5SuwiLbDa0zSpkPuqKT3cZ7FmT43A+Q9NGL1Wjk/O85WSsOdscVObAnVMsIbFyAV528M3MWiRwNa
U2zB31zVZYqicF60sXRo0QzadOwNsn6TgQlUepeLpzOe7youskPX/IPLF7Rx4J5AucRxHrBtWyVd
0VnFh8tjhq1v8NJ+0tKyS7p9vMvYFgHRytDvsOIR7V2qOEgPh+70i71Iw5i8ca295CKc2yoRXA+F
sbeQqgCwTmBymgrTp2kXIIty8+PKZE04/SJ9lbCxJiMKC/9JB7pqOJsHMyCarC5Y+J/aPaAemuGG
vaaaunOQZJTWU2JiRu+Vj7e3z2CA773oXmWxMXRXRBxSZ7N+qwlBHzCkor5oivh5OR+HLOZIqoIv
i/lq4ZEfdRUhjG91QkZOQUPIaT6XTf/SMI+czaNnxNkmpQxGyJwX+CEujyyM+T88yZDAm6w3Hu4h
uNXjZT1oqqg0KF1O07bYvFuzvj/VJMPhYxxZRzbhNQxG/I4teIwQ9KCl6/26Eppp/5Wrnfik6IhF
4IL7nY/4dJo4opk77rvYSj6n2GzQL5h+ErkxRrhL/7dfVI2WDher1CoEQGrOvX5BoxELFTDmqOiG
8fht2lbg7pdjGPDqngvAVy8Ft23/8qyg0yJFSkvfseNYqJ1c99mbLzFITSqkP/0vMMAKdOwNy0kK
fffAmsCnSILsLzn7ctVEcKTmcnLrUoMmuEbnG9a5RoB3Yg7KQry/svON547jKoj63D4Ouau1TW7n
PrkbwbJTcJcmTkrN4HdealdBsTdP+GWdzI597mLd9Pa/n3NuY2WG1EBnr7GcIu1h/vb98G6d0ubS
qNxbvTuXzQqIUW/njLFAj4SGqc2ahvprUkt0iZ66UI9tfgIrOz2EIYl9nxQ5h185gqVPcGVi2CfH
hp0m3XK/fZXSzxodkoMVWTRYDMZlXdAh/GQUN47ar4HdUwpTT7gUfRKG1xERWxergD8tT1Prw/m2
2YL4CyqGibov2Sj1YZvBGmaatBMAK8Mx2rcBIZOf2K2Dg6aM9kBp4+R+Tju16waz/H/4l19JYE1q
Oj4Soo67Yg0v9XYK8lLHco34iiTzUR+2Lwjz4mCt1du5IGQrO2yl/fkJkA4OaQoiwdqB7asjpxE4
2QXHlRR9DTOuDtEUWSceSYXK+5kjy7MTfvGM3T2DH7vFl4Zub7USNoObgvNOJ+4id32Iuytw5zlM
vLU952JXdOu0WQZvw+To3/OmJTVMewH/A1eH0d2Lk/LCcz5z2DO/faTNu0rHCDLYvfvj9TON3IzS
G9tC93aBY1LfJBAZJTQxu86QfKkF93U7D7G+7jPGJ7N3H8xvrr+1r9ckf/w3Ua3PKSjhcv5abD6z
MQJNwZ3rp9wFw77l8RXhXnNMsDM6oKYZYbQ8eLSPlcnj2jkuueFXMoDTYcEshV92TcexYHprP4dx
hbUgyvCeVMSEapw6zaxtdXXaK+JiO1cnjFImt08Ey/fMvBPrHITT9dcrNgLjz4Ky4YzZx4Fd0ZLR
73ZMbWqGPWffIkgg3DSWQduQbSwiPhik+8HhYe4kv8u/xLze7+0y+jJkWfub4o0K78dqOvYuNP8G
vwtdfXvIHpHJ6TcaofEAaQKa0C/WXqobPYCxZASOcthhFadFwgKbAJhq/+XgzpYwDeEG61BI/WFi
NP0dU5zmsyeLwd6StGseURDR07e2EVBpyqodzq1XXlmtzsUoiAHywHEUudCdZk5djQfW917xyl5I
IB8sJKp4ZVpp7X9M2HzNqSAQHEShaDjQr9/0H6zmNqgkC318rUjEET5+LwtlGnkGuN3sYVcsl099
39l2XdkDz2R0uT4s086vB8nmlJtMxi71gYp4/qcBAp7CsCylY41DeBMZlJJk8pwN0z7pamBoruNP
33WwSdW3RjaXK6yMMyZTzvfUZ4ihLYBzSIlrAu9cwjb3N98+sgOC6t3Nd3GB06johXUzHBNV+WUN
rNOC3khSLTr7RRYOmRojRYsKJ2fv4qkp25lAiu4gN6SdiUaH+tCRIyksRSAL9qV5KoK/hYKdpBZw
EcyPmfUGfuykaEmw9VDzTb3JqzW8MGf7ewsKq2Wj5cIB2Nyo90hCIIAzP+QqMgRr56YQKfayEsPV
dSDI3v/VmqQ/x9HVZm1oKu82Kpq+Jn5mMP21vbPK8LD28KettDyJeug8+KaLVC+1kL/719clo2Gv
tdDNpX2BJOXvagFsfg3ooT0366QXHnCxVTdBkmY7xTmbkBiEilWioOyUvYFRanA1cWK7b4kTZXSA
69oUIxAVXVkOEwo6aB6Xjc8E5rfIX6rfZ6vzBD4tDeGK/X3iMGY1MrfInmN0x+xHAiIayz++Iw09
8RuKF0t6TBhbZAckf1MJIxWDi4RRugatTA4XonyVDsrwso4l6hAXBrD+fx187h2nimSJcLuOd2Bs
sjuUL4fPo0pVtukOuuOUShFaMwcM7t+NR2bw1kCk+6ymq9RAuzEJ689Oo3xktSYwa7X5rR1eJrvd
Oaz5q+ORj5rhAox9UxYn63h2eEDaEMFj91gOj6INUN9LeeS56J94n4wJG0Q0RYJHgo5fahFoF/FN
RHWlQ+LNmRXk6Zl2LAkirS4cgI2woA1RGvd5OcNl2lSmQY5iWH79tafKtEntVNL6OM4V3ZhRXvU8
8w/kXPCqR2mAiXiJ1uKJCFRmhRAVMizQNzeG2OXY6aRIHzdXZUXR2qcR9gXd9FXXl57ScAzufNAK
Al8iUTSADF9zrK0PpDnZ80CwL4qmhGiIPJmOJYb0MVpS2bKjEUC/2j6K/cnqWc0QKXwL3Wipo1h+
YXK6fDos/kgzfqMrw9UlZXzPXWlrczhpcz04wGhJRFOB7sLVd8F8GsxfVNXWqt/30As5sw2hxHr8
YxZTq3XiDuA9HTBJXMF/jkekU0dDLh/mlCcPtwe8nkD0cXPm+KM/XbHSKlxsOijn0T9rKpKLztRJ
HMJ+jqpPE+JCISPnW0+u1B91mH5VSPWsm727cNPf40qva2oYa7S3/CeNyQmklcVLIzYH9GPB4fqt
mow99YbAwGrx8Dge2/cUFgdNrOfuXfCRaLtQ0BGdEqeoJ4TrmwyVGTR68c9ZanB7VaKhkTi6uJqJ
yLDlOu1ei8puvFawm6yLiyEbsSwipQbosHFjQNg5CcwAACIplfWsJx8zXZ46h1O0M5K/Wa0yHgBT
4vzQrzjPBP0X/KsNcdFuZ1Z+XAw9ZXmpjLcSQMdDdksqqkZX4zhru7aDt1W6uqAq+tnxm7VgQvbX
16yV2KNmclSTDUqtEyHwThLoZvPo7chQ8FbGWIDadKF9xKbFpBnU3IRscjci3b9uv/ZpIxHaowFt
lrPOdHIJWfHKQHwaPniahPV6eQezzskEzm8puBZ8N/z2sv4yon7RdBA600kTSwBA4rpxBktIBa25
4e+7XoSOWjjjLvzhTs/+fpVOsfn9iyd0VZfNm+xeCSWcNqIqbz/VrtXin+rp+5Eg8OuDIG+heYiO
9FztLnfrBiU8nRnQ3gikX7oUHmgSdwb8P0+cyieWn+Q+qX415JUEBHB+g0XtWLvKxydvxauD5pbs
VG3gAHrqdUrpZDkHFB5pwuLaX7AhlsDPrKZg95GKIeU/TSRGH/zd3spltNMOZweFJu6YEowj75su
PhCNfJjbKrE1edEichmOu3Y9nnOKKQ7XgxrMuaJBjR/+og4u2H/cVVlZ6SiXw6ia+Ze+JHAqNY+p
DyQSLDvOsbLJB8YVW0dCrnpYlsta1Q62AHtp9BwUxJ7m4C4FlOh8uAYkArOThUEjRN3nn8EivZJf
k1om11YWu+oOhjO4vmN9BZlfdCjgVomeNAxImdkInJoSpe5QKvTvjh3sOojJouGTFnZAQ0h5+0vK
sWnOhj4NtfCMKUeDBrRIpRMaYP7vMeO5743ik0nfo0Y0EBmGC2xIVk8EQ2049+d9LFNBrSf2nX/G
7YmL1xZVwKMjqA7XCreytSO7rSylJePMrLoWSK4nm5TAhGBpsd1CNgbwqg+XMB552+AD8Z2BAP1z
zy0o9LuzjYqpkJGPQ7NKFBrw95PiMU+1u/OMwrL/nIUmc6AQYTu06sr5SnI6lYJcVN5lGPQNnSPy
o393oCdZ/g8kt6182DXy/+22ctQMKyiN1PMsVgXdPEoKDnPpfQwop1CfdMYEDhR43ucSD9KZkLa0
u/LHE9sbhgaR0ipbSNqX1uL8IjCdg8K5uayNn8FeH0ztIT9dqM4DDnwDMFGGEuqqgfPdKLe3az0K
sl9ejWMe6zvcdX6kt1PW8i0MXYvNUNO3iQ55QwsqbH41LmBkMre7HsfaQlYghFlkNc++YMy+9HFy
hzw6sNzHPQ8c1t1Zv8X0sCQHB1fcJ2tBc0Jp9u/auBLkQ+81MfjHk9dXHUR9Gol+0mqGGGBqgDSx
j1s2f1cMqlU9Z5TR/ZxfEeR5h++zye1lQICcXQ/AKc+HM5nyGgEXPi9NIKbSMA7oAlPwaD3xE5q6
rKE9hvKHZrS4lO7RP6CoEyaUdEJeStcDGbOc8aWncbh23X2dgXuLxRPwKUS5FLW+CmWDqBP0jG2a
0u4BRZEUALLDkHxYfIeKB6rIs7GFKksnLK9cBx7qrEZ3UIVjqNAN1HtAQrRUYV3usDktDfyT5KSX
67Y5XBLohPGIu/PkOlSgL0SP00CoxmqEYemNkt7lK/tPccfawtFN9VDjndPmbiB2EK0pCiUdSLjz
CwgKGlmUJC/T11NsmBq9xapjRARDDgOm9cTwKo0KXeukL8EoeVeA4RIGj3F4qIrnsxF+UeX1okhL
rEb5LzLKYvgEneMTRSEbv1HaFIaUC5AhAKY83RXx8SzI0oNybx0EOSjb/h+YJF5HXIacdcelU98k
uvt02O2dQoylSuQ3P1QoUE7sTGj/uze6s6tX5PEL7ull7+F2IzKMU1mZ1DGi63sxSNQxr77h4927
F+TopmIhyqRMSSRVdk2RoqK1ZuCbFqyGGlldeyTHkcFZWkSk3I2AJJp/KMjjDBPTSCgkPpmk1n/R
1BgD+rYnaz1ZdyQGPnymMn7yUK/70GPVc4P6HmZWrVhRlvHnzwJkpWa1uctelUN5Kqj81fZT1bhl
YJULLBEIjCyF2+cToGxSLOPTE7TpOj8ebqfN/oZ0P4BxhBybS37Qrb3fLOusxXBOjmp+VcnyCAUr
V+IMGU2vwPHYsIeBS43Jiy4g/KyKQWhR4PttBdVYN81MPd5BURb3I2x8qLkmWXmFlJAWJ6So8/nM
8fdQCyrILS3M0KttufqnfeZ4Z6ZhWXJyCTlelCpfUITL7VKkZGku0HuxQWlbS170XsBT4aku5k22
i6ETFuoIRPmr3Jam2mJRBL6WaQdw7H9XZj7ABlhp/l7KasxEyUG9vZrFiQqRo5Mu6mlP7K9Vi/hT
mooU8RWnGyEK7Bp/0EzyLigTeD1ot6BK91WhY+1W0AeumJ23iAt8ocrkOZr08+ck5rOMgCCf9rxO
dVDU0woZVNb+2mMNFVeHD6+o8k+zwyXViNDfJILTC5J+SYXts5mSeEtD3nJ0CU7VqcTgO7FAc35o
NMz880FV15zGk9qn/jPhSo8peeS0Lh1wWwmKOoG4Ybds3RBUK/F/mA1lkgm84DqAc3BfnOsDQHJN
0tpeb6H3g1n8kxQL+KKitdKrkUAmKTFHE1Kg3hI2bIe8GAsB6KNcKsoNj1DQuj16vLPdgiGfljH7
T4tW8y2nCL+7OZHXyA3PRrnLa37mePhZhl24rZQpMz5fD1ZPq3iW9h+hg6RuKOXhiHoukQpqHup9
Z/ymQ6kMuMxBC+J8ukZKd3j7sWBdtuXO4aFLMPjYeNPGI3K0HdgfAMM92wq3qMeg5W8KV1nuzMZ0
3LrDUOggk/VTew1Mezj0YwEM/eYkpWv5t5akyZ/bNzxapFlzoNalrYFnWNQqpK24uMl3STaCYcLh
Kuvr0xKtpC1vx5XQYbAc+bVYqt9krtWxzliWGQ0gGRjL3nl9yzNi9mJgpKpEqk45eviZM/UZIjSn
3zZOf0UkEC/eurhxVUAx4ZipU1PcLB9qSzoCMRfQ3K34AqjM5MJnI1v7LTscqjZsnNAGYyFCacqb
KcVL3VzSg8NXRKzFn0iyGQoPxH/L80cShf1Vto5RcJ3tQBcSkoGJLmUZ9ugXGB17AU66IzfJInxm
Gr9qcmyKE1q9ASa9YD/wOCc+kDMJn3PDvjdP8SRtFBJd02GUv8sGDqxdlaNsnhRIRaxugzb/Jn9J
gSptTiB2mFJVbtT6w99YYpbfMvuJl7D+3pJU+qdqR4p21p8DIeRVDi17vnwBHh/oEyiuoyWHNsFB
2VOgm+Ra7UjiRGHpXltaOQQIXbIXenEbgiimBJcVpZ5Uim1sKKzhS19/2LVc9GDfTK+gr7TSWRzt
P1ML44ujD5zJtDNWObz9f2kOe4368oMUdsKLRzS53EwUgTVB8+5E3EECqGE9ZzYGAaUr1UfLp5Xy
1VvEv7IHheSorl46fK1DptrfsyT8Tsu6REUrP3tTcFYnKADdv9wroqS8mWLqN6W00Pi6Lhql9L1e
3n+GFcjeS2qLRdAmN4+qhu8sviAMRPhRyensvVSP2gFwyZvJLRSc/BZ7JLNhtXhmPb5Z6+oSDbyo
Ss5/Z5vSmXm2oSQbMeP1KnAJis9iDQwW+xQXO2pjnriUs5gKyxYjEDoB0lJSkD4zlouN7/sRaEwb
VVEqyawOGTDCq2jqC3Fe+7NeC+N2PbvitMo4Wrt2VPRFbUKsGhrBqzILGkr7OYhHb2cbBjycrfql
O3YW9sQwOdZ+GyVrDmB1j9z3+y5d/x/QyzxgQvOeijXZIZ6/63RxP50MxMI0m4vfSQDWiN2BL5Kp
BC+miOVpa32tguxOCGJ1fq/dNLJ+DQYRoWOjDZuoAQhgtV/lr+y7w8OEdRtB9vdNZYOinrQPbGZH
I5oM1GrQj8oGIyfhRbCb2AjY/DUupG36NLq3ATrsXkxFVnjxmNS4oveg7vHgAGnZ4yaWtzyn55+b
AlCL/LuFh1aquycI/py4HWsdOZDLrI2HvYoes0lFPgto3tpAL9A3pJU06nK0cjRn5Px+myNli2Qz
szSaynwaDtpkoQ92FdjUs4jm0MHoCriPqv17eSl7u7Ebiq+5p99/eJJyKAwMDvw9RS0VORwolLNo
nZZa8uKzzMpEYACUhEEf/QbHoKUOx7Km0vLu/ZJv4wG33C61C5dP5DlDnY6f3BZ0xITdLAKmO5WQ
nG+jQDJsYCv+Yc/EOVn1TU0/H8Hss4nGhFsLFp1TXRAu72OZomFtgcQbdvCCuxA2VgRzUI2NxFYd
WlshwcpdPS9l2R55WrkzkvqwaZXujKdixdYoNwqmFB6rh+goisO3qqRh8F0tUduhpfe7UsJdRaoT
BrMzqOdXNDwJeJlmoMx1kEWkeB9d/pkzi1ZiyT3GFuRggEna6ZQvdfT5AKc2EtenuBiQR6BBN/Ch
sPNFw+kjU0kGKGJW7/BPDF53k+hQS1IObXrazXGhfWZLgZacEX4Ko29ubvxWXcmJrdqbvSib558k
kUZS9QNUyjBEVmc8SZhwkwePzJXl5rVpBJSs9BnB6O10DbFOnyxQmoISjp/lq5FBNJrHS9ebtI9G
zhn3Pq74NGEwJZhTQp+UkYZbtHUZ0hlsYsnD3+pRrdjd3daxcXxj06GmQyO51aGeliQ/RvSL5nVU
uh+MSExG4/Lx44fqCoW93jbYUL76Ai/w2IwKr9MhsjuDgGMGBZoLLPPVbupByV+wb/5EKSEYF8vu
VtOEpnOdWCg3DdjmN6sh7M2vU2tR5uh8+uRAkhzMJSms8cdPxdmdW1ThfM0UlP6SHIwcXHQ3Zi99
Gsvm9/E4OpHgTMqJxPUcvbaxhJxyJLOQqAyycbkl+hFMcAci2mm6mR6h5eN0Xvng4b9RWcqbruO0
QojYOmTnWaKbSSNwVU63w6QvMk24rwARmz4NeJRB7fEv+bQzZhFu0FDbonjPbpbtSRwtUd4zHvsP
XrBvUP3Nc4KK9Boam3lVZA05xLX6Xyx1LCRH3pRaldXxHNbuu62ilYhFX70KpNSjwEXp0rBVwcxv
vKEqaySOsia6L9OVHch0xHsI0caR8cAUG3uPok99mEbJAtVc1pyAhsJ1L6sV2dCUaR6BpenXqqey
Uywfi/MSVtGRK04Jo6LM1njfgDGvjwmmJcYBPsFw03m2S+WN8X60hnbDVM86n2DrFpvm5LJHvyDt
Oo3qpM/7TALo8vjrnjYRhMc4hDV8OE24JvhhVJdp1vTN6dTy60uuN+ToAiPj85EytiV3jEXlafag
tspE5ioj8+mE1gvbHfxRAUhBsxNrxXXewiPabbjvp/oEoTdu/eylEbo44AKTEKfCv2T5DR4S9ESK
6yheNjtkODjgA8j7x71y83FifUBIRp8yFq6bQTuUfO8yB3b5I3PwvHgBwD+Cq9EqjnQ8UOf2aHV5
YyJBa6ZkTAMQDLPBLQxXhROcoj7EOKvmVlImUwOR7OfF6z8bmGI6Y2s3u6sUiLN/kNwdeSafuzoi
uWL4ca762Mab8Vs2+T7EJDTh90gKF0ChqRuGOV0Ws2eAmBGO2JmuISkl0wrTJ0Kh5fAIZnD/Uw5o
XJfq0THGjH5j7LN/9I86c8hUdOM40RWnHX6BvIpNeYaSRH0oAPuIH0PW+mfgNz5r2OD1Ui4LM7j6
0RwRrq4OJNK8YEk/o/yzOLiEv4GhXhmAei3o8HGjXvWM8iA8KE0KogTH6jRWrTQEzR00sahoHrNe
BQ0GIF6fOfv57CipjZj74Lz4sBpFKRiUF5z7f1seTMJsUe5hs78vHvb25fk70WrcFayjMJwVT+tr
w5SNuLWT+Kp46OP+3QxAzCsOVT+bDboUGHVYUCCOj38Jozi7jriqAPHt8TuLmiO3Csv5Oj6zKKuh
mMuDoKStI6+weaL6O8pwsCUJArcqovVhpP/MSdWisDD6uGbayFuTWRHMBHyisiBuAH+X7wLJYwIj
3yQj9F8/LYwYn1HiR8Y91tS41ikE0ATolfnGewieHbN4r8MpsgIhbwP+GdO+Rsk5/xAGhro7SwHm
ELW/upHelgerY81P+k09D/XC1D9ED+vNrffJSskKOfLUoZOaP3B16adbBHNhTk06CUQqqtaLsHwm
+C+q23yfo2HYHm7wWJRra8DRWRTahokTlc9pDkRFdDgwzfZ9vKUwSDO9sMdboY7pprDosalzeI9M
ht+ggxA88jhFrFZ2wODqOpkHnE0jl5fHcyMX7B0r+BKhnhLpiEDexo3HS+fhJILRIlVODYwM7elb
0mf7dAnHTSnHh53p0ngIzPvq3aCioYkNAoLbjDggUnvck6wVn1UrTy9hA6iIot/lhbCm7KcgI28U
JxDY38KXhdErO01/bZkTfn//ivyrhzkNtcZc6R8HSoce+4JwhnhGLWdlAgm0FEH6dQXfJOaQZ5Mb
fXNgaRmteJg1SkkLPJlYq3CaxRyYsGS3Sds0vmFxk5glGTI0lDvdwxfyc5KQ9wO956QVgyfj1J3L
S0902DqKDYnauxcfeEkclMhjaGtP+26GFD7ok1VaL0dLQEFmv9dt7cnv6S7AeOt9LEdiLP8EC9BG
eZb/fle4fx97a4FO+I3hFLzdH3WKzwovhHoIMdGFN8uCyHibjq93GetdS1TaxYWX2af0z0O29R7a
7pQYIR8qlBDgZidDmtYqs21WR88yH8F+vKNxz/z5VblQvG95XJwX27vzea37M/9dHF45a/tE5C4C
NTk0EELaU3mAnjsllr7gEeriuR7xJKqcn//pdjc8DM/ZWhbgip5DlSVdXlEZNVDbNOS8uqobikIF
K6CJJGmXWvrD3A6OFjc0T0Y8bitsVpiqQvNgL0ZEtySTBZwemor8K1kKoTK7bE4426B7XAaZJZE3
KID+R8RBkpCLUD5oGCK27/vyopqCvbrFAuz75hWxSJg6KboQ6V5GG6AkykLf2Cl9qcvHKZZFKNlw
V3iI4ms7lKEtJTyVredbFKZZiO7En6pj4iBpoP4NjFKCT5y2glQG7BC5spMFzJaW3ej1vrmxTUgh
jFM7HbvfnlFcebxGG9pQN8bA8ujt1SYSYtcfOyHm85ND105vRE+bMYTTwckMzfYHGwd5K6YXBYri
A0y4WilGCeCXvXU4lSn+E+LJHmbNUs8vUAa2vlrJVREy1Jo/ey26xUHLQd1ErM7Zl5e40ZGnS1SN
xwXK0ICPbqjJs0YhZMVKUzg+t2OMjjrGWIntdHmOyzs8OeyK0JPa6A2VHQ/7Yor83F+IbgNuwRwZ
TOCjmkSi3ZytKChJBYt6yeN3fUaxS9AlxPzNooArrkzbDUhDKT5VeBEv3JVqesdbSGdvTphsTt/k
zUGs/jxLQ8toPSPF6my+rg6iDQNLsSXIaOE2Ot9ObOhpCvvIMSW/RMA7SlCrfWZZpMWEj0m47Vx+
a1nvVBc0vT6r2hi42e0+c5yM+scrCryr27S1mxDKqhP7CIfasW72xXe9uuuWEaWcMggaEDuQHk51
b54Fw7TRQB/45F6lNpTckBzRVksSFuNgEo+mUHxZaqe/ZvqX5tiGQbqGtkVpRjeMrfzhGej0TxcH
o9p/RD2GhNjU02pcVzoO/bqkEEL5hG9SCh32YVC1Xs51aEh6n31VWCcKcpJsRkw3RDuPUDmKxL2y
GRvFa7sMqemhDR+RA2GjKMCO2C1bqDElq9yMyoakIoUlxMPgf3Uly+CWYpV0AspxPoVd3Y0wsI4T
Gje6r0q8MLss/1M8v8pM8z8WEFg3xkTDZc2WzQBGbufnyld9eIHIftSIfjfWbdsUopbnmAv6GqmN
4rFYDUg9fladPvv/jBD1vKh1aL8XNoYZ4tFPJx3MM/3mtntDIf2yu3kbI3Rtmnh83tyxvB0ASr0b
4CpA21qT+Fo7wj71tLpobxwFePME2vli/YTWX6qHKN5kuV08mqLVbARP8vJvpZHhZSRxcSv6EepY
C2GlJQ65I3QBFMhpUSqRLVxWmBQMn33RzFoB8NBfuwuaZOHqDywDoEr+SAjPhzdCCxQsffKVaBef
zI78AK8mzeGeqGw0wN0l2Sf2xSL0A2HjCJziRJnyVholePK2v4fXyIAvevxFqhTXeVq457yPtvLT
MGMa4P5jaRmmA3ZQLjD5J/d67yWjen05oBgysYmfF7iAFAPvhKC3L3tdngW3ToiM2CP1FWyetTT/
oOPu8Vrrwk1E3oy2d02r7wmQawDppbfyAP8mobNNInkuUjJfqvULoCSlVWYawwPhyV/4ucgbivb6
frtIBhwKj9zrz9v88XfleY2X3b7eG/u53TW88Vca2vdN8MDyh3MJmYMC0Bmhu5hTBaxDrX7uJ2oC
P66ihBs9qVqeveGL9PhH6dsSP6O2oWRIw9BgfMR1vuzs7pewKK2Q+lVi7LW0P6Soh77w9X+pxsv3
6MkuamZsTjhy06Zrc7/7wa6kqRwpjPwylnnoH38ggt+QYgS67VpGtKL7QO7SJV0mImjxVAT6LK/w
+NB29VAg4BHICOF06ByAKgQjBIz11FvtpCo8RgGI0FsFeDAiVOiVmXKT7vokTQTKQr6O7PlOtYa/
aK67d8sAaDedvcTxl2RvX12GqyYgs0mksj4WISWJgeq44Wsna/rVvEAZx/itFJBRUhSNNumpj7mc
hPu5dUPiVWSGkeUgwqT8Qo9QxBJt6Jy8T0FYA65SLmPn6t0QBJpzEOyOfwnqy3gTguT2iwiDIAls
/vcoioQhg0m5g3qzXOz39qYHK0mlIr9JTOvEulFBosh8r3Rys2QDicbSPt6aigSHt88R80hvjFHS
YSh+N2SPBRmTdf+z4njMfYUcuYutBopWlBUEwRUWjM9x8QO1AMbZD2toQo0abPJhOhfSdLrZeJra
QLO9TVXCFpIaFu2rSiq9Xb8SOs0ZyzvGmCOLF9CTrMkG9eG+ovcSJkW3vXJoIsBePDde8lJETicL
fgSmYT/a3GsMmjUt96927KcXVTBLN6S2VD8Ik2Yk8qjqtmlQ60vNIhjf10o5NWbB7VTiDfF0qy7K
owpIwN6rt+rxrRkpV9UhbdKG+Cg7THGgVTUPjZ7lCFVnWK8ycGeMzUWu9SusoV2gwaRCi3xYgG9m
6quXF4S+tnSQu9yTvqdlhiHO/uxdTVxLAdeNZB/J4NIJzRVzRvJtfCk/zPgNvo/x/vafewB30VlB
RkJy7JQti5sMUvwSsCFKVAvi82ZvgVeu2khHC5Kr2Lo916i9W3K2Ppt7L2398g6CpndzWe5rwYqO
cIzfwfzyL/g7jB4QjzvSTh4eGjebzXC8J1rPa4KIqK7mG3XFzvq4v3rVWUU8VmektqlFrygjYf6K
ZiyqVVDRQ9zZVZabaQ7pweQpvbrmRzczZeX8AJ3PgCzhUzDY3Mxq8uTJNpkLD20A/D1dhq5D0C5h
4VkonOQRC2uiQzTkwpmBWjHSMw9NBfrB/d5tZyBQY04bqhyZrmlQoRdJW2rMs8OHsciGIY1tonnn
fdBHrN9mWfDGHElrAaNI4ZF093wBeUNCALCLNITyrDUUErlTBapC9WjtgwBf0vRoTqPM+6Jpd6Tw
rwLSTgfbsMNJkVPS4QfP4S7m54IonKrHBEe2L08iS4Eag1hhsWVXsGIbFu3k7jzoSZpEjn0C6dF3
fjRPJgWUNFp81ORPDuiPwDmG0Rju5oPYUe18F2Ux1BFkRFn+jRdA3EXcDbEcdUGYbLhV7Ndnx57s
OahwTR5tj2jxWMJ1avyw2VTEzulmfeK9TjNTZQyWrIHtj52Pme2Xy/gP6iL/VmzXTHiR4Y9lqQIB
GYhMzcxJT6z5tG3WYQ50T2ylb7XCyx1tWGp8IaHkuO8YJ+eVhUYjuUwLOUNye0dMhCmzOdAM4dGs
xOVIElIeiAWWVX4PLhjrWDcCnhAWBTNEI7ItwEn7HGOHFZuPh2PHhToZzVGFKka5mPgVgMWeyqMr
73tnpAxLMxb5P6OpOeJpcceJBsIvDrYHzairhmS93pFtsIxvMFM35ruXu2RPYt0IfrTOYKk8Ek49
MpfKG2Eel/wrm84Q+xRaoSm0v4oHCzIiiM4ttIfPKpQJCdGpwThHd85AgAFDVQkJ89aV2O0c2Q1I
yReNeu1KehmKTc1QqUqiOh9oKBSGKmlLtQFiMhLatadF0fnsRok9tl+1xhfi5ntK3aFnY6Cy8U+o
vWE7CUXGsVJ504BKfXAG2xr2AtYz+4Z8HdLnpBuIL1kiIw2J/RAZ+lFgUXJHLNbnrMyJnZKhExGZ
P5QNmmiQPTVxVuSzOUUMwvlBnvzVCLFpDRzosDtyrLL/mxvS0oj7M0xINlPY9vDSvwyxhLBRiw/t
p80UTmB+Js3QBgNqeaJ1XRyLDMD8rwhu0YcMEZyO4EEPFoK+G2PxqXoBI//Kyc+RVVvjSIeU1j4R
xsySb/ApSS/QNNWhgLdZ8oGav/LkmaxclkW+Z1v+CvN3YNSoRcs2qRqipCFcEjKRcRS5cVw8EOha
z6LMCifPSjV/eI/PzteU8Pmf7TuPiWd+DtdJAiMSfCavUCkSWCWoZNMlOEN9s7E3LDkX+CMgVxyb
9jOSSvczeKrJrY6W9n34/8tHKJ7BrI0bmfHBxlfPeywPWIoNjZ8VdJBQf5X/pbN8hvYRQ6wbVEP2
Yo3Dnc7v/NEdITUf6ah6I/q9giUnO4IeTZtv51GMqs4kUUU4Y2PFceyHpNwOcBKR6p0yWBG59fym
QTRRUGLQpF+gdCmcucrb2UOjIus2mpPlSrxSS6XK+SWn6LQq0uDZjdy5zy5oiKilfuRD/Z6HjM5P
sj/qYmiiRhmn5HESDrNB/PzbIzDXouDjv9rHI0Mg46BdwH2G1INol89MjniWc133hGxIIGdLyO9g
vftAArX7QvpNhTtOwnVZ/Uktegv8GDJVJk0AZELKWvugLSVgtGzXa6G4F0+1GKv28zhSFQFeViqo
b1p54ZvUL2teNUPsXgCr+dAEuBE9v71Xk/8g1WQsipfgjHuE0Lon7vM71kznJ8/wepv4AY8/KbKE
e7owF42o4aI7mKgFIiYRcyFBBdAokn4PwB0/lTIuJAMgdMiuKrfadRr6lDy395578vLeIZb2jp4z
7cx93DxS4HefZ8SnaGPDFLqVt8KODMWgFc24sM/QxHmm7sE5r0siKkWe/jvuL6laeWXKx9wIfGu2
8LRo4vvrn3r1yRb32L+v9Jpm6UP8wN0lzuXeS8sVL8HE3wTL8Q+UjCFKOdoG0doelWgxe15ReuuD
9IAc5SfDeGmb2HJ52PkbZ0DZeY5clz4dJ4HIJHzjinID5nPSSBMhpDDrFduKrBzeng05VnGeoclW
F7xDn/70+GGj18xgcnvC5AtW2xfoHc5Nu4LWN70B4R+o3fyr4at4TFQSukaOzF0RwZhCTLN9nnlv
M6FbdJt+zKr2nWXwUC5yPRy7xkv5H/y4r2N0HE7J/fvogJjlhBSMAfXvpBYqPWKs/NLGAl5IocnQ
KA/B7EVEc4GDkNqQuhij3TYO0dTpSiEj2LVwq/J2/S3kH97d1got/6vhJldbXzwUfzvcBj+H1RJ4
j6/1i3vHRqfORz5Fka6YEuKlODwOWkDSZNIGEupExG3s04jo88ywPkChjYVHr9on8Zp1RrBk7a23
U6GPYBm7ozk0pYqF2KrM+QBXMA8DmSkZbULEBIC51SeorV+2kVZbSHsdzwBhnJpfINdTJEf1z6sl
t8PW+mrtrSylAWYSnlFOx/dJ2Mqi+5o3ppcJnUq7YPXnnv1mEGNIEOSMDgF+8ggNBEs+5wGwdRrJ
KY50oKxQx3NNZH1vMj3ZxOzg7OAAmV26aznKA8a9Izzcvr46x6TbcgCP8aieGNoJCXjF5le0RcvJ
WcySSxtVbudzoP9tz65UGCa2LPOnDfcOqs0OYKl+osm1pD5eoLdPvLpLyySi5BefHUnOVx2d+75K
3lunZXlccaVDRy7qNVBS6kEkJUm7Vp8b1pHzHxrOYOj0+KUhonnsDmM3JR2kdsnu8tpKAvCGidn4
mhVTi7sUUObajAJA/Th0bxqN4WzFVoVgIPM1CmAKfsZVYomYrEG/O/k30FXq9eiZeEITeqTasQKH
UHy+/prrJGOTeNhtSxl/LktTPQUGCnh/imFa/SdOAHTDxSgvePyn/X9YEXp+9YRZuG1D47f9CqOr
UoZGZttVPmwClIj582Rp6LJItwGY2w7rzehJdhgb4MhM0DWRPmmAquUYP+DNxDoKy+pGR8ckWLho
6OZLSJyDm6BK33PfY4APSGiBHTkXo81I51cdp8gtgVEK1PbOTcqRYbBim6BX7mf8KbotIqYkWppW
sTHBi8rNDQ8FbfporMG8xsqdLKIeBu8YF43lWeIS7Dikwi+N4kz8iiCn6z95jmHAL0lg/0svFaG+
1I9PLcR1esIEDv9Cl+li/H3UGE3+/Wl/efLaI2azKvSI/1W6fv38MVFFRrPzlmej2zJHtfYt9s8m
kJQwTGob1dHoGhYSoZPgdn8YVGZi8fnw06JoGlWIOG8Xas0pzqcE7l4OxW7OKGeuS6O/lSk1PxiB
KukNPgV3HgxzwGlD0oX9fWNnUeXTZ7/p7hufINYHT9XAptRarheCf/0UDhdxDoirSfkU/wBQBGWe
J4lpH0cxssCeXuNB/WxPo3wgh7/lD9kxF8tdbDTaWPInV3NgBjUJ8eZz61ZiMr0Q8qGBBUrhHOpY
YMLwrvurn3S6DO8ZZvy5HsUQabD6iDwVZUiQ8FF3m7WYFNK2RLKD2ENrCrMWRMXO1ENPSWqK4FHx
6lJsMGQX+rbMOsa4boiBEk0s8YEV177RgNQ+lQhH/PlVpnD7oupmRZoG29XJz32AAATIGkQs/SdV
q78f3MJoel/QxMOi98Go8idmxJhm2c9APZW06q2lr1krOABF2WUJK1LBsYtN5vwvyjcPLUaXzbv4
NMEgkFmz1Bif/4LG5DVUTn5Ibr5kyl7wvlV7cp41tAbNC6UeOtWLAseqkVYRNpXmQ7tc918vvxAG
DFu4CxTj9rr8ZxLbdpgKRwrxFygvW5vMuc9rE9O3HV2I+dwYTYViJLocZkHOVzET7YStUUmfXQSw
Udgv3c0eRPhaFziD4AXYLbyZWVN2fa5hYosq7xAC9Y2dUS/Ji56kW2tm6eZHBtz9MLRgVcKvKELG
WhILGRceKas1nWwDBHlCO3326H7o/MBUk97Vt/JIYLK1JdXFcO17W4/1DbcpBmh/I4nUtMqsunRn
ziWZsRgAAL7eGzZSQKk+xnUJiMUvjdAJsU0i3Drrgf1YThkmeNA9Xm5MlZJTlOS4NAmUihawRugd
8mjQV9AvTPIWDXmwHS9UzgdM0XGTnlw89aSGRNGfNwS0ehsQw076zgNc3AUyHNE8N0+nc/zvcP+/
7RGm0IIfz+g4T8ZjOgY/YN6bJ4RlaBnk9D8Y3AoccKfgf2axYC+CJiHpT5XM9ItW59RVhCUz5KX5
QPxFgm17TIi/1rso2L54Kwk4dQSV1O3wJ9wr+ENK5raf12paPqbFbA/1KKvHMKiWJbha5F9JGUbO
n5C6TRZVl902/E9npDEKq7LUc8I345NSBFB1X9qn8sqxjtueYgFcGldIigsJ0p0KpU/IRd0I2vts
zbqRCKILhCgvZSxCxFXVrQc90nR14XoktUzaz+UvFfdnUej7CyFJXSAw0NMbHGTY/P/wCGjLMXG9
WVWT05i9EIddnc4Z6Kiaq1dY8He1KHA3zX1MkpGf69miX+qh87+PnzUe4GmnHDwU9OH9HWo4lpWy
GACLg5DfYhd//4nmNbdKU6LngfFJzKqr6vq5C/Wyboz4hD+Lm2sBi6ITjRBKn0eNSDrMpVtVmnZH
bcumX8K2IakLqjsgrmVSN3PANjcFaVt4VNr7YA/x5+bdudxuiUnGPbnnsn/gRUb6vu08odSdJldK
mxRgftZ9dfqKMc/lkI1/FskFI13ALfHtiMOQIkQrJrPt/46ziisW82IhMFpNrnlz96/UmetAWiie
Te8RY1ypqMpgHiyVaccC6STYnnWUbC+eE3mN8Q3Ov+3DVpw+kSj5T+Ozlr7vQPr3CVlOY94OgHXk
zzm02OJ14J9lKoFLBJjCsplOalNdxA1CCwpA7CsBV0P6Wl58NCZe39VHsieuZHZDFMy76aytnaM/
1B60OUWV/fmZSMa+pBYgPS77yyynp18ySZz3NjHGBYKtVnspIUYynpB1dvm+rrx4Ty8HtaXXcY+T
ZObDly9jyB7Vb61dzfXPNkd6xaqtpC7Ixjo7ptpZGlHaip4ltVg11T/rPpuMvfVXyqiX4UZaOWkN
ZpLjZ9hmxs6A7AEZ8bLXmRKOKcfclux/FHHjUQImmLF+r7DBIMUDkjuJENaJ1Nv3Zo9O/50yy3Sa
x6D8THxied2XEfBrkrsJnyfOnwapHwp05K/wRbyEDvyapUiEYaKskl0PQxH+pgHKHEfg4L7h5cqT
8L0lW5J0ujXacNXpPPuHlhlc0CS/7wFIwlW/IakF0Lv4vU469JtO01B+UYAfdFqn+pjF5UphO84I
P1MyKsaxDETRJsfH8W+KQZUmvjQx4FrPoU2soFojIDThvmkuvlcUbEQq6LnAv2srkm68sCa0fjBD
GaQE/lOZZ5nZiY5Fy9IVw4bAb7VNSCRB4l+FPdY/kUzDVYpMQlHzVXd/lh57isKR6IkLwA6CUNmA
BlB6DWy0F37hujODPizFS+pI910cX5Zu6WBqOFZRLh8jqANKvnUDqMj1eNWUGWoFNgJbV4PGK7WG
cetAsP7/Hg7rwAzXt/9a/i26yI4TLVvtpMCHMKGCxd1VeaIiT1tTngq05v0HIR0uuVnUDwqpL0cg
ZJg5/wudFYIdnrao/Ce9WjTWTac4Bxg2VBj/Dxn/LbiYlZL7OhuP+nKXuAI3CPJ3lUeQlgv4jlho
13v5Sxpx2e3WRhGM3JtHA1Rpke4MJYeLSFKsWskCZFQdRGAc1WlPOUpFNoRgbaIchfzFIrEJepYb
8PyFFO/sI+L45+RYOtcvXqw3tTWLPJ8eQDysjSdgIJHirCwenIxeV6SSmhai0Izbpu+8b1b8z41Z
rhRzAnn+6HXFI8OCpUF9cfKROrULKweiUk8uq9NnWbk0NrGl84DtFFi92txxte5qAs3tdbME5SRb
17u1TuK4JlW9rEdTXVwDFnwZRlRlbieOfjCthDY9s2pXRaOoL2QwORsaHiB2rEqecd6RVy0hnQpi
U2VjaW9k7MC5kbWeZ+NRoO6bOeNf+PdZPqN6dQoPSR/pRmewdXMiBC9DY7kmILkjzO0ukNJAc7NQ
2NlUMzsq06Yml9cZekBiqV+Yvbz2AdFMVO+39Kb+LWVuDkDs+WywFNfMWkbzgRcb2mYxYZWdRcsz
Sub10vuqCNmeZIn7jAwN0rz3KmVQErRU4rKijIHpybszTjlgXYZPhHL2beS6vLkAdy97jHejvI7e
04O0M4aUkqf/NZ7+OP4IyFV0DDd8oVO8EkQ5OPty/LpWuFvwhQtk7v7yuID76WNvKby6aZu8hhc8
o25l3W/LSQIDr2LRQQM6+Hv7HXUv0sioAXs3N1dx7AYudxnWsgXYKGk6o8bXEvg2/4Swlt/+aBZ1
0nRU/raOHA/rtZZJvfKxY+A97Du80FueAC590EjH2SG2/fJgaTirZERudvJNxcMP6cQLWDheyvg6
dAWzDCJIQwJ2e4lzsP0yrW9E+0jGxmZways02sDQjtQamj3nAzR2W9g9AD1v9xo02Z7BW4LgmGkY
Kewo6lvueL+FQNd3ivAsGJl7y8Af/7Dz8zdtqi6nw/hKQ1REiH50/V6jTvGxnDOnec0L+yrYWtZD
bvFbASUtfTKiBrgLo2ea0v2YOp1WFmErAfijzdK5hqVzmZVwSxNwajuUnFERuWdAb280wch4U+wG
rLbnRgiwth5Z6YnM5/1wFVnb4574MH+kmlsY06dV/TpvSbTUWEcBOV3mpdrjWHxNYhPImnu+zdJg
El1zIrEvxWlTejqMdxsRTooRwJFYSOMb7TmHt2edXKVEAhaYbBT/3dnuiboK7q3e9WInJJ7KQqSE
gVhbYDxS7NAk14/ezL2GEF5HFxBnIo6ttTJ62kHWOhzTa49ikPVNnjChqrWp26GlLaVy7HVqz+gu
bWupFALOaoWWQG8SQA3Af62WgaOrc3Eb4Llcm8B+CNSdTp41+/DfQZP+3tKqGKm2HUJO65sjyosg
UccUNU5uTOaEAIg1cd+y9OBsHjhUNKY/c61iWJOPEXLnVT62Q3/P/lHq1yzGgRD3crYvRMOK90y9
sCSS/X3taeCL2wIF0mWcKMm5A68R3vupn/seGePA0WVB9VChCAgDx/F15TSAV5ESNvdsieyc9Zoc
qPT+rkYubDd66g1ScvMiCkHs2mNR5S61KqBsrTDAYjCW0aYygCSm+0Z4frFTK7yHRwRHvOn0HJez
GhPzMV1EAY4+lpjj1g2FPonm3G8zDmqf2Wfw/NuvbXJ999QTMq3kgBXigY3e52eBrZVxAqxsObZt
r53u645G5PyUI2edsI+e1j3sZLeDHGRz7lfU3KPeRP2pK6jN96iuAWhFFfHTAxHB6TVYdEsMg+F/
MhNQawzZlqNZ5wWgMUopgf0K7gaHq3hGrJzN7JE3P7+jEuf/OLe20eqRUVN+FXfBd0xsbqD9E0/5
VaTnXEzfzQG/pU58WAlRclrssCpadJ2z9U2QA8/fR9S8/aiX7paHUfRCs6D5fZo9CjIsvC8pldTa
iIOubTEV8BYvMUvo82aoOETRfVdzcy9qlSo37ImCPMBmI0okFIG/kAOkoNIBI+8anyO0RRYH04A8
VniYVwqWa6brb1F2Od2ZmFCjkX+b8xok6/vWIVzCdUOoO02TAdO8j1aGPMWNULHeuk45Iwijsm7x
kcoWYP79S68gAhLcnQvOwSYFX4a4hC1W6Y6Hmraex9Re5FPhUSJGfI9CnMi27LKlbCTeEoJz9Rql
fXEULidd96J/8HXXjuIejGz4hxLDCuHMt1b9Hf8l33hZa1mjb5dDMF3ggCDC17VYbqSnF/Q6nVwZ
J4qWooy4DE34hi7XWmXrYNYtYce46ZodIA8rBq5WqdG9js/CITRzyFazBonS6/8UXdI4tKgbu0L9
jKTggA792VzQVoYKsDAJMwF60MTPaxRqzCbo/wwk4XICV/VRYwcfDIFkhB92x14Ezq1K3s1j8zwN
B3HF+asbEpMUQr+i0Pe/0B23Z5xo8SwXomLB+6RBsJGl/LNaeIR/fi88dNxJFCldoCtfFqsY2w3f
WGEDxL9jcKs7MORjUOyt0MeUEChCr/5Ndaxww74lV6XsFHbtoDbd+7P5s8QtCUlnxtkewFICelm1
ZxpfUY72u57+isgl56X3MyMEkN1yG4HkasQt7TX+AMSxssEOe26FHkUKMMmUsePEeS/qet6aso3b
sxMfwpAAzX9QPVdtYlugda8RtycaRrRXLY9bQMgKByXYu8KxB/0x7o9wTAumsT8Y10qOGMsJgV5g
7UKFV0Y1jtDWANoJOyt+v6SYuNx71GKV9mEWPmXCUbTSGlh9QYnLe9NPXHpx2Vv+oYjfVv1CPq49
1GN+iKKcSB41hqPpiVQYXdU5t5Zyp+Rr+jk/ctvuCGc+8jTbM/q1GrwJEmygi4Ah1+3Bu3wNbSx7
s+j2epsz6HrM3QTP0bDC6rqhYNrknKpNo6eBbaJlld1DVUPMPfiYeGMk6tFSq8bn0WN/vH+oAjxX
kEjnYXYReYI/RpkZsRnpTqh2tW1cGnqyLOCRSb1Yv0dNnb66h8yNaAaUJKC9ChLZZ2n+EA61X5n1
QTb5yHbh2TALi4P7SIuvqxnHSQXkkVmYaxqttK7vf3QUY4/i6D8B60Zcn6IjLHN/VgngGfhw1DAt
2FtYhS9xULL/gD8Lwfq+fhMQdhNm8E6uVQBoY2k8jjGvLL1rRv3s2eYcORb3FB1UjCbkA6atogct
Hxu2UM0xNXZm1G+icb856myZ6lAuiRpRfYjj6ubR7UW4lZnFk3QW4De7B8L1msUdEseGP6/BEjUF
R9kotdIdKr7VgOoxvD1r/3Cp9C86zZb9/FwlGk9uq9scmMzT85SCxWtrrRAmJ7rTNq0awupO8I8d
DcihgJkJtGQoMEjE6StytITs7+Fv3emc9v0tO0O5Er84CdVGstqbS8P7cK/3wVfAJyXW8qgN+z5u
C5YPxrTfe4hVHo7R3XCJlN7h9JuCQDFyWSFrDI4K38ERBwfAdGxgZqlfrWwEL1ikyAPrPjVIt53V
LwdKL5v3QnnOfIovDfV7gVpzJrcP2RTAkBcrZpfGxP7kpzdYG5JML9zMJvPEQOZ+YVFzNpdWiHb9
AkVcIEfjUgw96fOio/n/9Zzb9ydJZyPb9TaNOqMTB9VacPAAiib61Soggauw2PNg91kjqBycTuCu
Y0QFZhEBgBPbYGLHFAzDt2cOd8nMhHBS9bto8zMokbnRH+Y5tYlgkybTJG4KB0CgfPrURiswtJXs
tRxZUD4xuvMXD5PA3BtGYdyWOYkxNL8ZadLsT1H/ciwfvvAQrgSGRj8/BDuKYzpt7zBm+7YFBK8x
n1LvFWkZiHq0bkEgbr/QLG0iWCv5nrVEGjWEoXcB6fZ33ye8KGqF7jDOURfBuDWhJYQ5QuAd7t1Q
XmwLrRe7YLUWyNl693XT/xpwRdMFBOgRI3tlR0wHv1N7hOyTBHTFVHHZMcxCRqj632NPe6gIJi8u
t8dSgy/1zyHeVk+8H6pyJ9wv8XR073XhjnprV3gjCJzAvMXHQD4O8F/8uEg42vpwwjCi2eVZrJ2B
fG+U++dCmAeJ7Ry6sXnEQtuxwgV700Ab66kPvxlh8Br5lQZHIYHbREtvoZykzaVP9ezpA1SVRl6t
4MpfkFzSnh/QP8zNPiKD9vGDWg/l2SfncRtDCBySO8KiYfwJqeHuQqqt0ct676gG52ADO43D4s4A
cQDLLhEPRfK7TRbqG/KPWxBEUFzRqE+j8ZPOTSkj5gcMn78+et1IUHu93VzfRCumNS+Ku/T9q9gf
Qh4VhQ18zUEVnZOvExjN2idlmVrDUtBcaHLid18hULQNbfiylXXnZuZSmQ/ITn72MnjQK+5GIEiv
w29tP4lq5S7WaGZoGZNHUeLAkzT08I+tCWoqgqTAO7+vrbZJMtYCar/tUB4u13MyueDn4hhy0rpE
rK2FL3i5Go16D2DVKHODdLalEa+Wu52heUlxNoQeeMZKxUu8Uic5C/TAYE+ety6tkS8y4wpHmAzs
HgpyZiNHVwPxyqR/z+svgr3R7Nb/l3atFFKnPjF+ysEAzBBuYmhEhq0En2QtLw+nvZfZHMxx4WpX
mFCpzaYltxS3AyYbH9d1vpQikkpInraXQtsb8S57AKVg83I1zYf+uOB7Ri9BBqAshN8wjj8bVIzE
cjRn0WzHrTWTLZyAp0n655c6VWPH9FfJnK2bwAlggjEzX311TPQIka+9bfBkLM9oI4ciYxjWNMqQ
Scz2Qbpk4fTWxaYOFUcASLYexNrJ88Vuy3aYb4j9ADPA4bhpcCAblaUQ/kNtV7FemAfZLbQIQ1Eg
VmxJCXxl+OJxDIuvga3LasyCbD0OXRiZ2vMT/K3I0MAlUPi8F7IdHpgT96E5fwkCKd46ugemtbUP
ykgHpC4Er/u2uLBqQREww9kuLLSpGbyapNTSLmJdhx/qk+hoXYHKH/dEpj+iBglQ1ZZ6q4HZ+0u+
TtgvVIcuD4DRmr54AHGH8eayBPM4d4dN5el+RoFfU49QDMR+c7UX95ZN6nP1dCk26v5skKYsXiDP
WD7qSpSB7GgUdWsbzvDDs718gwGU3yLf0f+iRMDNZJo45ymkfwBOWYGvM2c7VMy2HACvO00crqpj
J+aOrfCqkzKw+VGMx0HxnLEPd1qWfA3CBRquPDMn0G7wWMDs1kg9f4X+kIoOHKLzv+DgvPP6bfhv
L+1StvMkFwYufpe+ymCv0BWdAW+Q4pIUOipYSby+9ZkK7t5ZktYtZrEd9DquJfx0+Od3RIxM3d3d
6mbFpwQd1+maMgwS/ocn9IEbANfTKjiqJtFGt9/ysu8qsxdoe/m4aCy1Xwynr4/HbuwA0qe1t46w
V3IEc3lQJssatAdJxSWOtgADzz8LNYIAwQLTqt+3owELrONtGlwEZ4SrrNlxTkwuM8bmB4KwcaSJ
JN2+NBWk+PHWEctbcwAlbDhB045KInAvOF2EihP89NpfgDfhBDQeQYR6WSaNCxdAeTK0mfrUNIEZ
VK4idA8eojwbQQPLeJb4qUfUvZcChygjyVLNCirfDBz2JOQs0ZVEBzW5YzQMW/8D1NP0RlzJv07d
hB4Bq3zkM021BIrj4bIMF91Nl3MKCweoMlxMNzung81RzkjLLlEUSokcU5z5EKZ7+cCOP90yVe57
YyPtBCaPAFXyezYtI7DcSel5/5JQYedS73KmKDH+s4l1t4suvfhOiLW/zdW0rRClHyjObzMlAhET
tNmP7uVMYPKKXR5ZHYN3HfncAI59y5v6s5HAkTFaS7NZQbKQYFzUlCI7sk2yNJtdJAHUm9IkPEk7
LsG0bgnIy97I5lYE3hddcsYDEzbYpOYzO0U544kMveOGjnzknNxEkTuT0D6ppG5klY+0rsFlmjYp
HMqvWwaET+PU9YiuDGZO0YjJhzH4FidF6FM1P899evhWqZ9kY/SEN2XFDJaMcZRPj2U8vy/pqo2r
MMsxBgg8nYkdDFytXj3z2hNdb98ZIQpeX55kq+n9sBmkrI5iBOy3SSmsq0KBG90NbUIY5uuWg6bl
oYQSji6TagYcKYAYklMAB6rR2k9AzWrFnfih1Ed5MQnF4VpFQD/aeUumPRlRSn6e/E2aIUAm6QzC
XUDpS8HacKkO3RJGBwqskFqsngZr7JytFT0/usEcc0aRQxarAnYim7kjEzmib6SgVp33DOWpVebO
B3xj92LKwRyQiu8BUEbirREyl0KJss1ZpXbcM6HaRkFVu/V6VqSTRjFdMIBdqd+XCStrDpVR9nfL
z0zWWVtv5frhiARmkHwzTWMVFiM3GazeUbpDPeb7WLjwW/UdHxvjoNQv6OUy5zW1b2jEB98QK8av
RLwK193lgsJ+hdDebR1la+P+URyWrG3ubrNSAg3xmnsQtfAChSkhGnFYUY2c7oCULs6ACJOLFATA
ACqb5IVNCWrPPqs1FnmLqvuTZh4JKpP80fupl7eWHVnMQ+EpMtLUTz+R5TcjWN5ZLbxu0GQqHGKc
gnGBK3fpiMhAP7wBcmKOLt5DbcqtEai9b3uT+h/wATADET9aLc78HLGxM6DRY9NDZYY5nfwGYbPt
epFhBQV2BTojWIurkItnXXBcR6RgHjIMUAf7/8+yb2bwXxR4gFwIJSGudh9yIm5AzF8v1SnAVEZQ
yA0BN4kA//fN7nX/0PXEz3wy3mFI8fWcllt/WkbU+BVATc/5wcbBoCJp42d+wtEEjizSSADV+CBb
eUilu5gzaNkCI7zKMG2K+pEXtOXlD7PqK1N1sVysCFYZMAM3Q7+XGkUMCQPZJVTWImJXq3YvwtaD
BYraIg3IZarS2spyLtI7B5KzEIdoMgwM1iLPK+Ya3IvW9443wALmIGaObN5vxRXjOZfxcEMfOXAY
PjeiSDo6ssP2WqYO1NgnnHr2Y6epzZP3TRJ7jQ9+lIL+2ZXGq3zS0urqhua5ZDFFd5HRT3WimsUW
2db9/lkhK0AkhZdw+RhUxq25lhAZmQOJ7Cq2FO+5cmiw8Hew6nJMROaOirIUh06+klzkO/WuUBmh
Lc8VeIfXP5n+UXZaj6chCaxxS0AJbe7/hLjwwx9MN3LVAiyEHLcBuetLWEliWGEDrxNHVC6sQMIu
MNkF8tT8AOnEum1bbXQuwxACXdwifSOM3SP7Ai2ri9E9D5fGcWuinTdwNZ1Bqw9hMXURV4d6FZLs
BiDRWgta+Fu2Pe8u5DAXJhmcPK6dDomXlMn5cq4Bvlm0WupuqCkh21iquv/Gbqf65Z2o83w/48M1
+mgQGh9w2LxRMhMITscizGKx1MT9Pp16KX8leAh0ex4yn3zoqaiJSnuDxCbb3hmJ15+lgrYLxVNq
XskV8GXAflS31hK2fwTwM78UQ/T7dZ64e1qXYSrb19upjzivUyUYj150IMYGn7NmTGhB6mUJcSEA
rn0WwOzmKAaSmQzJdTk7fA65ElsjlDGvJnF3cG7D1/QTiV77r7y8JkjSh0cMowXvMroIWiWnSYLs
4nB+7XL2hG2OU+0GVCZBs8yq9FAXnTQ3XHiS+Gmg/TsfyZpX0jDRAVxB2a8jYuywpIUaW4jPo2Pj
D/tRUbWlfTP/9okbnLTIn76Kw5wYLi//S5ui77/Tdu02GF/Xr4rxPhwkCBEY5yVjtfpzb7UIDTB/
BUJgO9LGqWD/87C2nDkNhciPW7dBjMvf0tow8Ty1shZ83yPj9EvPZGDZ+rZsX8XpN/TUSokTO2oz
SgFz/5wn8mcfKZTSWFPbpP/O8qUhHHOCsJN0CbLOooPCYxeFgHc/g6ndpZo5hL8ElEBbZRTg3L1p
pRu08tUGjKtiFf4MC1KYFfhKzUqrk+hql4OyXEENW/IrQM8VIrT6Wc9xrV9ixXXSfgGAwF/sk6JD
9KmRXVrOZNYLg0T7aq2193YDJ2tOLjj1hAYAAxSb1mQ1CzFPDDfEBspo4Tq7vDFLM3qmWMEazUpK
GiQwVP/tq8uucHU9jpraVn/xhnCte7qD17dzVI4cFKdPiaXtDnuP1Ix7Ai9ZNpsUvPUcUge2ZS6j
rLALbc6IG4QDf0SpdKosjl9Y97wsGn6V+VMPgToDHgQzogN+RtpuydkApsS2Mn15aYyCoKhXdu2H
m4WIqdWTUEmEEivJBLr0yqjeFhu1VgNcHQayEA+kkfov5X7JjsNl/8EaIFCwJRDJkHOmLOmlLoxw
jR7hp2gaVT4l39JB3RsIoPSLA0Sd0vOgDSxI8AMMgem2fKqHU1P3jreOBJ09rKgJLePYW7MYtEt2
lr348Vf7Q6sDSLXb5y53bKM0m5xRlCWM+68allQV9c1eSU16Xi169e83dAzwTJJMd/09gTtxZyRK
2y1tT6d/4zKoPcPePcT7veBE690n/blkVKqBeiZKZbCdr2Fr6Hb7F2kwUiCxGUKOSj+4hy6uD/zH
ZvVUMIopoBpcJ0037/1iSSZXQmrhzRQks9fjwVS5Dy3AWeaFo2qfAvsYbUZd+bNdxGz7od2IDOqZ
U043XXl92GcINxtatdqLEjQTULbc2QIgwxq4zLhAjuRgoC8BGnX+cdhWq7dCmzOTGgnktX6BlXI7
iLPXkp5U2vsLgFYXuqyY3PQq76CmNHBl88f9hFrVN6jzh9ZcIG4jRhgGiI/tG6x8PR+7mmt/b4qH
RhI4nRZrSzmvjQaV0ZLvKfiUqbRcIZELk4L6wDnHmP81niVdVQv+mp1/w3l1yyuJjEbArPJUmImL
VOlKQbVrY7IzMA3tGrvNBJ1fw6WOi31WeVO6ynUSu0u3A17YpJBDuvezyRjbzUtC57hHhpB/hmOn
zqu/nFDiEIXKj0bC3JR0zALNkCZRieOKL76s9WZiOz9KC4CnsM4c5K2RwrjAtItt+XE9AV51mTLr
eLYOGS3+OM/HrpBeUus+n4xd0OKCZjc2j7l9ia2d9DVlgKkkMRDPWyCZlG0dT6ZbQKu8UmhO8d0C
fsuucbZIwRD51XQDGWL2M0fozpbIWhi3lOxqYWCb57ixCOmCYiAe+ScFp/s+ucEVXOfWEUvnZatP
JdtLRo4VWAICpSavZ4Vk+G5bXG8jlY4+Hv9/tck7Vd8SPmj+xVEJQ7hmSdhwvEgQpylo4qDFu4gr
/Ldfc0q/i5iADZWNHHxzISbhQEXc49z4pDD8LuYP/T9aOn30lNv7WUglYXvAnsYTiLvF+AW3XVm3
hdAV/w4ASUWJ9QPQLf6AujhEVVtmFkNxE1/TeAW6TlMTDQokfu6e3ZSAIkuKVQcJyQXuUKhaQiIn
3+zzkWCKA5u+vL9bWCSDEZ2JlWex60E5Cc4jIW0To1fZS1OY8Rye1uuZz9ZueIX6/0nHLwO/wma7
3aiwGTYADgoS8YYmNFoAy+moqiwxL2oU9uwS9mNtj4QGdac2XeqwRDzou/HBFcxoHEFOkWHNPmiQ
DtTxl/fUmCL/0HIsZdDOKauj7Q2Uh1UvveIGO9879limGD/ijLonP3z5fAovA2Pe+wAcJQ83ztbL
mNMBJA0xTKP2pqO0YvBhEcF7lKA6dCrTUaCPDRlX5NCFW9c1swC4uPicitGnqThoihDyYNamditZ
tHQmYwVm79g4dbD/U6MsGKKIoEdiWwbzWByDvn9MtJebKzYzUo6VlFQPsnYJJI2cSzHfS94gExZY
7G43zQlu9UB6A7p4ttyfC/7Ve8PaJGSrl0ZF001pb0DFHV9HUKliDVOL/HmMk4woFnetUnBI1Vqo
xfyUkqvnZjSOe79wRSKcYMQryWovrNEhmNTvTvc1XRk89R43pAp+6ZxgOYkzDCpG6z5OcFcqxsgG
Dw4X3rTsVnM6EgNCnZRfMFSsui70KDleCpzTZtReQd7SShP/6GaAMtiunAMi1R0+3GzjOK/s9USZ
VLyMxP8bizAiuQqwbWlBcrRAoT0kB0Bgvooe9RhzK/dmFiVVxTeONDxKMS458fiaYq6ds8ICTGQN
p0lgJyfP75QqJXng2qJUjLF7Tl1e0Asq1Q15dYNLD2zuWQVTRere9Ct9TZiEMHEKsOdEpLkNKcKz
RaEhdZA54jrVANDFdE17nPJQt7wde/MCKSGe9diW1wuknz+sdAhgm3GLn+sgPSTCz7wap75bRids
C+1XwL8U0hq+y8EuG7zWmJVOiEbOcbK8idpiKBQKd1K+Hbw+2nQWBsrwtxuU5Ex+VT7k5uhE1840
zFqiSMgzX6dyxAlEt6fybiGZf2+mH1xtfhuXRABBpoedXY9dcSGJeLvQZWgblrBntvUHJtuCe9Ve
+dFw15ngjRK0mcfkJPsdfunfwYb80ZRm4IHpYJqvkTu/PHPiSh7Ino/6KzXEKKankPoC51mvPgVC
L8HM4xKc4O5YswT+Jc01H/EPOqW8Wrc4oM0gNOvql6ay1YxsYlwPieYgQ8Pt1HpB/o1X0Ag/Bucs
hj6k3oTIa2qtsX2SHjs6N16P5vckbs0BSj+VQEnkTkqrqTunVNW0BBR7AIyFY9CVclEal3oAri8Z
/ZuVil1X/zxqsBeeb8uUWJpbFEaf235zbDwuDBaYan2fhqs5pH50Az/nhbfI+CIAO42mAFdytoKA
yzTZcBrlqqNzqAqcKr66Yf9OefVZofpBb2RCqVEG2Ec0sHy7w1pfCSPkonkEtCdHx0Y4kfgyBrIz
7BWCToWr/ggrUiYyxSa41a/jXK0QCNOYG3GcyZZmxryC59jR/Mt2qgpzv4Q355lwylDa2Omcnp1Q
FNo60iloFQ0q7PcDRhzDAXGd1OY711K/NZ/fRJVnzdqAQXUbqywarmaf69yGvBJWq4EJj5OHU4nE
aCVq5Ar7jnIymQSo5g2qD/qZqT3Y4xfZOZTvTKp3ZiqgxtdCmR0PioP5sbP+JSCvK1RCfLVVh552
sdtPsGN7sNta+4cSOei63/CYfoKE5EI2OAvnIS9LneJo3KMTxQze/Opb6GITRhFK7y0L95PY9qy5
gRblveJP2+sZGYD5xTJqXuP+pozrKmEOyPkQPoIhnzu0HVPp8KcNya5lO0QVdrpi10DzhD1wii2m
r0Gm/pCtmNyWpZWmqO42LlQuIMe/M36n+7ETycnjUK9/vNnuoyQzYWEssTMIM7DXImEfPVk3IyHo
YbmgIutrqMG2ULaG9aNfMR4ujkiq+Evv8TEZ3c7OgQGa/G7avfhUtLMRnGXJw2YjI9MMz5ktHc5X
aqdDHgg0UQjWFEbTVD2bRnYPSl0aWDC9DoAG37XI11G7kA42MnY5HRxRMb2xTRQaxa8S/ClZaM+8
YEUarlMvCXi7rpPaE4lTWlPvJ2Y/I6WRXlYmRhaRGmwnXO36QOgIpynlDGCS8/lbVCUTTMnNl5zb
nyaTzf12z+HjEDuEy/cMHIC9kdyIkxcgqrCgUWShK3StfGYdhDeqFWvEW5sEDcOGKgXAOVRroulT
+VIg0wUgRR2QASCeFUGlWLYGJjIuXQugiJyg4l2+nBrGNp78eGpILIyLGb5DF5h8nFvU+qZOE3OS
Or/FjuPPwBv2U5I8wrE8/PVORjC2hTiXCi8uQ9Jy0JiWvVcLemvdsR8t36dqIq03MCS3CGfH6dnX
sqIaMACrAtSEJZcLFNIzzNzsK1anFv66Bu/JN16h2mMjxIRlK+gaakVeoqgqwxYB0l8lnveOI20M
1m+LELf600AJxAs5Fv1rM1/tiLEMbGVEz8F3tzzTW/7ed1qAWM4shR7fd/lyGv/FdpANcfzq96RK
yM1DObBcRiSok2IMLAZfNRfArfcllegnJ24OllqSQw2rOZkq3o5xJqDanXJiG21cNVxv/laK5COy
gUOtBE3TtjabpNw3MuI0U6H8VufWwIBlHQjbfirYG1oTaMhyqw+nSRUkypaSp3rHlaWKStoFYNUn
ji9MUHsNlMVqJBg9InW2a5/CgD6aCbHiE/Wb1xLOZRk5xq+GeAm86PhAEv+yO64IDvupv+w0J5n1
o+0anUGRoKxNKc6mV1xd+RbQC9Rmc/ouOh8buVhLasZf+kxktvvF3zPxEA3klcoD2CUwdwBPYJJT
9EYsN5vna7wa9P7H6gz2jpNIM3REw95aJaIPVRG9m3+lbv8PnS82SYqKy23hqP0Lvu4AxCyU6Vsy
+SVBsJ/n524yKlrTJ1KYb0TGZE1i4rDNB42rlu77SL1QONt2G02PGeeg52dHDdVqnLUz5e3J2KW7
vGKz6hniXu8gizJ6swEBh9c+OBm/uBee2w+Qvr20SahVF2t+6H24LiYZPkbgOT0w7jvOm9er4wzT
TNIKAtFJXPWi2F8Gg/fI0Ku4tjjRR8D66VaGAOT07KBsbZH+vOsZHud58BvosEdLNuNCRwNRG6Ju
cHy4o6oDXcnqSUMdTa1TD3E/8OqXPZ9AfENWA26l7oWJpTKXzf4fO7solcQvtE/VCFNPaiX+Lgh6
oHTjRIprbiEsSUd3DnWNxPKQx1nrw/ew2grMHR+i5rwwwFXynr4CDKlNn/0/aq3JOJv8CPvvch7W
2l4QH7IAD8upUWUFwZJJnXoJk/6+zhkuIEszaaRKFYeyjhE+KQVZtDkqUazi9Cgk3RuyCQR4z0vY
KAhrO04QOJ6LwKYv8umPnF6bOKHO4H7QUFVOhKP+Wt7o0xvoiBFnFyGZGRXzlMVJYUdV93KelAyP
YDaor6uZm+ko9vSgtza/PZTRXU28cSN/2xFacDHDG4I+6lQwaP6AS6KIErVqk70WiE0Ci6UcXeIU
N1SlHrIFO+DcnDxl53wjzsdHLJ8c5Dy8b33H7X5b9+CmcFyjr0nKKCv4nYgLUg83AgDkiPiHZMiy
DCvv+rx/jxHowhFyrjkcUu3aR/mAdgMz1l9TmyM9MsNL4goxsJU82L/JP1Fwofrmq0BYLOpRb2HT
jGPMb2ACx42wq/DTZdYTNLHTBGTJJ2w06LaZ4CEWnWYtSulm2PMVrpcbIwanL721vPaiHKPBlyOm
wjpadUgjeL1z/rcqsnEySTdLYevh7n0dtjBzThjl0on8sPRbZ9Ep1HYYpKUS3/dazL/66vAAyW8k
9WUJHA6Ml+ilmaypyDqyYQM7He6mYwLRtzuyDZ4TSWacxUxpKYaMWynvCiL0TbRcYHlZVfivx+ux
DE3inKBTF85jnZM0W+/zlzA0LxS1zoozTml58A43Li3FD9Fryqda/ePsViKiZNUKmIm/0EuLu4zl
7Wq2jYTj1xb7/f28IklQxElZeS1cyi98VbhDatE/l8EYLHTiInXOH0FVkvMF6wXjRppUlp01mFR1
eH4ROUSy/Pgni+F25Du8wiuWYXkSFDEElTs1+Fh1eBvPrhRrYmeRS3bZ48LJySNmMULRgP8K7cNA
3BgTPdHlHDCmWXBHIhdDDOf+XVvauzXhyZLJ0vMgaclHibNSri2ksggbA0a0UmFEglfAYYTrD/QV
YAHApUsmgWHqPtmN5NJrtJBGfwVkUwMUxYYk+P9uct18sO1XBYMkZR/147mdHg2oJw/rQt9YxMIv
wj8rnVDO42hBQb3dZdfjFGPrH/Dr8wQKgwaixiBmi+fr4KacmM+aXyrZMpjNdpPGbF7d4SsAVM5S
qhmPEz+eB9wYhQrAGNMCyI+Pf4g0/RyXFQddolqoJkEkA3PBvIQ0GLDBZ7ic4lEJKm1hscko8ARJ
+F3he9iYE7QTeda+EHNAVOdb8dCZUzMpGbR+oi52vLKVLcqOYJ2v8x3ifA+kz3/1ZoC0OwIJGpkx
ALyrut+GiF872gOaphF643hY7HONQjfD0pkhrXuO8UahO50j+/EFq0Lw6wE23j6Urj9fOTHYb8rI
sVSSCX5JL13DX9IYba4/igiEHiFcD3GHI0YKJ9JJdzvurz5vMHKwOOzjxKDEfhLKIBo6jtyuBO9V
c7nRszb7EtD3uQK3DXFZoRyOETGvmXp9ql9mM8fCWb/sG/HljD2ZYHY5fOEuQguitAxXSUM8saES
sm926m18IdE48wrs6xp0rbX1KZT03vyfKaBGq4F4iS8wiHrXZi2m2u0Iky56kcaeNRtotlW2dABj
lEeElxKbi2I16hc/9hJGwPZkZFIIGIiXFHd00wKBE6Upn4oxIrA+qc8MAxXSFUqEeuUyrn8f2ab1
8AffVV4zNqrXkKzUqt+x4LotbR1f4hjiGXmxWTkh0f8P35zHtlSbTEzEDQA8XpJQ3iaOznBP5bvz
ULko+74mNLpOQhwXyby6l87Bm1Ex3+iF3aTxVErtfs+lyzhC0bnNX4KEfzEUQeo11KEm0nclaoR6
1Bzdt0vujDpEvFWNYJf+3kseOxgfKI2nPAXqZd3ZW+PuHrl86LmRDBSCddeGbiq+PQy+LWAntR+G
bAU0G0vMl9bCzgMqNx8k04R9kVCQQnzXrWYTlRrRJxMFUF5eMzn8msuV3cC2b7q8cH/dPCvNOnqq
iMwgxcyWRYZnMyirgaP2EoPgeoXPNZQcofQ5YEQhpxZbNrlegKSfRNpMRrbqLGQrBRIQJJiSjAN3
WGSp9dy5v6/4MOfqsrwGXmk1HEKeGGIDUpDlRiQiiVeZ/x4SVoooQo4HhL0m8aXajO7SGn3WRX4V
4pBDUlV5AamE2X8Fa9NANVfiZNQoxNW3wYAiXejifo7K9Gm8QAcBT1j5fHwTqbxHiXaDD47vLm/w
uBngnoda+DbPeJ5LlgTiH83AYQKfmQyNQrtlofpSwbVmWKJUKQMoQOLTE+mfBroMIFiy8mZRm3gf
nRR5ojvW5wWvjODXroMiodx41tUEIs5GLP+gK8h4eU3aSWPeJ+kqPic75VWYXliBEUmH5y6MyWa4
F2nvNMl/3sIDYGkCTzaFn0oCIhyBYM1NNam89Uno5zJJ8q95Zt5IC48absW5Ikvzf2is4sSA1769
M3Oc3FEEZOl7xIl3OTju1l8WEMSlB5r9CYaRaOVjw9eCetV3fbgro2rQ8hD3F8eo8Cn7cM7UO4J7
Mj23kMqOP3uhHuIHb8dt03rkewhmgvfdschnt6eT9Ooou1dkqRnWnVb1FHpDb8SQ06JYjPA3xexE
p6HrEfyEQ7f5np78P4uCdWPtC7XHNU3N0B8KRRdNMN1vjFD15U7Lyj0vJSVhssh40LhPBR8YgjL4
5TRhi9wRurLnz9yXc8QQaS9YuHNmUPB+9QJUEVFuyN85DgsL8YGDxZw10qZMMrQODWYK/mKJdP8U
PpVIEEbDWxcAIAFulDOn5Bnfd3kCWMFp2dv4ec3B0Xkp/2xxYwbHhYY2TrR2hNzwom8hBwXN3/4y
J3cvB1z+Ljp2KLk8r/e1e3M5AnL/RdtVbM6RBk6px2AJprI6CQ13IgWO8Tb3w0H14OMyYX9z5tr2
x0mbRNiVP7LRHXcOeCuSyDkCn5vkkKABmZ7PzsQqz1aG0YhvNjfbrmleCBAiu+p9cSbVo8OOfr8j
oq6KPQt5cf6EPYCWbAEl1Bpi4QpWwNEM8a29lCtNK4Ew4h/S3/Mb1V7T8dOYkBj6stZMJqO6ZT92
5yC5/cV7ByGJBDcsElvbSEVwv1/I2+W6oxvF8zgI2Vhl4ce1TTpE2/cyJwk0lRiteYPMMyLGGjvf
wVBcJyyiOBfRNm3RE5kXtZz/5q2Yo1RvhOFdpB7+d1E71KYLyEX9/2HhT6TI47ZsAZlFo/kDD98S
nFdRquFl2u2Dabxxww3A54ZwI/uGFlnS1cK+3SSHaTaB4ZQs3iAG9yFrp99acPd5uHTZ+uEQz+9I
YMNdFOI5w6FvG+r/FY6MuN8sagg8RdLKyV/HO/+BBkNYaacY1fC+yF0C07lVayR1XgDW9UjCnkvQ
dDSBg9Rn6TK/bI/khxCmvNU+aeHjW0JYLwLhbpCdzcvk8nZnQrQdCKTXjOLO14lDdJfpxk80nl+l
QDEkKcPxNo+WkHkb/3rqZv/Ezyb6VkHi00NtBuTOe/1v1FnmqCMXcTCf7fHOSIuwgwiL57fDapo+
ipTJKUgKgjMalFuo+a7TuCemsjESKmsLbDggUhaxCKHPukyaGXRNb/LNvbRo/ZZlDDblhvhkvjAn
KDsyBS/F7jum204tHPi1P8sBTnNcqNpJnJhMOfTai/oGPKG5vV5ji+QKRFbH94l081voawdIiXQ7
CjBWUl9EAl/beA4+CpRj5dyedipzxcQ7q6hyoac8e1ent8KgXkcTCPSo7TABCR4YwsDDTaIZbnlv
IINUjf6pSvLd2QCJ1ODpuNAJyttAHAmXv7k2CtU+es92O45cHEO8YnEbW3TxnV9KhigOxFTAUycm
wq9RAcJIykHE2OXNAz482uJGy+POtpdsFyLoXoQCwZoUSa1Zwx4+SbwqqQPcv8/Ou/9NVHxYG6xy
CWsv4uTmiH3sx0ffSKkuZeRZK6/qoUcSu1UX+hCz/MJ6AHUuCbXCzxGiVdTuPgP/RRkrrmjpmTAO
NxVi69v0e+6VUZ5rVwQIN/7YVGAYOA84ps3XnXFm2XGOZJK0N1N/tVUOpv6yfQEuCRqYmCNTFJGW
EiSDyHFus4W2Z8lB/Y7Eeb9YLioXjoVy6wV6SA08QSZ1Ok3O1+1VgTC5n7imehscaoEQ55QcIMhG
Ec5XyTkDdFSnNPrQTMt5zRIQ/oqUL6eX8sxuQmU4+a0IDlPiHsDYpi69C5/wZQyh7SE4CFT5goQr
kwFrTp/aiuYuCRQVQbmTqp7S0U59EYo3n8BaWbdH4o/ROrm8DciCfLsWeE/UpEcrtrgzvk4lhMH/
T9b9mwRgaNVDadNHFLULKNz0eh7io81PGIkpNoDbJo4I2m49PNG7JMqOS0rFGFvmOetE8UEOQ8eu
KplhMOSUht3cUNSgg83v2sdVJMC6xoLfNRmbCKrRy9wH0Ic6XY1ocBcVP3s7nlHhB35W/sIlsQcj
LbNT7oaJoq+NrIhsWQcNBfzvmccIBBBcdKydigPeaz94LF28MlxWHe0xkBnLy2GRHODAa3/DsYZH
lW6WP+qq4ceDrI5s/AHFLdr/0axbIYA0e+mhQ9CSjIO7S6GPqRmLSesdGdEOKVbsSgwKP6hfFJeC
Lk0jg9l0a6AnoUHnqx/Xy59tgEAB6UOcSCw2ehKmvXaPy+dd5IqxtDe/T7fmbFYnHQBYFqLtcPFA
ZOwyE2S21Eujf13SmZApyfDmtbLCcy7VHY7+JAgG2huEwZoZ0sl7Y+Ln7GzGIepWB/QHGy0PQN6r
qmxtEMIYBBkuDHitpbkYePozvdLtQj6+srRhNEJgSJd1te4nFPsCO4DeImF0WbWyr0/noeLGZVJb
8FepVbHJF9wK4vjMXLrmTnvGnmWRmNxH9BkmxkUlrE5/6oZPTj3xa55xD5zuthkgUC5G1J3c3YuP
SmRqXllRyEks+OgY2cVFQxTNZ0bXlc9yKByNr+47Nkb1XgzZhUNFE3LMsj8NtO9Bl5V02NlKoV+n
wR+KGdDfbuDTxd/wag/0THI/NTab6UA6J92BM2tbPzRFBQrPIfnmBQ99JzSGhHTlh0ctgH9i0dnk
xqYDF9JYRAXC8wPvr5ciWeB0P+kqW8vaq40Lfir0zVG+ku69fc0GGTFPYXA/0lVkXh9OIs1/c6ee
PdlzRb0RbVTPckx8C4ZH3TiULoPEwIjufZnYayAcGYB5vNrvHbokKb6RZ1IBvR6qzeMFB5wO/YWJ
Isy1jjzEoEygbPEW++aMyvQ8kww4O32vzxWafrfRqkyXqqkeQvptZMZkq8HpXDYFPd/4Ot6hv2P+
d5yawauFLxd8h18Y3h6tx2+xI1hH8ox6secF0GN2j+fxCaWqo+zqYdL1VWFlDB1VOMG/NmKp0h3x
mICC8ANg9wQF8ftkXGSbCiay/L7vVtmm4EO/s8K8ZsQf5PW+hhRrSiZ4NWsn6fvZ/3HpTMDGf2jS
sFB6GUL2HjpBbi9KRYuRfW+gEGJb6Isr80aEhmfOVCCmv7flz6fKtnViLGrsBzbrD+JXNn4Y//EF
saAGbDtinIfId2cL1IY4qJvAGj4pAh/oob3we9QUp7gFhFMqmwwDO8CxGQJkxIY2S17SmDvtQUzj
ok/BZOQg2CGIy1fZfbneQi4D7YjP9ME/glQbi3eNyvWPPf3U5koUd7WAf8FLdCv7td1g7/HlAOJ+
7GtY7CWPE1bHX1AwyjsIhSKjfxf3m4jgeBidcXeb/ZgPSlenxwPn59DW7j3C6YBkh/1/nn4ZG2dh
7UY4og5vdB35RSEvkkhrF17o9OqkK+IQmIya28BDSXyb2rUuimh7CpHASGJUNMV41dUjkAdR9XXL
rVXOKRytL5JVRMaf41imdN80bIxhq2y7InBD6efAGhqA8kQGDtEoE3CK7I7FCDnzpxeLKcZQiaSP
BRTfEmQi55m9Beg7bWS0Xr+Lm8u2ZY4kFdLoYVnFLHK72QJcBx1TlrYpCzoHnTNunbPPN5INNIi8
BsSEh0odTU0LIrdKZAyIAsuUpx+f+bj0IjX4nrZvFFi8CxrScBVeTo3mbk/nomxAu8/M6JKnE7ve
G9pRD7BcMJhZH7PGGxBz1TyfraZ7as2+X7zl1BYWzyQhJALQiWOm+DTKKGlPl6WP5b3LmBln4hWK
PYgh2OunipDLCAOwDeKKn5sCLz45m1YyYG+oIpkySMZWEy9ET5CMjbisP31SjNkciY14RY42QtcK
TJWW1pIMMNErED1qdO9voSIvsM9Mt6Ea+brqPlsHWwEjjRuMD2cmLA3IB+YGz7mYbSWKLaoet86M
KDky0NwP218tRcclYdkiIM4wlETUOdjw5EVMvm7Iv4wLPKwbu1fdVGs9y67LT8oV1sRffvD6bvcn
yz6ehYskNlrjwbIDBBiAgSPDbiPm++PnQjDxnBcElJsOgp21VTXZ1abrpZQhBiQkfJQnbYXnLZK7
iNLLvL/Jz+zCPbcmusMJYKyeUrR7olDilehksnQELMjX6g0pUMMJVxe0x/Jn2K3RDfuyDOyHPj6z
FmSKg+MrvB/J2BGhpqsuGnweuV8csbem82yNEacWtX3XsLH/02UeKftdvlOrz6gcQaCpcSv3yyPD
NbLbfkG+lHwdZiUG4j3v5GBsgIaWs5bTkFuJPP3jVtX56hCMmSrO8C9VKZRF6EpksB959TjLUgVm
gxuaWYzh4xLU3W3xBzwxT/eBkouMY2qk6L0xE95VveAqr1TlBIOUUX0Mc7rYqYtV+xm16qmmP1Dc
UiyzVuIO/MPNdxdjeD1UW6WWnVMHbrJQnEEUZ/CaQHbgQeLwIGAOyvhtTS2Jttt0HSMaYQIoWKFQ
XLLtXmS/nhVhzVLNIVp3d4glcH1bUOs6KD3DfILAD7WbhKfHIUDknAZTMmtHiW0KEJUI141ZYOa9
MOBYmjmeapSUTerNgFrvgXdTGIgpCYMoRg5BYt1QBuhjDd1lEywj9yZdePVReT89EnI0FAul6jpS
kuHgjj2SmzBA/aaO9r158rRZi8ojqifJKedcfJc18wFql0BjTWoJ8hhksXv/Voq9Ck5hR2PIMN5/
R3esmElkKcBG5ez9LmUIDzgGb/BJEFaJ2C58TVRDAbMyP8Y8OOBYVK9o8cAWlqxtRb9S7fF1dtVi
yEetWfj2ZFN2+Q0sEQI4LN/pGuzi2qEN3o0W0ahHF1lgMrJMDTq2hYIM8xFpYgnjie0okbtTY/S/
JvuTsNqs1WH86Oo2kc468gUH2xGb4I+3jkJUpRN3xoonjxtQiGcxdZxSurKSbRMSTfSk5ZYikVLF
SqWEVlB88rJzUq8CWDgsZPZbI/woS36PQMBanBegc3UIxvsG6TIZD6XmeEg2YBAi7kfD0Hej9ZpK
dkERHMkOdN51NY+XjG24gDYvkiZQLnKehLTJhvFr30yi7ojOcaZQR+Xj+ma5i+VeDtMXulqtJO6q
L/E1pHpGIOlqjGFf7QetMwAQ+o0fv37Uysp0/NdGvvZP2vZGkCNjctwlxcns0Kd8amFngI4prAfI
9KDOylMedZNNvKNBgGb7hIVVexyY80nY5vHlQb62jU3enU85u3VgwR4Xkie1Eqw8FQAeaAilhqtF
znH0iAd/FCjoFb6Rxkt4ZcdwA48z5lJXKLbmtMkCW4+1WiOlQplcJXgdhGwzLw3Q3HD09TMHdG08
lgUj/K50fsueOAXq6t4mAWE9jU8+bihmTK5qdmf2F7/PQwckV9T13HKbXGTsZvPFnXq/nwCO2uAs
n9bCSPtFHLfRFU8cYH/wMrR8jcdmLgO4P0wQOZawbYHxa7bMph8vdmW1ke7/kfBCAH2vzt62K7Er
TRxd+jeWsLjR34DQX2xagtYVuuXdxshaVO3rC/L9Z6TEMxhUsN3h+7WGq1M98TpshClB4otZtcIO
1Q9o9t7WoK2tPKfQ9KCTx4WvegRetvWOETkM1sA7gezSP6CCjIX4NZbc6N46jvFuwOsWsPJgGoxk
MRAKn4srXoTSaR8Q1uF75wsAi6NiHdICKzNQoKH0qqF443rSUf4m9C8kjrRQXw3ELtG0eapFGMaq
xxnvxFfUHz8PfJ9o8k438oedTdKLIPQa44jyT8a7AyWCJMRgq9TH0ZXb3WQhfJw/U2wMKZjhnTTD
G/NoqdtL3+4dSoDIDmlcgVJeiSvTNTeTvzRlj9lTBuTBzT9eNpbFGXnHIO7jP/EOT1LLzqfxYJKV
vQP9b40Wg4g4wEa2ERVDL+XTGYOMStsPGlA2DDL9vfH1nN4YVaPvP1zgyGg93Yimv3Znr46GFg0m
1zZ0PsPeqHd9ZkEosRDzzAaVfAPGA98niwfmA6pk1vP2t+jW47PnPTTP6Lr1yrSoDcUMFAtclm2C
H9n6cfGiwiBrDseq2Y8JDQY2DXMtlhdImOMuSe0q57xfkTnE50FLhEIU4eeHUIl/DiU1gvbhMLyi
gnMV5v038RDGPKWOMNKeUqyzyLlaGeCmuwWVdEDelX4BoYRozyI9+fS2AKB58grgE0NTlS6Cto3n
db8gy1z9nr2zZ7cm2ydXGHHftBgESk7S9QWAcS9bhi7HJ0WVXhO0A7CDRWs/EPalcxMWnl3LGkt3
GsnAAgEjMfWPBeltbWR0gBxYoj1vhkyDaDmxMAoKBETir18tSAHRwtzc8ehzhsWzlEjg2/V/fOFR
UWsdx+5LU+aCga3m8YqBKMFJYLty2mSn2NhBGzBt7QOIx0qdJI8EQf8euzUFbTM7LZ8pEr2Oac1B
KYmt3ef3TnSPVWYBzaOYVBbr0RT4prJA6CIRAfjzZeDHElRb5J4C/YDQlQQ+7dRuuK+EomxiPyeO
9jAvGo8EnAYjbUq4WLp3w5GeVH8cX6FpbarlULHas8uG+2OYQwqIpSm5FriBqnXNvuUDnGFl9PWY
g/XVgXLFcxrZCfDaTCy4wOkXZW97pyr3rrTKBYVRKdZYSfwagEq/E7Ut5ncsmLBWRCPHl5cisl9c
r7CXyZXu2g3fHfRIHJqGAY00YGIt4lZyiwOzhPzlpTyZgqXYmbSxhbRC5dIrkVbu9yqGyyv+k/pc
LTI6XE0XfriLPnIGJszjYC8DJf5E7RNavukDpTaDgvVMQoLuRM3DMsL6jc/KgSwvm5xJJiL90Ow+
uUjOOWOrDNYZkCLidb5o6UNWEnwm2ar6I3BzOvmOch6xT760ZZ2N5SohCWkoHJTsnyYZ/ZjdnxTa
yRAxOqnuslUeSN3ki2Y6ey+HTkoeaED2T7QAdpETtWhF0g5F/rFP7+loUTJR16HnmnzTCs7Cq47H
ws1tnC21N416Wf/Gi41fNySMiBdTUTHSTirsnjtWNvfCZy3ClTaWzabac6oJ/VgLFbvc+57/8Hlz
/YnVQP0D5hWdmW/AmY6j9xZSeoGbanIfXuYy3tC8PSG8UsbSAzTr+INvs7XVA2CuL0NiAvYNAIw0
8hktz0FRGqzTUijHeCszFmvkHrTJQRIJnrZLo9ShBEoyVSyGCRbM03SplDa5sFLnfg/b3Mzbxl+B
+XH7soW33ICY8755KJaGmuOEjt7u+I4FHGdV28TFnOv5prxTqe2/ZvMRSWuLhVgC89uUT/BrFLHq
XTl+Mo1RR+vLaeKV5UZ4nwKjgFQWw+wpZpIZbGwfPHVNI5DoZyKqxcSGkNvf7IyM7FKUk3NUNe46
Ob1TJS4mIzuXV5XJABOH54AGsf0ZyH269jYcFXlga6Jin5wTaxMXdBaGR3y2+dL3bU3D457782gI
j00q4vs7zb6qPxYfjkgGRd8n0q/156j7moCv5Fx4m96AnVA83b7Dbuy4VICZfBoBgZQtcV1gSOVl
pkIP5aVRnKJ3PxA1lbjXK3OnzBIlHGiYOsbI4aVKF3w0zxolLxe99yezv/phEITVZNu3Qjfrnyxm
UMr5V724bfzSACmflS12voXaU82mrIv3kgumfB7foGwsvn73HHp8tO3nxB1zPybviU6jzo+fC4b2
CLw3usclJBeV2uyTecHXoNIIHS4KjzzzWBwZGdSSXNsHOTByzFT6AIUrUzr6BsY4sMxc3zDjdCra
l0Bw8AETt3vQ90qA6Gu3HokY9yL7t3+0XExsO0g6Fzu5QqN4oJ1SUmnl8N4N4AbqiNkKW9+APFjF
b8BUlQ8BglYeoxkHUarI/aBXYSlO3dma21jfNigd0kaDnmIp5c7f55i7AtcVmQKbL4uEuqzzDyBJ
n3k1W3/+WLHPeW86w3dIIWNftG/51ffNOcVD/E/QmiVNlqAOxFE/yXs/y8UbogJqXP9BmyLixt01
he88XJjtOTzd8QxH/Nz8elSedgDGrB+uokqbbsNI90dvpCBFESOP/2kh7RZvTDnhjMzkVJ4qHMO4
83BpqgiLwryyvE9SR1eMDQQrXSj0bfTg8YL23KHc7Pcgxbe8FgtrGH5JuSlo6snD3dH6VjzjpIsO
Q3gt9UEft1KZFOANEEEVeSTjvc6YsymSNkjsJl1Oy0dBnKO82/bOGoHEWz86AN0oX1hOHwtl1cD1
q+i0/WXRAdDixjNmJjdPMW8xQpaRReV4vo4wGhSRFC+hiuChECzaKgMO57MoRPqD2Sy98AYHi2VC
hG38ixnIfR9N9zmoAcGKyBg2ZiE1odM5S2Yu1VHE96LoWmhIgZaDd79VvN5ls0w+asteFqXWZogQ
POSnWx0c0inDPqbwQOuwK+94boE6WP/SYltVOf9aITA3/jVu/dxmgC/yntswtYKvokX+v6x/ZeBM
FPQh1dM1pJpf8Cw20iPaGS4Rm7loQAoDODuSR5ZMjYLvA/BtXfSwBjj3jENXBVJgkrjcjZjSi2Jv
fuU+76VTsrOuCSDumApRf/WoaalWza2CDkANvssbgY2ZOEExt57UwCesRtbTvBDZ/Rci/8vqwDv9
7Rg+s6K4+NeBnVcb97pcysg5ndA6BUNSP5RZ7ITFOwMWMLFKLgpjKm+m+D/9b87drctqqHjS/rzE
BFuSjQEfqIQbrhDSOAGz5mvtImsf+jAp7G7s8yZU/tv+2jcssWz/KCCbboVgnTzjI8E3G5YxZmTa
CrX/tJ3T+g4WezgGVr0uKermB0DX7PEpZA7ww+mPsKajaDKrDUgRvrSc8PK0+ORByIFxnbMi6rEp
dxWoKPL/QL+GOxmDeksV+YMumZcxK4AP6VAk96KcDSN5Hz20QOVxFhP96sXCa5U73Moheo1/qYgd
mPATT0dR6qrwUqMb+b81nIH8V1HMf3I0388GZQg6UQWZ/T2W5Ik64O/ahH8n09OY8u0WqNAMl5wh
+rIumtTuxL4QpG+T8oF4acqT9C/hWTV9Pa9RbrACdLJforro3qzBVv+ciFWnC4Z7WHazVdGtST9X
gdPqcl1zgVugedhAIWRLYO97h6aam0uzF4XbKkptywaSnu5nR8afXPMEm6buTAn/Q/KSEcBEdzep
EbbrOOtQzqp83EVotd28FsIWUB3xR8Ac4+uqu+8+4g6KxVRS5Q02M96efy2GlM4krNe6FLxdTBNi
2Ont9CNQbEMRHG0KyUJJvwRcBCFYWsld4ei58uqAX7yceZzhtkpENUW+4FQk0yz4i2s67lHJKNVt
TpbhUUXXXY2bMjb1bMah3gthYRoQIhMffw6af7OxsXuENHyHTXhK8+68V2641rEYWf0o/LthD7np
yqgVt2Tyj/Cqfhpt5BBGBqTVBO7ZMd+m3I6f3DL+oQPgcUKRRkiY7hizYVfCBsu1P0EmvTUueCBt
LzsnjIMuDBtmwk47mi9eohTGYEvObgU6ChjJXGIGZRctdLlB3+PiiGQxyU2Ztb/MBSW/ZczGA5eQ
IYR13E33hJ3EpRkTgcxgsUdm+9O3KYscV70zAU4PiE7SQmG8bJj6AUZY/Ccn+/bZ6h2619fTCprL
mONO+eqJBgB0Y8MWNhgWxA9qKVhnFulSPEMx8ZqAnQ4+dAhSXVPFhaE2y8Ek00Rann9Wo/XK6PXg
nINr8rj67eEiilm6WdueWQG8wvoClP+9r1xd0rVEiV59ItOIzjiPdl1ZfqopXOjePQEXSQsToMyD
fse2BlYa0T/El7e/N9+HgbNMmFPKIWKaE1GV/e5Z+JkdsSLvtDq/ZhaIdJg24U1gZ+loAIGjPFn8
z6lAQSCtQaoGDyuITaE6hHwpEYy19EvgCFhjSK1SpxfS2QZSnAR451r/HsKNK68kYwSb0uhu2R79
TS6O8Td6LRzD+FhmmGS+uf92antyhonY3X7l1alEV5zbdk2XQ6+EA4UbCYr/OJe46akc19m8eheA
78gHOcUgdoMBcKpvzkj/QWPaNrzhZU05w1iVwrStCAYbCMA5I3eusBbOVjWGz0jWb6sTLGp+mGQN
SNqwpbY2RM/dhVCFbcewe44RXoyvEbO+DHjWR+CbxgCQ5RXznWlapzDo9cbn940YnseRgO02ajaq
846pNX/bTV32xQtZkXNwlwANDs1oAFiPvwoXdSG2tE10bB0nOLulNcb7+vt9c81w2Ty4rNFGBR+J
ZYXR7X7f+lGIRsFCmwpZPPhjHOevemcRFymeSIFIVe1JA0IwCsQdSHC63nQoWOPPrXgVLDd8ys6H
wYyh4szKe8JL1ity919r4MgfAIpCn5+26jXLR6fZGVOCFq1tUAfbJHA7lIVa08f41htxH7SDxr/H
1coiOhZtcDgqRmVRv3SeJ49dw+nyBcGJXwECciLvziyNyhZr9Ecb6H5YHQtKk1amBwy0mZd6o65J
2Od9REsJV8eX1y3e5sL6YS46xLc5GVVvrWNf+GeVMH1+FbKoxjmufcT2SCjU3Ar7b2Zpvzr1yLkN
5d87qllFcl97uxmmYEXzzcDe+/dHksZijvM6UUFCD++fAjoXPfLTGvx05s34SDscnIDLKVETgQrR
vmLYls4gXXkhBQZwwCbHLM6VCHC3DNNY94OWKsdrrEOGNmwUdVxsS2LQYZnxL2e9Ahh5GlEh56XG
HDJtkiCX65mB75jr3EeWFr+rrlUcCa6KjX7iU1617ACnUnmdcJxyBB/CiXWOYAPdF/QRNvqN0Ces
M6x9UGKOpevKCYbLj9HJYHE248ccRJ+hG9hmr06gG9Idm/sfv7VXXDU0uDl8/7UaeV3rHJsINO27
N83nhCHhb8Gja++vPL9BGTlGa2ddVgqgjTwoQ4vGMtIDHOJVVhte6qySX6GCSI0G8a3UwU1eWps/
nQ+xEL4cY8b8+wKTU6JhXfV1rS2srJsXEc2AE/cNh/E4UgI0SuEJglrrl/NlmERjD007vp54ghHD
mWfov7KbDhg8fUp0w0SZJ3ALSsF568fQ2DBOFCc9WTlL/GTQkkPTKudLObZ4hTxhvJY2xcN6AYVF
t6qwUQh97hc/FnVagCkx924qqp9v9pmtkZgaDM6OzTIY5lCyy/Npg72CE9FntSrPad9RV0YHbRXp
0/qKFAowvu9Pz2K6PC0V35ZWmFsdthsJidXMWNUgOCNTqVyvfsLlWh2uHwpqQw+0crd+Cwi2g80s
EU+gs9oj2g/iiY4dt8f7anmdpk2AGzmJPJfghyEjjZFXJEq6VaEQDk6lyByFiYcHP4tO0eVxNVAh
8FxWw/0OFo7pEhF5syeLxb4ydnrW4DtbjgsaGD45KXFN1GWqYxdTo37D6rAP9mo4IsX/8IdTKb1u
jGZ6r85hRH9xiGXIRVVD9Qn0PL9L3Ic4ChFOTyJdiXCfx/u7IXPlj+B7A3f7eUQNl0OaAjrVufuw
pdg6PgXfVHAWELEMzQsLBFO3hR0f3vlnO1BkPqXC/5stkW0SMVn1SO837sVcwsgn73rCWs2Oytg6
zJD1vhMLAh7qCMOgFqT+x39uqHKKkWXe6dJggnpwrV3SJxJ5L/YDQmz0+WZwmhZpwVM84DE6ONpN
w3KPCu+a0MDQ6qDVm+BLsl1xeFDZutiEnlv/28DXhgGBl4yd4dpjWh9+BdC+nkCEp9xyGSfHcptq
fJevlZ/WuEC6ZyvetJxBbEC2HJvSsnF3WfBayQhrwROuNMfa3NaMbmWOE7NltrAzcGWDwN+WIRv8
c3g1ivFwk5w8EPvu9ffTkRlOV2x14uhnT5P7KQm/66QGdsucMMleKWu3GdFSxy7ZUoRHhFLDCxmJ
MC7wVQmsRQ1nQPQWtLc8/mF0uTduqrnrrI6evi4eJ0p20mVHL7U8KgblfsewSpEWT4eyB++MNyoR
lsQ5MVcI1iI1HgFsv3s28Sd3QgLJHAjTinuFkyBYzXKD+RRmhk35y/5xVdDhDm9E+NoWDMOOardv
bfiUzoXyBM0rfegf4Qo3wk47NRE/cUuy3jmb480ewCkf2Xp00yCQg/Rq5qC5PxFz4hZ6fX6VyLHY
msEG36S7q+kiU41kQ9IndN6s9sHvAbpfhQ5rzozoxxO0e2dIPHbzt2SX3ZzIJxmLkM1thZyNSuk3
3rOcW7jXFpi48oiPJHim90oZwLGdsWquCiwpZmj8G9b0xNLCsabEBcHE1njITuwISoGtCgSK9UJN
3892I5VKb2DwzQ4ZErxQ0LZJvAMREXK9WASP+Vf0Ru96LV6kSR93YXV7OfpXmTvYu2eQcfLFP0cK
ft4JlM3NaYJO7v7BYlz6rwF6FQ1HnbF7a9BrCQOFPyx/wFIzLEEKdxfHwsMyaAaVrR3m7Ly7zqnd
/EDheYz0b6J949tMq0jzgB0nrFNVfEHE5Uz9V7LhngTDVgNPbAC1lCUy5JLH0zbRGhZnrwchHfpB
DoM1O5J1W0CKlf7Wh3IuDSkWSHu1St1vl3fXZ1bjEB31pfn5sQeSXwM1F/bUW2aHlnAc7a4VBv5q
J4im91PyH0bHmhE+Sf9pHBc2uN/6TZlfn8ULK2l+HHS6F1nebMfqqMAlzEA3nBI0OtC6t+pTZE6k
vw8PlxzmFIZPT0RVc6yFGLwQIMGjxRZwLiOCBX9Gdyf51f8diCCwkg40d5/j8O2EfF0yUc9F4dCl
V5ZHBdvZAeH6Rq/BWE02uoNPpjbqZ5aTEsgLu9WrDexoP60+gzlL/zrmN1goOOAHUhGqgo72OsLu
DyWfKMDSNLWgBp1W3cmzyq22YZz8mscULpWOdgqfEvJVrfiCM+R2ULUHXZwhKhvoIKlwUX9OEje0
D0LbeGmORgw84m4i0/vO33+f4QrDsdnEaL9rUlhzts6NN/kbeIGBQ5pfzYJRPyMCsZMOcvTZTY3A
t/ZFJalw888qVPMWpdqz8z+kuMsqFlQ0wFmwvN+TJRAFurXL0ha/eR8vGTHE7Q5j9qYjQRA4LePq
iQsL1GihTL5tpA70qbVwbtr/x39g4OMqAXso2QQwaOduVRdczSI9JXfd5Z7SaFUgHRCGh9cgWSIn
ADrGW8sBXJ8L+vtWPGTvK4Di5hKgLEi2TJrO04zbFt6GNTm98o8lKK0xD/s3MgfEaM4lTn2fUkcj
suZLVVHDcHix6bfKUyoz5NumN+Un5ay8/iMoNJmp3S7mcTrqoIAAqvxyqv/D2SPfQlEHin1Wr01l
RrpASRbQutQNTja+xqibsD/dZRNPtfPDp6Yvil4VneHZAHhhdnCjAwwh81R8AL94fwdCVHNXI/E3
ugKek3bU6qjSa88Jsf/SU+t24d+f26HwKXfiXNyyvw4B9tLul9AvqtSHmltOQqvXinSvfsYdmoJQ
C8oonC9OkQUrhO2pgml/l0d+rXVssoHwuly0vxrNYw4z15/3Q8LnAV0oxBeO5ydQ2wrQQRW58W0g
accWUfg/pR9khsHtrj5BMuoMEifKhP6dnwV+Z+Dfjg+o83U+0cpt6fRdrerKqfNYuH8H/TiS1tj4
A8wbsgXBacy0e8W9q6WJUBVgY/p8eeAjP7WWjAbfMNDFh8/46v2B8NcQqs5EBHpI+PXRp34eiSdM
oDvp0eL0UJg6f3oDrD1QLPLSi0WQ42gW+TXXHo/L2zA+5KIXXuJLzsdpkTEe6P/dnwUz1cT+vpB9
OaJfotLnlgn+ZSf/CafmT7MBipLSKMfWvi9p8X/IjdC6V33uD8kFc7RrP9nrJLD0Vn25P77VWOEv
ubEtN1kB+/CAghRD2QjIn+8v4KUcBrJJsEdos8u+mKxPupZOFdNzMNbg35DRAgOYuez915RV00Km
CGGS20j3Q1Q+F3VhcIeZ0LYs+cNh9rkyFD2pGznk+dNXnrpz+1pzJzCuhWN96U7EU3Bvf9qviw1e
3glYjxAFn9tDbdlfIonnaD5fSoBhcU5hZx5h2kHMGBEgSlBqMpOzrONPyySDul0CFNRpkmlYppR7
5M1ap4+uCa1Ujakxc11bEGseV1DC1Rmn9Nwh3x5FlZdKlSNu6oA5INnOU9zLhg2hCJpx30wKWz1U
OOOozZZZ90sCfqHs+b4J4EoqW0ebpIije7m2IwHLvlB+ORn1tXlv4wmNow3aBI30A8i9B9u8yM2V
WQsufqDXFa3PoEso6RqZF7+yFRjGEbPGdzPDLzBTqrgI5sbt00Xq2D2Qc5B+kNkXRzTP4Ji//F9I
DwnMEX7adTPVbh2aD9mb82mT0Sp41QDsY5EJA7gMd6ocwX4XpoSnz9XUZtRJZ4ZOBNMIZ1BSDrms
QcKW4JVHegP4U5Ore2EvsdJneY2gIeZPAq4dIgQ0ppiqjGpjtx6s7RNklrLJvafcT9H7/ZlpyNt7
BErQnhHXppuRRvUsEULkLhdvYulXkdVZB8ighoWssFx4iR1fJ17k4rLyZZze89faDys80RoKG9FM
lpeNBOdUeT7e0YGjkUOCvQ3jcdIqMN1qTReoX09jzaro1jH++C7pOBzpAc+lbiMjTo5W21nnfkFt
4fnjhTDibJs3spBPi5QuaY6Ss+CVTvlxhxtvcl/btSA3yg47HaUNqLx19tRgULy+yNPW+LbfzCS5
0K3SJfqg0BJ99tw2fVufl/MomVxyLgrTTLocLB27eJNBVps/bCzlXZgmf/gkHvEFuoX2ni59+l7p
QFSGt5MPtRCo4cmDUcCwGsziBWGcg0FyMX44rWYstknoLPvmAU6fezyCvwfdCGFTKH9IO/n0wJ2o
q2Yqj2TUFNwPZnEHBgYfHnBgiWHbrrvmFGGeamrIzSobwq5QpfoiKEOrgbfyqcTOxoMs5DQfgQFU
oDENVjtw2u09vX9zGIutyWV3dqn5JqkuhVlenKXkhWdy8kz3ACXD9HVvoP2qlZ7Ov82qwrJxy+Z5
u36F2hSaxhdPFk6W8XZ2roup4Wp1vaNQfOJrHUaVSsiI/kNgK6KnnUZ6VZctLbtmUVLzKWRQ/VsY
AqF0hIYNwKih1WE9zbP29Sua8IZNBialYPK3m1x4uyN+p8y4Wpmzb74baKNAEK2doeXODriDn4KP
WwY+npeQ3m7JffaotIEpA9qo8EuikmrTaxLG3KsB/rnP3woKtsZ5ZyzFTNlv44dQqkJi2ZH0vc1W
uaFY7YJ92WClyVrDfIJGkkqrNJsOaOTgSZYNaVkmzFXyAhUuFf7udtIO3DnyGj6LZn5IVjhQ7zHU
kJRrm/pCdCzm6VlMip2FZvDiIBIDra3/z/CyH33lQqvVIP+qJteVrMG8oKp4Yln9G7Q3kvSpadsk
qTJXAKhze4co1MGY6EcDCr4eFGBRlJ6anwDzu6g7TexQb8PS830vIeXpdmtPauKl0+YPTRGCUKo8
1LEk93qzvW3Ue/9tW58tg2tbjT0WCyG9kir+Zs3LnWjauFx6vMa0S0u3yPj54kY4sIKpbHlHbxP7
7+nAIba2V2jzGvrc8Mmifx2S3NtT/nbHuZt9+FQUvVyCPt5e6McBSry1mwUmob6OaqMMghbzU7rR
lbSPG9EhmbnROi6EbgpaQYItL5GeUuvdAQKzDaGZAuIOWF+6xbKdvqW6Cf4/Lt9DdZPlxIMYj5VW
G7XAVM+oU3hic2cnT/rKB0J54EC4/QSDnT04zLIXbztNAqHUuEpIOgg90pWrM3ymecuffE620bS5
vx/y9NUKGe5p2I9YwPBdXo/oevSfSxs3BUXd93xsT5HzfrstqOApci2MjyGAHTwGCaLv+ve4XMut
DfjkIKB36CFQ8PLJH85xW99Kgje89pKTfFfRJPaqUJ0UN/gkRi9ATEso10Y7cmMDtN2Y8YqYM/k7
4/0DX6s3PFvBpJiVNPP54Ou/AUN20S24JxDFKRNMH/ANqVTOvfsSGTT6izmy+KAM4lNBXgtgx77z
0oyWkzWzJE4S95fLZfy5TYEPrShAyAsmlDgLd4ZGJXK3qhJHiAWCAYzEoRAA/JGqR5DIQgN2xzF1
exUi+pW04w6q8+gWXvWAP4iFaawwDxGWTe6SbJU3u+VmHmakqBdCuvyfgsCGWoJFpkXdWwFowgsP
51JC8rtOpNynijhlvYdYUoo8hSzSTml6jH+tR0k8TMw5vIcu3IVzwkyHyteIsWxKeepRSSfKlz+G
r21lNjrJ9soZBi6dZxGhOxbKHt2VsOzdK9ZGBzvVN24y68gNt/Y4x25y2VQ85HoJrkFDi9LC5wXN
9bsxL18+GEEK6LZKUYU+IW84k2E6BHItKNAaCPvsOFYPqjqIZmA19P8MKUJnJdx6k+uoH6Zq80pC
n6E4rD9M4u96Qa8eRN1zkIdhnjEySdIQIDyB15XpdzGOFhFTpuVoy9octlT4GyYLzCtq6o2W2MSX
khiQkP+Ie1up8PPI+3lwJdsMIwgbq0fV9N/ua1XB06Dj66b8I1Prcy9WZESujhZqDSCJY8KnU18X
LnXMhMm/LEOTlyLwXpuNQxvpX77/Cb47JX63tnMJHNLtoqKsATtit9xwPSLfLuu+kEzc01+U7JLP
immDeNpJlweoP3pWBq1L7Pj/oKBUTDPMy3bq+rbsLcgU9DFzblzHPAubehnvpCR3bdA4DaLEPiXs
We8R6C2aO0YMPWzFgyOXT7UK0Fo4P/6Hr4wPSjep6eDEnsMghjb3T829hG2R3B6nZ/UVWCJ8KiKZ
NwPH43RY5FUj06CIKyBBIP6DTPKxqX4BDvjayeO8fouBkuTthzyqb67X6DbEC+WiS+H4xpX64Y8Z
E01HYcdz/Jr9yuJrjIvvCheQmz6J1cWC+JyIBRbq4u5k7R7NpqAw9NjSKhiVun8v19zGqrpECdlF
UH+WyMk13SVkPrPaq9YJlNXIgR+NyShaLEjK1XXAIn48lXRL1v7TqmY7ixJzXOkzH0Umon/A0Xn1
R5auBTSRPvWVCJ2YujjM5iB10tn36C2Kq27THgwiEEVEh5DdfbQxAEPLgOTckSfe8zmRbrdEBR5l
JiQPu6Uj/Xu/lIVy0qcBNu8sAhe+qCguZI2Fi7CLA0RrEDkSxppSoVqnWnOpojCvM5SDN+VxRJ5W
P2zLyLCXm/b41lF8lw1G+WSP/z6cbjCi8yjMmFG/CmKxyoS3gs8S92mFnGBN60/BKB54BcikUOMu
aiKy1mxuX3WDLeqPdKu4DxuEzwqzTqNY6XP4cABkoEVYm7mmueiQTiM5MGRg30a2pOXFmBAj7TNH
QlTpSD31MCnMKSiMlhpGNLDlBwXsqU6s3n3UEL25DFv88NHWH1Sum3dB/+G4z7Wwt3UuCeEclW4P
pvQSfz3qvMwD9NWkvIvw+jxKdkxtJD0Dpq/7m1n1xYv9wWw5LPCBW9VSMS+o03k5beNtuaXd6nsc
87gVjlqt+9A2WtmXctVbR4v7YiUpMgS0aIx+y+IWbd6copamaU7aCKyAFtqtJsVr+9NjvroZOpmw
toTmNQSoc/F4agKvs1rL348YLBOlayGroZhFJ9QOi++vl9Pbh4gU3gM6xTDAISrH1v6Pq7PGutn7
KRuWumfoT7aIWTsvp72sQO7unH2MuW6wL6DKGZ6impeilw6oXKCIJL/fneMINSGmaSWx1+/MpQzu
TrmuyuaLHRA7mLEMcO+OlkJ1eFDAXC+3wdlDCohJ2r3eFb+eAx7oZB8yfuFIhW1+RjmaQRs+6tRS
D5tQkbWGHwsClXw/WOZ/RZK/72evfdbziboMZL4zb3SWz9Q15Wh4Ex44N4vBWw6qNAL1NSo57qsp
Ai1e4ya5Z4cPyVeGGimVSPee6S/fobGoVQMqABOCUQ1eGnquXyu/5FMOR/k5bQDul/tu9ax9ga62
RgJHxMYAnx3UVNqMTHY787J6s/xzzottAGIBlCvkpYIAjp5w3rsoUDwUnSNKADu6XhScTnMYtijn
HfXvu/UfSvI3I4Y9vMBkHjD9L5Iguwuh2lTYFkbz2jeCHAxVRDSvomURXp4YDyX9KOORDsxKlZHX
UwEskrMvSEq1cA3hmvvG7mwcttz+o2BMPvTftQ9dfCgGJnl/xK5TAM3rVD5QdxDCFsHhc53ZQ4e7
FnWNyh6sThQTUwZvlChF2TeZFdxC6igIi6zBWYW0AVmtK8m6QYa9Uh0Zh5PrN/6aTB6ed0FfMH/d
qEwc6BCcHXdwTfRYFOJoIJniFn4+oahQLYJJ/rCR3CxEF+Htlz2Pd9hWxHyWV9upkAD8JtiPC0oB
qNzg2yrlDNcyadrTa3n0I1SK0heyZK5PY7pzKqoBYu2oXknIBdRoMhTqitGJA6TLmBVWbWPB78Do
BRED42XIuEbBMzBTJTYaOXrxGABdGmx3xIyHeapsgIzNYaUyfz29t94gQL7e9HOjnvQXCzRsoEc/
/bQ+YjDv1hxnPdmbWs1flGqcaet8p47CLqSWM5VQzv/SxfEXi3y34/PrepZ9yFkvRF4U1D5aydzR
M/pybiEr8o/PxbVFsJNO+ScT/1/Q536t2Od8r2KD+rBdFjFgIjlwN0KHUj/qqlqy0tWchsVfJVNf
YeTLE1aEy8gx+9matM6uRwAiPZ+lUk6JyLaFZxO34voRxXvT6fXhRs+LPfJHNA34OUh7JXE1jqXO
XettO3GgA3kFZsN/6G3jCDiqnsuBBfBKuS8j6qqa6o9zCvV4VlY0yd4gag6z88yW+Mv9uoCbf/GN
jp1h2Erm/t9Ip56mGPCuFfVw/YMpki0ghQo3i7vdvsl3BoA41x/K5uFpe2ae2r/61bZXRe5YZhpF
gH6cm/7kYc6zOeq7R29sBtVfp8OzmetTjzClrM5h2DsYc4L5oqvc07GltLXjeispt0oVSOFOb2gY
4EFPnCT/GaI6Fan5N4KFJb/ihYlspxNXNEilDWaI4bUYYdJXlfFOdPJeuhvApiGKNB93sF6ifujS
JDY0McJ65iuR3ZFaQ+BMEzxZRywI8JXE+xLuZyOceUht/TT30/L+qjdR4uu1y0p946VHhYo+xVm7
9aOCRppguzWdTY/sLA0MORqqKeIgK9v7jp3R6T3wHteDR215Ub04vYdeU0WxxgnB/uFd719jgQT/
isBcgnd/dfa96FLpwZRYwIVZzJcJUWTBryKgEPNqw6Fep9cZkhFVJonam9eIRKSWcxpuAMEolW8E
URmQUbQnXC/4qA+rBJCaJIZIaIrc3fGyRQfseIx9JQX3qxIUjTur3H+h4u6RgdwPo58/nFSJsaIV
GUPy5xKYkOJg327YDcxN1d3laU1jdv0v19OaLuINGShpfVSCXUHXaelglbL+akT3oUQMBE8WlKXI
Q1F/VTQgQtRulkuFl60NHsQQpNg5qDvkCip7GH5WpqM8x0/325mUYOzzdsVGN2iXrgbYjRUVce4j
LvzHoTcOLm0lvGDkNHEf78tmSJbZGM4mJiZTGknDER8qrp0zd3xL6yQFCKPDYM+kV/KjnFMWjWTb
dlEH+QPE2INCf5drVp+9kveYJVZDDxKq5Nywq/cym9dMNv16jDzcnnQSQotWKA3R5HXOUD8pqFkV
PcfOFLM+CHVyw8ep5K33oJiCtZkIGAW4kakzPEiq02hc+ddaPNoY736rzNcig+IYnJOmv8T0wS6Q
uLtKVxqMDJWHhxkuKWskGfxOb/EpaRubK3azYq9h+ZjI/R8v1gw4BvCImYE9ojBrhgx05C91Bb7+
fzUUJCWr0SU47YUtkiYcQkZEXxEHIYeAUJgPwP+gM0G4TIPCKIkxzFgZ9MRMo/HJNsEcKYc7u5rf
iJjN5RyzC+7rUYK/fyfE4hE1FSLraMcY9e0fkmB/HIjtHKqmiSTT1h1chZtpZsnYc2vTSubWOdlB
sBd5bdLiVRRqI0vzcdHO19AhQO+PcsdBLlgyz3mu7hAC6iQvlLj205xhwayLkmG5+6lkKvs22eJN
lL9+uwipMTgKKtQtzD4l2yVot3pvU0hEbnO5ia1EmyO+MVUuf/B/6ArcEtpF8LgEL82lMvVf+S1l
1qSSTEkZHXPQaHiw0FvJJs1562pP9WPif0RAOb46Qi6NbcbJj0hbf3L3sm5qe1AfLAMhkuiG9+a5
3QGKym/P4XG4KDHOmZ+xiuTTmomLZzFuBn0L1fTtooYfgGmRBZLLjd5yyzWzTFhpvvTjOfbuegAh
udQCYiAddzygYmq699MIqaH/alOhNQWbQ9YIqLQfj3ZvlgCBnXNQSyU3p7wIueCuQ/I9too5CFBP
DRHl0B7HZZ7nqQ8J409ED9dLbVBDYZKkKtq6PhFQFyw1Dfc1FAO/gRv0DqyWeNKbY5+IsiEZAi97
IXIV0ZGavfxWMeqiovhHnWt8BCPHqkLZb/4xF5uhl+5CWYltmieNxnttG25YQGSyKRUiKcC5BLkP
Evk5znYFdGlImf2UnGbJwvp0KxWUIxm4hnrDeAZvHHsA6fZKHInurYHJpR1FjyMi5pmodWPJE80l
88rCRELTRdiIOwJBX4pQJmw6K+ZGela4Zjq5ZRAv4Up5XNkNnocNPmAYsJnP7uzsvY2t7KxtGiBP
k7EI2DWOHeTjJ+YqUygkqprN/mhv8qiqNuFW0rs/OSrxcJLdLhon900nbkCOwoiUpnH0qCYNaO3S
ber0NRz06oabz2eac5bbtnvfUbvFvqc+E0LIb8P8tUMxO+ofW2/cLoWNky2aocyWPDDMsTLfjXHX
npfhhJ9jzdxJzTS+6JuN04mtoSBVEisX4v60z3DtxhkGKvrcCEOFjy18YlLXQKRtABUJ6FZhlf+W
bAzrVMIlePI/os2BfgXv+00PAERYFG/4U4BO9y5QDcMAZvok32oHaAmnBlpRzCNe6a3jBWWEUROc
m8KcKJLFjlpTAYeFlXgJq6y/DJ2l2p5vZ4QiWWj3gAdFNmvtey4TvwJC/E4dDj4vb5nKgxMllnPV
qB4MzxGfwp++8Csbm7EwWuVRhQmsmcQTLZyBxIaYKDH91wA2NY+AoslRtcWBkshBzm+mLO7SVZax
hwNv0LK0Gurmp8rAx70Dl3fSRMBHmypPg0qrAe8YGqX0KSjJY+1j+pB/ztd3h1+6yQnKBAa45b11
HXnUSNFBp0cJ1YNRtLF7cPDJHchJKLZf8MmqvJgyWehqMeEp6kNPQLI5wytgu4b5nc7XlDrZobJA
nNVn09qBje4UtXO7sT2aKikgtBKKg/VssFFUzB4cEJCeobpSBDJoguE9rBTo9MwQN1JlHn/eCLop
nQQRG2jHI4E5jSa2ZSw2WsJHtMe/3gFa6R8RI/dNX26Zp7R09FFPMwIM//xmxwBJIUuAikyZd0Su
V/AIGtWZdYyoZu2bmh14/WJCrbUUQT5bs+KcniNsR2x5G2WbKy4npDUsAKcuPD5mCiMAdWBzx3BD
lhTghI5SsVGPKm/Oa8Ai8yhY3ONdJyseUeFgvdEPD302sX2OkXK+WzUjSa/QhCx1eYRx4xwpC49n
jWHLM2KxKKP8u4q2hZIeBstNik5wBDZowKTuSPHBFXJWw2U8dtsUf3Gkl7+IajObL343TmtF7HTH
yQV0ukKvdenIMbumDCPMPogoCbYa0hZPy0VbTuPsPj9foh4JVl+C89dUtQwAWynjwL5mQwIrAB57
jloHUARVItMV6eyzqpT5pmQLta8p56vqK9bmL1i84RQnfWCc5R0mbKz8wE0iXcYaGJQjWdWw0ttA
jD90g635emgEFYAqoTBEyy8K14jMYaX/HPNcHvPHgiKct6wQ91diBF24uJWpQ7CocMaSTanvrhr1
vO8dOon/nrjqeil1FmzsGX0yQwK3PgVrKDWwLo/4YFS7eYVmRqK+9Vrqlq1lTiDQnAGcQtvLWuo4
Q1u/6/STrD6/o1qI5djeqtyhVE+zbLMn08LPMSQ5xg/YXkJzwlVK5K8rOZ/qD6ub/nP9ycshYoNk
1AYyzdLCTvUWxSETxo+Tlg22eoMddomSYORVywfw33dU9d41hF+xYEnGfi9KlblS0mfizTWXaWm1
ksw9NVg4wldh8MnPnShfkFhQypGGXB20MPBjCI9/DYcBPtP6wDgXaAaf0iDgua/K2194CNdLg9w3
BIbUvLNAOlzdRkZAOMeyVCPFLWQ4JdrytKE+Kbk1K+87lkjUqcSzWwOnNXjOxAf4nfKUKM2gv0wo
qbHcxwPLzciimNtpdmDxz/Xu/H+c1MsCD2hqH9q8/LewMcoERahWWYbX5OmjgpJLmTaHwIBH8+GH
OJEj5yHK+w4g+fodArv55jJi5IkA/I9pOwvUEO2F1Lj7OOBcDhBAvAxdTwUqF0cZYoBwYQq/D8K5
zRhhnyBfyeFW9ik0cWi2fZ2JSonD2wvrqcU9ajfjE79SM+g6XEB47YY6l8MJKMD7l2m5e9XHIUII
uZHnnDqn1Xd/mTqUMGesAXK48s3GWHlgiYQ3NVAsigRKtbMZGRmwnkWCVhOfDaYDMW0CyIQwTP6H
/T2R0kPwj67/T5/a4XEc2+Qa7lO9pab74ZrcWzQNp3pwgjatKM7OMhHpJm7HKeq20lSnVfDnpYuH
Zl29bNiS28GcsRfPBbnaCh0K0fEZMcUiMTnqqZntEACBQIZWSMGxuAuKgQZ7s3MrDdfcCd73cDG2
kdF19RMiJeD+Fxq9jFKrzH/WelF0kUg0roj5vsAOuhy2vKLXoNcTleHZuhcrGmsyz/d5a7A7L5h2
OkcACmRcS6v7yaH1s4ieWYgceQTejwV0ECdaxGxDBVCkJtYi9m63aiohqXISFaCpr+2o7IZdgfC2
wIy3bpM37TKSC6CLyoqRDVgunYClLRJ+0csuU1ltbCpOhnNvjAOtscH6oAxa/kda7zBHXdqBVaEA
a2YUpi41dpmb3tOZ1b/IVjCVEn2erFOGYVWfp1ZJgAQ+bt/5UlU6HJcHrCQr8usXMx3rCsuxt0M+
bW5rc3YUB2CjJTdyXW0OTjFKK9t2G3JK5W+d4lPjdVtukAeRRH4qinvHBM419fdvIJnRNHwdpcj/
0XqCW+EiDqpbZZ2zco9osnVp+UgBRG8o1QTHR2i9uXcTfOL4KQ8V07kOh3aRmgjdskPszp40yP+t
mP41L+smKfo7eAnPwJNuAN7G1tgXVLzZN6ZGeiicP4DUIdeNl3gP9iK3MkQbRv6GIVGmvJqA4R2M
CECjHG7s2oTree7YM2MPfiuestYZh21a0k1XefxPM2GP0K+Q3Ldz60tX0yDdPUbCoS8R9vlG7gmU
bHaqjMNI4p6e0pB/lqoYtV6GYN80JTQtMOi8fkElM7nj8x1W718b8YzTuR//+pKz1gw4hATT6+7C
r9vmCVsBfeiEYXCbahDFN/Fehqng7KI56ZDt+hogWcwLLfOpq++/O9Fb2htEE1HASJa7TQBW7rPh
9gmfjZYKdSbUQgC2ZRnWnoYBsd9M/Q58xyq1V5T1tiUjKfoqI6grnCpUXnI8IT6agrgV4iMYj29x
4FapxE9fDsUuA5gO0mW2mb3cHaG64NgCMn3R7Xh2L4mUC41RmsgCvcODt1cZ60PUbeWKGZ/kFs92
LRvX1whwawNu8UVklHS+gCVPY/ernNkiupIjoIgMRDyvrQ7JJ8ST0NTyaF2jiV9nBMQFVLrzLkAc
ghbgPFodNytr+mxENvxeW789gEUmUwr9WdH3v1rw3U+ELA5y+1fF/lWQDbY7LDA4VQFwh5g3BvRT
RDe8cuOOSltCUCZ/4GoV90mx3yl7qD1skQ8ddSzuqKv3GLT0Wnd/OaqtrjoM8BvMDd5xWBl8ccLu
XtXTTu+IxLZR1dQG5qFwk/8tikjA26CIj1gCA3QMcp1frz9beeG5fxvlTFCma/yV8fLanRWRC54e
fg9ZBOxnsaGFKH8DQ0eqUTpO7IUkIWSNkNmq5mmKk6ysmYhsdqxD7aPgTVnLpNn6n5Nc9GXIb695
Cf5KTgbTnzlE4TiHuF8sglMnKE+Xsay9GCz+NDgIiuI/0lh/IhYlSx1qejaSBVtT9Au/o12EU4jr
3UptPzKpPKpVz8dRQncqD0QBCxSE+6OvIef2I03JMHrtpyEefzr6Zd49EVy8FNq12gGZ6BnT3pgA
aGCjj3Kc2hnY8oMwHgiuzFrsUjfqSGtputo7OaATEIg7Ez6VpOrXi4YmoXiMJUjSAdnCgaB0IOcr
zGI1e5Bh6Q8MNme/i4tjbdND4uokKqqRA/Sa+ZHej7YeksSzTR4S4Y7Pww1XRM8dgCUCHRRBtpBT
MvgzSri9fXExMMGARc4I9MXvw5gue/Z/rPDnsoi4worMY/BlIDS0PPAfmDt/0hGZPYAXZ+mK4zer
/B+M4w5p6+Qs/CRUiKwChv+wNgsK+4Bk6KbgyMJ3W+FHc2gy//pJJD8vcWjSPwNfOSpPEqzV9OSs
XFFDQ7M1o+NIrATfIaSEyfJpy9o8uKT6PrmHSYiDoSzR+b74mxkvzVYj8uxtm6QrvIEDc69bwSnV
VYqLfxkhRNqrJhxZfE2CF5nylg5VyDL0dOKA0Jry5SIe99wrlAknj6LsFCnI8k+9XM5rtN4mCXkX
nXBv5vd1Fw3wg0qae5FJOO04ODuA2Ws6kf+JOGigOwbOsiS2dqSkXQWg5e33AobJQVRtWhzgyERA
drNROnVKvyIaLTSvxpk2bVQbKx9fmgy14Xvngp/85oiLEGva2webgeodKmPo3Z5IMWIm+SkDsDM5
NXc1ePXttd0zb7C5RqfHPD9/sizN/xdjLKHsQtqnxTp1tPB6LiBTysa7qOesqdlJLUHFx4L0dvXj
4yyh8xurMxzRpge/g7x02ZehLRJLN+5PimkDFKaSkmz2yLA8/EhP3DneECn0aeZhUeS/Icj2+kAg
5e3gm3l/Vwp/RtUw/Wf+bp4MT60zgGcHaisYacar+cm+9hPgpDl18uuAP0PGXkX1WvWYNS4OngOf
+u4jJ4B2C2XdJ5lmR1CJIdKMrIUc7u0MdeSG/AhwKPAW5TenyFaSAJxMkNw46r6izSWV5Kqxg/tZ
XfDYAJ625HgtJC/Pk1qCkuYNTlWKjmWxwgCkLLuNfrcc+9xSGwEOsKLuk3/Jt5fEGxzMDxFBvTjL
76Hz10pH/HVmpcPZBJDraRU53xlXPu3nI7o1IpG2hP6pumBaxKFFihVQrnR2NhC0VanuFNYvGI8f
N9Zx1dVTZk1qLNBmpd6xyYcoZlf+AmANMVsQsqvQj92XTU0DYrI7PRtxO5wSxrs0YEpH+oqwy4u9
oM9J3OWrAdbwrc3hRNqDQ3nH/V7wUu3Zon9l3PlKqCvmDf28ovTpNZxH2Yl1UCKk5RUrlbukMBfC
0xJGWonta5z+7QwP/P/I+wDpVfwBPsG6uM0GpKcgX0S7DDNNWfrvocovINJo8GZCl3V33u4hginB
DE1joJUhm8gCfQArJPKVAu63ETlmei9bI7zTPcsi+DgXfYwC2jQ1OmlKnH7UJz6itRwaopKQi2tB
xamVf5Bz7/tOS2Zigo3kvLaLYDffUywEXDMkhtSUNevTJGWGXgCXzjo9wgcKwy5KHxWFS7wzlI/T
xo2YU7cQ4sY98JTTnreLUXnHTUNSyaBcvOdgkIyGryPrBUBdJk6RH54YsLJhUyAGpgnvX83eLOpn
G6I6khX2zwQzD98YRhrYzwebd9vQdDIyp53aI4eshG7x32/51/yBndwc5+SbzT94ISkiJQpur5nN
NN3K/MTk4IjeJhAkh9iik9ewEqNTrfVDkpTy5ui6yEwvo2c/yG3Zpcxrx0AEpWrzK4BuU9Oo4OFR
3KBFv9WS7kM7A0Mo6EbihvR9T9FrvkL22Zo+V43AXaEOHo4edFARB3QQgfhhACYFflzrb/b/eCbB
L6A9fUAUlbMRHcgpC7F33M5weOqHOy9S4ZPw2p1jcI7aPd5GkeCRJvlKZ9MDrM0CvJUdfMzVWZkL
8kynASWjPupl2htlShqSshz8J0iwPDf2ybWILHtdHs5KK0JKKaJv5HgOf6OXn+px0C5XqzPOBiDM
rnW4PkAZz5EFb+rv/jSh5k3uBrS7LknoV78JE4JWOzgnyHJSlr8bARaDJnRa6oFVYdXyBjfJVmcB
LSVPFGBayF+Y+0I+tkyqUNvd42yvaeaU9GkXzNeiG2e8eViIoSCYF0OgcoCl8YpwDjZsWhWwUcM4
pNOwmH6CqTJfihDh0Af7aOwrgipMkUkdpb9OBNU8IRj1xwarJy3ouBTD74EwGMG9sfuMgQLQek4l
o3IKCyu87LUMqhOBFUMBRzXa0n9Zf+c2yKv4/8Dkzap6GIknLtMnk2abJtwE0axZC8cEuDDEbqVH
1rmbhV5lAdq3XXSffjsB5FVoU5dNnQq8Im6IGI7pPOlT+sF8aToeu9mSexJqkTAePQyWi8J61qaE
ue/8bBuVV/UZziO11O10GscPe/177PCJMIO9VOkE06HVZ/83wbao8lLl/gQIMBFAytrIh+a7ofhR
D/HU/MLaTHDwfyXhYGDd9FMWbGj0AlOWB6LZqzHZixtc0QsSqm7AdUaLJE45KRoPXPnVHOCI706n
4ePKl2Q95shSHgJpXidMuedRWn6ix+fON5bVF0vb8NBlmzGNeSNZzjmTYrLHV8j8/6pfAWrQ2su2
bxt9JFn4LPegojpinkw5kIvOl+CPavWnJQLezC8mpaTvtq72yOH4lhjbFFGnzw/HlVdH9bAzn2Hq
sNMXRaBXaWlGradIBOpztPO2n3VgFzGbJlOIfxl6T6e1vDHVlj3J6h6kVdJlG5QNd1YqeVnm7dBH
/NVDxZXj69LNOQd3DP/8BAU8NEhlhQKtEIwgleMm6UxD2BaHUjg0kkvbGb/3GTHJNVScQleDPtfO
OdoMuKY10LflUt5pTOPXlbwARNyysVDD3BSWiTjqhjFFHy6VMXN0kQRqN0J22wqP3r3hpNVJ8YwJ
6KKwcpmQml912r34TcSjyBIapUGusZucRL862cwC1B15sb9i0HjZ7HlsVtKVOBrCq5uAzg6F3mA6
dW+0+RcTbhtGnPHavcKSnt+WnyYcadF4rHq5dKyeblgWtbkWYV3mwVP6bYnc3p8Pdvt+gpTPDPZz
1yGj1PBHUJO3WSn2isDt0h6Bsiln5ivNxlUu3mJGK1JEH5fMPpcoIuFiR7MEcxYxunUzwxxjJJTT
B4VUpoS8h6r4rOq72C3CYYPyd5EoXuWn3pMDp9zFMxNkFMig0IQTVKCUUtGvJQkzcyB/FKE7B68Q
pcqGEHn2r1iVtXaFipQkadUQcBY8C9nQ87wurafo3DP7BvXFkFB1Rx0blvnJQtqSpDs1tvxS9As8
jkPPAOfapcdGsEGTxfDQroUBPIglX7ogLFC5z4qPa+b2wOOVsjX1fLoFHWu2Y70rpRPYTf0asu/K
Nuq2fpydlmN0ZYiCt9JX9lAZ1jrAedAHALeTF08mZPqLbrcPP90f/bR7LiC9gUuKrGOpRqL5qwDs
sMDKZUzsNsQoLkm9bnMwqFmhocwzDdEVED9P+Ph15soqABovMvS5teDeCfnQ1ffrSCrUqX0+ahk5
5/kjQB3nymuC39O/8OF4dJosaEesBVI4Gm8Rx6l8PIyfFzaoE+dcB9Ctmbvcl/KmXZnzM7geUxvJ
df5sIgTlpef7wnWrjzpn28KhzX92uwNp0FMuoKdJ0CfTcyHLwhJsgGN8ORhx/8BWwWr6QLszwI42
8U7Neog97DiFXBtFNOt15QVBDH2GHB95PiV+9wxGWeRXKVyqPvUA7zskyBuw6mm5hMNC47Ge2Q2s
wtRozfn5bHyYS9gJAOZfugsMxjvbtj7OXSPEAhilEhN+q/KvJeFW3ZXWqibNdkDd8r8ZsNfVRMJe
JtNzqoLFmrUSknt/YvvMyTqej8wprzzbhTpjykOsGUT1qiKFjDtZZSWTHOo64ZWGSh3wB9XKzocy
zBJfycTqBoAghFudDpDQDz2KKhcYlriI56/aLf3LCKNUU5giYQ9TxnjMM7TLfol872fx+QUkaiDi
23lulJKhq0iBGt9GK04yXZ70JN03S9/7z+usD9CV+j5MBZ6kDtce0fsLxzecJ32MV/acH44Q67oM
J2ocfZlk6gfyRcMxXMROclZtK+K68rMUt9N2ibLIu76dGhP8MiGChmhn97X0hwXTm9WaSSUC1Tkd
T3jrB/+rsxzY5mQ2veYiHRUZIdVXxpm8ZVGI0PrrJ/H4XbCF2ouXOF22dOKo7nhmjrCbRWgsAFZ7
dWbJsoxZBh/eYECw8ohle3s5yF8P3CINAbAtNueN33n+mtrVk/J11NzRxgEvcPUy3nwHTtioR2kT
/kg2KcY+uOpBRUp0Am6D2/j2FLU4tMbYeKXTYJhv6OTAfxFM/KJRyPFXBZX7L8cUn8sd9SJryyPd
UWCsEv8y1epOZDRi8netcC0eVDFONOlFAGXPuLf8Gvo1bubpwV+Bqh39GOHwruBSCgLQc+gAdahj
7/9V5u/8kPJYnLknr3xc21p/H1h+fsH5+ph4IPt1GopIcAlAVVg4MGeR2hsw4VeH0EXja0Zi2HYw
fzG6yxUeFwjPI2YrMgEPWNNGyhOIM56jeFIqZKYteDwmTa8MmvhBWxOVpEMvS3SeXkJB+bc8+K98
dw3F/EXxZ/dKqLxQb6pRuDyWqTyd0PWmz9OQ2k8IApleOOrYjZNaZWl47zkPiBeODkWzMMkHLS1u
RzgfxA3SRFPGtWU7WiCvYNoQQan8+6dc8v8yiZvMCNU1xdWHhwXi7y2EpS7BTT1xkU/VamU7jVvl
IE4CbhBkQkq92/8nYnJ1SsnfK5TV7N/UJ1uGGWK8OjqSJEdmjEA2W8VHI+Tqut0JxZu8Dryhrg67
G0q10Isx3C/RQZc/72/IVbWRDfUATHbACJVoIyNABnMG2NFcUx9AXJLjGbKFKP4C5J5se+QZSrHW
8m4jisOFOO3/gDLvA0GKSFtcYiACbSeONDNeddcJ9dvVq4WEgvfEKNs7q3BUfsr+LBLTLg5IENyy
n+SWAxUY8P+Cryzhh8vurykJ0ZVhXbcFHkDxGCpy0i8yPvDidJ8RoGxxJfnHbQRLP19YT2zok4+H
5+HBAUEpQoszkEjKG3XEDAD0yZBbGnz+lh5X01wVO+CX3wYglw/bCFTKZJQrgYv/qrPoxlKqm9wG
LIT4hkvqDAtrLU6TCw91HDulObwcx0Vko1V4MAQ7CpwP7pm9zlsFhgwJobDi7HfqcTIgldyPf7b/
aTICEKYCz3LucepOYWLSq+3F4PG0kefgZZeToJJ6aBqcYbe9n656wpnlbxZ+rDsG/bTQwTsCo1a4
A0ABi34al+3Svr3/uTzqE1m2f0sFI0X8YB0tDfk4ZUc4AadYi8kdm4hckvwYW6f7YY5P6N8ZiH3U
zE/8NSgvm8svzv5ppxyw7C8eMZFo5ZWHFwIc73v00TaCQEJOUj0hD1AzBDtOdigPYC/ngW7kflOs
+TQVhLNMlV+r8bvGGpV2Z8jnKHPRSXAPdNQZJzfS4lqdgJQIHmJzLjVgqpgtNBVfYLFcpFcJIzyR
sB0//EfC3RM1pvLDet2iXdMwTFACzWSq6lH898gg8nUmWvB6MMcYTBFIr8hA7ivtyFMPelV/b8xQ
cWUiWpdzAivRHiAXP/d8cjEFm34rohvOoXPKAvBp1M5u97MuQFDag2jslS4/ZBCUGUbp8s+ozWf/
SIMcr5jbG0LZyKiYlParmcPWEVvUW+aiX6ceQ2l8uW8udMVsdaa2G+aLB4Wj++tg4RECTQSTmMpn
/9oMaNnhtFlXAG5KkjA4UDA0BE5+dvI6EmneWVL0wLhsfpL3JWic9vAdhn7ShT3188Czf5uI+VrJ
r6k+n1uWo5ogCr0sPmhi4KW4RiwWgZ2i/G5tji65Z00uHH/mlQzK7YDJzncv+EY5RhaIvPKkKwrZ
4mDZVe1lS6ZnFVsO2pX+u3nU8Yv63EOdvUsTEyYFR9guKTFf2Ik6YEgWpEl/qegRAJjmhuu7qlmD
ZAjcbfMWwdpxVV4wun4ZSSpmAOjyb8wkSS1b9N+ssj/42HCgGrKCzicPIWqTNcMZoHw1oQEJp3em
U2E8vNpQ8tKcPh93jM6s3vMs9DM0WCp6MRwh11VPm9AFIvVrVbTXDy5DvEayoJVLKXUjJ3U/XzG6
HsYz9drgFrlmIu2WOl27juQkq/ZDzLARMZ9pjewcNrlX89g1rTtsvGdIZ5TCW/B3MnlQlIq08zuj
33Dm4MoMQn4muUqTII30si/1mbqaKnvZWK+Reyy2xmI2zeM4+7NRQf2U+x/DC2gxX9tC2wyii9iN
snD+06GQ03LMR+XQcWUJpZ5RZkga1bDlr4MFmdcXOyGn7PmKZqTTeCoSs3TSeDJfirmfL7fCd3xx
iCE0MP7J20kQKahqJLavEnVgxVgUog9Klxk20g5OzsWdDljLO91VnpP2jJynLplw2qn3KRBVRVOk
1yASH9C8HI1v+oQDLFkL7QvuC+ddnjPhg6ngsJLVnrQHIOxt2xRyOSrv9yTXwqvBlPLADIaiw9bo
JQjRqWAfXUxN95PTzT0H42IkZrxXikgOnDGz5SLBfJJFjLm5X+ngbz1bgwnfREaKwp4a6WjnK9fB
VUmT6VetH3fUVEItsFJR2NhQEZI5yKhx+jT4YQ76UApueU3CDjIQ29L6yJtooXJWEqgh2EVR0Wy7
NdMjwMiahgnrDQ6SRPsndz+hXSL6l2ChzHXUGtYc3IfFqcmL7l8n5aYpqZb4xpBTVZS7B7iexYS5
jw5+YZPpPJBjbsP/o7u3X5+0onCHoXjtfxfU635BBqfI4jipYcekok1iAfOzzgcwTkVtFi1DQMwc
mXTdvQ7Scg3pDmmjUOZaN3IQ43Dh1FV/TOSXF1W1C+S2Pw2RyXbAh+RmXYYOlVvuKOqXagx742Q0
dGvuhkSbL7M3BsYImXNS590HmZZj52eBRcZiAeliF0tHDzMa1fR6co7aGEt6z4j0ROq5IUntQ3Qr
5m3E2UfMogCbcQ8KCKmH7CKHHuf+Y250xcJMHSJCftqHqcpgIgfRngyItJBGsUMJJ5wtt8UsYROJ
/zcyjpuhBGY2gbPUfmhSHsp31zUyvCxByuHTGfJO54WHOfNq0pO/Adp1BKbAxIYwqm7z7XEWasMT
JvZxgkyVRJ+PJy9DqG6SbDUnL8kLHgjj71cWf3iCTxaJ2lrPT+paltMNSZKfE0b9LzX5jU0VAhyu
OO3u216dqvLqBaT7V40OFrHO1xNpRtibZEOhNRa8/Lq0Ndc1ZoF1ZAZe2uv3Wn4Eblc6JuvwXqVr
lKkzTk7ClYV3sEK+UkaVaLrAB1DMbueH2lDcfQBg+kTf+adlimfeAzTNPT1VWXUUvwgdYV9Ebe1e
W1JuEQ7uA0BVhgK+tWxP++7bmVKzoi5uREpY/js4iikZPdgpPJU5JgAkoTiaMVOot39iDAkO26p/
SATybqc1Ow22Clu593/NhLROCmr3LEZd7QmwvbJrndM6TJjTcj48ysJYMxk/COYagDCgA3dD+Oje
Il4NGjSSgUwOZFAczsRCMr2PwE8OtWeozgEmXXr4PQiTu3Jiu/xBXzQza0kWMUDe7gG8ECiNbUlI
s8Lbt0hgTybQhn2DUhdZaHAy9H7KCuRL5UKxkGdMpBsuEA0g7Fsc0oenk4IH39VaQCRJawMuXdM+
8u6jmZ4hv2VPw7JQX8tahI5bejsAxPbJY68AS0nGDJtg2gDVgymWMkKDwlxKMe3hpG/IL5pOWOHN
Y3jpqoLLiMoMIeOSn8WgEe8BUnb6vOBpKPX8ysyf/R32jMxys4cwfYDcIra8ZuyTrcimTrVvKyJ1
9cJ44+zxznmyKqe1NmalUA0yAnAjUGlkbze+Uq2bYLAWyXB4sG3DEJHIevhfC1Mz6/n9ajHRRPB/
e0KPBRfDu5h+7NLfh0OJ1fZ2qym0FIKQ8WqJKhdScasYOwh2T1Pugp0diLGgsqvtZ+7oxr+NWIbt
ijlR0lRJZuyUx0fdAtVTCYKB4UO2Rr1IU4cvBmH3DAic+5zOaKnxbQY/Bcx11ityqR9VXs53o9cX
1nRE7eYHpEbDA8LkpEkErEizZJ8msX4AOZTESEOhRye8rgRGNZ1aK5fa+WXxhqGojCZxaAtbBNSI
iqXt66xwVsYzGrax/h373Cr3APrbhZLI9pk9vhVDmI70JKS/znDmyHkLeoYNQ9jnCSn+B0Oc+OpD
iFwf4RMEJ4nKM9/Ltae/kOjDtc0HkibUuhstgRZktlNcYOpEqUpfOB8rTvf1ETi4m9SmDq1vK0CU
fDQmrod8G5IU4DHtpbrSO0gr/bwUPQQauQdaS3lRPCUeL9pgEMkuUJMTgPI+mkyNQSk1T+gL7u+P
DZSyj09nTYnPoY6UkyU6NQN4u5uz7VhvB1jTv3p8h8Pkmh17xzvDZmEMarBYgaYtLFfw//gI6fBF
zqrTm3Shf6OzPjnpmWeeJYj/Wp9FFjvhSXpq42o6hCp4gG6hX0wKwwED/m+prqPlYrS7lG77lBhn
p4jNMVNNN9nDA9cMHUZoBV1DaC1T0A/mPzuCnI58hvn7UkWP2x6scXFStQvrb0enekAqS5zXmROu
gbzykPV/9yObFK/saqCQz4uBzhiNrSS1jfHst/aauKJlE+pOHhjUCrWyqWrwH66b+40TWQuB7bcS
njgbLuQ/3tQ95sAHzygLaMCdoeRXPQXDOXy9a9u99LFfSwJnVE3wOyDdZwS0kKYGcZvt9+aJ92Ff
byIlx+I1xH2w03h8o8Z3ZwN73bEM+WzYRzDCTIgAa1Er1atsel6CCqQUC4benabD5dBtSzqmy1/0
lsbfovvQd09Xb4eA32UrpslN2vhh0pahE74es75fm7xkv7dGuETeWAUaDR6lMxrGQdlu1DtUWiUF
BAWWVXY8q0LAvzvazhYyuR54+UIDzAME45LeUT/mB+fQfG/6dseq8sIEVffyBF+RVRCwQ1PDBkeh
oiq320HFlA3Ge6aYfAkVj9a0c1uzCFQCkGxP2s6cqCXJ7B2R79sLjfJM3LCjZ6J2Tra44pUlVzcE
JfT3BdK1qYtPJsX1fZdj3Ganoz69VOjfWXYUsOzEg21Fez+qsuYg05+0Ykw1E/kSeghIkISwl+BN
EkJGUIaOGrj0yeg1cImcM7AjaWNA/lZSg2OEUVes41deHwI36kjgIbylsiPpIjhSC/TtjaSF5RVa
1kWhTgPDtleMgEzUMNJ1Sk4Tmzp0E0T+mjokL1d7f7cTEl6k+rAGjmVDGuNq05hKxaLVWIBgae4O
7JFIk3SI1Py2p7l8QJYc66ZZ1UQeriorZrbutv9t8UDaz4Rn4pKjrOCt1cCBmrQwIq2qpAta2xzc
i8IbMeiWdhmyCzpXSeDyMGfjjJdmp99/5nKYbgYcxizGxXLf2D27vEG5dGDk1OjMknf3hjsOGI2w
+wdLUpAeKxH8Vj3BLaDAsUnU4pRjI2c95rnO+nOLIGLPIO1eGP3/NCcqeLLef2V7ta+jHYTujJJo
FB0Sjb+Mamj8NxQ0Dx0zG99ghjLWconXcZQGrM8TA/fX1lDIgVU8AStY9bOzo5MmbaMy6MRt0Ts8
5BbkVabKoMOu8CRWSe2hOGE/44e2jT+lJW8+e9mOF3iQm+tI+Enh59niT9ZxokpBvVKWpv5Ey6Ng
EsDfrPXSZLvNKZfZCkkmYEg+12s6i/U479pOamcncHg7A6AE80HSbUO4TFzY4iSLNqcdHLF1f9oq
+OsCl3/3NiFjjQfWaUeJNxwCfyw+DFPFvych+3gczdaJqMO3T5aujtfQ4rPpW1yeEvFaHLHEGePN
WQU17LpCpy0eJ5Pa+l1WiDP4K16h3/jQVe7oTHEZw7l1QaCgwSe3eN3WVGngH0FXDEFjpczQHwEB
m87qj5SCIGAiyQ7RzAcE+2Xj3U6H6O8NjpKz5ViQoOTNApxfxj2kLm2hv+4oGr99MLKMFo8ihW3k
eFn3Bxd6V9QQ0Eqco4DYuwmAcAR3mYnGQJdFTmfCpwpSyQ1HDoBMskjrI6PMzlDvdUvrvCvgQVIr
MCLrhURJE46jR8OX8tXW+l51vpQLNnf/2Jf3EWmOwmvkMmo6c0ZnhwzKPcOdKuTNYTYqZZfwc3B6
oYGLksAueV1wD+IycKogKO4i2g1vbLPKcU1AP/LqK3sWLLstAeA+BbRM/lU4AK0DzBoLWqQthTEN
OgP1kpfEnZYm/B6f4SAfFeVhDYluv3QCotqvsh3tH//8LDBXlhni6xDhsb764xSrWNchogKfaChG
rGtjwEN0KSUScmxov/52WdWStAozwblkRjhPt1HsQlbbzftlJC+INxT86db6YbcdW4A9qcawbsz0
1Cc0v+bk2uUk+8SToIvUu6hyoNj3ijVWfq4vsRM3dg7CHHQtIYEx00RDFr1eng185pvHNKKSRB/Q
3f0rZ9joa3CBBYc72uIKWuOUUfKQ0YQla9lHyhj6kVXLttA6lXkp1drCaNI9PgWFy5LU+CIJYA95
bDPCV6pJYQTmL2qYtfbrm8+66FeHvMHAfSn5S0iTYjgLSJzfrpSGb08YAqGiKN/CHERF3weSHL4V
ccyJxGjwDEaw32RiPaGE9eaPUb3tvXyA3Wcn7Qk92tKod912tT4w9PUqciIourgLhRs3FydA5aI3
Jw70SjgOtMNhH9cRv2BhKiOMgTpYWu6xUkozWRVDuIbL0sPkt+Pg5jzlOTFyJtQKc6Zj128uWq+i
FuQq5/z926AwSyyeQj71yyww8ytLkS0gI+i4y1ViDFdmrhL9N2dpZo91Vzk+3eKff71jiGYOyKKu
4kKVsue706nb9dKw8umBbnQlb15PxYSJ0LM++ceIIgf7algU0+Jz/UJbmzWM+EXPwry9Is3TIRnw
cguiqFJ/1VXEozzQeBFFtMw0hVVg6Mu7PVruuzMNQOTiiIfUfGCcGpmdEg8jhrxL+BAZ4tJPF79+
4IxKFy/1heejto/YjfRfpXSGuTfbkfMwCTu0R7NKDcrFx3lIEM8zgGY3c6plcfToy+Zf9396wrNg
RRFX83E48Ibcu2BMnWZprMVgL30HrhynYta7/sKmP5FCLzCswpGtWazbn4gPamyduYVW6q+oBuM6
6rHekiCGmgDoe4bf0BxfAib7b7YywgciWx5yqg9rj2vxNWmMybuozU/J2FTSrgWIlIpwvQybQS6r
zyYwGU19C+1d+eIH68xp9JaM/BQ/agvvJLnn7QO4Z1rRAT6jmrWsk02hIHJOShN4EQ2HyG2sFh5B
Md5pxXwB0P+qn1hOQRrsroQOmUBjYQuJVm8Pj0338itfEwcbaWL5HnyygM8pggaE3IgCx+urdfqz
sm/jBAadKbq4aV6wq/fDY933zOFYeTktrOhzT7IWBOVkl79Xv0Nb69DzQ0VBD6uxkKSeXcrVXZEF
tnrNM49LBWCc7M+jh/74fw1ficJ87NlQfGnb/pclKqTP0M+tTRVJO/y5jlt7062YxkzM6526Q3CY
BEmVKvpQiSXN5uBiuK/OpGmiL4cFgaO+mWwmrw5q+t37K4WJq0r9z8q6Qjp+dSJ7h3R0tWdDOYhq
iMBYENbvs9KJx3iuklUbYEz7yjyE/8FJ1YSiBOW+5zZ2WNTGLYK4ozqIAheOr3FPLEtnri6r8SDc
ZVsjP7rsL4fURnaUdqWEzxIrACDo6OmZjmqvEWnBejS6ZScK24A2/mtFCMXhgNBj+csSpm16r2Me
5m82pzWopuS4KG2IKUsLjrS1RMU6NVO9Dq++KnaomUAdE7LfCYXU3e4P442RlnCyUiNuEozptea9
8fRMIT0PLu3nHObWqNBSFIyoqz+X6Mg4nM+dlUu11GLNG7Xwtkm8CCUAZ28yPBN9XuUEkVkRVkY6
6bYrXfOjPptRAO2f03QrbvgJyolEEDXL50x07cphbXL5n23l/pr+sD6WtKLSo0QP9Zya8w4OGL2k
AQj07Zm+lNwshMqPEcybZYgoPbvnzGStrwnkZg2EhrRAOy1/y/WKKmKFfA1DsarhEXCtxvcrecIU
82BUUp9wL9Ge9rwYIKDx9AKpJVt4wppQXKwgnBBLkk2Hu5H12swYPTXq4xkN4k9yQFYANw+f5qIp
iNrfYCFy6LMD77Ad0oWplcF1VPIFxN0m7u/PZk/+ZNOYpJlFesWC411yR9jgkP/4Mvsu6AwC6fmV
VuUGltumwvuienaGMSclz7CvaosW8nFm7I0UdXqO9zJbJGfKEpfMHLBeTKrEh0xb7ojOT307Cp92
8/Ubu6Y25YPyFPFP0Ui+sKYmXjUfp+tNuAdIONeP8f9Z2psx8JS9gDlMFfLyhqM3nwsvxThoL6fN
DQsY2TRqjFpxt6WKQzBd3YKnzYFFPkJiNMsz3Z+KnDgbFP47AcqgbQwqtHxwfUcnaq2nZpkk4Rqg
T6sJXzEXwlQL8BBJEP/sJIlY38uAFr8dq0uv67NC7FJ8FU5KZx50+jjK0QcTSPqaFhmBxKktbhr3
yt/hVfp8KV0O6/srVgO3OCYvKKNdkTqKqBtgRwG82AwFhGDCzAo+d1yl22G8ETrGJ/vgLlUrYxU/
m4S7pCN5bUroXnZTvf/4G5Z1APLzLcSKyZ+FREUh4J7fhl0Vp6phXUUvCIq/nHiaBEWj006D/iFk
BSp94WSkPwPoRrWmgUXs2dPdvQ/dCK12CVVvEXF9CyTPFrqif0XaLkA4USEnuhv5xq+NBBUhbXyh
BEmG/UZBUrguLh+vnntNFp7gilIMbPiJ3Zgni1afbvEKvP1uptx3NDao3r0xhkmmp2o0HrVu8Q0e
3qdBpbRTp8VWNHHQugQ6lF+1Cl1ZcEgpjgUQpNSelxl69bjFKSKx86i+/YSAXOJe2G8i0p794rpu
KMpZa3ufXZcaM7GhNIp+bFreE/KGzFnq5dNdwBUNXJzHQH670A/YKAVm3FtH+Qdu2ErkUJTT6Ch3
LqQNy0jveezbgTTrO7p8dl+gvAeu2dHcu4WzXH8BSGuYytzzNFYG8XEjAs+zCBrs6hIv8JV+S9x6
1bglKTJuqRmPzimHDUHXRqVS9QxqBiMUWJ4ALYaYjBsgtR2nWDNzcaOngwNPJzxCC1+Suv5SUER7
q3LZ0LGxn2mIimXB//9kfVto54OQu0RXy4gULs6DosCgqLaqSbWmsZKRlLw3GAUca+kzxDpPbGQj
MRwuHtZaU9tmFGWVHQ8DJmml2/oppzme01iYEfpDVdUxjMBzz5OsjO4+qrFb6OJJ5ps9L9Rb19H4
QjmQTxUh4tf0fweZZ+XkqdU9G4OszuhQlY6catPUi3Ugz6Kf5MXf/Cg8+17FWR1TXtKYjGnH4dIf
WPVo1meHbMKBk++9hZJs/9TD04udxgjl8ascXaqGbcP41s2Z8KCA0e8yU0xsqYP/mqFbhdQvaHCB
hw/oDvONRGbG28Qn2OMEkZsRqaR2kIb+2tJRbpV1nkKRZ129nUgFIXW/TvmcjIGaSJ66tNHghk0b
NNDPCj8SdRma7r0y97xtDIugrBAuBafKtVSEBFqGK9Ua+9l9SoO+Y/3S+AyQBUoDxS8yvJlYAqlY
rR6Q3jD1SgccEY5dzmF6JUlFB/O8Vre5lv1aIQNTnpI00GsYRyz8q7njCtCnW0CUNHhK/+fXdX25
G5Kl0crsL04SvQAGaWlugnzjZS35OVwUKYxpDyqYc8Jjx9afSbCDDzJ1kWy3DBKTtq3b5HsFqa5S
xYLebhbZ8OOqmR6iDtAdjuHI2/Y4YTRJOkB75ECDSmMM9pTOZXB4jDe3PmYS3M5PAIQwB/Fv0O9z
TQhitHX+MDflIFf2ogrmojzatTF67sMI//hQlBL4PrnycWdf4VFh1nO4SNuCzv0iEiSsnoUkt55E
ukDn8uf3JrjliTkk4oCJDZoU78LiTxaUfwNK9xZ9k+tZvV8wBIMXNYKGov2fDxVm11FY7sLdZBkB
k13kZlzAY8hwiaWMACXJRXHJNGHubxkUrq4cMfCKN3fgUymGIULXMo/ogGKzHzwhHRLD1lcLnyTi
WQHph1SK4UpFeGG7ttiwdzVN7um/k5Gj8gzsiV7iqZT0plIg3Z0IKiAwZVBF+q3FnCUWSr0FBUu9
ltMJdEmuhd2V4rpkbPkY5y3RE+hkTjVrzvfdJTpv48JRLJIQtycUyZNk/HVx4v7goVznusDkJrU0
dAXXv8jjPnuOXvSQmYjlN4HhBr/ubupmg/uM9HDXMzoNu6lS8vU5L4XsUcbbPMkPyQqdMBlZdtxo
Y40T5d8MCudl/gppotaQHu3eAwZ1xKn9hqs4q/iADTgf4umTsY2PoFwURQ3nH5zNU92phBM021xx
gCs36mGPALeAVLfsqBiU/AxBmPakPdc63chFF4dTjz6j8sPtMuemSj/i5D/BrFfPf/Rc3QVCTlh8
j2neyaDcsgpSvnnfvE765kZ2HJaSN33dbP2JbI6bfM2bgi8yE32pGGIHpYe9LxPB+gSP+chtlE6t
jUe7NkvG9TaXKgi7itABDAQKhomujnvkPqRzNX6ck7IKT70mP/HzpV/5CQXIRm3rjzMrMWw2sHoe
W50/czkugQPbI3O+3MoyzrWCErlgF+TEHFrVCfWyWexm3Jsg8J+AFuzqNa+6ug/icFriXbkqgOGC
tbA64bTJlm3PDOy55SAdQBsmH8wjMTpjvKTQ3FGiEv/T2c/smJNUPMjv64aohnROQSJdLr9RDenI
Z8PDAGTF/c95pyobLwBsa+sE1ZFqQ656mRDwe+K+hQ4ylPUBrnIzZAgaZQn06S865EUoytWIcVnk
+g2L1A8qLkjf8mL2//A3G1CfEQ7q9ILb0T4xMoM+HokJH3Hm0QucXCsqQUKdn7ypXUYjBaUGay6w
xK4KHWKAJcrG0YHa6rFzcQ3tagGu5hCBVWoDz0RGvByXK444WXkIuRLS5BYe/TPmT5tnzdzVCoJ9
yoHPbPa/Q1stYhje5z6S1IrNJdx1Tpgfqv9yaeDx9SIIFw/M/OnD7VXXu5z9PlMBYcouIUKy8a89
HgfT6Nc6pf3N1LxfcBIfEmaaH3v00eFjK+7/OulFgGajAFrsmzgQf0bQOsI1gkHY2WvT/6pj8Rxw
t4bqWxAgISy2r/yOfHqOvHpANPPPgW9hy8gkCgoUFtK3AOG8JFnpAQ5YUCylggelMrxbhc6APBf5
st/nVYvfFRtRPHX90JU+uUIz5hTWArOturNmj5UTEFGYnaEFqJXuYjgKP2XWr1DmxmHI5BtcSqqq
t26QyGCOLmME6xPRw60G1JRu0CJKqUVMGogHSgbHI/SbWCDdSZwlFDdW/N7ntitqdEsb9cP3Ylvx
KEoVzEd2g6YedXS+CdShhGPb4EHwoUOZl36Se7rtH+P1tI9w766ZjhZKXSzAexsSJyJMMdtRZePN
hm5jRWHypvILIKbtyRYgLXZjJZd0OzHs9kIGsOFtG6WC61xlVDQVVKBa2KsAD1JleecW7m4ICkKF
2hBn1oo9iJ28pREH9oD/sXAcVJC7fQEJ/FwLyrd018ZjOhs6Iq9UxdmhwbnqcamphIc2kBazrAiM
dXMpUzmAhQk+bOiK4GA3TbRhL1kWaq7HQyfedkmZEdtaqhuT//bpXUocXPjXCpItkjsAWJQ5MLlL
wRNmSJx5NqftiVTpc0OPb/KY6Hb4oqLDKmohNscGNsQdHlXS8e8/vrFHYGFexLA5r9hlNqUv/tTL
1sJuxDTm4drVn2ki/5O60fFd32Xh8HWNYnOcK7W0bXBjU5eH0zsqBgRHGTa3aVl6zkAnim7+57c/
F+g5QUTRGO41bevy8W/bQywgmNKz/CqHVAobWI2tNJlYhgJ6gNujpFmFTbG8SSTrzwfEH4UZKlLL
CzzoKB9OXcO051uwpvL4z5YYe8udZLROPYaOYbg307QEx+2ffa8kFPFsdZHy9M4lBM80RUrh30i/
E6QOAf0X1LhJ6YOS31/ujr28yxYZxiSoWxyv1bbEEaFyiNRSixBFuutCrIzMIi1sWQ1hAsQb9J9z
onblk6j+7zgs0XQsqnfn2KTcfJDeGogADjmYdBkp2BU5Mv7+LAz/K1LV61DdcQFHuU97mYXRtbUf
Eu3sf+vzIyIHTDkadsKqLc/CmS9Sw0vptZLCUEYRA91QCzrwGC4UzEJh0r7yXF6+FWDdgygnoXfx
BtMUOi9vWghj8TbG/t2JPQ67P/GrHrn4PAmNDMX8ErjXv5eVi0NIxYm37/zWWNI647qRWto5gEEq
febcUHNJgJQ16taMLUnvBm8BaKBKVps2Afzdwgk7QlcKtOeEe9hcdpTsP9MIrPgYHrD/SsKQYeje
dEJLH+Twa5lhsJ2w8QGv8htAFHn7D3ylcnKnKpskaZvWsd8dFP3Y4wAtuVuRAnIox8iG1IuXcaPO
VgDlxaEv8T5n8d743gix9FJMLM5qPHQA8Z+L13n/pL0bkTCk9G3jHr02af+esEk3T1sy0Q/z/qbp
v6IDzSaSDzCcR3HPyep+x1p+SCRlhFc3XDUbaRTkPQfTIM+CMLAlh3mmnLgOnb1mudXMRdb6PQb5
A4Z7OX9yfa5JiqTriHShwu8Fqcp4hfO37OWJQa1KWesuhb3wns6vtDOoTfmYpz81hPcICu6RljoM
eX5PtqYR+IZzNBCiuxroaszRGvGSajp2SZKoU988YIwFPw+lxhYkige6lsVmTacDBodKO1UZ0gfp
z8+e6TKn3oTRmZMv2FxT5L+PsZSvPXJ98eqG5bjC19Bn0E3hsAZen3DbCAVAM+5eEUTkzuX7Jk7e
5TTA4D5kPoNUT6LcFhK3Kd/vNXTfM6ofLJZBPd9pjmULAtZl7l/qREoZLa7CJT6srCDfYOBXcVFJ
4Oo7HNYHoz+QwdTvLmIJlDfJhHtEOWgGunSILGhRk4AvxfMYUa8H2HfDh45DV1CtTAodJbKMXGug
oGHoGdJ9MTi8xLbMHYMocVNv9AdWFURKemINNLzJpKDBNd89686rZ0z1qoK9bHjD0Tvi+k7D0h6L
fhFP7J0R1EKbfZHDWEcD+v1Es/uef+AGwfjviwR0O9sITHesib8KtjUhnEnlrSxnprrpfAAbo09p
wWvxhu6UOGOGszsWTC7YRg12u2TLAGKxLmcBXtZRY3T+ivd7/HkhjXiAczY8dSokgel1ShkYtnq+
RModNBSp4h7iqHl3YcspalmH3FnGMJsFZhOkU8O64d6WAFHJw0CdTOZjZcEhYA4oDiGD9NJXAAzw
qR0EnLTmge44LkJkYZnjNrewvdxiBzpX6pQInJX6XD0zwmM0jI+JJS3XFgIMOcvYYjd/Wi8go768
RZZDOj+ByLWjLpytJ/QsfMvpH7neJ8YV3B9MMjK2+sLL8h2AUCAWmvhrA4ATBCX78JZG1dxfXuy7
19z5zCcMQ2WG6fM+nPSbR3kUX7XdQA4GaxWQgOlVOCGBwlqT1nzK8Sdp9f/XyfZbvY1EhiM8KBN8
2ieOHwF+iLseMAA9SmDpTz65EQ8JOivhkDGXGAqACj3ycl7OtiBEMnTn8J6xirqdG96GSnF0sHzd
5OjnwrlX36jO4i9dkzQLnB3abhCpqA3hkgkjL8cMBECyHx/IeQl4tgel67HUc/OUqxHyYBAegsbz
cR1pZ8f8grdHi5DEvncLTagQ1eN3Br8eV9dTARE0ZXhbJdRrTowDoWPfqcfQGz+ouLTq8sAl1+25
qnLjhGoNs1Ag4MO53UESBGx+5njTq81MBEJ1SD3SD/ctyjHenh3UPZ1aaYyBagiwG9A0tv2CioJX
M7hh62tHSR3OIPvfV2RLsZ9Q985Fxp8+oflmxzk7S/RCF6QcFbeGP4UY4VVL9V6BJHP2iazw590u
NogmObzH3TnKB2WddpvjG4SiTLN/JR9nmtjQHhfR6NtDSf93+4xZBrODyrzcx1EJx+iOVWH793S2
EfTGTOW0VHQRHeq3uy8IE000eBoPmHha7vgHtWDIzOk9er9Jp5Yb5Gp18bePfKCVSVHD+/FD1a2B
4OdCOROZcogBwvOQxokrq0bZbzTKvfdMTRdllzK+F6EH7e0bdLc8kKcE3jEb43f/kALJAl3iMdV5
igsRpzjZj0nTl8h66nNt5tD20N1W3ovcnVmvr7xNtEIEfa98T+3q/vhkee+vVwW34FWALr5oBIyS
XluGINHWr8rFeZEWQ68vHcaHzGZ/U1h4YhLoSqwMJEJPoDdQB7EmvSOiw0GWLGpzjfKFL9pKZvlp
gRP1kI7XO8EgnbfNHbb2/BiX0ohfWYf4Kj0oNc0fzbAMGpI1kBCdnfEPxgBRvjU8qMohPSP2rSuE
LJi6O75tmMT3kVn8IV6qYzdRVqvw2m3OsIMQiyCNze17hkbwXsuCNR/22ipF/1oZhdJAD7iBPge+
9KsOHRTrrkzsjlTV7X5ZALm3oWAxNglvqwbJxKSeX/gojf4Xw6SnjUD32wEzispnK5bCKREGtZ/6
2eQWQ6I3yNcuTB74sIE43kAI8GfKo3Gpi080kbOvQkNQYHxx/bq6lwaaC+C5ZFDS49rA+vkuBMm5
vkVs/qlZD25dLwT0RGQzwCUz+0zYk60VqK/wtNWrwERPEsfyQd/vII5qufDJ+jeoxTXawKncnfF/
SPJHuTlWxV4Ll8vXINS7Gw3czbtiu19qJdTSz163A1Y8hwOxMEm0qc3tp1VqLnwxStRXk7egCRHm
Zdp8CZNb7CPG+/sFEGMnMbMqIgF59nMK6DzVM73CAG35mpN7Ua1PmJBpJfes+i/8J4QlYf5cKRrJ
1UPc1UcxTM1QEqOlpWS0tOkWA61mtxj7Q4f93jPAogKnnMJqLqDYfvqvgKzy0g4oxqQkTPeWvM2o
dyJ0CN/ppPrAhTbuxxwYzSLywjevWE5+FVPwsYCLT+BPXs0tEg9EE3qB0iEY0SnaVrL6TYMiz/KR
f79ms+QAoJ5uWGwoYCnod0L3epYh7zrfIcAs0pTLllRB33Qq0DYTnttlA7AcThKI0bYgDWcclDAD
TqPljIx6bPYGvpN6WnzZRXcKXqBHJOs53CuTDbf9Bb2oDaSWV4gIUFXsyLw0gCJdldmHKbQq6wwq
yfBXETvqa7V3N6turI3gvEwk7HXBPskxKr0j7Ffd3XLbJiKHrebT/0Y9cpVsyXBR4/X/MloGu3zL
keAyByzyZ+Fl50a5WyJTnosmBBBfoDNSiYfuNpVoBFlMEX8xSvWEVb80b1QIZOdXmbow5fko8NxZ
SJEu7jqcNipz6cuQBQFmOtxZJEhJHNgFkdEQoTai0MwVbSyyEOMKlGaxC9Hg1kgxT1VQmuWTyEp6
/ewT5HEdUxdgegLOhFqX2ZE+Pi5xYjeub/83MMnf5ucTBdhRvGjsIiOPf3MCD1dTil2vbtJ8jAAP
OP1C3H7+O8QLm2h0ixULxqmjsdQbbsO34mkasRpQaxPstJ1yxSFRSfoEuqDnaMXrLKDGdpzslcmy
6qMreE7RrcufbhedxjlBgraFPC5syIqQ/mWP208VGw9AU+bUXFrWkK1g7Mrf1d6opvHxmdSi6snO
WvrfyDulK62qHOTRFg6HqLEDawjMLhbnr9xzDruLjy+rCvOa9p4lQcZ0xYUpHDQgnPBkLG8GSBq1
BMEvwyc8H5APo6FwHnsR4GIqFdiKxdiV9d8mEKL8UwVP0A5SfFl8/TPN1dNXe07jNyv/FhTCUxzI
/XeK+xt/r2umVScuiA3ofuZAwH7ppfVXq5jbm7MfgrJnnwJQp7j7hyaUpImH77AbeUVNNJ90GnvO
F+M5FUZJ15rJRt3KhGlaTFnqVFecxL8YH7uIL/Gp/8b9c+j7yw72R8tglJCc53KB0nCJRuhMLh/R
TZk6+SxseZeWCjM4FsSw4CxMACXHV/ysoSs1JDcWvKAdtpPKgq3u+n1NoSEcRP8qA0/mwXVrhWT2
jWLxiZIKmRfMjNpO2GacLyycKZ+ObA63xTP/+sHtvInwisppFuSJzO4F/PIBg/6FtnaWIPTO7Gd8
ESZAU/fwzS4mLXsUphxKiJ74nm/YlXv8hE7Ahv2cnCQUcq1LRZ+I9W3kCca9Uv1dU1gROTVWRvem
yjd/jM1o2/Nlzfh3ymNQXNxngue1StNAzyAAEwLyiUbZbmMRjk+8EvCp1vTwe/jzbxn5saJMyJKY
dVyXJuZkWC1yI0t9yfu232ygX/Z/zAKVrd3s4wBGW8SJSeR8i5jbrj+vDrSexXzjfLhiCowITW3b
VlxSLFRhUeZBI4oX787aAXFKMU+49yZLhksrbbzccW2/lwFXaro7I/hbh4LHmlZnwoUJUu4tAS/Z
VbbRWSQep7YAb+19zAtlZIPEgWrkRrQtqtd07I50kU8KQyRAXwgbQnRCNGV4Zh3iaHoLzwAVcWgV
NyhDyo8tJq1O9ks7M6Ur8GlmHY3u16wCIZbQ83aF9sOSsS3Tm9sc6O/ptSr9uytQrJY2yZbVMt+l
NblHfm1MA87Xi8dkUbLSL8VsqY0tHbBaZSEtlRmL6tYUEN0li3IUa+U5QswJcbtrevuR3graS4fe
uZTihAIgGTpk4g2E6m9GPS2AOXrhqZVuRHByas1Qm0Y0gDNmYBg3kWSK7LD+jrJw/tCEmxTaDONe
xNdDUYhZBbujQuANRDrMDrpR7Yyto5Z5eRvcUVinEoZiFvzAqCG5g2jwfzZcoWwFMg6iaGB3UuRa
EgrDHc4+LOsHi5ZPF1JOASi6mEoS7ZTs/XvUIt2hZS+cT1niCoSgP0SlO1rBN4MXFqRjIsVyalUn
y5lXc18kdSQrS3OucfJov7aXxsdRcfCiwefa9Lyz3RgUPmvbpNVKjw0MWULh9pikuZ/lG5at2Enf
0GwWXdwPd19mE5lDdFn0YfQMb+YuCg38j2YRESd4yhhcAFJ+DC2jKUfwFX+AKciKuDRY8+CQXnxY
IA4PgKlZUnTVsvevGQWVniZsThhNGvfO98BdLgvMxaOyZO5eQooE/sHoqN7B96Aeff7sUNvoLyje
Dcpp2KcKD1257LIM/Swc970AsGhtjOT8D4pySu6BvvCM6SUkaUgUFCyes81Lz8S+4FeYMv9jjO6/
nCv+nspWygahCLe3Q+I47yeijhMjQ6FEAmtkK3as5e6ZJ3RSwzFfY/E+B99xSWSgMxQCLUI101Ca
J7XijW0bQJeg1aAGdY6UQmFEMhpPRClfwXW3xDlAEckceTUXkZalaW33UJoxXJfWAZOUkQgAwskH
bQzCAWBY4EQmqdoKGcUZvzkO36kCzGWWq1bfJEKcI5C8F8VcRfQy6Nek27ljtH/zpGGC7iqynepe
IECMo7vbqurL0vhcfLstgOUf00KZLJKZF5Vt0wpzAg30bQgJZQVc7cFfxbYMnBiZ0f9rUzMaCzvr
3k+mcFgEkuayWFN4w4mdK7IA1YSN3/KPQ4aZ1nBjA1cG8B+ae+Efi54neav3xAkkUiIc79DGptBh
MuKV2Sgwjrt0mX1BKh1Lj1KP2Iq2T+NnadiMViHAmBB75ZKSGa/Mz2r1sKozAlTxMzKYChB9g3/P
e641x4P4GzVQHWIPo/fbwUNl3W6pUa8+8nBYm4it751ykMBrg/1vPCf+y8axD+2HsWMGg0glY2Xp
EiwxElf4QuIq6xX88RhzyyQsRI28wQD7HKrPf2C4vqjmng1DLTW4ujK/5bVLdMMET3EFxzVu8PEC
gGCzbHVhdcAZSwCtF83jF36ryZ2zP6jPF3jQCWAWWMV4WW3l3L/35sUh5XohZibEkPQ9TFCG6vBr
MUEcjiHylPahfawYxiACLLktR8gdE656D33i/rLxRnuVsIEYpe9JXOZ7rK2Q6BcH8xpIEKLOR1TC
LogRW0gN/+ykPm/SUgKixxcvdJP7ET6gSFV52of2XKNNRGA/Q1WcCHpCWgj1NxlLytIBeBxKURIx
fm0E3CrM+EhQu9xOPQMD54KCWPQDr6I1FkzHG0yzAT3EPwenblyHMX5QkodGY78CX8lMbw+Hj02v
FemK3Aqv9jZTfTlzBqaUrvG1MBQ+etO7fOodr5Gi/ixGz+cssHFqMe91SpBQOZrWRmka27Xmo1rm
e0gfW60J3SGc442WeuaCuaINbl0+87JN/jELwJ9mV/TN0oKyqTJWUaHf2MGIegjDbnjCU3m92CMw
nQowRDpn/KQJlUXD2V7qKrHSX0vrYCuxCtcoSPs2HnCxveKhwsanqshn0ihzJYRlRI2hrKLR3VfL
i6RL2m7F3m78oQxQhR+hTVZy3ov044h2fCVzCrnmslieGlNx/4G7mnKe5Qa2fs+x9Fke/Xagoxhh
RcWwftbuaNjQEVPL7KWbT0BjbFRkfRQPBEiwB45XWVfI/3pEVNCIV+LHPLwOZtATGcGb7N4T7E8c
chlLxp44g1DOqE/8fV+Yv0lrirKYlUS1mYgMwZ+TUpC4inAX1AFqJCQo9xdlRtGe+KSVQKjqAVoZ
kEbbXpjcXrF8exkjvqlBF+SpT4S2NbKrG2EeffKPjCYqG+t04PTnJiYuC5M/kIzjOe9fTIGCeOTT
1GJFxU4vn5rSPvLCeq8tL42mGlrYc2Ipqdv+o5RExsFFPk7tAweh4CXrdjShrQAHEFQnjshK9VY6
x6hBRdxl5dnJVgg+J+MqWWMYSAf9icNxLuBjrZwpWrnhrvqS4aXA6NdEtdTuhpym0kiYNivG2aXq
ePoK5dhbt+ejyaw8CAQZZqGNe2GsAii07/SevIiz4J0b4ByQA9JxOH1SrsVYeRI1vrj7SAssNTia
9emWSJeiBb7wJGJyqxJBimZjIDUScOA4PEWFf8AD6TKgLB1mK/qLDv/DChho9W8lcSZvNG2v+3io
H+gGFZitduTRNK9y+VU4oNdv9csVAMIL1pxPYx8t6wOS6vb7Q26pEZ3IqsSy4l0lGDzClIzvwnCU
wrVptBr3tMkLtv92MVYIrgi6bmHrCO6LzGEQTzr7kSqxSG5/yKJIDlzENS5twixvlbVmAEVOWQBs
B2hfpqFPf1jKlR9GH4rNkp3YrZzXAnS3K657UAYmNc3nej+R7NdxatvEWVGnRiYA9igHDL8ooFok
v9U5iQhpN7vXH9jLSz8b45i0T1HCsaj82SbPyx5ICNdAOTRfCOuutQb8LiDrLZTvKaPe6Li44v0y
x9F5SjGcZb477AAKgtLOV2T2gR4BUNXndJg1h5L672qebMmmobwZD1LWK7HUvazwG1xLKe2vU39Q
rpht+8rm3omtKIGaaetkkFaOgpSktjnhBs1NbHSHokCBOesur0cRMzRmk/74Qgr3MyS4PPChMqWw
nIiZUmt0GmPzWoJIHL2/VzgZFVxFq3I5DDJ8ze0COX+ntEZSkIn1VxRlIoiTLJeTMORMcvL5cIqP
sNhkwM20rxnj0L8nDxNwbOSARrHBfonJDe80esld0QDVTzb2HUA8cNUZGWOPNaOBRmOQl4AmS3gV
+KtebE1Lhe+J+zjKqcUtnEV8Y7pe7FJE/MRI0V5ElexAxKCLcfU+5hYajlTdMB1ohvEM5r02IP2C
4KSyHGEEgmFs1agogCKo6tgFjjCN6aPo18s2C4LU1bReqz1jjim7kbu3Oez7V+PAaX67A2Zguu9N
cIZyBhpaUPqtqNd8TsGLOoiJglu3OF3eSiqMA15CmbXrIok+HH9xNuSjubZhcuMGiwFe/PL34ei7
sNIdpliZQql/f223j+9elheH9IaGjbYEmJQ1IE11TUX63Oq4S5AXnPzteVhRxZeFyQS60bLbGa6F
ecv0KY1fh4wswaMtlFiFP7v2DZtg700llgTVQVGAJf/ritMLZSPvLkGNhVkZ1puL/weHsC0wsSdO
Af4qC1vQ1J+uEQdcXw1dz4ibdBMJoghVh713reHZc6cCzvoJcf8BgZ9+brrSkn+mn/Do3cLOyPuJ
6vRWXiajpCLYnneEI1U4Z6s27+Yk/go5wBQCxjVZn6BEXRmJgwhNFH14EKePmYPdkAOZUIYCi15+
6jZl/b98RHOdLUWy3j41eyW5S26spPt1GGfnEkL0JqmLjdizYQeKWPpau/QElH2YbabiLye09wXV
K/1nooM365JgRb8T6qXX4kJO3br1425z6m+9TFR+r/coVqKig81jk98JFoFxo4egiiWkzXurjkdi
mjBYvy1Ns/SDEo0q6L/k/T3ue1b+E18bg9zNWNPcf1DWZdimYAvChMBmVHMk5W+46ygaaXLvcoUl
pBNniJG52gWz6XdsyLFXopTnDpeCi6ZvYM4pe4rqx+0tofd51RVgYQ9SwhJg630N7xFXbBEuGO1m
uMmgMY8n4kFCde9w1tDsX6tWXb8LkvtdPipE6p4xTpRh+ZmXDnAmmGur1YOMRGzgFvvz7vBk0y0O
4c5kwxSLWWvb8dkHVDnvDWWb0GMoe/vYgNf30+p++stFrkLsifTeDnKON9eZBZvVOMRCiMBYkWGq
FA2itFXLnUP2eyyN/Cu0DkHsrfLhMlW0WPEVuiSdzcRc9cFmqhGI9OBR2aWZvOVtO2imPkYwUn3P
B/2V1P/z3dnit8IUhi2TrRJIe7SQ3pli5NBVYOq3pF9MhLxxRqSbA+xXMvglzIWB+xgAW+hapzkh
+uj1If6OrpyuCU09LLqI2LayUkFWEWjgkLq+k36BFtFJVaniTas7J3kqNDpNzKeVUhhE9F7lnv2p
OnSCBwC1N5jnEjrYhGuMt1u/CpqCIftdzvu+bWQx65ykn/7C/V6c8MLxUIJSxudLL/PoaC5Mf/HS
pQLW+Vz/ScqYHabnWC7QU51EU6ZuADHPGk51ObF+OJfz7fsjcC9cnwMAhWVqvxq6PCMYCUJdLkSc
+HQgKY+uhFA5F5NG62usmBe1CCKQeitE6/Mdlbq6AVCULb4likQ6zcZr95JqZWUvyU3t3277gsKt
aJ8BOhrXXVCERVoiZzDoXT/zX7ICGe1AVpC3Mfsn1p6W0VkbiSv+aX5pcg7iFyEZxLMlLGJyF4F6
hiF6PNAcKNgNac+/Ve7sedfs78rHaZ6dlzEDAMyLqvr4sAk+qtfDvr81Ea3iXmQAMtZ3OhwUFvAF
1pKxrKBNVi2hVsKpl4c5z9udV3xuemroAM6d3C1tO/Kp4RVA+FJ0FbbAC+9uVA6sDyqY8x9/kApp
qAAlUq37cV6dxvyj7Rn/aOIkQKamVKs2j/UQRA+fWsniEZT+oPMs7em53jDf+kLQzUheTln437EG
qV1ZdosREJwQ9aH4g3Ge63qexOLOFDpinuyE0gK+eTpqJp8pbFJTecg4Ql7XbcZ0b+o+2yevHXmL
knPtTAjkHIEre3EEBidzdWPIaOzJc26sNJJCzZbQaanW7ZZAr5qWIQ2AoRegyqD62PWFxJkRdoEw
dSZyAF3tm/64Mpg3qvPQf2FQdn+HpjYUOdFClM1tafGJ3DrOC98KBfXxUDihKSZT6uwJp1y7biCz
RU2ikLzp/lMP5escFDnx1jUABPhtE3qQCT//mCPD4BJ4jBt+hFPoP+Qf1hNfc3bsQ8znZQuyjBYN
dXdCqSpW7Se9z3OugRn7U27B+u+OfSr3WBi3mgEIY/Ni4bvc77vdC2RrCf1ar53lOroUwRK5ASWd
zkHJzVnKeF+WNT4oIu3zOjzaP+InzIA2RbRG1w97QUePSeUMQy/UykFuw8Wg8pgpaeK+Hoz0r1OX
/KghIggARaxXH6UW5uM86G2PA1tUElvf9MDctb6Af1HquzaPHLrAEjmzxnpWKnLT1IEZeTqkm0OD
DS2OrnGs1HHCXx1IFGEu30Bzi0Xe5T2J7iZLvxODHPAG8G67BFhASkX/LrHYNFwhXrI31r5Oloas
CXEv1Vu6m3OvNUfUsU5PoneMZQZPPw0ShZihePKGelqcScoLLTjwTjnH0buTelTrSZDcn+QZvRxQ
iuYfiXtF/vuE7dZWqxLaa6RylI4h5KSk+NZL5p16VrIRgFqt4aHnWdZb5wGaeMxUI3fuzeEpH66M
M4LE5KdLnydRiZHNkIFsL1ZPHjHvedbV/G0GLw1Ia40fJvg8oiH6AW7iF6KnlilByxSA+5PYWLI8
5kbDrvmRRcqPvWdZbq6lC45WZ5lmV/gbz07ymXjTvuekPmGEVyXv2Q264vLn40R98t1Apq9dTpe8
OUE9qaupcrpejR2i0WwyW8KN2Qx4SoOMPf8tLZqnqFy6kbmbugmXSvYAki6/63AOv401N120E3Fi
dy/J3qRpMVu3vcZiEzbJbAwipUm8x3tsfbVcnmz26h/8Ie8c5o0XRJBGMdOWmT1ckfzXKkQN/1d9
tFraZE6YqGHMMyceYcT4y9djOgPtTz8qFNKriVZSOualAcMZ75KeToMl2Me4TDWr20N/dMrCDShE
hXhiomZmrZyHo7ZTP3jPatZLGeC5ZniykV2jFJmVTmf8JrYpLk47EC8Jm0NKGGbWhdAZ99BkYb29
5T8DwVE+ji4WHq8Yu0cPUvE/+l/vvJEIuHIkl66+sFJJT5Gz3X5kWRSR6xI6/kYO3T+t6alzKr+I
XVZ489nqWCgodJLgFJNcqXWGTwzHpOMpKCkFfRS+M8s5pll4qJS1AagGTL3b859Iez0207DteG83
x2v/QPRa9TaWq4y32glvUeWv08MNgCs+N6hLb7vrnaYbX3oPq4ybJyv2PWnr+LMdrA956DawiiWJ
RkufJfJp3uJ6ij7PfwJQzuo+E0T39JVjM1/3+6SAnuFnuKh5vEoUKJzSOI+zOU8xBtPR6xQbSD/k
yaTJv08tt389rv3Wr1ttz7wUcbRgd4WOVawh/qz8HZi7cwlk7lb6HJxSqnUQCqT0BPu1rmcbjHVu
jFrjLtIU2RCtCoFSJP1G7ruB1NX51Z/NfFCUjr8B0jJA3ZHDjZncWUMcCiod2RtCQfMDdGnZ7eHV
U4LLLOIjklT0DfRKvtgsTcLsSzBj7oHy600YjOj85l0u+bQD4BfpfuzhmPpZJTmFAzT7dnhWC/XN
X+0SEJcRRc+vnyfWPyZmNlqT2t4AqZJcgy8MKv0RcYQGsi2wqbMb4h/LpY9CyZCM11HxwgW1jUjk
jGy1aDbwS2hO2R00pqNM886edXg5U0EDV6MeC3vMok0jbXSNVWnDniZtwFswW9blFk70xQ7LWiiI
dN/1UPUVtApJKNDTGNTfL8SOj6BD11ZOpC9Ghe9Vb16WeD5ZHceteoOx5N8VsnMj25G6SsJix/au
M2UHUt2vQza4Co9zZeSAv2xbMmfXEpf8yNSQ0A0bg89Ke/vHrIG2JAy4NkbK25ogdnWi9fQZcurF
3xl1xEE6vs+sJ6bc9SLJ2moWRC7xjD0zZGsLOMd7NkORTXSv4qPzbAUwsjVLugL6VCrbbghb2/DK
Jnv0qFxj4vVS4fmr9dEEe1EWxxzju5jsxvBs00Hf+Ozbu06pyEK29NrIz/Wn06Jlxl5NNEdVrmig
qmFx4dBqydH57vYXYCmES9y7QHZ/JGy5TWbrlcbSBm/Q017Jq5rSZ+1kpTokfE4A8kyjwLw5aGIR
VbFE5758lUoP0txHRf+qmyGg0GUB8Xsg21Db58LKxmuyDH405ajJaiV7e5dbmlWje25Bf00dFIuB
eSfkCNko5eHhit5qajwg2NQB2WwWu6SnsUBJu1dKIooTZU73Q3pq2Ygi/dABZj8L58lXrsBkqVrB
BAI8AeIsSknG06FfrvF5UbuGB8jxpVThbzok9LP+kbqPfY2eFLM6HQRApe621lDgUr/NR8p6ujyg
GsxNcTqHfDSzrDUimQ2mjR50A2VRBatRh8xDyF3ooY72izvIeU6AxTujZtLz2LR4GDFE6x+IUslv
0wwCp5wpyps9cBICr3FwCKyLBHuvNcUK6Pu/iViatXTDh9kneycy2KMkX8TdL8isFv47FjVNm464
EhbdMYNvbyqjkyEzVpoCewJP6AZTl4ZHUqd94e+Ht7NRDtxj3P4uFOHpbsd116hMWeTZfku6pXfK
k6NuzArgpVXOFd7+J47cjpQ++riulk2JMzh9n6Y+NX7P3WKE08MPj6NY4M5t0dX+fYcKEFbt6IHt
8U0qevqW6vW/EK5WH/JYnWWQw6lZdZ/V5cOCt+0sv5GDT6zjxZDK3bWI+i8CsgsqM5fNKkxqzi11
6N0FHVx6KL1o5BOqi37aaqWRZk/KfBBmOqJh/yU/BEP+3bduSAkQdrBb61fJ3lC2frrCzl4E/EKA
R+ahFvqvwrnbI3XQ7CHCcpplhPA+ERIvFU+seCQPYPt6JRdCYAiWXPAAv93t7c8QzGx5L8xE2EmL
LJRCh58rh4jpWHFSdwSJg7KTYEshoACLjO7Y7VDX91igCxvwSM3J7UUgEnDElMWl0E2ycK7867Et
6WRzZSU62CE3Abeb1NRMR5htuh0T4Y5U2EmdYQvBnWloVhHRt2Wr8FBE/r06r1IuSqOUWmbvsk09
bOrm+T3HOTO0+/+nkNyQyvpQzZ7RcccNiVqgfrOoNAjTC9VUP0m4ZN4WK8taP/y42vBU+iKN7Xp2
uym3YB7dOQMZY1ZNFsXIXz7bUHOgtl0Pt8XdxUZrO1UeJGyDRPmsQfDEZzJUGWBAV9PwIq1c0mst
VDDrtq1ZshXRrVLwwvAi8xZnHN7TuvqThCuWD3mZ7WYg4nAtXGLQ36ylIFgPkRFGcdKZFRdr8lYx
2Ma84delGRTP8xBrVqxIiwcM/RM+sir6zHRmGmuWxKfTtv4IhMj3Ee2htEjHNzdsvcHFirgcH1vB
wzgtwNIFvpCd9oF4oyW8+4J161XMXeMZRurhbkoKTwd3x5SRgjVTU53tTVgVEKFzLqn1YfG9/8ma
IHErbqoB277mY+U+yOgMysy65vJBAnz/+V5XLKJiJtc62O3E6xHYhWMT1QjgU4qSrLAMwTP9kIrJ
BQFCOfORoPObk1HivTYf1UordiRmg8i2XU0NJX501FlY0XAH20+gPF1zVwtpu1vLVe2mZtW7zUia
OYNyHzAoop/SykYxWNA0KS6TwfrWAlU3g4TOCWjr1a3DCGDIYFGIG1rA4Yf2ariXHcbcqvcoHYjy
6bUD2f5rtoMMKoOkwn82ef6vAh3ahoonmmYcBwsk8cef8CDtuY4ebS4xR7AV7UayxwuDq7Sx5oqB
LSqq6jrbzXdCazRKdvZYFZT7SygkMEgZFhi5hd7UvolyXgjgcfcyR8NGUgZjrStvcOBZ0JDuMySe
Vlyggjo6nWbgJ4u/XAbXMlEjb9cDslvtVTN28Lgsepny8TigEmibxSHd46d/CDizIaKa3wcNd5hj
+pCVxaNQoEDVYA2CfEGCi7ivzBrcaR5oo1lUrFDxzmEMXv0BAphI26ljWD78KrXRKzJo/M5Iiuis
0f8yIkMjuO371UbaVGbNRhdB/vetiBE2hevTSOUNua/cePOTz0T1CU0ZQOsTKyztrGYI2Qjv3hUJ
p+xzDyqwAZXezYW/XmI8Ps5Gqi+6+o/UuNBl1/66jSwUeqXcD9wR4ou7/pG6e/UB96clDdB+y2nc
M2ht9EV+DJYr4ST7sE/78WMsTmHc6pYpEyLRKiCRLFDt9lmN1KU3ea0/YHquR22VclucHgvQRn4X
WVuKJ79DP7ogXxV8du4ElSFe2wM1oMaPGl/d96zF7+2VXi61SQrWae5GPSqOQKR0+X1C362i0SaQ
1vIEZw8qN2kicXFc/7uRlPNZHsHyrKQMTL3+E3ntDl+ciab+s61cLx14thU911CRcysmTfkkQQKN
I1NWU6Em2fnN7xj5C0B5oKkWUfvPcNEoMuRgSImMLgB7HM33EdBm68Mdpe/8uFypNjUO+B+i0HG2
hT5GAhu2BpQNm2BMTSKLnlK+Hqm4Jsmjuxvbi7aHTm0HXhPCiKQOipw1IOnOXiJbhcH7o5LtVRP4
umJNePSp2bnyx3jdaFnb8ozRQFlARp2s3xHepojYzTfMmxEMoP9HSZ5hy6h+7pJ6waLDJ/e7y2EL
I1bAjSAufC2AD31qNFUBgqjjyPXp2DDabwqvDYoEKe5whzRnXj5/pWbwvxuAL4yPrXt66oovESzn
w3JVT7t+9FmlYtQ7zoZVgjyfXvWfUj2biYFGbeq8TnNDPpS1jtOH8ZokW6FEyLxeJ8/+LxyLq/tQ
GB3nl7W0fEgsidKLNGE5+Vne6VYrrtwE0XTlDVyaNXUeCZ9bY5SYuQxbia72NBnsrnr++uXjsWZb
JVUQrUZv/8uC+1TSfujFOn/ArB60E3OePwiDdNse42wtN4BGXRSH4noMieNBDIHm2BAHTsjDCgMG
yCctcr7Imsp9RHUfvcjajSQJ1I7+VHWWdPozyobs4RYii8Krqzmuu60bD4dsLiZ5bhPkr9fjoU5/
CqdCzDu7idi8fNRaWF6NpST7WQin4W12PgfYfd4HIc0fK+8pBeQ1AGKTdAVuvtQTwXj0JMmmaRut
M3+VU2QGooA0r0eqWuDyC22kV6MKVbVwLvXnLJ/nMJ/8HZ3zs7eO9gDsztfGUeFWV5Hb5zS9A/Uh
8OOSVk2HgrtkLxuCAxEDiiQgr3iUHGykwbslwt1fbr4qbmzM291B0zsuZrc9y26wGvk9NjeVTSqb
hrHg7rRY1se/+heuEYr/JC7JP/oAA7LPhgQ9dH5CGoMxFwZkighycZNSh9sOG74cHmhajaTgZ1Tl
9qbdAA52iLtYW7ZsSsSIiMYP1ZKzlsFXpzyLLTtfHaBLpbOy7tRT2bTrykc8EpQSKFtGnR4mMMS+
0WmoEGatSZTVUDRRiqlh7sgLTaScjdWnJoWbsS+ik5op4SAyiNd72TNPqfxkywx+d5NK8mgEIVy6
zLcus7e7JRzd9KYgMrPe8x1CJk/nnTp5ey++D9cr2OadhGUUIWAxt3N69AE6PkhjWbLCLL3eMtY+
9KngSeiYYDIfWLuoJcWSWc8ujPftWRHRrE6zyR7CIF9CO+F3KRtZiXdIx4RZ4ym5Q7h9/sxgsBLK
e3GtxlDcSwMoZ/IGy/w2HG7MuZ6OHokXzLhavW7blxRdh/T0EstXvQ6OD13T+nQLNy0LAwC4jRdQ
k6LpD1NNPvhuBWAb+QvjBXvAs2c2lgFLf/DYFVStVIaVIoJAy4e0kWawv3pw0jURracXYHO6rYoC
LRuq5bkf20B8XqMSOXMeQDAc0jaockQBYm2kxEyDFvduLlBaElYRsBerhbW5jgx4gs5mQBaiR9aB
TzGltuUrQ2SwdN/2MVpPs3bCEa8xzVD2G9Sfku6fbzEFFi3szFBAfgFVaCwtG81JIdsT/OD4h9Ii
y8R83dFcnEUQh2t7PJPLeg6F86tspGjhKdqOfeuzTbFXyLa5suQ3xHnAfK9hhL/w3Fyyivgz5V+E
YHALOTGhazTYsTcuHZeOtghxw8X0jVYkCg8UCHnBQdVJw7oJNswhqBpQGfl8YGwN21BmBYoMfUhI
Tm1tiyGGnIrruiXS3Go89effjBGjX9aAyOeu6SZvCBPOP70s4I/y12WTz8/rs9vEustAh8eMJ2Uo
TTwVV6+fnCFA6ELJX5Zj2QNmnCDK6sIkRq74DAt9wIqEgzcJkGeO0TRVXtkYyUsEJyGR2BiEQGag
F5lvpHHD8JU8EUuYP0VSdKI+BdWg3nJn2eEKIzTclxpJWgVXYF5nEIsdUfZfdUODesmt9/Exuv6C
8ejY3W/vxKRt7lEaQErktePb6UGVk7nZgNSJD69jEtAooMS/S0G9XwRRt0xFhbSQckUFyuHn9y2j
rq/lLO224Iv4ByJRadUztgCRApB5hUrZeU3JgzdndYl0F/V2Ixws/jgXHOwner/B9caMTZgbRUTC
VW2I53HhfDfq5k22YiKbyMSqW40AlclKDid8d9jHplo3CCB47cLf0Mh5FX/NHVFekfkOXitgp9+5
Z5Ktt0RYYhwyuvCoWp9088lu4RfPocFFbQq8L8E4WQWLh0+nMEs4fy2vzGnVeq86+XlimFMT6Qsa
/d/bHw70L2gbzdqBt5gQt6puqrG2O+kKhjvev8+w1bGV5RKdQhZifSUdo/MoMI5zhHT9VmmMfkle
apDC7g2qPUmNO7ZVXjPz9bWNA2rHaz42aFGYjCWJ8C25iZw7Xzb5uZKb4o56qUN/cXza0Ehjor+N
FLgNqSGjg/yNUO5LRMd/8whvhgtLJRDl+NpYOTBBO9HTWAC+Ca/b7AGdx4r6/iLcd0Gj+sLavXr2
rSQQJZit599ByKYwSsrkKGS6t0rWxAxc3t86s9tN7v39OSOMeKIvUi3EOb2OxaQM6mQ+F9YZSmQm
PMDBt3dRgyhidzxa1iuq+reMsWiptoq7UwaqioLyuxWL+Kbp38ocOhs8o1TgQ5KtNdYvx/kZT5AL
8XxTmjyLQxoBRwRkgFvdVwEJ3d1bLLoCEmQpQxr+7Y1qEt9h4nndqvPyHZc+dUnjwtxbsqDowcT5
C2u/njHMZVECdN5n5PCP6GZ9H78ZZe3dNjUthN1+0Zrz725Yjwt3uG8HqdRN/yDx0L/uGEGHie3l
ff6EoYm1CON9DrEDTv2xtlCXuRfwN5VbP9M4CTxUmeo/qPmzsqfTNCJF6OC4VtW+wCN5nVMKkbms
BoTddjZ3iU+r5kUVlw6/G4aR01quhh9Uxv44VzFVvIpNNWJc/Zj+6EZSoANPgJNY22zhCPK174rO
mXx56M4IyhzMsBNTQ8tUjF9zrc50OSJngn4PHTfxFZxjqQPWM4yFQtS//Hd5HXU2j1A1e5cUMxnS
buzJFNecab8SFC7Y1OdGbvGyZ2S8FNRFOoKKfOnqClCmcKwdg+D75MYbAd+9aDKJZ/BgMJCdWUKc
vO8xokcjtA6s/ZaXwV/hClo1lDx/Ytqza53oo7B+OFJHL5GZG/Y0UoOrz2lYMv2thKTC8xOvtx8e
D3KA3W4x//nLNKiI9XhK2ECdFRv1NG3CwSMLUhCWhP44v/21ytTyKcaBfd9KjreUeAIb4dgrEZ75
7OZL3ma0WM6Iq9QG2gpSbnJo0aogMM+hTAzP8nSZl7bfsVDYK1119ME2bsv5FzBYJ8baIcAXxXmq
BDeYA37bxYnB783uwrzs8+lvmIFegbh0+3y/+MS1WPUBZVyqLZm/orWawhvKTUSvkNBEw6ReZIzq
i09EAo5hh7p7nMPElvZQ3Y2yj9T6HcGgqq+yi2NHaM1nUHKbNNdwQxgm6Fzn2z0+VZ5abovyp1dA
sEQYoM1PQF5iIHx1a+SBwJqsIpd0kYg2GlhsHWqZaQk8rQeP5nl00anklh2fZZySBRh9WYI6W2XK
lux0TqBS7Q/CdxIHHcQEqIi1LhrYZr62LpGAtGLqjXiaovVoF2OUFQkxhkxWGFL7u3iXeryDE+Z2
BeCtjKiQjQYbnwXfUgTR9xCRCt30SmKyU861qmWiyuTbDs2MXyar0K51ZTwgmdoFh2RaBYSUgMvF
9J3oj/UTPhmBaL52JToN1BKJwfX25Sd5C6kkEjfCvR+afsrdEfIXSHvUSWzh8eqx2MPXKdKhz9D1
rZqSw0UjI5+46Ki2n6cD0HiVzOmoElEPiiqWgl9Jm+XneUoA050xVOm+HP60TB0Db4x1OSX8ehQh
dH9ME8SA+eSeCBZSzLsADLzJB8LkJuf//X9yJ4sf1RUNeJXuhTQRPP9JeeJr27YgB97C32Bppl+T
y1FPrSnKil3LqhdshxjOjsMfKX9kIUG3sMBO7ysvZGHDmMZDrgd85bJTniyY9t3ynf2iC446LxzS
VJiH8XWpLw6sPgsOxJdajsJkY5oYKG5l4HjEKc86SZBkp+IpoeH2wJ5q49Q1uTDD3myf/Msz280X
ARBcfrf7qtb5ZLZwtmtqRSRXkIFnlzU16CDXUTrqp0f4FqThNYIhF/0ELKC2kOxwTpg35um7AgOM
4vkC6Sscaw1v7uxLvrpnAPzC48OpyaprbWTdYWCQtezKQVdAqpbTKGFtTvCataDSj3ZBV9xD4peB
d8QsgCDrHrRRSa2HKvuJOihKsE3k0LGKGE2XD/+4g7Dj9sF9xeQc8G4O3xngjiN+W/+aEblap3Ub
T+KyH6e7KxhGuXlzRfdLzWCVGxihPtO/FPNGrdFihb5IudP+u5kc8EgrGY3lcsjXTDT7e3pDAleB
P6WVVDxF/Z/i6iHUl7BHzc55RRehfeI34spIsQ9wNfC1SyXEkb1dPZuHPEULzHx4voxw+ARFkkhA
/GXeiQv6dCaCVaH28UfX46kWNvVoEuk9e52WQfAfI0nsYE75b2wnvHUt7B/WsrC1vBkODHJnleWp
bWd5Dl4U0TgJCCNO5BtjXKnnIoLne1Y0gtjeD8QMdFId0p1FuUUhSX4zCel+HHK0TXSStpCmUsRn
yGXRAU2wagov59VvBnbM/kiCCjXy34Hd5M01T2mxlJQo77dZSJx8s/7G9KJ7VRhmKDEeRTssv1xG
64hQ8Uv/3UBiyEmmyzswR7RO3lbpOTMzia5ZlkJ1JmKgDa5zLtNYcoAuRsGbBaAuTny0g6t9P9Xo
EZ4FgTD+bzDkbPfjiZWi6c+7OdaVBUMSiiDTsqUKQpVWwlZRd1AEPzE8w6miAmDDAp9+EcHAg+Dn
QnpwmcMLpFBYrge7BTCvkfQtWuSm2FFwfkJSDQe/Z/xxmsWiD2WK2o87Z53z9McIn27aGTziLAGq
RBiZ0/HLi1SC5auHVJW3I4MzSQnuomU8uY9/7MowS74fkDTDkKBJ53ri9fvo9dHWJumfL6UqmMur
NeB5Lkf91qTRscHTHOUzHR8MJHXmfVjjuM5wS1c0Kt0CSkbzo/UsB57y/qYxFlxTeloV+dgMQ3ly
owhnEBopIZ7ToE6IIuoRkeoM4mGoCpZ4q3v/MrotpK0Uf5GC09VykG9yhdDY97kuplrG9NJEs7qW
w+6hOhc/1Citw0FpLG0NdAh4yP5ulRwGbzVwZ0cClj9Zqe2PeIehAAmxwj4R+70eqZmmEKNNwfE5
d6l93kwMSHC/SCs7t2/vCKx6CqlhkpdlfIjfvh6UyLmuTEWm+X9o+fzMR0/iU0A+gTdz8b/mJKXS
DdKPu0CV+wJ7P+VJYu40AqkQG/imQnNuU2JIg9J87uOV3rL0hshZvpDXtjoPu/57OinoL9us5xMj
XOX1uG5syY0Ypc/RAIkdLZ99rNNxMm9OVTyP1Ap/ZkXjzVZLcVXs3VfB9WweTb+fsgq0W2cfcVXI
+t/UkgKV5EHKPsl7Dt11c4UkkCIEwbH+Wgqs46UCpUUz6P4qsPpibMuw7GJfBA/a4aGXP71kmjqi
5DJCyln3MTOf41X67Ir2Z+juk8yoxJKyf1aGeIyhZHHWv0Gyhu5bV2sKtXQypLmS9OIJ4uVxQ4tj
XqtYowZnO/T2d2NOh6xuiOYc0Vh8Kgp9xGneYeu/3swyQoROyvQRJ+r02Cnt8GYcu9h1GLFba3Yn
vk5iJwnBATvRghZ5UAuQqKuGpt2HQB/3K0EbOU6AJVeihGFckIM/519fsBv37Xc/e462l9q00ssl
1ekLgSltcI8K8+s+ajumI+2NQxqv4ll7Bb96ftWp1YtbxAcrfp5ua/xK32eSQO4BCsVcM98oiAPG
CO7vGXTOpYAt373NW5uZXQQr1WTUVHcEtcrqkCVjvCixjDoFaHOdnbRhcD21LZM7cSaBlvxSmcJG
RYzIiV03sc3vAn/mz/aBidMGncNzVR9FRWaJOupcEn41KVpzaqRMZLO3p7YlBztYKRkWK4Ob0/qh
i0/oTPqq527yUc+NOU4A/+cMgfUEUJNCMBfaoKIgawowTVKCq8ZKzuXSO13GyBdehr3fyo9eHYEV
FGbQ+Eu6dupRF1ha3cA4C7HuGXrEmfN8KxuXtRIkGBPVMO39xyBSl+pxwGnsw5QnkS3rkC7GPFHS
lucY0iMtggElFZMFGLFxnXn/Fan7cpzJZE9Sw0MDsWXWfnwpp01Wd0D/WPONWaAYcIArVEaLPtIE
56G9DlW7nMJ84soS0LmMc0O/BqWripjtd825BpHolH8cs3GGOjKoE/H5F0mBvBUND1dCQA3R+bcQ
aX2YGSfx7wF5xBR+P8+D78u9aExVZcXlvRgsd1VkSQhd4aIlLAhjA+hOsMLZXxiL25hqRyCEFWhc
PcRq5JFYXhBTPTlL2XwoOZO0MnqA8DiGqvKHkMqlSDOkVEL4Khwp+uSBSKkh6gNW4ymMkDTUFwyD
cHiP7Eqv9kljP0djaLUC1sqow74hsIzX7dniZKmBxn6pFdElRcqPHYPC256XgGc98eNVk2CTorCG
jnJjRAyg4K1OL6mDDimwlXpJDqIjAW7utY5DImC6sFz0rQAl+Pg+/wlY0nQf2w62wMclxhWJ2V7C
fB8VicTOHyN/Slk3bdqSkrjfg7dt1NzkCJEColyH5vgdpQ/y9ygrn62xSEEyY1daJWnr+sYAjg75
tZ9C9hwAhD9eeBwknvFAhyhjiuRiaG0JSVQRStEMMP3dtgBJS94+bcEt/4Ti3834hAcLIxNeFegV
PxRFYrGYHwNrkLF5QRHmT88GjwYvsQqW9ONrch+mlWGqqln0CsQw3HSyr0EJag/6PCuaD/g07CPc
JWnwXNj6+khuyjGSaQ9//3iYl5JTdBudETges60RwvTjdgjG/q+sgQHnYAU/4/zcxhAg1tmph0GT
GTSsDlR7AWF0J27Ss3mkV2QAZTzI9teGZjuJdLQtuMNdKZ2dAlXpw+ucEHdDsz8EbP/CUeG8vsYr
DwF3NoYZKAyjkJwVurgmZkLmGHaCaPAstdL0KC8WVZOfHcTdKq655nArOB27LLniuiBxTjT7RNt3
+3NhObTxaFmbVIqPaJly84pAWT5iFu3otq8HnQyLrV5iGI9zl7odcowuESwdPZWXfYrkc0kd4fZT
p9f3ZMp7erYwAoQTDXWq5hyFXRK3MtMxwgIT6qzBTQTPRJyxX2B16rMogYwPcK05oEnlFJMWaUyw
n/1Y45ek2QAu2eU2zqtCLWhQGB10S1zhD1E06/YizKNatZqHnx4AO32M5GLT44ktFmRWf23B5H2/
L10aRG4MAyOUjpAMmGksfl2ReDohGYom83v8VNjOXwJdWFZI+Pq44NV8DEbiA+yNjAnsvd6mH55G
7mZpassZ6puBm2XrV8o6pW61Xyk/6OEFbSN7G4Ym2zvAtWBuHvdvV8Ev5eMcw4DLU6ukY+KoCDt0
eoaoq1L41yExnf395/AcHucP2QCtXhu7+Gzk47dLherM60gx4ZB1uuYsFtbVvB/I3qk2vvIvq9SA
7jmeBpMjZUP5GBPN1Qb7s+URbXjnkxht28+8kDc+YJ7n7il8czBjq4ldQs/dw4SbiJra31ZzOXVT
eKDnI9j9KKGtCJI4Qie1xgSXj+UfbrLvhu4+pvyZqfQdM5p5hN3UQgklafsfGk47DWKMpC7wStOL
Bmw6qOSv7zZCIOKx/yatobeBbPY7qhbznjINBOhFAGgOAg2P9LGNLxH3ctkmCnw2+jZKiBMS5nR5
mUJh2sMB2J4CqIT3dzB9JLoEHnSDkjoVqLOOpaqn63lFZ4/aejWEUvglaQNsnBAZcjVHd5u7ZFML
qwNINk7W+ltn895Q5lFuhEpIA2LVYgORjOoPoaEUhXB+2Pddx63VvslS3UqkOnXY9LkaO3OpoN8s
zwe9aa4sZHXnUKq3gStX/I5K/Klntn+KkWKfi1/5JChGIsoWdajPUGpk8FsN2dEXS3BXpLn5yFf6
HtDa+vQnk2umRhnxs4m1yV/b22yzFOGHFE/xb7iDmKu4z8faRX3DVNypM9M4IxIVbrP/thEU4TEI
AcmZpKrfjoc5WDZ8mFZ3tTdwqoCWUGjw93OADimj8Zm5IZ4yc/L9HUbRpZWwHF37RlP1JFXatyzX
RXqJxPJawXyRL9zoV8IHx8Fsj6cOlN1sev0U++ruBOCg5skH2cB4vWhRq5unThgoPEvMNFmNs7GF
0DX1LZUewcBwDjluD4cUMfurg1+y5nJ8VJvyMcbY8yK6BjDnJZBEAKfuZz7uLJRFJeiODdKMG4dn
04XBTUitEfwABrAVS5+/h2ciLF+3rOLJjUPsuZNczN2yYWrT7OdvQaY25O13kRLSJVwDdiAfN75B
X/fOGOO58breLotqM9owvoYt1oh8qRC63K1KYgml2gkahxQZ1oeho3CFIW3axNvrQYzY3MywWOz1
HshJ1IWhz0dNbuXVsRpzKLmQcS7ur17M3RaXQqCYx72E6Vxjt0xP9L8QegGpXWRlbQ5vt87V94xy
1TrPR9EApMNW3wOgPERoAL2r82JBBsXAzaOo2b1Cc79tff+9kB+kxMUxT15k1Av62CIJTvoY2V8O
U1eDZ35Zf4VNRw3/ovq7K/nLbhkcMxPMJYl9SjxzuaBdH4VoO3yvp60mZSNLiSQ4NG0hclfBCPkW
hPIPdA3zE3brL5vmM3hIkNzSzhtr2bUo80oYrAP/WVWovlWVQvCnnMZxfKvNtTO1r3XGrSpu40tL
q9TKHp6Bp1mxZq8WHkmoE35z+mZ+rx7OuEmVunih0RSdupxqyZJQF5lM8rViAvpuLf5nDgZr/Nai
9iMmy+Zs+acatCExdyzl2Gces9AmQsSg+4EEPTiS/UwDdterIyJB+8sxFkISro4vf5S6HuKlRK36
FmpI8RAqcRFBzMIGGDIYdI2CLAFExgN724D5W5zHjEztpIxmj0DZM+vw31SKTsp7Cxcvhd8Rinqr
YUf6t8iAfVIUjcBw3touZkLj80h5k01t5F2yLKkGLn8g16fMM1LqXP24D48ogAXXpnDfDrWMa597
YBXY+LesSIPkzZbUQqQchTF9pzdSl1wIVO7EWOH+NvLM7EP/iKUA0+KiQ25qIcoK/8ljAQ/Q/Pjr
hG1BKnULJPMjZzXBs/HPPBuENEvro0mplie/tpLkT5jT2nO2jLcRWLWTBS8dc+RSSf5I8D3iEuic
5JPNgCfaH11Qi1un4zRIg2k8yQYQIbEMmxfSVQ/SwytA0D5Hx+Z1MyiALeB93TBW91aV2rc+U+Tk
xvzIfiK+fDKwboSxrlACS+roo3q/5L53tSo4lTbb9rMkeTd6mP625SvZvhh2vb1guHmA/h3TeUUS
SvvtM/tB33ub+4MIpWHYJDKtGcrmY/Z5Kl4Ewgm0/L612+5b5CUBHy4RMYzrQk9Ptx+VLZZGhw9E
k4oBDqwu8giqQPc9E16a7L8qhbIVSa6Lfd76b2IuF1X6HduiwjqJFBSIRp4I2UaY2YYASfYcv+BD
m+FQBqsosQYCJZtrMDi6kK70tG5shQ5JpyjEJdL/Dr3qe+UJS2+pKlL4AlwmqTVxeCdGUVeltptS
tMz0I5Ia06vxKHb3Vd2Baq2/5KxICqnL/obJ9p+Jpya0k15PZXXqCgTI8Sfa6r7VBT4FtWQYpwgt
wtmT4v5178pQYpZOgnBwb4BiEAuak7zY7E9HR1D4A5OabdjmgnutZd4Zm5NzpGVzF2IEPd9lwWVl
T6CJoXcSfnU6R2fxXk2oyx/V7r/X8mukQdC45+6fPF2KGOT5hALIOMoSwJ1Cx3KJ2x4MIByZDXB7
NlWIGa+KwvxWzdTKyO/yTgzcPIHbzG2MDHt9SM4/99J8OOz7QJONSO/fCI0J35WtbnL2DnVisj6C
r2Too0Ck+jIqHpY9BbEmby+aEkvOe3oqjsyjuzbhDe1kEQFOvLlE9Y+n+VjGt13J5nVcjCu4RHzM
pHdHcNbyzhNzt/qdYutJ4EBXySFnP0zb/plPFS5EbeCn761dZ/VGw9gc5Jx4bn6BVDiPi9RZVCxz
F16qAtGzn2G+TEAWvpRJbQf/A7nPhmhRAE5oErL4fyo5pcJegg+EmiC6F270cJm8jBf7BL0uxaKt
9BmLwZLAD0SGkzBa3fpjkL5VZA8HdaOv1Q1M7yCky3WcHRxCbvUUTzFIkUEvLIrTf6jVvQtNP7/5
je7uUgkJsWbgg3MuoLBsB2I+UAFA5Hsm5hoOC9sW7RFU/Ei7237xncXBl22xv0spa2pch0eLoBpL
3yZxWiqnFRRzZuRQxv/ESlFb0SUKehh+NiKPbWu5srOzS5+pxsgri6jfClaTiC/a/Dufxa7HxWmk
haaFjUKR/8ov8ArrrfZPAZtnYM+55+DUn8pLQoC/94amBzVM/1/+8EU52cnPLATHPQdHt/G1CLXL
yVNm2Jwf6GkC3VDFNtMbSuS3ZhDHxUksJN62B8tVgANkxa2ZU7kjUkOVrNU55pIW8khvDfQUiSTp
CN4/5P/cS28mBjQwvE3JxeMcrv3aDUkX0pdcbiucbfW7QIvT06Vfwoy/rZbvEC2gje4JmSqyP0uP
euReE99FT0afJPPXSJpDYPKzllcLPS3/AR6bHEMJla2/2ghjKSuts97KAbsT6bonRSQrcbk5tagA
9XVOSX1srx954uPOGI80eqaYXlU1uk5WADDexiodfrl+9E8sLR1EBb3tsQoDfhrbYAoCxzfyovjt
oSDOZG6Sej2+3Rui3DfVQT96XefbpFhTPTX5YuSLGHM7IpyEd04cb7VHm46WtdrmOGGjejDI6XUZ
5hNER7hX20upRiyR/QWvqFdhA8lKmA1E5ahO3x9ZTqIeABzwRcU2TTxYsbse9w1LnwDme2cnxQBw
kyPRtMxjGWAUWJuGldC7Tvffq+lMYdkEyXSGn7AjuKlSt56hcmzuwH6QKHRA/0kRihCBgG+RqfkZ
bgv+g0+aRrStEvtQCi/+P5V00IFAr5iZ3WWdumj7Wo0jybSqUYMkkP7OgGz3nLjEYIYkEe8k0io4
Z3qJyVKM7w35PYTFrp8EOIbnnaOL1czJD5n5Hifu1BJ5drmmhIXuHbLs25p0wyt+ZwZ64j4DED+r
vI54duwYEit6SkCZzR4NsUMdR70Q7FyWFLgJc+dq/jZpxw3MmICWFyBJ39AZiZDthuwUQgFNG/ZI
I+awVYL3s1Bqnd0ayEAkbW4GTPGoob4I5kFMx9C+oxFir2EjBsuaRg8md4AsbwQoMGEMP5m0luh1
bRpD14LWFef3ggIxgE4tfwDaaUVnChmSXX7u+IDy+nUTJxUzuFsqx0WLh42kbClpkhhGkZTSCSGE
VAKc72wVKREhU1yns15M6CXfUb+JyIoVL/kTP508xzdI+CmrBGnKkxmsoN3HExQWXGv7gEXrIlf+
37C+xLhZfI1QMe+nLjw7XyXM/30YmosNQozRMeQnWGY6rWd4KcRMgP+q2yBAC3QpMO5Wngme3yu2
C6fIMxwbVQubaE8K/5ehXM4JokVW5ptEqna4niwYNrYzfKhrU7ymXnUI+yJGhy5K9TzXhQ4Ddcjp
+Q+T0I9o24IeLxJ1Yy2DZdagH0vlrvK/OeemECflHeGBcqh0NyYw9cuif/JZrHHMJTZ7hU23aIpF
gBnHi5JEdUpftZWKdhRL6PQNeY46LxZxRlLx6Hky1xUzOpqiH2I+PsCQgDL9WzXfivR1OhnL3aa9
tem8OnnX45K2Emr2tBVZzO/91y2YAR00eTeOcUhDuXkCgBqNPCwih7ookutZnAbqSsKZa6FqIrzu
QUFHkNV5nhIUuODFeaXIdnGhTuI7X9Lo00vUKzXXFkwH89Bu6kuoTvYLnvY4ZwtilppbPKQyJnwM
a3bfavBkxIBbn7sSUsJLmGbInua40A/MlDweUAiujPX6Pqw90pmc6IGzwjTkvqHEgd7ux6G0yj3i
/XHiBrqk6JNZrh0ZooU0+4f7Ml3lcYbpkA6H1P3Oow8ksJRVm4+HRuJmVyM4pLB8bx2Lx9+O+JXz
aNozlUbnWSxeIUJ/w2XTy8acRhyfTWQJuu4L1s72QnTiQKV7V2onDUw4ElZmPYrNWgo6PCylktpm
aLwSZqHTFZbeQWHGR+D5ehd0N/feSxFHK96J8FX4WMB9EB234jX02KX4S2UdGStg6kUpbObXC9da
HhIk9cFDKosJmVTMusG+Quy+UXR9Uo4IZ5GVz+Nt1CYwO0X4eN450nMWhirjWbUjQXBUZtTVT2vt
2W1zeiD6MLz85/r+MPcyrn79qlobfXFjFJqwjJdQWG9r0WOF1lAsyoPVUuhoOMmq+SoXMJuXBCbS
PdQvAeIUMF8HPzb6tJh76T/4wBQoRWyKsMrn565C0dAtpAP0WQWfDHToQ0wSMzd0a1i03KgSUeoH
Ih6R5aFz82rALo+s1ntnmt6pm3rPDhw9T+FVghW5t7m+58b4iA0g30fyvB8Hj5U7Mspjt01eAZoW
HqvV4QzhQTbF1d7EfUXzGoj+6hUo6AtSD7tFM9UFxrNaJvlJpa3Xrk+I8i++rK2MiHvy+C5uCad0
UxoxWKHQwsH1+e31gwL9JqlhGgnitoai+dUXpbOuuz9W0mpbgTsh8rkgdQJ9RQqqyqbQlTgud5k8
Wxe29ThaT/ioP1N91v1L21pl/7vOfUrrCNGvO81/7sOuj4fxL+sZ1D9hN/1KzNFSJtDEfMwf8Eo6
vsGL48zUy1Q46DwxY56m4HjdfQ1WAHotO371XAKdNOdMFwgWoTAxnzhX831pO9npqJNI/V32YBXK
bK+oEPRk2F0vhQZgv/qEWoWYFGmbFF6uLIm0i/uZKZlAhRDENrshElfh1+tVZKNyXbwGKMUb/63R
k+I92pcovCyMYMnKDe4Z4BMb0rok08Tq0RSxxReZ7tWJR0q/zS7fxoVHVpTc/qzaig2JcTYCDVzW
uaru9W7CINrb8VToH0PHuRQ1hez0VTXQXjsn8nTAlS4gjNVf8PALCF691LBbCoLU1V9VueSewpXs
CZ/96spyBK2j3KSbOghnRMuKyZ+FzniLlVRA/QXHzNJAj6gVF/Z2nYE+q8HhUYlorX8Ytv3K0y8Z
YrKBW7mzdX97J9tz2WdgXjoFZSqtlLYtrV/mihbYMk2BsktZGBnZLpw4BT4cn1JCuzuuqEYgBH9w
C2IrU3R5f7IFoXEoHqd6Nk+reFGpqBjU01GJ2gkoWQYnf4z6lGIkZdW6dBB1uiSG7tMcMdQV589s
CYHJ4zEuT7BcUKj5Agv3sFYlRKEQBT+3ex4USSMo9D60gCdYtP5Rwjbj3MOegO92faGCNOaGgOWW
PaEu38xadlbLCUcIr5Y73IkmwYTuVwXIBg2Iy4XzjXJ4NqvkPsfz6F4NBQFc2vONGvvMYph/Lgf3
o3Zl50lvyXTlr1+Xz7eMP7iJvADKvcffvQ6MUEWBQF3exJVJipBEVmBGequMmwcu9Jw1CNBUPbJk
gO71JxX/ysYzK9NV/6RduWJ/en0h8D9lkBNTEUZWjAA9BhOofvKLwl27uOkmldGviv45VItAknET
GXq4vCTW5TekMJ3gzwyvCzDca6Ra3Vz9AsXRCotw8vS3PBTSZclgtJnBoPmtmbK/nkrxUQEx6aZn
vFqJ4RF71DoXZ5t60p9d+KyKLRgpXcDFuSjEvQ5isDsqmio+obdUgQJWsZTS1P1+ZnJv0+QOjjzQ
SXB6rUIHZE9KgUAguryp3bQf3pQ9rIMYWR5TkHEGw58sah1mcUpOEX41CbuCayZCeFOLGcwtuCsi
/qX67HeFW4STrTrdL9hEGwSOpdRA3x63asfaQdgqjr29vJTwIQBfDPDtdB0c5w/LZSqIQurpxrua
ViAm377MBTLbrmlCmz4vWLjzeQITfrzKATqoypin+s78Ah6Jq+qVFG6aveHZimYY4MZV+nr6GoSr
8Dn9qqukkX++76ZwiK4ScO4ak8Z5I8Kmr5j1FPxdkD8DE2dPFmOu2T9zm2pRRDdkE8XOd4RMXrfT
4OCEM6b8Nlqm6sXu7l5yffO85AdjzhCxI4Z62BhkdbtyJim4NOkBJZYlMuoXlwX0CRhbUFJJIp4S
nCRGA6jEzRScmRHkP0++2AyLccS8ZUAEen8ZK2tMTxOWPgZ/8as3RveDTgsExJHIr0Rnx9brX1BR
i+kbL41YrP3Bfqv+lqkOM3RhxOwHzxkDP3sisWwWeTINzcVi3Hq5seMeVNfuaI8eSNTLdgg5xIV8
/9QH8L9x7L2pDCj9t8+VJwlBlTln6jfMyNqPW++iKJAbD6kogOgZo14HC6YnMr5BqepEs40+P2V8
g5xfK86UPjJs6mJNyZhE0u9ptNn55ssX1OQPgSYVozYdUgMg0FiR0cGmJgX/MLQOpc+yIz7P6aJ3
QZq9szFl39JUx3FnXCXKV4qUto82leTZ5BXqddTSOGVctvsHQ3UnYo60KLBSr53L/RsMXuzApl7n
B1zUoBdC0XvI9rUX9WvwwCetgwqsXpnlO6nNYUTz0FPZr8xpdAmtLUoZsDOPVgkBCeDDFio+kCAF
2ImdVSLcM9jrdaYDCHaLkJ8TH5V4eyOxkSX/AsPt+UUv8roBlvZ949BCx7MUz5eJuRVJJGoJPewF
ZWeXC/J4+3k8fyJIVqmHDTY5KuGJUQoBHy8FJUH+43kAK8xlOA0MutvdXf14dUVp+kayvP3CY6XJ
jGN949FacXHE41yrJFBMk0Q3/tWihmwENgQwlShmccxbJJAxDdIhNpp7WgdpO52iSzf5xecS1zA5
u8rKa/yeorYpF/WzQDMRnbU5somuaBlczkMqfHVecHUVZpwYtS5bDyJt6yfiGknIYPczP+lsDCu8
UheWS0HWOIYvB5h8tmPqLAQwjYUbLsP3iq1JMbrrXLzphvGszOid9KMcM9xqtaLsFPqjfN6+IY4u
GqvahegOJYDRFouYtTWYK962ylne/AFYCSiE73423POJ5D+I59uBVm/brurJOh2JcCCxkwfGxuOL
hEW8MFTcIU5AA6QHry4iG/egB1qJwpzfVm8ZlAHy5k6dYSOUNCIy1arNJxyy+FbiFU+wmCjf+7mb
Qax7qatCpdNSyi/nA6O7rKmKSFvOmPXIoLaHIwtzjaKEAWvwQDo/yf3L6OIpndRzjQqNPlmss/L3
vK+kMK70E7RQPjd0ySFcZ+G3whcBpGFkh38HLA+oSx8/IgGXqEl2PiqlQjL1RwToRfGTLNtI/aSD
EPeEEhbu32pGz0lgCSkz4zmNFWs35qf8wI/u4bkYrUBQXtDHAje0vgpIHzUNtCwsig3PVlqUa7GN
UX5e61g0zRIQbNmxz/go3ARaOT2qjYobRoxgc4i976rUXaMuRbrb+lezL6D7lfwYfxejoyupsV+s
fPMdUulZRVLQekstYgHHLq/jkq+Ju2OmSqexeFH+8sIQPMbMicyVkn5cKHz//2+0O7UEU0wc1eoU
0Ky04QuZUvSLleofjYP9VNkhudf8NH68l7ZXIdSpuUDYyIdx4QptgqmaJmxt1f7q4xEnqWFApTcm
cfOBb+co3Wn57zJZktH6yYRqv7vqPgqsefv3U3R3QhgZI8NW6yYc1CM7kQRi1ZxMemyQp3itzdpY
+x5vTQrIBKMN0mIwh1uqaRL8woO89VFrhPi19nyj1nLnqNO6DdbggHfQeAljf6q4phbzJB1RE5ZT
PAJ1MtefCx/rzGI8ydRnNvVRSfQ6LzW351wppaUoRaA+dGmNqSI1mpEV27B4/eGqZJsDoliEst5y
+/B+i1yALLyH/3WbF1KSK/bE+Tln8uu9PjCDyotce0aD8AjfGzqEbw6sks1KFqQOeyQf4PrO9vrf
DXHL/3rB78N51vBDak7Kb4yTuHfMhmwQ8xaatLThfpwt97RJZjtpfKIqqhg5RbCCRidUooXPryh5
lWxjdtcKHaqg5TrAHE36Jy9ZM7Y5z9zpYw3OvOYE4lPMN3PVThc/bJvVXW5KgIVhsXwvNS74oOsr
ErsQ5NF/yFbDNcGKfK3u8ecAIpIoYoviiPQJIN2nCVP79VEUFqQv6x4aZZdf7AVsYVqa/2J2DGLX
tK/0PZ4bRGYb4nHH7JjFVbYd0MbYuJXM9me+WldlC7qDt3riyEbNIMm17cl8C2HEHGzI1sV3U0Fn
G4zkBUv1qdSLi3pze/w6IIzN+NaN9VNAiBUXGzHCEp7g3vjD0IwQhaJFBntQsu/4YfCHwNi1GYiQ
qETawtYUQ1TD9/PRCywqYuO+mJBua4b4fJe6gX8YUI/lnQ8Lj6lCcmEMX76P+Fb++n0cm/Ilo+2r
XFS+3rVW1hb4dVhCrdBrAjXb9hHBj393945zhWG6+dnwK7jCR64hTTqnBzhOqJcWVG6Lz4gmHgwO
palm4LON5xFwux6jC6vg7rBntA488xyy6iLKDecdfko7fthSTlJSlxYAlAZfoshSpN+uFN3ae02b
0K//p0/Gp76/v0OPU3wDCkKZmKEdqVWuHPTOMErj6lqEfsfWMQTFHR4yuEmiBmRxnbNpAMXOclKz
G2VP6nEUzoWUUW2mf00Pw0hQfiSX9N3nvRdETJLk/NqvVFixoA58RWa8ZJoTbg3JEszinwrEo6FC
sDR4fWJTs2vi6JEMiYUM8cnIOIpZbDrSg/H3/63y13f+1rCm7MDSblSXRvJrSF8f1ho3ECggMuFC
70tfUc9kJQQzOqj1Kv2pAtqJsKllrnj++2dBkRa+uVJQWmABmITkp7qEOugLBJUtfQmURHjLlNHT
KW11FbLlyhkHXgSR6ELpFbE3AZGT+2eEuBH7iOiRJLUMKoUdLMMgBEMSbBbper3+EfFxFMswpENQ
H/2wERr+wunDrcSKFwvUN1GUMUofuynXarcyH5+zwQi/PSm2tVJeiZ+qB83rLkBoTbBtVZ3et/pI
uCO1B7w+LKMclNeegzcXMskm+5GQTRCFcHSR5IYUtWOhQ8IjD0YJ8i8su1QYqUrEYwpeXsKMB+JT
iP9+AMvA6viWvM0O67XWkTMmoHMiNbG0i5CVC8TDIJyC0JLSJvrole8x66IACM+qYaX1Y5HUHaqh
TGE6DhnX2GLIMEtjYgvN6rZ2oWMNaRZnsYNbwhkv4fh6J8Ztyr2fap3vY5TLLSSuo2SGdMvFwnSh
Xn9DjJimD9DmKWYz1yCZ5K0XJmY/5YGsjip7Dx/uOCzWMrUJQKvt3oba3jqh6TUUm4vuxSijh+hk
VWDn+t35hAuopzS7y+OAf2iF2F0/OHUYX1Beem/oKIgrWd4Eq1tvmHVMzBKPqyVX5ymmC04afR97
dQdNU9j2azdTJBahmBRMwhVmN2QQheiaq9o/b5mNJsg5C5sZtUDbkwhdxnsi8Y62NmXJSYh7nKlQ
4WR5Bn+7Zt8ZsS1mGTiRRNfohCuW/nWoCebZU6hnpe9kV4j949M0dP7jid9v+K0SBjblPUCWWztt
FMh6p/u5vL2bgO035GasZYD2EKovzw2y8u6CaFoCaRuHIYlMTQH9Sjaqqhpg2PsrECA1/ru6xpyg
egrwJGcsmD6G8icbo316XkaKL7zMblWJoxXSbHKxwh1h+Y3QqrcFyR4ZkcOJ6ZCy7UfTgayiKdMJ
TpR5B57NZsqFbmS42tEaIajahbb/shKLJQ7RAY1jaRNDKPnz4K8lEqSqtnHYzQzT3Ns07hEfiFJR
G4H7Eoj8UjYlOouqyAGqla12aslJujP+MhGwuGkzRyCmuWzxWVIFjq5oxQ15Si93hpHV7mPh3SYj
J+LJVlC8THv7oTZupM2Ys1s9Tqwk8mRWDzhhztSxnUl4aheggrkFXXO4FsAxNdczWl+3qyxMJ6bS
w8RhwZWJOGvCFrvt4PmYy5NqC7e7P693wLJ58Q9RGK/B1iTfUbIoueMMAxnh0HTBkITHyr/Z21Fq
B38owrOx6KxQRWCcVBMFh7mQM4y5ThybryJ0gASEqBIZx+ig5I5BrQQ8PbyEf3C6306Gj0bABrUZ
krjqXmxtTW5sztZWro41qkCWhK2Z5W5MNtD6R/wOQSXSAWnOgCE7Sjam9UCkyVymih893lrMOjOx
i9sqJVM+N07bsUyUXOLAYycI3PZfmXdWTs+FbFhfOY4MKhEERTBI+mTOYpqnzR/pRC/9OVtme2AH
WJqan60EknmlGToWnNWuSzqVoc03b26Qsbq70NFnEcJrl0jXIKulDQoANIaxYOZfPJRBpDwH9OyB
xs2oPB/gJwXkDJ0U6xsNXJJJQGF1yBRM6Gqs8nYuSlSq3GFe5nV2TNZc7xqcPMfHWr5eri8NCV7X
jbxedxFiYvcheAhZ29b/DPuJUHLdT3DAKJKdW8t0nqEGfnsecAcxy0QLyrWjEP154J/vJ0z9WZ5W
p01ZoNzCVV4CCkP+lWw5DbcldLZTJNIhlMkDgybwldcNNeT4txQ0uj5oazmnOWsZBFG45gQtQnjX
Eb41fdle/349LhmJpqOVh172/JfAGgM1yEltLwc8lPU9/dT8nehn/5xpzYrkl4LHOaX+1IizEQAy
a7OGbB8ABiDw9Qw+YrtptRmDDQdE4F4+KaTaCQT0OiNHzGrs6DWKKX5uOapDWWv0xuyCzrQ6FvsD
go9yL7SObUjrYwL9m0W5pVjmRhyasVQZKAdvVNs+cLtR537ZI9WdymmMkv+hnzgj664umXZzqOto
aj4ReYrIwVV+IU5nZRlLrYWcWYaWwSNQluXU4jcyE5kgLSwmVh2MzZSNhF3QF6/e75Vk0lNPNJYj
2C/EpLvJltv0L1g+kSWwMhXs+srEy5YdjS1nUtfh7dOgkZJF+ePujEktzQFmab1AjrwdF4cD2g8a
s/yLD8DbyiLferMiw2+F0koYnJyTtJUD0QhvsHpQSA37poO2tT79LGguv6smYlgCOMK3Xkpgk+xv
qoowqRn1R/UjAU2QTH1Z6TMSIyzta4zlKaaBlTCKW5H08Kr68NrVYPCCFJ6Hj8tadkbCYjXurMaX
Ho694FMiocewqdNX23ns8/jBRzXUGqHMwzzNgFN1e3Phr4j5zcQFBEssB+ZUTY0p614T1EVP1qDg
0kX0gIi4ZO5VVJUxivambE0OzTNjgs0vzdvr3iQCYcwBpqLfiuZLYOTntlmEfpcTI/4vZBFY2Awo
uB+TzL6Oa0pAYWoQ7PpT/pZHSJBa9/uIGh3j5zGbskPXB5G6Hx0yRDu/wa5uPOZ9RuNyJF7EmVf8
lCx+fuhs0PyuOENP9MCW52WePZwYZgvaf6ulvt5wMnk8WsT6LS1JZUcMVx76sH2K7ZWX6h32LYOg
068ND0lrosuHS38f+QEXZA8qdiJT/RBfQ/9vNb62dKe2c85XsHKRVqtFBixzbij6eBf+6UcxvYkq
tO3q/DV7hIAWfkYnEl0HHwc6nOCKCJc8IyrQu0aUm5fWglvZbIJsXds+HD0cPSjw7bvl4BUR15/i
qjP9epXOR6Y4iyTlqAi+y6/e2HrWQUSxocqiEP2zR+q7Bgr6WcI8CDhEv8XxnYzh81TwhaT3hiLv
0r4l2604Xqnglt8Ng3RtJwsWtkH0YgWllHEZjuHEcI9T/UnbEemRDLqwh4h+MvnpcTubfeK5lO1u
A4usmUWOcEBrfXkDOWDhuE0g3g3eM7XCG8UhefhDRrXnaj+zU05dD6LMscYDfewlRbtSMy235Cjx
Y2/aH4mNCffNPpPFiztngh0RktFGfvydhbcGLJ1JhucyGLSC1aaMun1yd1CmTDOSoSYQZKNWblmf
OsqNgf7TZ8CVAVmfFE4KljDYV50zTywoYFJmwDhSFk1az8DtKCfbBRH94Q4D90tMsmjWnpRXHWar
fwlDHQUZ9DsnwApu0fdXxpHANeeh9eggUQW5GafMtfgqsXRnVYCvuh9lAFBioyfqjZdAhIHgexSt
3MYiu3qI1FDxJsavmHzC4kRNEs6KNpKPpK3chGcP7II/jdPdgEhXck6fF9nuByMasPDaqJl/+8Dg
URaKOnmIkMZvCAeprH1kx1ptDS9enJcW1Fig4QH6QvEm2fGiaBO8YxNn4zxhl53tOZnYUHTwzu1q
noHO1dw1tnPO/hEa4bTEXGHJrPa2ZD+MplAIJaYO6EcrPJVMgiOcRWPTktuA65I4ATVtE+Jt1WBg
nL5Xv/DKN0gamoF4D+P1E1sBm5bk/o7Md83Ji0geATNWu4+wh8+ygBuuH762F2iXd6MwF0F1BGdI
P8vh7aqPsLb6U5Ivq6943VzVuulaWrKRbmDthSF/eHiJmqhMOkxFH45yXKreHqiQLklH/wTf7uYH
OdP5LYT9xH0SkI/nLM4818xkGuVTYbuaKVixXN5hwvJy2I3wyMyoaEpig5/zAgHQszvj228Wk+y1
3nfo5ANcr5bTKjp9cTQTUAaoCEd3zJ8BXw3+hCk9dAf3bLWPAoUy6Hcq78Y9Xpovoy2dpL+e85/4
kkdkDcqKVT0aBqdYnQxWGvNzHs4YjiiHSMNr6GvdO4x1HkDLUqnm9kX4Mv7+gxEy7Gdh4D/SAQ4l
bghPbCNASBGZ5ctTs2Bk3DSyqARwl3JwU/Td4w4Qa2Ktmwmv9jHMCowEvTQtfuIvmgdRyt6MfeuV
1ei2fZ8220kCGN7fh6VLWCM+juEIww9o3bBy8/79LqyJEZ2LyefFV1KSSpBRm9pmugB1tpRYOlQ9
hoPRbXyl2NFjwPQv1Nd4b6oFpQ95lC1mFpxZnbiuG/PQOktZbVt6yVqBL+BGPhWdCYSUOpy0BBRE
jqPz+h0mi6N+wB5GfFlrBriDG7PfeAZc9GPnvOrSogCkkUklbQiyLJuvaXrX+xeAZHVt3MhPIgfi
s6kmsvHyp3I0J/DtA3XIwTO/G65wh36fF0Og8OwICMr58VLV7OAtttGSUAYsxIUhpD3uXuuwP9gM
Fd4cleOFPckPjOvqPep425iYeai8oBhGEU4QFYIYKI5voy/H36LPM+1T/t3ISVtOim0t6bnVTNl4
HRK8E8foMRn48bxB/+GdUeOWfbhJNmE0rvMudzC/BdL/poUFUxUR5L3cafUHGbhOhChPWal6W289
1tV1GZxvroWLVU7ptm5CoWtJGz85oZJAjWfKXcXbMtx/NT1ZbnkfvW18t0fpM7zK5kdbAe66Cu7d
gKK7Osy+9QNHeol9M3QffiHrdI03wtN8FcrD0um9B1YZtRokSueLt9iE4HZYzBS/ggrdMn+wke0i
fU8JBojxJdRC4toJWJLzZBHdQq0xUMWGZzjYA8kYz+GEJUBQPf3PPJ3zKhK5g4NEXZn0qnwD02OA
ouS6a+HA9iiq30VfQQ/zlW+t1HRmCuJClhxw3JVjQkZJm2RWvxhbTgSBTT2ZB1pAalJs+ApZxBVX
s2AyUG6OIUI+qBnmnuZHB68sezIgjOxPC8RCq/KQvvxAmCVXyUfoNts5bUmpIeA4Tbj8r+AJAYwj
1gdSXNx5oWRy8QHLCYOt/xG+bzPnHVs43FNaWbK0XgDDmQ67sZv+E0PH1rqdsbPV3L08pLhPjWyH
5ShW4TsMO3KX3QGPC+rRFkDzISjVcBUG74cFc76WUbvl5fT/OZ1bcO2ngJ5tNKl9PhjgamqPR2U1
dv8H3UvTPhA/F4chTzFaLQWGJkFtZWNo6swNbxJ1rN42ZCNSbRRzSpsbTEfI8CfgHkMFziRQikQD
w4Jq2vOMAMcyrEG7vOShjOXHu3+KxiDI8qe8XxwmzbPKmqBpyJA6StNnL0hPWyz1SP9kS1plfoD1
c076S+Ub+pkmqf8l22sfw+FvZmZDXih0JnwZ5HND7o+Y5imDPBgrktXYaK1viw2h809tznP3eKrA
7t6Y/vN9VnLJqGoSbvXrrv5etQd79cQQcuMr2KG47qrPAcCuX8BFtGliVR6IMgXPhPARCA1sWtjf
L6kBFh3+p07nVUwBxaNyWCbbFMNaidfIEAGpdT1q6wG1Rn+vcqpOkyGMKmkDmLEq6bcRNBKihXOX
PIgHt8XYV8oxs/Kn4CdOV2ssptVrifrqymteRLZvhP66BEDcuCz9pXnRBo0vfDS88fbQW9vJpqho
0hk8s+r13Y6oYPey+q+O+pOUowRP+RIYRpfUeTapzn1LTM0VWNQXN4XXkBvmJyo29q0ZyRzLA1ND
5HqEsi2ZdXpVLupSYDWR6WshgJzYziiqbAIN9kdILAKi/JjZNLqmCX4uHzNCZpNCpVA4qEn9LYBC
R31qc+3HzgfKrP0g6+koBM34WMs180VCmpO6MOYl1vwUXdpISQErM4w2zUJKIdSS+4XnNtKo1lYP
xAfqtKdwNtdaArVH3F3af6lGkrM1Bb5BZfwBUwLuHlcvjVkTbCq6bfZFvKeOo065STVRWofquCZm
xbF0eVpmw1Vu1xnu2uZagseg8+Imtg6gb1cYt9SUmLZwXNjPgZQPlQvPPgu7BtfX0GqLBCvN5BPH
Nk/DKtnK6AYpO37kkLPYG1inehTY9zdJAokhMcwhANtoMnCjgCtA24cxtgYDrcN70lfiEhZ1yGiH
mHSrfjQASptW8GySQQpK1hH0bn5blLb5HDPa1sjLdC/PGi1Bz7NxGnIEFq/9zGRuYPGj3D+9SIG+
EuEjLDkQcFPJdEl7MXoLS67UZjrL5OXEISmp5gLpLKYIq6C8gEAD0bDJlIB6XBP7PrTA8YmAPiih
9JcJtxZVakut0We/Q4YyKgThQhALbNcX6yQmosTMYD43L4x2gYpJrCtiYAfSjffgMbedx0ZQH4Mi
VW5hB7jXBM3E7LNXSIm37VA8/94ATE9DT3DmCQqzBarms1j4UzkbisZ0orUXa2oald9Lr5sykf00
A02iHEtNDMCf9zGXhfaSvBqx/00xnfwR5uVrAOSPEIWnWIjCGoE6hIvZDBijpzkr3GmE54oqjmxp
pXk5F3czRxen8P+xn49Xq7uMYvqRF/occ6rdzrwyVOSIY/XRvhA97tw90ulPNxqmUGsyY2iD3kvW
S5NCQv7/FkuxcwDR/6VuVwAYVstaQF7gX/GjmO0dkx0c0t7GPvMjrW+KtzDeABWOo7hj4znEK3yM
qvLoD6NEmYgq3z02G2cHNR6B/jETi2ygQ5bHQyFSSsiK/QibVO7vkUAJqhTk0Y6vR2KY9qLIl6Bb
Aw5ycEgloPs6yXPOH5uu8N5AFK4YDFeWC57++pe8KhHZtvDwlc2rFGkFNNmGRasqiNK+WpZFaar1
qoF3NUQm8eaE5Q8Ml4H56cF8DJX7CL+Bk7GkgukNF+1ejA0Ac4cIlGBE7yQrXnQTjFtECDZrQrYN
50cQEyR4UaDrCFoAmW/ZWkZS0ZiwDrCXCZOgK1H+l4FCs3yJEf1UwTtThfd9bd25RqxP5KQN4hbd
Fbzmpho/BzgpwPJIdi+zwN6I7Y4CxENKhEfY5w7LvqG+zTD9/wFotgLv3Uo56LsYUoafh15N1ChA
nbeRNBmsOdCEVy4zttA9joqs3ckZi1CP2hDKfinaqNgQgDZZ+uz24siqeosJsEe0Xc7529qdexF5
9NS6cY63D665+Dut9C2G3Q0kQknBxO53rkJcxGYpBP9GHWs4AmS9OQVzvpt08Fqr20UwRPqIupVG
f/BcJOj3iUcM2Thp3oKhF7vVHv4J0JcPfAt9O7ntVH8bQHxDOzglPO9mLmDKtmArEEW/PtfWGfzb
Zi4jotKoU7WyQqG1V3updQguCPPPuRn09exNq6774SgY4Q13oeaHia9K7yjybejkfBZtpUIdENTL
f9gEOjLWY2ex14tsAAjR4ItA8DhyAiVaiQJOwHN5A9jAr5A6N26qUkrjj5oiGlxfky9UPLwMmvio
t+vQ/Qa1kXAFZlk4adih8iebiD7+E0dUFKr4Hy8ePAP/MLfVUbrzwCotvhYP213LmFfBAXldAgeU
SYmiGIujOkO/+vOxMAG8Q5rdbxiwaUB9A7lPjJIg72qw5iR8AzZfaquhmuq1XWFFPEJ4Xl9aE5KA
SJyF8z/TEy5e1q2GGdND/S/Ih2GWsidYWwSmLoH8ibJAp3Hxqb+rP5gUzXjgwfYaCQh8rKe8w+E8
18b2eyeRdx5+FH2CEDmodk+EcxVVSdqVzEqif6HByQ8FBktmfBckVB46nPmnThZP50y6CbPono9d
95RGsrgMgCYwVkYAhLNcrQQqNUloFyy+MIzKt0ye0hCGLjDqgtolHT6Z6BsDaMRWlUdgVeJO8e34
N4DaEso4vcPsAhblXOj+SBVcWSMZKMwxjpbBiuNKsnMxK4Ydu8QWONneFGaFfGfmHTISnPxYA0je
BppjVH2ZeZfHmm6rpu5fKJKXIwCu9wOtu6DSVdJsEw70gCOUXv0JMaoyECMILON1sr0AWnuDHZCt
UbAX+Hva/vwaq1HDrKUcgRWCSRRpj3BmrwwpMOTO2UlwS7m9LbV22IA1zseJhakdrW2Xi9CegbYf
JzvJY+/LQ37qusANJNXlhwawma1ZWpfXd/dAQ5M3ViG8bK8E8lFMiBzNk8QszQn1Y+sfU3yIvp/j
Z5Cjyre8nJL0wDUei+/o2BRMtdU61RcdFXSiJunmTJvjq+655uwMILSzFY0n+/kmCDjOxous7i1f
NYbUQwjijc5PLbZwyOxf1maur0J71JDZ+V7zUXB7I1yBkD6yeA9G6N/W27z/IgtOUWOAN7JUeXMN
YmcuvgtkTHUcVfCdXXWZ/cPKU2nEgT9afK1LhNGw30JLNcmCB8WDPp7DuEtLcES0J7Tj/6nrx0Kx
A6O+ZpNa/hTmp38l+2/J9kxruf+z3w2rF/TzzrmqTBtvqpuWkKESEx1oIwMjm/tyXIYZXGqvkLVD
OifJySkrrkFoz4dpm1hVdV5QHH1BZ7JyBQ8usgRdQ8cl+uTOWIi34VUJw8fKkYhvfdVlG3e0/VMO
FjhRHlBnhW8VxkGPV+wfvq6/gmcBrE8fK0uh/qf++nNzrEVH/Lp+f636z8akiH0pZUayfI+1orOJ
EtwiCGqTml9dWsGGcXSydEjABp8R27pP6MkKR8brPdjHA5nlrAGcW3p96XidVdh+Ay73VdvQyINV
uED5TeSJ40bL8BV6C9KJkoWgiIsJGZURtplJXYacp27pe2gH+0K2XLOEB5D0BgrSxZizbDPFdNkU
0398jGM9pdcKNo38SsLRgF16KKp8yPRwGWdjHgs19jtGgqkmynQl9wRpJUvSjDsjUuM8TCBA3zLi
mIox2R4CxjaA1HlfxUC8GtxU0gCXcbv2IUXrTIKPqRXxQs26thsTQSODyEtfJ52KxNoa0ayDpxFp
lXbfdC/MIQRiTwc2tX04nzxyX5SZLhi+oJBJj33X4X5+8RiCd1jTSqyHWDLzLJo+JgH+bF598c6R
sVowv1OJYJLrR34Kh3/KgyMeNOTh0ElOFaLHC/91+9USZUn0bz/FFoVrZY0UaDKfA8pNGaven777
lKRIdXoZTEq4B+Hf7/ubj+VbY1yXRf70iQWge4kcEhuRNskmR6BFj0pPXyAXOiKLovvoN6COquQ/
ZRI3xEm7HMsAwwu/Octm7OqywRADZY847NBkXmK8eS/o2kWc8JxswiLwG9Mftti/9Xb9bHvG+R12
66SVmJWxadiPLygQwHdXs/fT3TGewjmUz4xtn9VfiHyIxvhCwe3JXP87q9czL5sltr8dxwNEQMfA
L1tGGQKziAaaDd7xcc2b2psq8zNXh7awniUY09DhByK5+L95tWB1C+J9v8yM+4S/RzlI6m011jQG
7TjJmnqlW08t9IjDDXZgfm6X0S4k/YO5NeBthecgMS4wr++fwvFx0zTLgHTJIcsS9EBubD5hKTm1
kYW+oCXSWP7zqYXX7o+8+at80d663blT9LiJFHZrdD/RWXg1Yl8ymC2KSaXNeUfqbOrKuIuglNhd
3b9WzMwwb2hAqg5mc4dOZHuiHrcb9RiF45lWXsqmjGsH1VmWyIu/Gk6F4eqB05BEM43rOI4F3enq
/Hh690Nx3civ1/JFn0eoqbctqatZi/L9yV4OSbQIvhpFtqA3HEYMiG0UzHu0obafDgJxoODBTxYo
ohef1AhFdxdUkvp26qM6q7uwYd3jR2NzMWfN1R3mCIMZy1bkWlbXa/RxzgiKRwbhcufMRlBDy6TW
H2/bp4ZvalnDBYS/MfBboj35YgUn4xhqSrjLeVWVDa54PE0i7/4+43tbWdUFoZzBr6Ne0D/jhBZ2
7/rKPjfnG5OjfZ3N3k0dgylt+CNj5O6mpAWu+/YXLE9LqVFFzO0XRvAXZfcSEJatE1RGrdQxs4S8
ghVCVFXfMOBz271MIbTwiX/tr9AG7jF3L0UqTbH2EmpZ9IVpCq1g7tKFHdSTTdi1eFzugQ6O65rF
IcsiacZLc/jbxOclMNpyTwU9E2Btcd9NQwdOf+e9RX7GTuqb1t6+OL+06cpdiYGPTulqH/9ozQ0x
0Gt5HKXAvk2c18nk793rUwc1VzGXXc4MgeE4aclpyreD0bXbexgoDjvJnef8rdw451sYB8QttbKs
sy3m9wiaQzzjtLaFCKnnAxfDVvoogmODIfAhtVDxMbu/v0r5AsLvbKVcKie4xlQgCNfjC+kMHRhh
quI6U0RptsIgUwTGhemi6ite09JNUbMyD1u2RHmL0R62zwYF8A/VcRAXS5f2PckEoaaKT2uuovM4
fZmP20ZQw/JEF0tzvz2pJbEMx0cb6TipIbn6ypqVmoTHU10ZgWmRaMGLvoTt744aPefH/1JylJbo
oMqQ8x1S6XBABzaIFrSSq62RdKS8DAvhGWATb9p2oGpq4zpPRXLRGS+/p0MrZRuGYGHR41TAU4fW
RFu/3t0RoW+22vGMD2aOfB6qwYUpYiL0LYtCPOSPhW4hyoYHII3Tcgm+yXkPF6mDZkb2ztOwU39P
lLrK0v0Vbv9gGt6EqOZ3VvMgHC5jdSOEpoOpH0dLfuzVwmqLlJCOJWRi70xFV9PpIsoCGKJII5rB
k7oLty0Qmtt9m4oOUNtwZWfYgp+Z5U/x1r14PYdOf8/46PeDosSWy/dh6NA3Irx88u3ujXoaMgva
j0Dunv5RP+y/6toBXdQpfhqYYmoubBm1ze6O8eSXtPpYAfRHOLrkIxIg2pEZi+wAo+3fhhNDKWB3
xaGTjIfQN+0XDZQH0l1GhSMnbTCBZ9hisYFdlMm19vbbrtEvJMcbflIEwceXdqYmacUlL7ALVarZ
+KCadOp2Y3SJppcRrqkgVrwvFRQDNUhwNcNcpB1h4F7TGo5pN14QkLYFNyiR+XDKV/A6/3fut0CZ
j79enTy/gC416KXBhaeWZoU4kjVdG6/QAbyg5aTrvV17VZ+Wn1jIDhNjNk0LH0JEZEGmjBtmlRow
vCbRTWTdIXeGZj6AaNHXoXFL2hqyWnqZj795yiqZTrl1RYbm9RnGTiA3qybSz42tb59DwLsrzoUX
Vcw5eHUiU8WGovGrXF8ln5uSbuDxY/ifFO89kYKP5oOghmb3rOd2WHCRl1LBqMcbPqLSyEcSIj5r
JWeuyk5lbLJCm0NIuxkQQXZsQhw6p3oXQ109UA8HjlLcOWvgSZ4oG4NQZpO71f3Cz7HwqOujNwL+
ZKZgntJ0XsSADdEVvP4J4LpadJUXeZC5swQaeOhFvC5lDZN27by07BuimM0GMxPsezKlGzAP1EeR
iPL2e/ovXS9CDL423yS/K3sme2Tfmqc+PLvmhg1dqU+a461eWy16XtdFcCZb6dBaIsZFnAgYyYVA
AvlylhkX7lWdlVJNwWbxU2kYSgZ4fFjMYlre25wM66KFqdG0D25p8d3RAktAGBrRmmXWW1I3vyaP
6EjPZlUW6/s22+AQg29oKCx/qm4wftPQUOXn2nJHMjFrsl+ONP3ZGLDlWPxkQC6Iz0IYFPESAZyS
Fri3wISauFZtGHRrGfx69/JnijIrLg8ZkGQ5OkNeLZ2guFXq4qMNX4SIkUzoU/a5LPqqM+KmMG28
BXZ/bcVCuwDm65MQLplvlMcMtkkYcRv6yG+R+sYCUoS9RRjJmixTPeCQshG7XrqWnK1QqSlUB7jl
z0CfIatFYbysHhzEXzg5qXqz8R5AtQcIb42ZVki/FMou3BHIQOumEJdIp2w8P9w4/wJi+CU2OGzR
kXXZvxPvGaesXyvcergBJusYD7+bL4CGHMGRpv+jOr3da7ygyvRYhNaB/1GP66afAIdm4gGA63vK
povzxQrDZuA+t68bNOBXdGoJ6B6RAfbGHKC+yrVVQCn5V+I1ixCgUU/sfPAlq0Uvxbk80Ecifmxr
hNlmo8urzYNdbJtePWLRM1MSrWOejLxB0tdKboCHZ/Wa9v2vassAZAPF00b2zBFrtmJLcGkPwIhq
+aGc0o960jsTxCfBildKEPY/zEab5Z2UFck/p2otbsSfrmKI2+8GI6Cwn8SqvYwXsKz2glE9xvTz
RN9AqlxQZbR20cdYiEslkIdgH1ACJwrCRwi3aBXhK3HyF5gneikFeDFbty2X87nSCq7W8FXjtrZ2
kKEQJelL04+Be6wFkY3VhPg491wiqBdgRW3UCw1hWfSfaw+LZFvWAZDACqrFFCFkek6Vh+r9P+z3
KNx82leFJ9S9vbWZUtHZ2MMGyfTDmeubooolgxJ/f1TX4nb9h3mdMPG6PQ3m4NqgkLaif5iYFg/H
TgjLsQapwgZoIqGyKLOFc/UcXEYvNiBVtEviIqVgHIPawfkMxHC9mj2E8+n2dbM1dx9hBnDkiNa+
6Lpd0ixC1wImfOBAYKRRIyY8bTM9HU6si4rRcY1jxFEekJwx62vH4RoCnbeZx14CRz+c4ZGfbGeE
cIEYlsxx22pKXNvIJYcGxX31jhVhqp2/7lrgEemHm8ZtQronkuHSsvJVDsrpmF+AKCSAGxUZiSM5
1KTHJ7viYoMD/8Uh2ggqkkRAPnqjyxYbAU9OvaRi8jCA5AfXwFEL2IQP2dgtoy456n9+GAglwyeq
bZmt+WX4Yd2NRWSMOdf1PPqQ10cGSwYdiGFgSt4EE4TKRjmcAMw1dfnyhMudfs8f/AK6Xt3iIpVd
2eiNy9A/4b0X8tOeslz1M/qXkPm3GPvFSe9l0nJ8SBxjZmag3fe0BNWc2MoYRTPJ+RvI04U52Q6n
8t4cFieXAV52XPk/bRjUCDNNCMz/CxpioXUXAetVecgbR+HsN3VGwoxvSPzlqTyFkOq/rQityKgm
W14jadMy5jSkM/cuHBfubycMMT+XNRQ3/yDOLc6WEPOhc9H+8izS2wRlW2gntC0qjZCpgbLH4MYk
wkllWaRqEnYPoimvrlp+BdJrslOpJZ4Vi88d83Th5rgCb+Sd4dKchAYsaLedxaMD4GbmsYY2pPqh
mIRrfYcLZ7SujB5uW/SZwyCqNX48t8DUcnjkYRVz9OieYepyQArT7atRRUlrpyyjUrBqftIhH5PS
OWyw8l+ovHrRQdiXZWHzP54ZaQRa2jbBq8r/ncHfnagQrp3Xxqj6xTLbvWq0vxESB3GeVZRkbcrV
4tCeC223G3NvZxCsLgPF2zjEcbobBBIf3UlkOWg4ZIVLE1MbtNw/kKoj2mrXeLxX6a6a8kKl+In0
M+T0QtiHfQTIbkjUUpuyTpGGnSxbkL4qT8tF9/KLY7TUNHjjcJ1lRhpQ9T75IS1taKujtDEPGcGj
uMc1N2eWNE1si1lBimRQo8CvjB+wN0iOdx7NMVfyfXCtwyWTeOhAL7dgg4HtIbtFw/WLu+ytUWFe
mgNmOhkQT8dtb25De6/5L8gWfG8y3Z+dg/W/+rG9FDznVgOEMg6raLhUqf11yjnkIV4xq46mTF7R
VlDpIRyIWXrDszABbl0zOre2T7f3vreBRRhkbaHGXHb8dIdBvFetjHCGhXOT5qFIginC0dUSk59i
4hgxrO53fA2zn9tjKZSB2ZTHHRogSXeUgenGw+LWZcyrPUdzxaWS1dd7S2CqiZyojIaSLRoCYQOx
UpU8MgjHUZjGQnzona/y06RXtCFOBI8G1Q8lJZH7wqP2zp4AwavGT2Sulya55tEyHDB+QUcJs4Su
TyaA14Hvduzu+ctLedhdrxGWjQl0EL8yh0MsD1tcHmdirdtrrTzqAmmgD1qi1fu7R+N+6tFK+CJC
kM4Gv9SZJfHkW9D2tfSXOMMxivotfSH5Rc6hURQWNI6ET9gk7/2yMd9um0QVSsY5odN5bJ3wj3Rg
mrtn5Y6683oMoDHXA4+W2BmG2C2BVY+fgKra8ogSR4rBxV/tgEp+7FzTVCQfGB59GSF/FvxR33ez
IJYYoxWYdefzykOsvJWTuAz6pwClZikEV6EF1KiQLRk8TCHchJ8ljX+SZPSU8pG2rR6lpovmtRyp
6HNUsD5XmiF9VJp5ruOf4SqORc5aIDXiBJ/J0V3qVn8KBZKbGEzlbh34S7eg79GEq5p4+w+uSqyK
vr+Kq6vlzkhSTEBM/vYkCjD/a34GWuys9ed0nNl8fQyNotxK2Kk7iEBnR0/SDIWkR5AepINx6R02
k9Kj4K10IUJCQbZcG/o5DSNcoiD2h3qgJ4BDgA5NkCovHJh+AJibh2lqrVIQ702H4l4IZztiyUhh
iWu0pQ8leBP0eTOUiTMLcW4ZaUTrqofiH4uHPDNJE+uoZnskiscqpw3k6Lgf+uMCzKpOb6FHGL6T
DBSe5L9CfP39cvS0KjgxWrjsR5/zmTppTn0NwG4SDkTNgPwF7+mRBYoEPNUTvdYpBZJILFi3ZCg7
/lGSQPpWRG8XRk6vwDIR/IfUPXpWI8bFPr3EvJ1lOdToo0eAfYjjosz/Clor/vQTKKUlPWZY/DIU
YISD9fnDpacnpDYGuzHGFOYvyh9pBpl1GrXCsIPoeKgJ7ZDdHjdwob425+aT92Ny/R9pAjmmtGBb
fObmsgVRYImRsUAFXZPxt4FYJvbUDg7GpCh1mu1yExAyG5/yVlevk1OzJrGYUGWVshb0VErFL0vI
gJN+BvhdW/mifCwDlmTgnXtM1jcOz1bp/ksrl27/23d88rJcp3/Atwfx7FDSM5scEErSJqTEtUup
LprzR6/Ui4+F28g0SVRW5tJQ/SOmj2wTuV2vhvTs1+NEeKgTdOz14KNd1DR8TkNE+2apcPU5bxEi
AkWfeIayGIaMw9iX2v1t2paIEaBSqzr2z2cRMlT1kd8ZzP6KzXEvumCIbEWm64kRtIT8H1NJGI3B
t6YQeff+TQfdLSggTVnjq2fmVHGre69wANxkTR67y7LWNYYRErENZoxBpyYDF12hCUqsZWPmGdzD
a2j2ep0WXgevYaDyn+Ha/QFe/xgiHj0CjJUzlGTA7UilAZ6yTh4H9JxkGTocu6hlP5b5Bp3RYlKh
Poi+FoABr9Fo0dI3jYl7gnLH/7H1gGPRcjnEJDSTt1wMFSwonKFx729+MDhy7zTPgqCcRjr7x1EE
24SGNK1f+74DXm94o1nluIKjWS6CymniuWNt9VbCrOpmFIXQbdjC2KrBWhAXc1u8n2e9HST8l63P
/vcUpc5M6/oglhy0FCGEYy6TS5tVXf2AuyLoP6X0h6WJIV2ndExUqjSg6zKyXuGgiALHKvuqr+A4
WxaBW1m2Thl14DA6QExFSGE4G2VcyC5c3KWTFjUWYVfrSLGQJEg52foQGlOcgVrai0InG8cmk20Y
syyzm46Tmr1Y+qLUYhvS8JKRyQQ8JrvyivVXUTMeFt9QhsgLuOqd1f0uIJFwzXWwnxKgmVC3BzSZ
rVJW3bBybyA+8sPhtB4b7Uo+J1GdWfmmFucGRWZ/+SbKfkhq80wYKl3uRJo68NB4C77l9dbPnkoD
3q5ZWwBKRM0fmFPoRvB3tnu0nNTfUVhrDIwL5x56dVbbwSB8JIu2mpAWSdTbzYT0AIlITD9eLCCP
9p88PqoIJ+7gZcX/7wu+vkdHC+Yzp1dHEzxcOjr9mltcVdE8CnjWlQ9vM872F5ndI2V7qliGBTTX
IwcHHaVLW10t2RttzeK01ZwqW8GinV958fu5JKcHJWDpuP4NJrsRhWi/hf6ZB0GQirjgw/0k3WgD
k4IWw3tnhZamy+FGTZv5o1gAe8h2l1+6BQODDHj0eBy75myZadr11Cs8mZI03DVSEgI1YZVh4kDU
pXo12tnGc8sy5YSXxSr/0vD0lPX9KcqyMmVHXoaY2jnlYpTAx8eIO3GcctpT0B7KNYLTzVXKDX/h
547qOS33WekQXTAn7W1+5zbScvnkNHzRd7bgk+W3m2Ipmmo8mhyBYk/0jTeRuw3a1MnyNXaLL9XK
j3g6Wm4lvf+7uUuGqOv9of8hkIHl/0yDe/p1YR1w+xGnr4DjjwraZgAAsE5leGGbq+jgq7tnsAkj
8WkKfonQaQz5sKplcsm498FGKpZ6aCj9ZMuYCCrQ7SmVWz3pjs0zdLS8dpURvzbsfI5OXriyDG1h
zPnMSeWY9BDU896076OXNOJ2VBzcPZTb0BlEIzHWHw6BsYO7oyJKsz1Jnh8/1c8G6xEREQrQNNHP
bd4HW/ciy56ZJ2KC9OLu8xC9KM2YjIrjpiZn1tf8EFHWrirryfjfpUA+LBUGnh1gZYjr+0cvItC9
UaUh7Vs0h2eVg5FHC2ovEbTQlQ5/Do0bQfaqucllOzSPDAzQTJml9cw4ED+0A1I0uVKSg05CHPIw
D7svU5KIH8ijkrPtk7rVMlcnx9LvpJf3nipLFYKkbWFaSu7zIyKc0RFy6xK+aODn1NE5gi7eBCtU
Ryh3pmziktFU6ooyPsHS5WuE04sKd8UYxvWGNg2JlhAyjO2ArnxOL0WKNI2QIXVXkvFslS1msd4f
JUYradHg6B3uT9gicmH0dyTUHBxvvRGhopVFx7lAuSRB9kHKoHNzUeKJem01RE3Im1m7agvqWUI0
RQzkCkHCD416ZGQT03CStUbaqZz7pVGS92Y0Zx9pv2RW25YNurTz7JIsb8zfyPwUCewIJbSBIjem
kEIyxWYnnif3I28ulJtkymIeNLH0BzJOMAs89bYbdRbEOWzEd4CPqpdl9cQanfhBYynr4WkOacM6
icPCp9It1y2qmlS0S3P5Zt++gLvkUwSgdZ04/i2bUIotDwbXuiqn6SfKQcP9OD7ZOoS9ZbaMKWCe
ae8tSx1M+vMh5sLdSjV0rQ6Ie013jj3ihuiy15uLAhEbHNzLB8eOYSGEpBiEhckfql4CvAjX4tVj
BWU0yVn/7A2bEBJw9K8GddoYAIinX8PGYTCGmsJQ5x/+i6aGw7J28Zi3BkHefbT12Ujji4bjKgOl
p5YnZ55hCa0H49TX+NeXJln9xMWk8DFrSRhApi9ugW8MQ4pXCTDv9DoGijz49sxXWggD+La1Nkot
bRb/SsOUlqjCrb5iT8UqQ6MVtuJlQGiDH3sv0CokOhzUHplM7z/BwxvPBZru8VHSzaEWfAhb6xro
2uYBsQPiglb2aXr+mxtr59Ey3rJyx3yk8i/l8E7mUt2JSn2TZXozBNFG1wiNIdS4rPNTwZ0aFd+P
nMXPXJ67AqFSuXcXqm/opHggFXz7JBlTIj9TbumG6BbutSy4A8LXFIHwIzI3uTwFgyPpqFHCgqul
AQLIYxLSCSl/f1xULK1Q1zWTfCSA32CY6UeJf57dUs1MmC/pz9BLQwNuT5LbY2ZJWFXXrP/Ib8eN
N9rg0LyNt50SINhrG3yGiGDYh71RPgfb02Bk2aoYRMaPfA1U5cd2O8pvUzPb+BWnyGs+U8Glaclw
sNRnAssxthl3kJFCDejgXuiYS78leorbyUIx/gxtkQlH2pyNwVW8Q+tSOmaXfTzu378R8fk2w6w6
FOIh3oQlgDZ2GM9MRnEPpVoeep9btjIswFg/AFm1QHp2JchxrQSxXgNiYOW1a+WY6KVxygwE0e2e
ALJ5Es7MEQIcHT4liWrb5vYbu0XsX6bhZh6/acRbJTBGOLxMaqngCI9NlLxL5urZyqEKD9vqE+g5
sJk7QVUuglya7BgAIruz5SDrwctT4LWU8Iwm1E23a4NP8kUbxwT3Dp8o4YujPxwLCkykzwgPzhIV
pV3A7vyLrHIURFUzDHbCwRElUXNHoq3DQIwR3MhJjbCuThTKXJDjk2hCCvUwLNysMLBhlYhls9Re
jKKJxZdte5nKGFIwJEFzw5kA8QsbER7WmA6VfwcSZ2+R3wxULPVH6+m8Az3jEgnaiobhrzsIMoAB
ZSp/z5+YrOlFjpjE5ZTqf1n2THecbKM+dl6NWvXLRqI79Zrta9VC7sPDzVDiBUizQ/xbg3iCAtbT
8Temo6usMRooW/+jD9iIh5ZGakHeL3MWKY59OP7aIqWrKmdC4N23+8jeMaGeaekThWeyhmOK8QlZ
vUw1w29B2Uut7tGWk/TFearqWBRaVMexagZ0oZBrI29ubHbEg9hrj/FvysfgKQXGtui4V1oO2Kog
/ubmAsC3L00IzoPW7X751LqZ2KM6bHxSoA5fZtGc14JiBEcQF9Np4fGwCmOHgc5/GVyZT//wD475
/i407tv1jx8KWgjljroXOljLuHkMlmYjNT/l36bZUwt9QQzjtW0SvULV+rBkA7IAs2+LlwFjU0QJ
Io6X64wJLeYACaktNdkYVTAxKcpr2XIT26eBkysM3EHcm7GJMm2SetEdm06HywQ/BDWdiito7ich
V8k2kOVqwH9b9ITrWuUrU6X5dhhVrB+b7LxNUecE12XO+ceMw5G4E+DZkSLPhjSde1Sff6+YzFKC
eSEsmjCqSfpoXfGrSDlpqsybZzleQ181fS9jcB1u/C+MDWOZjNuJlWHbb04XWsXaeKzjCRqkZQhu
A7GxeLrike9dDzJGkOVrhHQ5vruy/5DBtx1/uB91dU33CbXpGuKqgLTA+iKLa65pG88W3ghgpXx2
CuE7e3tizRQymQ85ygXZjwyM7r5bmvE/rUe94YcpCgOjkqNlr6M1phuhuqEdzRZbElXFnEEusFe4
x0eTexqGRACdmypVX8BIp0I/rry3LvzH5DECffi1DB8zNLdgOYhQRyKEdlfnDJMiwqV2PMM3dA0u
9vGaZkOKAQ68hRihT/rbPs5SDx0GhYUB9YpaP8Kh794hI5vPNNAVvPVuki+fsRM+8OSqINI0VdDN
Z6GTeRhTtnc98p7ZTv9N8n6tIHFrrvmhV7McQnr6/M+8G5gS8fa/+DS2mhE7bDCSG5oWHB/w5smP
kj43EFkwdBAejFyiPxVvo7Rh4snjnjWJ9DdrWuxhvoempPXULJTVuEQIT5TJdSG5dhJu8WunCW40
rtKbHjEtJcAkko+yAcLook07qT9xIV3FFUmXOz4061+0/T4MLsiftZgGS1NBm8OuvJl7HxwChKmo
lcpP1oi3QKA4XC45B9Qramd5WWbBld/IQ1wLZ8hVe9TPpC1+SthtnZTAgIE8XSbKd/IbyALPQs0U
ClIXAtUn/VZwUOW6d/qSDqY+lvmD3Y+um5Iim/ZCM/XVjG7Zf1V3iXDcliDQs1RI34xMbIsM6x1q
TvL2K3KdEV2uaaa91wbBiw3Yrmoo/ck7ZCB8NU82AP2ehoZvwGa0F+7uXsifPRc3HZI+x2Cmuwc4
c/+R+w4BOtUFylBmMd6QC+I51n/jne9F22swwnwVKR8iw26vJoZrSr+AQbejVXxMF0M1gfisGk97
cSNiAP8LadvpOkNGahymsEm087izx4JjTeCXHZ09/irKFy5fHAw9HxVIC4joZy3bkyU+WVmi+9lj
hy3Bv1/Xq3FKdzW9eEHNM7dSZd7jKLZHMRIWpuVAk51OOe0oRzt+S3cAEf+6o5X+ax4OPjXGU7mn
kRMgvmsQ8DcxLRlZEA3K/U4utp9TVW3IlDjbDsFa4P4Mb2qD+VC94NSGRAo2HeY6FL0Ll/G6dSJ+
icm6wVe5Dta3XwIMGnxsnASlSW6HA51/GGY0tsKTTDD/Y3U4K2AVqSYyBwzbw6mcwXUgcuGry1ZK
/EbFzktAeD7eKky8LALpcyLHYvhNEm9jMYEUMgZq4CqCrbqhWrJlE4DQcNlOIHFbaQBSgi3JU/Bs
82wk8lD8Ow5zXZ0w21AWtteK6idkYQDcnE6fsUGzrMx4BGCm5MqeNq0/7ThzJrXDF3Xe2hm1u2WX
FqnmapBg67RWInxjKA65NWDEER0/lmrL9LG5ypPcEtz9nRnZy1qzlEUnAKAfnF0vmw60fjWUMWmF
o73JAkt2Hi5GW0B9cCpOTgxi6bKdeKz3FJqLDoKvDmc8iQrEKtZZLUZh3kTkCoeIq90TFDyO6V+h
ngOyXnATXciAzBmeF+ofVjIa14HRL5SuVSu1uizk92LlOKAF3wn07Vzcda8esvOeY0nY6XUynjOL
W35cLypdve/fF7wYybV/q0TC2dg1+eHHalynM2T20R/m7zobh9dn2ux7eMJM+ZaMl6SSLXRfnYjk
nm/chVdx3e80cEJ06u31VXnqlZdHqWhf+Yvzw2FDWfF9V0PlqujzcrljGO9C4jY8fTW3/1fnwKCQ
PmDIzvYZALwe3HECyLcO+lWqL0ImIXwv6+YiGjT28Tp8mmdVYe5U6pfprC0oTiM6MtYQBDSLkxXB
BmwfLIFTStnEH1cPVjui+VhmSlFHO/ud+ZTLwYjjDVJSzCv/sLkYb/RjhD9LSkBFccCLCvAGRHJS
xQ66SeTxhjBUeMURncRMXdImlmkMZuIs97tYfJQlHAXlmAq6azKh7oqIVQbDwruYNWjogUonXOKx
Xv9ha2TVLYf6spyDbLRK14IFXcPspMmb6CQU2UuGVRE9kOK7wWP9TIdGOXCDsf/rtEnQFBScImGC
qUJa+dBUFKQQzH/GhUK2QkLmJTnq8P06uLmo/rkXCdqCq83mDQdAkb8YPiC3lrcSM/3pk20fEpyQ
pvHpGIbCbg6wl03I0Rgc4I2FxqetHeevuEQ6J8YnQeTNk2vCPKfMDiQku1o1C1R6Dw4Aa7xlnqZW
uPI+IwyvXkumpsW04ioWtv/ntZmEN3B+eK95L+Mfd4hrYj50d0N35XuNdELGxjqb0ssOvfDE5H/r
A1R4NclyOjGALjyc+ahfv6ecTkvfhERfU0ORLQ8vl0CJY9S9NlZnUr9qJbgthVSFLPUj/BkkVYRN
p2vzXTAYbqkHA8KIhxymH8CsXgpZZHV9auEHMfLz+OVbSaO0GtmWFikeMMddRn9u7tKP11RT/NtG
tWNJiMyUJkXL8McsjOdeymGY37viXtAMWj3Eagc4DBVjFc488I/NU5fsOiuORGvnM4co09z8Kw55
nGVexDXSQ3cbS0FiPZAFl3WEVUClhN/E//IB9B6T2Bs1iMtA5shPc73UW2uqm9aIbom6Pw5Fhv5v
xd1lkGf40Zi19p6ZHqi32YV151HTxcdexc7TJLFZUnc4sQA+DvfQApO8RgHb4h4DMA/3qCebKjv0
Bgr0mzbUjrRnjCt9FDoz7zESXxQvjZdKRr6rZGD+ePbxuj74PCcppvH1LeOrxXFLEecFsgeq2jRz
VdmEPzEonY7Paz9BYajMCnYNgOoLR1g1iTyzpTNog14NCpRw27pZVMQUbYeItJISHgYon+4UzbWI
3YiqEUqtCxyQMuBzCRglkLJtgfKmlacaKK4j9Hst11/96uKOH6BqYZDvzisbVo7A/pJtyPTXsWek
R1Rb4E05tRK7KHvr23WIIXR3VacN+AYFmSusmPqds4G16dBHJQ4xSIegAC85JzWwS2I3ngqbJMM7
520RCPcrZUeOSA03k4b4okeckoQ0cf1GdO8tdMKvQPTG7OIEE1iklom/fNpQL0pQvFOmhlBQ6oDL
mHJ0S6NscB2PVnlhQwOhKhrqlvRsbf5hsUJXHVFhbO8K9gwoOZtQtM87MJ1j0CeHsDRML8NQPv+1
MdugCdX1T5sEbrcF/YrEL1yADppztz9XDIpR9laJ1jeZIw1hp9PNnWRlPyYQWlKgctrTe3+1WZ54
hoWZQ6MeK+r6mjXK3wv2RflldV/6i13X+yATjnVA5WKbbd2HG8vpOD56/kN1gN4byFDX81RqVyJn
M+RzzsoQQVHPzkHuu1nMLWNwjVxt93sfbUGzsu/JaN9Te1K6hTHFKjJA11EVv9oNIeG274Fjz521
+ZniSuyW0OPYtP7ZZFStxHFCWXZd2ZdiZAHfLFjmtHSLz7idkuJDCyPEnjY9JVciO+llejpRVEUs
3eOUkbYC0NZulT2Z7QS4wqCVsdks3cW+PZDUGN8A5i3cn+wvkvON8K1o33drzmeGZ21+aca3CywC
nO8elJwpNQlp2kZ18/r5uEbHMc4EbyDhIicgWRrbxZ6h5q/LH1pu5kOq28ZHhYCG42GSphbHeQB6
nR9T+60HlIwvSjw8wmL84j3zePZFQB0w4lXOolhZMUbqUprk9KHHz5YVagcTHvf17oD2bhZ292+3
cpjskjQslAlBGZE8+BWSRrvGupTzxJOWv13chyIRQBF/3w3AuWfdMzjR5rKI8N1Q8J4xsAmSyCVC
VlNJFLhI/X6QVJgVVE1ngWC8Wkoszjk1GB0faINuMZ6X/sNgs5tOWE2CjI9jkebps8AAw+Rq/GMH
r+Tx7Zuq10+eOA1Z4ecmBTFiqncQCQkLLqAZsNmiE9oHlv0yYcGAGnrNZLMYOVmpoOD0t4+JRXJH
ONqpsHxOxALjlHQ42s9RlhzWEt24bbMtft6AsHdHKxWtBb1DuJ3j5/N0URdBQrLE72o0e9A8jzrs
eS/pXev3g8uubRraFVSsOKwq110N0dpluxGXNhYpEm/4dm7MRzeioC/0fngi/4CEIZf4uAaxlP7M
LZMa+ZJOlFoSuXk6/pn6MFoFgPJYLr2Iz8UluBEmZrGFWfjaMlDNMuvs1IIr5KBHhVPtminF+/ln
h2+E42ZeHI75HC9Z8gbNNLlwirAgt0bgAAI1q4xfHysAu/Nz06oUn4YGbj/NQnFCPA1v1dPiALOg
TuYSMTLkeiAHe0+G+MQcubTgcYSCXghs0gqL8EIH0yqLDKb+7fqvkmgu4/asL6DtY6R+LrZRBorw
6Pq7mGdjCwYEgm2FbuuymvPlffTTUuD0inl3KSL+cI0OJzI4sFSWumyAe7m3sIXIalItgNXq+Y7L
boHe6XhWaD2p5lmMd5kTqNIUxUE21coVPSsiYyA42hhAUJ0o8VIOhiU5Qt+9xGNiy/Ka5QneeWRo
WtfrizYFd6wXz57SY3ZEIaLdC2SS/w2fl2Imv/V0hpA2kBOy1AVmwTR5oiDteAIzw1Ud2pq2/iAp
ZiTyB06zexjnZ/7AsXrMATDaaB0AZk7ruqjAL1cpa4cp4zpw2g6y5RQW3PGKSCzx/p6B/eKTsfgK
oZgbb5kfoy4paiCNo/Bbg5wQy7G0AkiBCJzlmAgXxnkFjVpPlDoRdyTFpQ+DbSXKHQCET8jZlzop
mQ6147A096ey346vU0bdpzzV/2eW6Mdl83r96UltTFFsE9Jkf56NljgQvZ3gcAoWhBK5ol11pv06
J0AcVCqz4aSjXkPuJyYqRfEHsTpjOMjvLTlWfiJvLi7OprCiE6b+EuPSoI0kZ/JL9Uz1MvXEAujG
2C5BA1fOyxeax81vDKZlTjpJ56S+KkATetJps0R+LnvvNMTW/3SS1VKjov5/rW2aAohhoPGN8btR
tZTXwVtjkXbxINn9pFafzlDrk7LNPZ6Ip2fVpoE6tHYnlL9rpn8bOGBSEIEIj5jju60XfrZe4kmv
WyzLn4RVC9vGnpHe7qwGij7YeK7jzjeV9X50xhkYvKPSxKCXaacLkPVIrdYrsuj8QemYuFshA02S
RsWgWR1fijOxyGeYWKBWBdnXl5LORah8Tpla/7tkci8fGv3Myf7nYdVsCPYyBiCvqAosm8Ol7i8R
Ax7aQ+aENc2V8Gbx8XESgoJXz2/YBm/O83FxznHJG5M+K87CI1UOODZQphoaVXteXe19HUt0QApD
nXRIRy92IMDw7FrnbOM4cP3IaDsj1wVeST2MK3jDI1nNRgO8T9WISgQE8if7nWg2aFDHA0LIxypQ
Ic3AHz7JlSA6pBnTldeQZ+s6HTuGXteFm8jw2A9WuLlAePqtMijEfQcUxnnfNZRPobCwdyd+5j9s
pkwpBDIY7Z5SYn7bOVgRbguBTLXfgzRXM2z50VjZRZW6mDzFXL33YoTquQ4AnmzA1wJmLoCkEMfF
nkYDwqzRZwh5trOqzAebKtcG/2Z9yW6trE/yYejwemHLTj1LKtRxAMNoibL6/rNLA6Xq+a+PmEB8
l6AQc/Gsl3o/IbjV+PIG22sO+fPnl0QHR1v+JHYx8XEi1T+zvYGcU3xf/jKfyYlX/9EOAFdcx+eC
fFSez7H3H1b4kPZl8p/HQv4gsAva7X0EQy3slZclbRGFjDaf24mZ2m/UzxF9WuB9UyJSWBljFJi3
Bk+tCBNRy4HMCSduF/ttyCcPAGZ8XmPokUPrAvcBaFYId8F/7t4botdExsS8UUWURsHnv4sJuYcR
6lIdtEfjmLS7KK122r3uX/1/X/K6KOcj7wDd+GJLp+nl0tFOjRm5I97E9z/Hk+9xeIurhpw4Q1Xl
xYLSDIRXVuCDTTNPQBJf4nTs3RpgysI28M4Ggg+3zHm1wRoifJFm2TDpRLCfFK66Y7nbLXiv9s/1
6Ul+lZhKerZMyhM5iJ+baWf3n8j0TJ5YB5gC05aaQ443wBvpRuXnFDz5QDZWG7ugxHP8eL8EXBLa
eErmn10JGVBrRIk5SYp8A/a4LI7tIVldxCAR9DNnrkQ2wL8MEZjm/8ooL8O1Z+l2gGWXEabhHlUA
tK7I+GRf0CiYivB2B5le586qPVn7wNeGcJq005BGMtd7OoWB39tVPWTUMJP8/3GkGgA9w21VF3Ha
KwLY4AdyLcqFKfn8cjudzeoML/q+96venLCRiQYO0yofZIx1HK0oqwZj3mF2oXWytthVZrmVBhb8
rskRI4ZKD+dyr1HBfANIFkWaIjfRgxO6OjAZ9k2JqctsEX0RNo8tFUT2cIzBPK+w1HJX5wmBYO1n
qQ9EWU2oCubTCdyUu3p8+j7JjL36rabgZelqk1iMAt/H53NobfCgL8qsduAKn0yu666TBeGua+EA
tvfVTNvNeKQXmAbcbw64TE4XvwVQvc1SoXQ051hybD1Lb1vjUCh3cZr7OYGAPU/DBXrktx9SU5Lv
rCCd3Z3bqbzz2KHVGf3Gca8GlmAQWVxHC3BfgsZS9oCexBwcb93Zh9DG1RoZaFDbP/oTsn5TKtzZ
gDUkrz8bc0Rua6PAPO7LHC/aRaf3K65Fq6noR/QuXTdL0cxZPVFnXzkzGQSux2B/sWBEASqdxouR
ACqX+3ep6g5A+VvzwZHLZQyd4afg5OVPcjY9iGG1DvzzgcRk6yURRQE5ii5rnLnEGC+JQ1Ca41OF
mvgH2+8ePdTfdW9ku6h+VsAOfJY2UvNdpRiYsy+Jv/+IAyS3lS8nkKaHjE8CZnwxYLUAQ1K8tT7P
dNNoxn76wMT6t8K2trPx6+0kYWYktPgR89UPBaEbQKl/6Um6wuNHf/pC7XQ+hnr3FJrD4gXVSpj2
QwObMGycj44dwsrdevwlg0hOBI5W7li4DOEZeQ3Iara0SpCUfQQ4NTjlPnYtI08gSXchaEADoAPq
w/EaH1vyh/6Xhq5I0YfLai2eSnZQe3Y1xRHno0avLLYaHMTiPEUdj6BNjhKanDyoXUDSkaQm1zTq
1j1IwgtbZCpEYCTUgjZu4urjpS5yXurGq6aF3gJ+pEfWSji/DHlEzGPzAI3SnCR4WNoHuz8UEhNa
itJNZ6ryOyozItY/VapTIKeA/U+8Ye03Fvt23iXXPSdvE9tRGzl9iPXvQsTkYzzPuRFHMGH74N5D
BnaWkzyT1BZwtntQ0YZG+zH+z02AxeKpn26TZ5LUv3rRu783aSVZ40GwY6OzBGcF6yT8pk0VKJmv
AdS7ZkvfUIa3sw7VMefDgOUObDMc8XiRLGS2uBNIlrpmNoijNFO0dQ0bAc2trUpjGeGW6084BoGK
JN/JhypZJZ6ZqVZM4eU15sJYABE8s+KD69M26IRqS5o9702P4ns+LMUmYeDWLdzyfkJlLDeTv3Jy
YJccS+zJSeYdcjFskpdilccYkH9PpvOn8AC6sC1cA93vIWDKgldxOZbtNioDEwvtBZOGghIPlNQF
o9rwCyc9E4kiVW8anCPN7uLGoYw9OPyj1hIYkHFWzZ9Tfqu/IKVIxldY2yvqle9h+uhyUX/+1TPl
VfDrbfqTF/ZQr5uck4OU63jFUNvzSeIhWeogPkGbYEChq2URziL1TJwubIvauyyqJGyRJQ7YdZGg
BxnIIhZETvxh21zUEkp8H12PBYhrjjjfN5uBJAcxWHzw7Sqp80yYdAuGqRFKZPcOHXZuz7tgn3k9
LxyG6eZhkqBqofHclqAeuZBPVRkR9BetlAVZkGN5jEMs5yUl4CpBPtvXBac97fP9SiUdtkVOMtcM
iBt+4OImzIr1LT/qiqggBAeMThBCQ6fqN8DVt8k4xFIbLuy8IIDcxH2DHiuvDhEDj2qlRMyBH3VR
5yEEE1lvz8QwLfcPj7ZA5KVjeXP6Lk+Rf5tnTFPnPTsGYkAp1Sn24uI0QrJoCzvHR2KB+YikEhO0
buPceQC/ym19fxzXJhhZ7ZDHETOysFG3LQvUmtXqpP5h4G5IbT0RBRV2++PFnXvJcoUil6lB6YED
Q5IFfRRvtn4nhnNnfTDdKX3N2dOdQX0m+ZF0X5W2fuZ2QiaYmABdzFY0Gt93tR3DLpXj881M0uDU
akNistmlIlC5WGAUCGomaBuX4V4t6HGl6iIcS29hre8XZDvnPeUqeE5shjBcs020QWMyc1pGhvrj
C9vechsiBJqL+9+lq49EgXInuqpxIrbMwZPtntrGHww+HC/s4zkYvy3oacjYhJVLchJgGOuFfEVd
ycKf/lYF0Lb9IKrBLZwrjlOWYeQ/CBNMVVF0YaWZjdro47X1K/qbH+eKi8dCMoQDcTmGwxwwPXeL
JtOfH8fXWtp2AiWAG5EmO7RUA3tMCrRiklIjxYCRfsKONXVAazbgIIMUQ4k72tDsslvhewoZbJmM
P8H+1Si6MiCSMjXKPj4IXVM7KLvkER4epMe0gj+mZjw9FUzmhspThlSU7+Dsz0jlSl4sXpIa8Fed
RjYObu/8+O1IhmRRKj4Wled/tZArbM4LX2uUvrrHTtzjyYpIILBrC/2BmjPqF/0tpdpx9bGEKcxh
rQhVZc4f47aCeUBF6NFMhgCM6b1scq3pYRACSwoeDI9CWpRHNMdszeMAetTRAKyH/61VyCTTfZNO
Y/2mQP/3MQsErW78aWEBfUlQKOCp6X3vsqVhymIm5yZq604VzohYbmk+MEBOt083P4SMbuvn0CI1
Gj88ec5hgwJqJJmPHZG4FkGT58K4igdnboIXtz7W6LM2SdxZ3Ed29at+gSPA2iMtKCOe98yRInGn
yIGlLy+UovdPEj04VCUYzAUjryst+fDy4pPoZA1QBBHQu3gIF2elNmPwfXla8aU5VAOG5r8vEAQy
8j/5E3F/huO4b94ev2Ziv39rcZ517CSt9/NpuvhA/yYSUcLELrngFn6ap6zfOWBcvpREfnO8LqYL
8uYA6XVFs6sa9nZ2Ji4UEsvsimmZ/8tGD9Tw0JzR+ymsdsQ1AqkWv1CU1Fa3gCBw6kaoSMtzFnMK
pAjBhnExIiHBJVRJGcDhF8zVWgODnKYrKL5ACMrX+78qghDVyV/J3qbAjWJ1HdhnIwb4hdZyJqSw
x4OpVv26lXgDxapdeUryn9CPGkl1yCq2useFFdNlt1T4rWzQvHUWhc4i70a3wDDosBXLTbZmQioh
5UwxVgeUUxAAK/LmelpsIr40N0654YkTBpPWRiKBZYdnag78Hy91sxe7wJmTf6aNq1EukvyEyqU3
X4ZJ901ITMLKP5LJWu6QsfaZCUGJcVaSD4QqGLjJzcg9b3IQOgD4Lwb7uF3BxLLtCL6wy31I997/
u9kC0zDmXc+k4mPdHhMQ3sf4xnZZYGSvp3y+S/iibhtrDAnYqsJyCt1pWYjjgCaHMUkcqLF9qNPb
uDqXkpqeU2ZkQSALQ30jDkbIy0h2A2G1pRJzdPkuIcisbvqcx2LffsFH+5dtmNN2O+R6QfiPFQpf
fDDrd6eqJtFLsgi1O2v8dResEDOM5YJTwB7/tFj3b/I9jjUcm6dDyNKtE1n11a3nj9erPWjWxB0Z
CeTwblrD6U0vxilPlCDBUM/8OZNvYYW3k+cdOS6jVTmYsaZijgwbbAcFfTTf5q6UNgeFtkLVkl84
W72Ddf3QhSFg06rO+AEJQ//apAKhPpJdX+pBz3cRcv/10KcOOYIYCqn1HkrGgFZqJY1OjyYVNKyw
sjCia9JK01el3C4K0mBKm9l9SbOQk7povWNo9ll4ri0UP7chuLZrLRFUPYY4+4vd+/kqT+efBc61
fTkdRChBSnQ887ZMYJMD2Rf+Qen7OQYmeFp6aAKQpqjdPrWSh8NFbW4Hf4hNtzBJ43UTKipFHuet
7BVhHODHUxMQsnYOW9yWqSormHGujlkDu1ZYqUzZE13HJnAfPUXPpBIZyGN1BuQfcNEWEqxR0lRV
aR+9kLdmIzMH03/dcn2OOS0wBvfcaUeMsav7RIJRjJAfSOC6wj4k1joIuFdwBh67KH22Y7UvMH1x
m5fdUjI1JVJns/5jWMuL23jbagehxTz0Gav47VvHisKf2MTW4rzjx6vUlY+MbRGwlx4M5hJCG44j
QI7w+mZe3S51Y8Zws+CXrZ/IWKLiykWjvzOPFc/el+z7DP8J3lqXIZ5GsL/KBmEvzKc/raOAc74U
+lpLh9c+S0TZpQ0pBdCQd4QHtOje5MrwB3tB4ZFNn5zILehOy3lhE2yIp0wDLcmfjL2jPtMk9Xut
CW+TfsBruODZ25dwzquAUhUuoH5qiAkT+FJE3DxCtijI3185iC2uNaAXrrNWoopN4JY3ng8jOM1M
gXgRXPo8bFygnfMLyNmzv6Jp5iVGHBC3ISqnZx36H+0ZX3+Fis0Nw9pO/2mSYnxxU1pUngPx/1uB
Sef308qVq1lHTxyFnaUzWsXNSafEXG71k4m/EKclykrnUDU6IDYOEG9zSN0tlg1KXumTp69pl7VG
CyTLN+qSg3/g03LnBk4sEeSHTW1fg2HvLBA4Xdqs77oelmrYqgvxr+kvhWDWRiTHNfffZ6cyt8tU
ddmhR8w8772+kDVkhy9Fwfeoba5/AwKPE1vyPuWawT3PtM5UtUf2BP588hxrFncGr4F0CjDavGCG
dnrEBOy09ka3I1fSD5PDPCoUxObHn4ClzD6/EMXJ+zKR0rvG/ELk1C0chTN9Ts9tHzDUIofYGBAH
vmYE7uUl1AC3+MAhuBtX502cwoXMdLteij3ajBJXnRBa1GgYteXdfgOzKZIBO9o5aFVXPSDspiJj
7/AQp5zfYWrWn/k8CQT2JpNx7Uavx9e9Vm5yTDF9Rsjc+w/ZLiQnOGk60H9pvxRMCmQIUO2J6iCB
9YvDV96Upjms82ZzmlLTukFXMe6ua5p4Rt40Y/dSt4uxuvgOgsBzin7ked8FXSHUhDSfCF2s88Ls
+L8fSOpstDBmFERRWRa2Q+CdBnx2/1Z2a9WRp410n+dYvaBzT192TiE7zKXLlJQJ2LOQJXIOMW1Q
fS2y9iAn+hbXGPxe+d3HW5lozbyXocrgjatoh0dXARIP+ygdg+4Zo5aSffg1J8D6lDImwIpPVtcZ
XA80yomfrJN7gj9P7QPXJqCuaaVAux/rS/DajLtWOQCNRNPcJL7clPXbE+cOWgeijUKAM8unEe9F
9xzXhzOpwnih9HD9Z9sVFmrDe/ytbWlHsrGciyAM8lK7Vt694OGlqxR8tKGy5EyU+aQTZc1KwYk/
Q3H+CNdoXWfrrpJDWKT8nC00zuPQYoGHv6t9x53VgHZ0B+/MEJJgqocdbqkW29c8NVPDsfFjpr0X
Y/6YlNR+Pp3+w9VNYpFEEXo0UzV+3i5K5S3ek+AwRgRwzEnKGj02CeDPFWs4pnz4eLVwRbEdsGGY
6zBacj329ZEbWrg8RCY7uyTura4nFOWuM1q21sA3ds3Pd9YO1/nrte8/MU8JitKHcTOMd7qEdnWa
/wiyRI1pQnacOshymU+k4C1pmHb4pZSV6EGH0/zz7HlNsRVFqvxnWJv0o8QI2A5V88Um5Ai4D/Xu
3k5y2tg5QmBzqRfThfQc8J1ouOzC6Xv2yqL56ySWPDWrGamQTiTzXVac1rgLMFg993E3gpyOUiho
Lx+Y1yhE6jdNNEztBUEGd3kdkmL31eeZNZodJsmnFS9cfNKI2fRujotk5uldWKrUzeZaQDv+RxgC
f6v0OgwPbJvPGfGq6rzW1n0Y2jGr4KZ5a0DiP8gRdL832ab59gjBWprvBq6lPj7Il6O0YzLPAAtZ
a6KprM8aWXi+le4x0uHTf9/n+FmT1CON0syPlC0kZ6TwtIfodolEVE6FdzTml3iFj4gTHZcz7T/y
/cfzxQg03bTfQrXvkApPdSDgaoZBmG8hiYH40cg3goJ43icPUvb/l+Us1zq5mHwtQ/dE1rlIk9+d
vCsSdL4PPLvAQxT4crxZJpM/UDDAyfjL8aWGtjHBIIlM5J/b8L/D3EkrSC4plKlMj1CCeB9O3Un2
CIYl4Vw0jcoilK11oxiL92jlM3GyOHbazCO4DALdxSIIVVizBRt4edWQxZ6+8RWUXrxezg0Pq3KH
uIfKWT2AxxtL/nXH3lZtUL0u4+qTFl47Wh0PDUkHBqtxD1UE36D5sSrasMkLg1pb02P+gaS4qJ3q
SCvfAgXxVUB65opSY78C7EfjaweF/ilCP7+mpuKwT+RfuJsQ6IDEMVb3Beb5Ev88ywgdq4/tUrB3
0z3QTbLKdWvb8TqNnZutX0Jy11pz3cxVb07giiH94yFsRMk+qYzNnEI94Q/++f26d2nV6jRroy8W
9C0h5RWlDms4REHry61TGBRUTSCN8ffYqsXQpsVU1tBGiQc/rnJn5FIPeWbLhmLiqM3fS+yX2DDX
XRIqOU4MAkex/je9VaKgJ4EPWYnx12GNLHF7jetmwU6Tarp0gx0XSnRZp+OUO0Dhgu+N7pxLiOWo
tcUkSEGO2Kj0fG8QjIeDvpHQ9vC9mY2DIuSKl2XDfoxVKcar+bPZTH3g0a/Ns6UBk9PNc9WKvFMF
RVKVTHmu9un7GMvtC5tiu5YbFB65o+7Nlk9yyWMChDvPEVvVhHdlWn/v6Uc2RZRCQUJYnh8GMQWO
3XDwZOy9dUcz6SZU3jvQvRQl9aDeQ7r/XpkIQ5SuTLq4SP2l0vlAbBCSO8JjsYYNxfUhT1WYEYrl
Z1VMv3mo9j9nrMeJpj4CFA8EZBD5/FkZmJUlz8A2P2f9m8lOdVjogEXZBhrlufhcbGjkzr0c6Jrx
/SZIaw14vEbgAohffF96mcVhivhLZxDOV1gRSSAuVngBc92DB+xgC1JIgoK+Zg3q3QCn3k2/93XZ
1Pq7+4z46H8IXE8c43vk1PEDigRYyWO0AwZAZJdICIka/Xzjd3lRRfyKKR5BdeKUtLLxu/qdENJn
jKqlAywphWHJdNjRhB9LyN8j2MZx6x9M5CcFz38F2mRvhPybBQ0Ygiq5mjv3BqAOjfr/aUZhKyB1
GTuxlmiGG1iqJQaE4v3uSiMsNtfrLqkJ/KOWgkxQdIATeGxFZmQwe4IUeT7BL1JyKWk412DrX6kS
4L5I1g9eLJnsbMTIaY2LWyY1hc7pAb/Diz6mTqSEIxhtjsHB6T0Nw8f/EGSXUvx8rCXadkuBF0Z+
4lXP/F2kbyqVjaEu3TrTfAo5QcgrBYnLryXQS98yhbq8NeVgAGiM3BdByYaSpTnAFa7jUGxLeOaS
QEpRt1kSD5hHS0oFs4hLRCbUXQHislDQQGXkdSkoTgxkVzFPOjXLRm2bGlVVSxW2x9TePDXEIWlq
zsdNxhSlP5qD4y6u07w6A17dPXnsRMknzcB7fivDuZgsyaQW7yOX1njX3j0tJKp5XQSnx4LMty2V
h96SjTfLtp3qyGYqzC1Z3BRqTNxRH7ThQx3n50kQIaPxlOipJ8IXwyIEujroXd+xYH1DYYk6vjCk
3NBR5qD+u2wCfPJCdsLa3QvLN5YOBzj8taqgbt1MLY96aAPDnL/CPjXjql8cgE+GXEmJBDqPaUvR
FmXB7OAO3kqOZni9hNpk2ZxNhTFI/300JhkjNPStcifpEvx0c15vxPIu4CIHf15dB3jodXcherqD
CsBnljRMGWX+3WJPXT5xIZMA4ZuHzhGNGi6rZOZHxOGx4z6Bsu6p/Fj0ZR5x0uZe2ZKD824Pxt6p
ST3Ex0UT6JChvSom2ZdF4gS4RQGGHowAUHO7Xf8qQqZcxwsFpPFibvNBodQIsOg0fDhJWoU/nP6P
jG+5k0d57CdgnPZs3mPAjUy5ITlKxZM+dtemFCe9l5lAOEwWgE87YR3ZDd9bczLtOJFKNJyclGdn
CsASzd8PBAQZ52QiNTMQ5YIREh8Iae9FPw8fLCrC9euxk3JfSrgiMTYqeaSb4eT4vU/hwqti5Hvw
13m7Gc9osZuRxJ3cV9bXypIlMPdX95i3CYuK90gaSNFhybjRY7bXNR5HjN2bPVxJOpXfHtrh9gxs
y1Wqb3Ur0rCDw7EQ7U9mAupnScYFwAFJVY8DFvMnJsb8pcqHiSTz9Xef3guyxFhwyNFfrjP26kZR
y/uAVHTBQp6FBNSlgHV8B1jQ2LnRv/3VOK/NeDE7YO6hpvpWgbNcMMzBinyhtdS8azDYobbgDrdv
gxpCzv+/CJuE03/NfyxbZ3o72r0VB6WO+l5+7ntaFeotP19/yB0K0UsdWK8yi0QCufCQVDJBFWGv
OqVEDlm3B7UjM1lvWO0TZqAP6gxwkDfa1+VEOUutE48eDDT4oG393ixiuTNenmsdXlJ17DNHBsgX
ZrMY0mNPizSGqt8XOdECAR5tEEriwf3koWjVimc/qK2E4XKGr37BTQI9quefAvZYEXnUce6a2JEW
eQKAQhL3rOlLEyRGpBTUkjtivOcnM5qu9oD4ckD/rmdMJpZ5lorAtpCPMp0Uy9k46ADgFZsqc+TW
mdW3ifyL9vsVftA2EvSf7/R/sRRBX8RaQutUY9Nx4miQWRzj3mwU075Y7ZWwmwFEwBEiSYyo6krC
CLZYJOYYaY0wuqk/AxGQEa8c8rh21DNwswFuUnWprWSSlMNsICYF4CGRWjmHelcgLVvwHo8qC14g
VqMZA00clwq6d4jqWZWyB1l9lXPFgCSfl+soPfq5l/hzVwbuii5ty5g7ASfG8wjiCslhOxu2b4oB
Q7T0uzId1Z94eZwySF2DfiJn4di6cuIJeG2JhroHZrjJ6yVnsuUiRjWLU3HZWEuRwjpHDfpKuRSB
YncZ5P45e1H5pZe4z6sJLqzj3NBb72kOVq+F6CWc18S14TT+1781wU9nVLUeV2ElwZQXUJoRCcIg
xbaJrj/C9huBdf2aTzkaRpegmDr1w9+jSt9QzrHJc+IjwFvxQtmvRe30TUufAwbWXDyL6N4orId/
S+hwk53W9ll6SNukTHjicGwRQY56zKRbEYVZ6w2zHe+47eNCsao2ki+NG8h3OSBQmtBTPbjm0pHe
znL2jM2WNQhFTgKCe6wNJsLbML0EeD/PXf+iuiRNWrjsP8oAxuszaqT4ZhhPoFSIYMObP6Nb8aaC
JogkyShDKymwNbEVzKiO2mWl7Fnzp+TehIuLsovfGHxEUbzLuS8ueeRfTEhps5oF3FKPqbZGFthY
z17+HPSwbTd/b5xrstIU4figjzmO9RjT3fd2cje+kiRzfBn+LtbHg7m1ff6XTLX3OjpaEn+i1bgO
1ZDLP0+MxypXpw289cH3g//6Df+A6PtE0hVbKOD12GLI1tv/cXBroOhaYslXqLwwpShS4cEZSRyL
0liklnNYmj6QXyOfhron99iCw5HyKu+Aanss2i+FuO9J7iDnOLJXbgU33F/Mk6qRpTimjkG5maQg
8fx8Fie+DUSY8w3NXPwyBtnlrZMgnVVF3weVcLYTgL80v7M04GxiElSRenq3w1WnZzy0dJqzDQmN
ijbWMhzGlJAKGShSGHPAmdeZc1kOC7eJgx9E6GEpOeYlyH62jQxUZfJEn0E7CNntlrwdS9yZsrlU
eXn4aSVOm0LWN3tuqbSDVmgnZDKNvPtVDDEO1NBvz4DrhFVRkjnzBvFNnhohPxXtDQ70Fhmy+AyF
odvPlGPATU8NnMVFiwwpPSJxka1mAlfP3Ze2ZGmrbWcv/a7zJWWXNhYLDIXmfys2UCAekTd6EVnC
ynWITaZfAr1jJCny9xFtlBCFt7K5xfA4dwwwMfCfKvklDSb59/O3TJT9ykFKXK3G6nhruYVQmqJv
oN+K3SAs0xRJ95Jtc3GBVN1CjdhBCDTtZXNoNM390Nj54LDyb6h84vi3ovKSDhRKYLlr7d04gN4I
ENeBdccWvlVdGky9yQNUkOeSxmUnTjCcr3fZSAi/Ny9O5sgY5hm3NtVeTL38mOzRDnyZHubjr6Z8
BdUyGbiqyAjg9UD82zvM8AgiT0nlM+ZnwLa5kJkgFp8szoECz0I6xKm5uhwXt8EL3zzESXL7qkcT
pLNdtyKmogOnMHgia9RxyRvgbtMMYGIQUm0KISzk2YsDM0wfMBaoVGOqCZIephMjqsaAhqOnraML
SgzWcmrsoOKV1UmbdNYR+hXn3XoCx6GlvRsv4lwfReQGu1USF7VZL9J1JmuV5xYbdzCYydIVMvsN
ICcWz7POxYufcF/4DpyXcPXbqMiyrfQe5UA7qb4sZe8ujYe6zJtHDzTu4KpZ8Tl/zaCoYiwgrQQc
EXc7TtFPH1YQdNzkCzso/3HbNUMk9lB5kodmdwcDZ18W1TaopTvp/x9lw8OiatUDdWNPdSo0RVD/
lV7+OXXPIxW008gGUoORQB8Eyn0oWFL37n233dFoey2fMpnF6m3bATL3g7OvfCpk4Tc5LElOVUiq
KCIfHT+2RB8yT4mxzAGcOotyu2fSql04iLiZiIdQ+W8QRae+6k5d01q5rZ5qvTabMwY6Pgd5fs9U
5+jWiDqrt8X9uCWUkgEVBe04ZPa1uZhaIWSzeohI3dFnsbiH4IEsR+tkN+xfdrrV0x4fj3AfICQe
oR1FwlZQaVOJ6LnSzI9nuwnaqfcwby1yRCqnjAF4Q0EVZD3AmnSf3FHrHtjw0eDYwSaZp2gUmW07
2mJhQ+Y3/SJZQ5VdRLoAOhbBGbnGPV8AX6+QwL7119DdAaW94D8mM514xJCCLp6fviKimwE3XWly
mJb12xFopplt5dRQDsQXXkeo6R5KB7Jo1x23l+2FtOg8EcCunZG/swzQLlOvgIawg7RRLf7R2e3F
ceXHFdiMdXK12b0viKjhRcqiY/e/Dn7GBc9HbtoRBar6DNMXLQjvZ90UNguF5duPCm6u7KTpixgP
4TPpNCQlT0jgBqyRbivF4Cw2vzLWL0EUAaUWooVyfAfXYKjKzY4BUIAU2/oHuQ9vFAqvQL82qZR8
upfpvBhQ4htKbzVNDg8MzwsvGcFJLmFj7JM9/Vh07FdvNmTx9hc3CD4UymVjGo0PilMSn+JiqVUn
rWINIIrH92MPYS7sCWarWiDDf6JbAtOyCLr+7RDpE2zmiCrQuRuOEbfaqIxHiYjR3WUcs5LXDGDc
Y0BiZrJ9qtoovAI5ku9LI/YMS2uANIup5wmjA+M9CHghVWpbVTn8EAy28pEXAqkEQTa/WXaMIUxk
EhCwep42KCESD+aaRbKSHi1ssYj/9bbAwN9EGBfK0IHuwO+j39SMz3DfvGeGKkTu62lRg75wVqzF
hK5jbVUm8+6bTt6r1ob+KhwCyxE8wQVd7RJN8vhtdS27GgFa47dIt7GTgZAEYZduQ5NM5pwvyAl8
KJYIvB9nL/ETdsBFx3GCIr2iIcFitIfBQOG6vkMmjGR5W1wAFPJ68pf1PiTHOG5Pf3BqosI6Gl+T
1IZBaueXBS+f0Av/rMqmjVBx5mN+sjCdCB2EvlGXZKmL2EXvOnvqiA6Kq3IbZGeKCLrkI3QCLi9t
T5kLdRnc2aBWY495F1FOGGI2PC1oMxYiZd69SYYaviK3GRfd55wWxFp8KDHFrHbC0gA+wi3hFb2M
QxvU3cxftksx1gqByZB3ka56s5e/mVuIeAyaQNMqcNzs4WlvxJxGoWhpSXBLpHOFjlKGrxr/X2+G
cTkab028rHQKeqrBsrY8cU+dPpEJQ02P8rQw5rlv1jfSZ56Ad+6PDXSpTOgkv5WyEj5jagJdMZQR
NaanWaboTooNKQVyEx+E1Ik1SmZ4OaSvVb+dxMCVIANeg5rC+MITEqyAhfwhAvOiw1D87kVtqFzQ
S+Dd5U3JgpEBlx60vroWbZNtdngMN7q8UuvEcxFOL6KHTxV4KR1rdVBrOUY/ZxZnJqd9GAcTftfJ
oF336oGLmUlCKAOAOKCaxtZENHxuAtcNguXMpiJk4v2uy1T25iAIR90XX9uZyQiKYcTEiK6JKNJP
ofsvFYcYKMcOt/7SKdpAhkqxjQ+m8VNC/+Yn6JqAXkxXQyTn4Ewpe+5OvV8XUOwoddXTKLA8BP9R
tRvr2BQdg0mnnj6KfzXgN9cH76J2riAtzSN8jHmjSiSWQ6WntAQuJNohiWRcignXBJXTk9dQ4SCP
Qbt1sPh44kkRjkOD5q2WfQxg0x89OSk3F+P4W0dhU1VTEa66J5JdKY+LFuoi/vcx01DKWcJT7axX
gm/0SpHv3XF5btZMbTv4pA9CwrDo7CuxeZt0TpDVQHURK17dvGaV6WtS42tNZQLz7YsRu7kUXKpI
L/CXfly4/g7pqz27ib3r2yaLEVsEzr9sngbAjJhGIF0T6GlTRNSHA1wuAXOoIcwhtXla/qPgJxvE
Snut3chJAb8ILYAOlGKh+KNZ/l+qvvfrxKnXnq1p/DbpeOrm3hqVQKj/ANLLGfWVsENu5Y8Yy9SE
jR4Jg3goq6IGVYRkfx2FzIzwXaDzw2WWKTHcUPSvit2LKekrtnVEOT1G+TO5LyWVQzAMhauFjX7g
Pm/0rBcYd9mo5yH4iCAbSb1+ZNebjUuDEWfnaO1kAKcIFwqtw72cJLY7MlYMTydgORMrLrLCIXYv
+sCR05wTVV4hBcsY7PdL+LyWS1YP1CcXunccfvAPXw1lg5eiNbRHHfr3Gnx7RjuZIS3z+U5Ej3Qt
/TJutQiP0xP5vggu6+H9r+kOWaxQ8sTcE2Omtt2uhDqz87Xus1G1ChEHJdUFzlQPIp1VE+IOfh+O
moPA/V+A9Xw7wJ0Q8jOFan5KwTJQRUBNxgDL9sf6cKFW4gwLRiiGEXodZb0Bm9pyALfKpgxVHH/+
YhD/ko+9tzy0ANBsImQRcBS1SZCb0Q44KHRZUavkPEy2SQXX6HPXeHdzvzSQkkFrgKwUDIjJHoG8
hsJ1l1L52F7HJVF3xr+2y3VU4IUaQMkuBoI10wDVM3BxAUo4esYciJB4Pj2xEpNjmlDISDJ/Ksh5
7QomjTUKAhyl5bRAL+m+/JAVPyVZWrU9HRPlCosu9i4Vs+TCdZOVeD6/cVES1xKeMJYj4CAs1mGQ
0CXnsp82Ay+Whtsu2/7OxzE45CVJi8lJ7lVoyYanJTMRc5I7OwZjJNjSrfDlbbze8tIiHBAj3tNk
sFX8k8VLlwS7ykr8H1nMegQ9OvCm6/nerd3J9TEjoHtg/Trg+HGlchFvGcYB3El6HWcLHsuT+pIt
v+muk4Ye8idgvSDTAWo9dmsTStjgT1lECWv1JCGKxE+WqdDnY5NMQV/YDt6mIZ4FkqvLAf8TcLYY
ZlX8hOvdg0APDof6paf4DWZjKsKW/yOk9fraGuC1eEA2npnqRWbWbT35T++WzPQAQ2mf9T37pChH
NyZzT5iuOMC1ZSSntY+h1melrSi1fmtX8Uht126YalVp8Y7o3UT+Cy8JytnxEk0z6pqirBzwLki6
CYYeJwgjpxarfHOPmde1uQAH2Ckte9NioVBJpZmocNk/ZJG4gREQ5yeKFQdVQYkOGCwBmNLjx2HK
DzPspRRfahorY7lhXwbp5491G7UChyHTTqkob4l8+GqfJDNTrZ+O7bToytH6QVKdXLk6r0p5UmbG
OPNrFQkw1waLpmmMgpW4H1VTWXo4WVc0xb12nDarox33gW+wDYGsLMo34HaLop844iJVuczoQhIF
BjtD4Fqt7MZXr0HRP6mgG0QDRjCecsqSfrq6SE3DfFevtp/8HaqLiNMiYiwy3SYl9zkFQLHgIcWm
m8iG7s8EPk/uaillwskZTCxFTfCJ0sMfqZaKJxn0ZEaoGA4WpHI7FxNu83dnXRK/HoCY357jnPjy
rZvarrEuJmujxiWAGqevO4tjbcF+aeKgrMjPLi00YGpaOKNAXQQ8XFT75oLhzmgOAF5S11H+0aOI
wYyPylmOdKSYMGaiSEbI74VeryaKWVUCkaG4a5Fyo3FkFcKE5kYKIkqhhXd5iROhjeKsqOTHl1jh
atG/x5RIAbly7urPjuMadSUKjXg8bGlcetpgFf0CIKjNX9kUoNEhHhsWiq3esAt7MZOarKK4FH8+
YwEznDJ2yOo4JsauDGEnKuDg39KhzukA5G57x2rPXruk6Xi8nQK6xmkqXKxjuay0HsGhsRmHubCL
XweXWI4cNxzyS5qeHFfaoqluQgcYUjZEgZqcI1bWA6DB1ll5Dm9Tb1UE4wBEmj1S6AZgdbNO+K3G
VHNDB4gJAXy8m2U478Zc2SEh/2ewogzM4zPV5vqxtPQsMN57U7ZIDkmli0yCj5broOESjGlO07YC
ehXbnfWM11kd4YpjscXEVWXpk6N5hGX4h30bH6+gMlEQpboYfyn3CXurZK9jJVKvbzvhJ8iYD0Lq
DeKfSjZnhyPNrZ/0RiUjJ5fJzU6iPa80Me9G0WD82LZztyWjxZPRPfuCNY36v36xES8HYAJT0a2X
7E9gIKCafeV/YlaqqdtY5ZZ9SpqeqacJ4Vf9n8R9c32egjNprFdODHX2AQYU3JTMARE3JHLcPlxX
PoD09RxwON5o1Ivbqot+Dq/x+xVfBRu8AUuSpDWda6IWU3sC1RbAck0elQiPoe6Ei2ipm19A/0cE
QyslDKO7yg0yZuPylbaIU+y59EeegP48AbCZZoYjEcOB/yRD6aAQBTQMftFH7/kZz5WUm7r6pPJC
W3xiMWeSvQyiZVCcF5FEL4rUn6JF71jvwSgopEhP5pY2BLWhVuE4wif9tPFbvKnePCKQJQLTEFia
3X2RX1QdxKB2n42XyLDGwVosIqLKMrI/zkUU9i7DBWAS22ZuZpCQozP2Knq5EDe2wTr8belBRj8x
TLETUFLsUYwa5LtmPoY+fgR2LIV2axnfSwn8WQZzKaUY1wrV43Icdh+/BIoOFgpexaLig4nsjY56
IXGCAJ2Qj3bgcAywgePTZeiV6/WHK16Ultw9SvpL6j3BKH0BwMvYmsO0TcobL8BNjuGKmGaWztSO
Qwxd9DBdRefOAQteUyDYeslWahDLJEBVz+E++KqEGESh83/84VOYC4SgGEv+u3RfLiEG3XIlKrrc
2DiFLtlCtpvDMSG2oeJsRrPAznM21xHMbj8ntAVWqvWE6HHEpUUuoupkJ7y89KY1qnfPjAK0wjVy
Y056H2SaW74/em+QuzbnxATA2VEP1zfz4g+rNPqOJllQxEjKRV4knY1ylmeOgF+bYwEzvSy/huod
bFeRmnhDHjXrRAMrm/GPTcmYpshi1DncveqV37EeZGmUsCYRzBaE2VNYcjvQ/lEEwwIQWUDWWc+y
T2yTSiE49Gu84EmYpKMhR4g+JGw/fgIcEdq9tA5ZudR7jXL4rDAZFJGy1KJJ4ABnei7EvOhDyhHD
Pgip6fPJWNj9Jae/jXASRfQbLo1wty+oXtqpRkECoC+L4EQBjVg1cvKN9lLTmBPW4Du5Cwd+7fqH
Ho2vax6EJ3jNEh1snRz3X4ZVXstB7NYYfrz93sAwlZCSqLdOyLTrvZwmVcTC16oGaFfu567UBqCm
GHTtb6L0pof1qqbPzPzlQSw+GWNPrPuDiEs1qjW+BINFQEAQm5jb4yDFd4vyxn7GZQsXM1k7UGRM
5V5PiLb4XMisWY/4X6ope+buZ2BNhdxXF/of3KVG3NAOgxHEyTkYA2u2D20D+NesXNQAf6tIqrGr
JM9SqlLitseLIEWMCcTv4LEEzUGUzNgrqWHCsESHnW75/BIJowWnGyOPwIT/rjwjzev4hVypo24z
iLSUGnLBRZYPTj1ItdJWcOfyGRRb8piogIq6KRiQTDHC8CKTCsBwQrBEFTkQXKREgn1+KMtev226
ZnfslZadf6wLKnhAkcTC4DFyDFhxxubIBIrKM2Os+eiivYRs4IG0evQg3UNR15v7q3JOrcUjz6BU
ZgilJDeOBLUg9Nc3boPyKKiVMyxJVuzJNJjmgJRyNptG0DSEEH9+BiLDnUmYxWn0t0PrMBzdCiWd
BAy0uaAFs2vkaKBW7EdMkf6WRZpYQxOjbMOSEOW7mZUOCWfFYkHcO0qLHHjuFwdVS7fcuQOqRbRm
k4F6iTFGqOeTGvIhkKW5FSi5zh9axA1nXLfBq547/YuQAbTmzNvfPbV+ySTOO6aNLLFuo5PtxRU9
fIoZyUb7FPrfcv3GhHx0HlM29403D65nbfrvf7CZiQXHl2RkKsILbpWie+ZLUYZ9UpFDSJST4QEt
s9ToFe7oPS6aNCw3R+Qhsu3Hp+KDTXdmHcMOvFCdvfYz6UgAErLBkgAszq0FQrEeYQoAdR0ay5zn
d5EX4i4Dyo6sRhkxPI5c6CvDEhbN9ghDQdYk6eqiV47U3+aS3BHspX8ygtiFzME2/btnNNjnvCX8
1x/WaXKBw3IUzlWpikN6V7h/IM81ZN49V03q7Gcr106gAqAXIFSr4SbVlB7AVeWcbn3GJi7DPE9j
L6Eyn+RHHZphoerg6gG4GzFa1j2AHwHWBXJbs/4JtGjLXlEDYTsFZxg8uVXQ+Vgxo0DgGI+BbEpE
IcEmE84hiUBMfxbmWNhsHpbNenNgX3ZNX9bMvxIIXWh93P3JEoY4LgpZ3rYa7KYZWi6MmUx9FJ5G
Jx7NN5FmUsIAKeFLEYEqUl2EBYE8D5YVtzrtVYgnPzrxdXoykdH4g6aNuCRYfVhxSLKo0ioC/Gt5
/Os9/ZV8SdEgzHJf2MdAEMLD+6y3D7KUrd1tCjlyF4ZPu0Vv+/2wCB1k85KEyRZfyPJuz4xQc5pZ
YeDcRiI37I0KHNa3OYbEuxibvQkJ7WNmWKjLCtRVyjX5/N9/J4iU3VHlg9WBv+SpHFjZUlnFDrT3
MDfcpoaRC+okkOce9kcKoRGFSxa7VA9bNBA6d6VhD3r5iSBmwLYv/BQ9syw1bPZSEuSAon83QTd4
rhHY6KjIGFCfRgOv60zoFAjKsr5NBT0nkKfgWzT3WSvZavLzvMpviZ53PDTscHJ6b0x6YiuiRYzn
zwrMP7omjC6HZu8Pe3bPOcDSBEwpghldPf8deXtq5cjGVRYnRbu7xb5du419knguMuHR7Ur2XY3l
m6JD56larF3DgkMbBwxTnhkH+5EHa42j8otrrgtM6J+BOPBQNZuMNp6KrXT0LOqqZyeCj+OWRiCM
larSOH4f2Sf6B5pi5u0OJoqXj+XNS/tVTCXdTnD2MBYEI2fDqPNybY1WMp1Rj4tohx/M1CQW1tNk
jX1BtGxqyLUTIxJniCFeH5dNV+R7cBdkbX0lZJCdB6cIxREL3CKq0fV7WVfq1SP+UL26yFudXCoJ
PooSF+PDzZvhLbCqIEUBgVSUhutjW+SIymSpcplFMVJcViUQ5mT+gXQZVM/dbmSVdjQPlbD4fy7Z
oHRMtr82vTWckO7yrWiQwHNZw/CAW2F5fyic37l41SMEGPQTckRnenNpLFShYnVJJcry7W3/hUbZ
Df86VeYjrFhJfvAX39WUcL/blnRNRG4PxFVIj1saW5xDztWJ3r3xfZ7IJoCHaxzOMxm4D12zh9ZL
EATsn7zA/dbfGaFk1VzDiTKxES5e6MWTMli6Gvj10YtdqpxmgIXcD8eVs8wfUw4Nz8R8KXsR1u1o
oa/9THYeGT1vuJp28HJiG1kRlkCHfieC3Ck9HbnoO2ErKTqaRdwojvPL5CjoIKy0ejAjBrL9TSyE
Zt2TeKrHiJd93me4NXgOUeZobxL2rSypLtgEu3gRFjZJefy7KK1CqhQFyCn/kNtjfG12x3GRtrmb
HNvv2oRfxo0vW7yXmNcHUzApcbg9oca2Gq3GS8XPCAg4/WCj9UD54hKNxI641BCZyVNEh/owkuf+
SBQycEgoTNKQnxEYNTjGGG4aj0pqt+egJwELyOZx/BchXbbyog3bEBLQu+59nePadN4wanUZuiFj
6elW5YKAZc7t+8Lpz2KeiZxWzXXYOCk5PAdzlTprrpGvq+nyUfQnDw6Epg6R22tUqXHHaFR0Wfkq
uRFfH0yOqVGh6ZSsx1I37Tnf0bEOyQdbfb2Qhu75xjdgcZULXTf88C+z6k8eKc6ntcTsu/qkvFMt
vRyToNqzgbbwSV8pt1rRMe859Djpd4gYan0zjtSt561PeSqX7yjTMwrcVFon2CIUESW6ExZyhnfC
3xHzvTBxyGsR8B6FCNlyuK0xLZv8i1rwCQMgMNAq69FGCkYvwqe7sm8sFRoK85gQIIHKQROh77Zm
T1QFBe4lVrhoD5PbZJlW5Ao3WoNXJPwkVgcB37ymavCxxKjFSaJoHY5GSHJfJSC2XNvvfaTtkA2K
XOpstCUX23GbD62BGXFwclBpbwucOWvg3irjeq+Z3AjCZWHe4Nx+qU7HeZOFMUHxFOzKuKNRbILr
dvnz6UCcxDw6g5bYy8w9KDLznd1WxI5E9S9Kba1lbi6TH9927tlXdK/wZOK1On28MPZozltmQbmP
h1YZir6WnlP+v53/uX4LI0x+BaPnz+X0B1aiNrjUQteHV7uiKxPR8/Q+SSJA70D2BM0WJ40+lGpL
HiAjyknfICPME/YL2kwF6JYuV+2L1rihqKPBcxAsWOCq/oaIUFDPCLjek0/CXt1Awnv6D66w9Xwd
aTutwrKeDx4OlkRtUm1iiKzAc9+6/3idZEjQtSTUqKi/9hVWYp+3CwRfT6o4+GHoyg1ARVTIjlEJ
4oE3xTKicfeiNiYmAvYlPycYi0pkgUP6l3IZ7HZN9L+rmR21ZHwNXzYLJRPL8tjfSqIVbEZq0hv7
qsq24EirOIRW95TY5PbX8W5ZuwtImM3cUJyagjOp4t5wihLxhcGYE/7bwe5GFYEbT5u1LgRkT//8
4pzpcNWzXfFsP30RSsdAGopAEvZjqAsN3BDwI9te7VSJqV3CMfGrtdcGsFqu0ZsJx202bovK3ooD
S2qNUxSjtQUpzDD2eqzxPHLpjpMVre/tyXrSznvbTEmBlku3DBw5WHFVnrSdZE3hTAI0VvRg6SEv
Mum/FqTgbHjWdpZ+RvuuuClQJBHZ+Gujolh8YQchoX+N7KAfFMo6XVyH32ByDFEOqJHG/yPqTrXp
0w1igHaBNatXL3bU0/kQenoN9eL22yQsrrtseoCf0pCB4maESzSvELfVfLSsVkGBNKj/G6Z5sy6t
7uP5b7CnA+kH0gjbaOWcK09P6NhClXTDCSx7hJazSEvjxj+4bc+NzobfLxBx6UsvFOvO6t5ZoaTN
3FR1spXQydvWOHmtSa7rucnFoSTfxVlzGcjvoFOzvR8ogxFHIWGdTnIiuv4MkyO2v8keGw3RXsXa
akKCdFg/O4/miX0rELFnk/0+GjL91IO6gC9iePtVPeAHp5O1D0noNgzMqDUOfGD9VwgEvH4JB+6e
zK5g7a6iUgylw60dHpjI9bMZH0oKzIjqbcLOToT9Bzusya2FMPCKZ3GVGAmE4d5k6O7Mn+/XJlWi
ZPLvLPoEN4F6CId55iLEuPTOPleOlT0ULfNu/GW0GRt3KNTdacpJrZVegtadVnCZodziupnnJ2Xy
Mq4W3SQld5WQvik7KUDYT4kPz7xXB/wyPgYPUjmlzYJrwpeKazynvewUqFr3wbs6e3yNIKcSXDC5
CResx4UCqvWGh+IedRl7iXJF1txuuzqrrnMkmn/Wo7igIAk5Fqnsb9nG58FReL2SBJcDsleEmh95
CDDo7+Gnutavh4EMdruxjODHq5WSxdX0iYgEaHrbeVmuIBGFLYUnIOHwOeHJXxCHBcCu0EGSGeeS
rOAdEmZh22+kxXxJFz92vB9iXMyzHZt7FGiUp3CC129FqZ8gUCKeunvam6l3+6hrcTOQ7b8zf6sa
0f3z7b3Cdl7jObagdRayUenAzRu132/LtbnKHeeZtMdAH2fP/5lRHQJTKSdYQHNa1upYj/2Xzfui
zespanmzreo22oziMNP49uB8oUKnkXJerRXsjSQ2htE6zAd9R3NANkkcRvi4SoefUcmMRcquZ+Tb
WDCu64kDbgaHZBE0pBW/H/HZjsBAwgw4vm6hIahc5pccs8WP4Rr04t232zu8td+0CNH3yDqe2Ft0
q16IepKg31EeJi79KPYqqeJJRXgmKm7rVQbCNzZt3gVvQT/PSNaMmCmrTMEtUvD+PwyvJlb1846T
16bVg+zAFTQsN35rLKlhnU5gORYi5BkXfsaJ5fdIwiZklgwzfsYibAvlgcK2+cn2kgT+Un+eNg1S
f+ika/zQtXpOPt/1R4TNZA4w5SXXcH7DpCi8+SkIFDChCgs8AGRmom0RsehiNXpgGL35/hiv3WV4
sxo/6lBdaLYAZEuldFUVfnMPJA0zcthTp8h7ks8LAa5YQtdM6/5iMLzRqMCHR5DxjAdZSMWneabU
/NtuATDcLCd4CBOG9DCppBR6PLDifc2Gsc0LahvBvrN3T7/stoM7mYmSctH1L1+Bg1mvLu3/GSs/
zEHMhx11MSB2zzs2+KJmaID+ZxTElZ3IPH2jvfiGVfiwp1avoEyiuPUNY0ywyAOyKccGmQy8LeZf
jlNPyJMfd1TsWj8EaM507U54Bb7YrM47YT0XCG++YdCtYIGLnoLpUfo4NhgkJr1aigJdVSaRsCpm
Q5cUv+ldCq2hQUsGYMPKHj3El5vR69Je7mdesZizcJVH/dLDkdsN6EanRY2kACaUQbulE++FkQUz
4LsLeV0clWJXv0RVMDy7J6xLkHXiKyOK+tpjZm61krxa85AWC63pUZ6X7dq2EaAF7EnhPYTesuJ7
ilKvSrAznMfB1leoj1uULctA+o7Ug/bIa5P73ohbFEukI+GcLRYW39zsdsUTEVu+btA2mrrChRgI
0T5vnOW7dlKq0WK4cBfBtb3FnD3Kv4NtbY0ZU7MVXmFLC1NF2DPya5N0u9Sbfs2L3qwqH5Ib2PFS
1x+nmfHb8BX3+WH3M9eTrcUWxSJHvC9Puck3Sj97yCUz5KTlPd2G9ga5ljWyt/7KmiaI0/djzDEM
nLXhoaBOp92zJTlmOfb05Ohd4pLt/ven/gdESS5h/A2MV7Pmq+XK/qRUvljKA9Aff28ETiToDXvv
s4WSLwsABDlM4HYnYlmGuYIrhlnGFsTdmRnCD+cKbSzOsG4to/xyD+RPMQpOAST/KAt5lJrGk2bK
Pki1Os+N38kIk9PVqyGdoPyEPOBsItI/yyzpCqPnW9PtOG7J9Vaui6eDWmsjCX6HfhggvZXpAw9t
QM5ZVqDjithcbLQUsimreQ2RPt7AP8EBPjFWjRuFuQ/nCIMLQSDf4vuKSacXTjk7xNnzqS94Ez0K
D2o1OwIHG6xSdAF2RXGKqJN8QqUEfsts6edj5BBxkhxLoKoWurvXKSdaJT83HyjG21UmdUotSAqf
ZLM0QyJtgiyYp6VGtYwVNDuP6Kfc/Mr8+ttqSFfJGYNkgJj9iADwOrb2tWiGBvKqRI1U+uDuOEnP
GU57RFD1jIvZlcYpoGJgOJ9nTEUhcjU3wvZo4yJlV7yGEghEKZiGV/ruh+FX55oJNP12ZmxMmI0L
JS4ZykquCk31upsXrClR3IZSEcII0zLTNvdHvi7mBSuGudBS8gpLtT9iMrvU/+qPs/a+hmE7P7aS
K613/c49xT2+tPvGWMU5Fue4Povi2ZcoERMd9dVtUVmXuLgy1XMxNiCl9G21vuUinIZmHk6cvP6r
ZHtUOBgdFMPaDtLed8RnTJM9mrO39ovOIUocDVYqIjFBFaev5Z0AjG7iI8C7C++ZI6Qt2Or+N9xE
/RNjhIRQRP1zH4ey9TFobxeCBriL4DeK0bqlYdvVSlAXDEKJ6oqpOP2PcN0hZ4YTO++H9+OBYiY8
QJAPuEJLqN1oOLKk8sH0ZFIVnHg2+Cs9ME7BLhGnkrDg1E31Q1F1p2FBtBKqD+pRaD3EdR2Gu0QI
vA8dEKKb3+JzZ9Sj27qB2yG1tB1fQedGRZRe0HgkymSISzucaEUxDCCvkb3jrSJpkNvC8G/cXh+s
gQt+SAHBGhJGOb3PjXj2MloDNQYxUx3xWhLj1FAIGnbpdkeZyKzIKufDFa14zD2FVPvbhE7YkD61
oHUDOygTDF+ZOXmhmIrakO6+yi196Dl0mbsZnNPscd7Do4s69VPO/g1SRxzhdBlLFNE6FAlTIFR+
Y+cjyBEJXyvSNoFwQpCEewkqAoNG0cVGZVfgVu9QNxCXD+OFGxXHh+93QMeI0FkmeScr8/sgmeUf
wLPuizP8Zbs2YOipxMLBXQfP/TXRJnAroY19XLiZLoVSlXjSwctNn1NPds37K9bPL8/yfpIgj2Fv
nbT2BTtTST6j2rqnqtoXkEEd23RkJtREDIbN5m73WxNrUhM8DIgys1JXd7W5EGJoh835FOIAhj/M
Rh0Dh/Taw5hW8dORs5gzJmoHZsUSTnRdh6xFdJzab7rGVWLhVv77TTxwQskdY6amTx3YNWzbfmCi
6lDBLXN0M6BkA1Ktnu6ZZo/UW+4W6dRC0GoaUsbK2RE8yojhv7zHfZ0qnLzCGPvFFtrEIE6Mqatv
kKR9EdIgxII8Ggt96XxGfs4uupBLE51zfHaz7Ug9WqAp210toqF+0RNi2M++5FYO4fghPZUmihVd
JecKpkiv8GlLT0UHWMj33RfCiHVqFWyesbQDMq4XuyAJbYFOlBBe0HBQBMBLk8JcunQ9SvXL5aFC
NEPZAqdHq6vS9XGHLHLFzPM2Phm7jGCnqKDKQKg1nzxmD3tWxG9/+JdJWP+Ib7lCvDXpQhtwTp4S
MwH4AXuSAy8LlMwkXV8u5cPchZd1VsIJRjKCg/5wO8SgFaBjeJj982iTgTBwAHyAYQ+B8mQckq21
2VP1SrbK1ja97ec94ejsVAsMX79K/jUHt/Fkw2BSDUgTeeIJpUi+UyKyXCj4+GJWY2FUSEeJxkTr
E2To46usJYSbcRGgu8kb2vO0WuhfmKFYJxEr12IKVWeO1H0et9/F7x3KSAZCMy9d7jMUSv7UNnEX
lDYF12Wm2tnuISIqVs6tWrvDt30oKtD8Ilkj/5+kfmlB2Nl0FkYpS9XeLBXQT/qykhDSE3hx/EWe
fNP2mQWiFRcWv9kEY0OppOUDlqZ6Pnx5kvkqhEtd2sduM6qqGxLvMJ1gzBwRsFquNRa4caabwvX8
3yEa+Ps48tkcvhm+l9u9xMMnBVNfAcRRHeO2IPV7reViSt9Y/bES55ofyS1Iw+FrvHWKLvt/9l1U
OEh6mBfaVhBePQNHWIRtZf85NHoEx86C4snsrt0SnglOuFPneVsmge9Uzg1YO1LtiNafSR3uNtt7
r7dSBgwxaBjc7GXCNLTQCeirO0TGCc2+xAAtNgv+XoXkHDGqfb5/JCOHpI4DGwV6xBcYpaRXN8lS
b60k5AVzWykqH4NNv8sgFaWj1a8Lye5GZxHAalfVLaUWuDLB7IDPwbBkrqpaoX5jA9jSMeFKc574
pfR2bYNiGScevAFLFt7xO6+mNaBTE1Ye1uVb9LwfmIfK7zW0RB1paIE8sngHaZT+Ae86i15qkWlk
GeUGjKg5kI+BUY6eZdX+96uDGWNENGepNnSySK7RHw2ugVjV89BrBvC+P73pP0BTR8PmCAEvR0BD
QiOYMhgyF5zUJJ3AlVDUoZ5laAkXIaOUbHbTQRz8zR6+RcCWS4BA0QviFVgUQFfl8aKslD8E44vW
wSp9nrSVYbhpg8GgJoG43r9uuT8pqj7imSbLMCojRs3NAF5XZ7UHtE5Np0nfFQd/ToY5d3ofDsWC
Nc6zImZ8x0uEi9nXRQSwFNsbziHvERp/OXkzhDTWD2soiVwU/bRYJSsT3FyP2noIxoLMMDLUPkxS
33yQCx2YbqH8G0f8YrrecYvfsiCopiJQFDj7zNFPRteoer9GgARnln8JCblJtc1AhGBbiiIazQcq
9QhLd7fBeCmCfSVipI1Gk43gT+9Q1sWfaHViPldBBfPOOAXdy2Vw/nqs1Mrk4/QNNG52WBwtb2rm
sBcMKe4Mg23LspZKI+zy73TSHdjVcEFaUszpvykSEXIihbklIqcm/hrqek5iQDxwVNPGoLKs/7tN
uNR9TeIYKKTGiSZXIPkZ/CWi6TvTwVNluqH1FlRNy4d01lIzKupthKizuvfYGQ5Xm4Sk8amUpLnM
fNgsLpiB7JP3J66gLhMCS8HkF1CpG7ljmJfaXUaOVT2Cm4rMh4YAx5ku3ZdbHtJQUu7PkzAW08AF
M1qZdz54o0cvNkx33YMXkDIdrcwY9JWNK7ZtFPfoZSD4rDvCUd0aVg3ZdTO7dNJoBOTtu4uPpZkr
9KEEA/g1eLNVutkBuUfMO9IHjREKVVgpRe03JD0AwPsKtebSVkKfw8CwYEdq0iUtglyN1ZcOUzAW
xC1ow5pbcsMuq7A7ZR3v/E4VyGkVgdbYgzW7CrUsIlwtmWivdG7PFJeDExDxReZm0oHoWuW7mV9d
r7ochmbNRTg+xTscOy4FsKI7k8bomuo/nNTMOTkKfnCslsCC+erKFOF92JB0pfuDwUVyHqBzsVzc
0QjtIrDXrCFXm4QJ3mMgb5ktwhaoDbg4laC08RRoBkCDIYKtR3Zsv3lkLnrYuSuN+RBJvauEO73E
nFDYguhPVMXOK35jDKvl61GJlGfSd6IFo8jC1nclelZbmBF1WKpcZKrHhWiqzu3A60uahLgBywXi
3roa2g9+JvX8aEbWYE3/8PYLi0sTGB4LOZT1gRw1o3QIHyQVp+X1dJTbaR8+TBCb1SjiLnZ2rwkV
2/M4jbanlwN+FB5dcog4vaGPxR+YlPRdffNbT8gmho8JD9yo6RNjJAk/WPwKsGtLhKFih1JHBfcx
PMFRhDo8vJ26ftuhoKsI5b0qK9go/e0az0p51Eisb15TZPApbiQjuqUxIzWwPOHAOZ/VieeA90fY
i8FNO/JI7TT4es7ciUXQT4FSZ+CCvyYgfTdXUfi4Kk6eM/ZiC//AWy2sN88nxRE/K/ngogy6jD6H
MBUQEBdUY51r8aM+vaheaOtsNCQA5Lw6+/ZP9Vc5mKF57v+wG46rcCCLWTKZ2e0esySQ/QVhAvvS
sdMygA7zr0/olCVXwgzltLm1x14LrZNNM803la6DS1pD6q8GrkFuiKwquy0yOig7o5PDdeC38zrq
0dqxOU/brIU/0CzVeWBlnHbdg2qTyxrwAi+LqK5AzXIOKaqhiSoLTU07jIMaq6vevfZxbdKC+90D
h9hHrmOcdeiy1H4HjRBGas7oj+JTmNCd+EiEAzV94jprjb4fFZ7oQ9ZjMALYbnPkN23zBVNRvipx
EXg4xmlv5nItXICMryqK/bVU+4yH/O5wujjNrPN0dHspurAb3TKg6XcaN7GuWlJcSYvfFRg7AyVy
b0cohRk0bPvoTAFfJ9ZVAi+qeekYsjh+ksDQgFgj4TMXvf9JKIjiIzq0xmhCFbAk8JCvpUERunc3
i8NAzRBWqSuel8e8FLyeb2WXy+ynztqZJq6qMFOZX86seC2o/a5UV6FRsOWeLrmYrdO4aSnq8/bG
cVXG0m+qUuHHlHbjj4rB2NpS2QtiVohvg1Hje0vINHydXHYbGtpePZbiZCumH8ugTF4NFGk9Z5NZ
yrxHtf/1skCN/u4i1Ntip/sjam03KtpZ/cmFPJenbVwD7CbWEIgUXp89/ATS9FGpA58Yw3ihPaMg
Auo0klHdi54xzyhdvV7ndGbk6KfAATcoVfDcZPI1tGkzIQH9fpvrG7VOGSoc8/7sm3Q3i+Dp0n2v
DyIbtat1nWgTc/DPK/ONpEj4f637qP+HAq/rBXimPkybEfhWsBRvYiDCEObMcQImWUGefT6m6Siy
+v6oJ1ohQCzlm/RbHMbA900SiQ4YRaO28C37A1bp2o7G1kyFjcIf1qoPZIMg2M++2jpHeQfZPBbI
TJBs9toDJTVrcP/AKUrO5GHsJ0m5r6ZRebZbDalzVUKI6D/u2QunEd4tpubRwYceoyezPCNPU7Mp
gKMzQUFojbKiSSRo1DO9xbAsNsoFmMbEwCSX6XGUo6bok6jiNcKERtAYTBd8pLMgrcJ9W08wz19l
nnq0ZsK+eESze26umWhbC7PFXqRXv6rNLBml0WVLdd5cCbKZO0Drb61bI89kMv0TiNxDAiGvnswB
9HvvOJAYs5wlYSDSyS+3S6zdr4rFubN9fzP1aoF1gLsGm0NHaSe0p+rPSQR09zM24xgRxJ9Y+N0f
YadjCZhdzLU7YCB1DuPUmOR9F4xTsFrRRy/NPvfI6x13oR/T7dv4oHHOfA6l3MXi6zWBRjXW89Mb
mQpt51soi9+4AR2WbA91eR/VWeKTKRLUKaA8bX4QXMIVoa1oH3Jis6b0kOQwqfToIfbo6DE3QY6c
9wMIdSqwV5VrNWndkdHnVl7n4vnm5JFRCThVnt+8k7GhcAptXwqSZmXk92CjLmom0v1wxOevJE1B
qHiMHmRf1xQJMCF8GwdJpfMzaHwWbA3xmULgwLa+Qw+bMenAQN1bbE3wIWSAzpnNA4yd7ajBBDy3
/Ir9tQWKqZUY1uRw9twpecLS4Jf6U52PLHDYhYk9ef7xQiZ6/SB2w8HMko7kc+knBg/lkuDM1oTG
QWW4cy/bzNw+MojyhQTcFnYoXlh1I92dSD+kBrsw1aCWimPx2//AC/f5v74TaqzO3EgwVVIJ9ktE
uXtxaLjyARspKpXKR7bQOuj1GX7ulY/89mlE6H/RLhN2CRLd5lMw6fVpdv70H2Rv03rgPB040VnF
cr+jbZ5CiTjmkddvjy7z/LFLd9dPr5N8Pj6W1CMWDU0q7GntPSwqPle4yUFRQDbUCH/HUOHwXdOC
RN1hr+G0YnrRd4AhIPs84eSesDbO7eXTwfvpt4F6F97cffxaRbxcZJeoBT1yTSYWkGB5eZMSSqig
lDf77RoptTsytNgKC3TPhdpZUFqKRMsKYwt72slVI02jRTTXI/6LTYQgvTC0YQDaCWSRgF768LU1
2GAUR7bODaDY0bYSyvu58GPlSMjsbDh286AYUfG1lQm/+Pp6xP7iYqS7r/EEkcQWDmp04LAJRHmc
FrHxXKPtFr/3MdSAMgo/vuItJgzyG/knwKNS3LcUAJT4ArT5P7YmTsRMmrmsI9NhhhT/Rk4hMwp3
vO8KM7xdacHU5jGJrNt3G4gkdFG9PbuBnZd+Oe7C5F/BprRfAqLhQf2LjDZ7BMEOWcspTZOtdgGk
N4N0jf27LkaQ0B/VfuKCEQuvvtFKo/SMhdM7kdZqs7hfV0DeB/cn+kUnvhu6dvuDW18W0BVuyVJL
f7Ad0EsU/yQiAaKKZSfhYjj5F7NCQ64Oi3p+bj9qMkg75hXOAUQScm6inRoJ0OJHMnFcx+G2fy4K
atbaXehZQy3ronHUAGrEiTn4/xE7KwVJmFE+Rhx450hq5yixzVj228zXSREdKfw7PrQaJgl5wCpE
347pBrtRQSLg53Hpb1ZkuYxtfZTSK+YHZbtlpM4qr7QKru7WfD+0BPUURqdhnF2nl4JL3ImlMQs+
Cc3Jxuz422eWxhmFgqBwsN5Ij82VcndaE1bpN2aJv7EwZgL13gTuoyU+8AgCVlJJGW5L14sCZvYj
9ThMf8J61ZmKOAwqfxQGM0IqR/+VQVd77WkLPx4VYNbHGbSxNeFjnwyDQUn+r5ToPwnAF62miZ68
2CoavdgepKU1mU0dYBfOTvCQTcVGUx8EY7/+qh2qhWJOWVcsR52IMmkPdzmV9aghWOj9cNUAw8B5
GoS+NkSJ6MMrJYnI7TUCqSj+I4rtj904VZTixoGEsq4ZK+ZawlLgy7SUZHlMGhGmkFE7pPVnEHHg
jOU78Y1yZr0s7A3ZK0Um3rda6LUjmZpizGiZzX6mkcS7rV9rgjhp6uGxiNpWBl1dGEGyH6Qf81ny
9jp254TzOQhuZIbRLU8KaguneWR86XtR30eJ6JfCooxiN4Gb4yNaiXTO+7lUW2cXnTUxMqemOXQj
908+0juu+NwAPxv/LAnQqzekWsTFNQLmGjFnPzKGAvMdK3h0kyrcwKm9lG6ftKKil1hQIe/7Qw1B
NQRo2+H3GA1DOof/uy7PCt41PJo1NPPOb+kwrfsrHKDEUpLzgQpx0YviDTRj5mfZS7f8mh6Q3W0U
PXOHYjQ0MnO2GoWhWJh0g6ll1r2ThbixK+AlUlJD6r4ev2zB2suS2W9MS+jEBG7jvCPvSASEAq00
rC0TOXDwQyjMiOvdFaEc02zUBu3qohwsQs/Bcb6AUuyc4b6zVaDAJPvswP5e9vXpjwWpK1KFTMjk
JncW8wfVt+UwZzGpWWoB+n0ozduwOj+8ZjGFYJUvXVMtUTIvzPNTxHKHmhoM3GGLtllDtAEEzeTs
1IoEHEsRGOd2IdBqGJZphoWCPPPVTDy0I9A5xf/1D0/bS+cnJKxeyPGlqDpn2w2TI7IN+fKyfz3U
8tRncgggnq7BBFxccfixi5aHmANPnNxGoITWBaOJJUX7HAsSgaExne26BHAYwDisvcVthQLF4pYO
KETKKP7ViUxNdwWGRMKHqVHhFDoGu5h2aZ6h2EhEl32DPiKQOx6OGVJGveA4gDhP1MKCBEYRIxcz
SfQPudA2eX1Z15J6ij/1KQs5UrzO7eCPOKKoOG8qorrLNFRVyNfloFRFjpw/0I0lH/ZA06GZcHIm
8k2sW0Cx2sT2B8yb9jGJvupHes/WPmKkdRXHeSM3zwQhDvD9X2ndx856k28aKVDu6fthf+UDlyoV
j7ussnQi7MCZ113xFQE9wu2lmY8SollHqNYz+7DdRi9rsyyTlwjfnORk0aFxSFdyCmBNO0p/uDF7
a49H3UGm8Aiq1WzE6IGbVuLPzXN0gdnBKrn5p0Vw0xVP4NJSID/gbL548i1tyZI5Bmv1NKzpd7jZ
R5K4siq3Phq0H2q3yfTLEjc/ZHxSoiYtSSYq1wlTC+wwnQmjPx6DvsxOWw0jnhzUcF+Ek2ibhXD5
/2sKpqnjDKLhQ+hViznjXoaGHSRZyCNZPL92Zd+AMyUV3xTvdy9bk6FAZt26Di0aT0cGWM/qMni6
mZR5dc9oxtaLQ9BSeEQwctQgu5xSKBEUIuYjvcRcnHCRW7Ih7X5Tk8Mz/s1Rc1Go3ewRl/AdfeRr
wdNQtoY5/qBiPg7aEjeV8YzPQVHuP5F9G56pTiRMNThpHCgOchDw9eAbDi4ezaLDuV5FqxO6zeo2
alt1i3HkOu0Eo/8Y8d+f6cigICvpJ9wU2bu+Xo5ykLDWEsIWWlQlnH15cTJfjpa6k/u2sZ1+Bh6H
LFA+sTy8eXf8503wL26XkdJcupOgRBgoOY/MujT9OKcXcSNqkeHwayqXwXCRzBLBUQb0u2yqaPzp
BQTVybof5e9HKDx9n5dGPtmQa+J5hILULw+zEIYr2uS+4QX2vs8V1t/cO8flsaXsVV5VSnO+/CtG
qQLxGExf+uPSTydYTYVcTHxPkrjyK26fjXEndkpGFMSn18ajtGuX6gnHBrWaXbwisSE6eDHLxiHE
PMEmLxqL8yr52uKE6sqtLJMp2T//qpS4stWObq7zx0NKQ439WsULbQJw3UpiPEw76GtquLZBRjvD
yArs93wkn0nxDnYYn+OJbAqtkwj+IiHpptKXm68QHoic8I2IhP3bCQyCWt0cBTI9VN5BfqpQPzgq
v+MeUNFW/9hdd5oWE206zTfZqQ/MWw77QYJcPr+Y71fY1zinYREEaNIRBE2qE3dRTpIVhJpuq598
iubHg32AIUWmQfORu8rTN2Ce4AUZYe5sgnxCeSPGy8i74rFvKI0CmA8B9aw58rv5hZloF70QZClJ
TenfISaDNtE1powOV7aEjXPKxLeOh6sFM5oonqR5bczo8AimXzAHFt3LxFPhjjGt1Xxoxt5gCpMY
OipIwed2usUS2jjS5M8hvcHHmEG/z+Yzz+z8VuOs3xAiBFW3OtvWZtoXPW6u5fCyX1Rhfr3CDABO
gF4DEzJvOFVLK1Y/jAPgbHfHLceSTjuaHMfNnTso3qCL54LjDS1HgHj1H6K4AIAL3dojEAzWBXY0
oejaJC6ameTxHoRuynppsp7wdOehWbNHGtl8Dd8zjEGcu9lvMiCaIX3at59yGjDi0iUWfQVEqnit
WWVz343BdhMoGuhlhpItK4GuWDKKQORNBMbqhNnPiWKx6jN0/zH+r3mr3jMT1lWnzO/xG05qcdWx
vzGeb/qP8c5SXd1v2xT4teAZ6O3cDjU4ZMQC6zyDj/IuKFUMQQBufs5h0qI9t+z6dXPdGHrDt/IB
SNR5VhCD7XaYmcWRRcNmyhOgUiTaOVxB8JhyQF0NjetpniAgWWkbTO91Igaubnadscct07osYuWP
ceuXMUOlgzM12n4c8CgjNQZqRR8GGa9P/aW8QctkuhMe4wy9/ynT6/O7uvqvCskgyMbj3693wzUx
jfsrq9Y+6IEkhKcTlp1oWBwhudCkNnmySN9JYvKbrP4KeFChSkZR0GEt9Hce/ov9cX1Kmyx8GMqI
r1feobjne2SYtQnqkiEX+WA/ka8WkxzkF+katJ1DSKXbletwSX6KYBOo7ijWCi7us3zvqW1JlBUb
f45WQDdiDz0h9wXXLb3VcAyyuPt42zGtYWzmtQlOT8UsQvptD1y2knF4qjvexawt32WbdL83QKKK
D1HJsac2ahucFV64alNVPJ93XjoZdEePhJpGc2bfT0ahv5dU1Y3+wdVQuTAl8U0fCDxO+opNI7M0
osS0YgCQLivuXGPntMjg/sne0ohZgahLxT061O9PWWUiK06psiEfsiiT5dcz/LL1CRuwbfgNgqNq
j/CaH4Az86q1Xwdlnoo79IBq39GCVaWXG9e3VeM+p8nLJDzWEqJ6BvfefSc695uV+eSHJGLafVVS
cS31vym8zyNefOvBiuF800D8um7Qa/s8Yxq0J1WJ50vrvi8EFsSM0KVJfO8zJwacG7cC0UCy0A0y
xq1vjbHiI1pnKlq33/MppklBVRJ/ivycclzmcvpNmLb4JIse3h8hGX8sn+KkJqqm++G40w2aQ4lq
mO8fsC01qj6at2vJVGJBUKa9PTy2UmstUhuY2mbQeT1oJQxXzQBKsPYt0Go+QBgmW0TDnEZuz/cZ
gUOZ/glZkRiEt7fe2X5bjIIJ5lOBKBLbivObjat0gUE7nHxjfviKqvfmo1y9YI/noTlw0PsRGv9k
Vm6N3He8F86LewDTr8PJPQOvZG7+iG3d8nIgG9vjgK6rA1OOe5PE0K7gRy0nRKpzrOAjeiCpw/5F
YAgVPL3Zv1c5lT9DcZZbEFPXiX355wDG+6k7RsVZcGja2sqT8Ua1ck7cm8Nseik6mGPATIOLvqNz
0tgT0ZoKg7wwrcv6FJNmieXfUeJKJS4463OmbE+ZGLx6Fv46nfsh1ZOb5BmFs4VhrVnKl8Yx0Sml
StfjUJX+Kk4NFipjOW8PcZ5LlqCWRhsaJD+vwuI7gczvAoj2RycJ3Cp0xvaW4DaR24txfy1+tlw8
9y/ptndVfUBlJGNGtsdbqPMQR0ZmFSzPqtnS7ITKdGigNOjuUc9DTSxuV0i+g8DA5U6WWUt22GCO
sKjA46jIsz6mO59OjAmMDib0B1fHjuz2gJCHabfp8HFmk/MJtk+jcv98AXygGXUudRTBsj7E6zr5
Ocz+9Bay+mHnh3hmkceN3SZYJk4T2VWvBd4RPg/xUxechgo+5NKsNNcAVZtd0NnzDrLEItAiypPX
T9fxzEJ4vGds3Xcu4hFFNR/CgBx+gCsU8guPsLY9KLqNlU40ns74gYiBd6WwUNjPKNynP6cnMJzo
rN3ni3hWucUJZJKMwjwycrxKr0Bo7Qg8tfefPkc8j8HeEabVGwLIlXLoJn68Vc5k2qAGSLRa+ZL6
0vJSRghMYANGuk5D9astN/SkWT0Vvy5tAer9gLCRMwKTA3C6/L5h/zaG1tIlJp/ATAXGC/tK/KJ4
E/IAt/sh/ZzpgWqv6XrkYPdBYgip027Xh1onfhDW1bCrTs+VPjDEghijF6sjsOLp1L/0a5cqMOUb
dK3zJCXvMfxRx/rnuh6fuxaXSSPIchgELDrsy3h78glUqQeJ9Mf9+2rLtdCr67YiIQoOifM/ADuF
rBLgpWdyGI0ctSXEpWvsD+ItKQv4mcPwIDQkqVzQ2q8DgPPv3R3yqHb/CnEynGXVrRjZ6vfmwJUw
Qm27p0nEZlv8CqCjH6nEW08Z4kYbKNY9ydpMqGQwDS6MoeiQXyFCRfV7i6dHJJ3hPABHQ2s1YEpY
fKXZYQbn+WGjCxU4bBdaErF+EpNQ1WQMCs5zUZCyU4mgTKPvClqIs4zCfkOYPFKXrz6/VDMus3Ps
X1oFJ8ZHaI/u8bCZLuDGyIbcd2HsykUQgHyAihDst8SJXqSCsUD6U6sbVRrujopqT7ICqm/XxATA
QULpOBRPvFHn4M4Qew9VfXIo2jqQj9HcIhfrrHuA3b2v5AEjgbpJrGymG5kmGGcdtCEjgbyWF4ML
dct2ChQKXcqzq3KIwJz1bUJA7d7hbQgqe4uDemsJ0gnHFozu5Q0TpfEv/kE7XYRBwgGbxecP0ku3
Hd27htDYu5W6Qu3N+/RI/cRUZ9xs6SQL8Gz7Dvt/fA9ZJkJWiNv5FL+99dARC8c0aDQ9jfQIgiV5
RK6LDPTISYJPvRAasIPs3BmrfWYqNCTM3LD/BmObXBBloDiHqRn5yA45Eo6OvnyY8L+uusPjLDYd
HXnUyWkMp3l2HR3SnZr3o+JbXU+s9XbTnLMII4/Wsl/lp8O+3Z6Tob8GrgVInghzm9tLX7mQctO/
mqCfsVcM16PdoKtfTMLqJ0bJjcdBxZAdf3pSlCFTwSJdQn1ks3ajjNhpPJchdXadQR0ooIc7Z3Ho
DfkwWAXE+80SVRE3t1VHpVe6f9+EmUFPlZaEvQFWyCPfXnR5swTUiDjBYLAZn/9iBCqws5GBg3at
QzggpvR++xZTIBwEYSJ7iuHZfvoL5lap1qk876CJ3kxyWfGo7Tts24rQN3mdwaAlBNk6sjK8Gpyu
7OCNq2nFJzPWuCq6lx5p1IkuRi3LP12WyaTVz4u8v3ErjvlOjtOhXvDY5flb7tryBnyvFj2DH0sS
t+v3KnlJWM3ejIy9bFzXvfzbsyOLuUlF5V9jXKFaYwDiPM0T6Zpp85XyuYEFSebNOAfAVXPAASiK
UngUWY94dqUhsM53C5hXLhcswzF536Bdf3vKIi50hHMuZNl85m/4/qBo984SK0k0SE2hT9eKBcDg
nZa4N4V9/7WKQGs838xET/WprrMIOu5daHkSJYNpSzFybeEluA+6OZo1Zi+dgxqltW07lZW+nvYz
/Ap1z25KA/ruKsKHhs/UC4cEeDij7z0Bqvzuuas4s6j/1I/EaKrV+nGZpyB3h+kHIHjQ40P/uK2k
9u7a+i4/Owi6hTcxbOl2gGMlK5n6/YFoyWxnXGI8wphFa+Bl9uLY0RGTawc52005PDbCIuNHGmWn
TEL71aUTj6qcjfjp5NVmF1MWSVqnH4TV/kcTrraXLNbD8ZP5vKCK8Pa1dvGuOHljTnoUTVQ2qDl1
2CXCJ1iMNjIrkd9bDslSv6WoEQ4xbSIoGeudbY9kuq4kpC05unGlsq/B/VnCht6kDrOef2LwvrAj
BsSsqfrPS5NW1WsSZ0vEa34I75JOzrVULM4yQm+5Ld266feuRE3O4ujoNY48T/MmhcKAL9wFCtXM
xhO4iRSnfqGNnaW+QzSOrfu1qvl7QhS4P1A57VTqcYqkGqrUxCGDhI8jImWNdD9TY+kTpck5OFuT
Ne3vCb2c6TkFvKkZXbpRoBWXnVqUcgNPzeMczaXGljydpv/mVpueWECbC9Uo83HeAAA0ldl70FZ9
nuK6O/QVfesCt+IYMHG27KQK6BCYCvVYOv9tdnTZ6V/QYLXYh2rVBHXJ95vmy//tMeUS9v+GwvEk
1vLlQJlVEtdBP4tDOuZW2fbVBmy3CXqRBt0Aw/v6Im4YgzoDlZ9oFdbH+DnveJPMmi8VWsymFzwS
GJj8eyP7H/mIGXD03SiBF3+yFKGqxGZjiHaCrLusOoSBkqR9cx4suTqk03n55/2GD+xZ4ym70Tqi
vzolaIACOJaYxcDObkjchvgnh0G86VzMFOq0QpM1bkr8S29egL2hfnpxr+h7sKY7IOgFojRIog6Q
cEDOnl4iO1hJkcpB6if55Rv94PZjIPEob/kEgO/7fA0tfDei+dG1YN2GOjCFMMPigZaEL5on2YOa
Nf9ay/oUfwW5up9c7RIl9fermXFjRRB04KIh1jcKLuiBCaSaAhhKghOJsd22vSE+wCwJOKgxAJtr
ssndembliamMtnraUWq0VcE60PFMXJF2wYeOcDcYVW1mJw3uXXc2S39J4nGHqbOko1FLZSDuBcXM
dKYPPRJHJQ7H+nPSX7BfO+DOfnHRnFqER+g98o+Do0q9IlNnZRnQO2NeOcVxgxJaAxOTD5E+of9h
tN41mlzM2LaWPEek8j4Do8mRbdCMYbfD0TmbOMhVPHNtoGhu2kYS+ClK4xsUq6hhqNIOsSWfVg5G
TAg7x9rDuIpNHw5EJbedgTF3hdDiADV7nAuQnWLgyX6Goo1NRx6T9QHcBgLhOjL8TzDV64ya7Qmh
iwSm2iAkh2p6OkZgrsLliqCplAN+CDCtC2IPZbHuncUqJsPhTcE08K4zFO8juWxYsHzcIlFLd+SK
IoURCiTLw3D3iATO+LALn7dbK03Rm7YSaQxINzLryBvqm6P5caKVzxhOWNM7M3JFiJQrymT3Z/EC
LBQ4/oizVt4VV7DprsN26xZATz72U3bz/z189nlvdAPIqyR+EEf/8UlBFHPmixQTEH9RjUk0v/hh
t23IjkuIHPafh1TxzO9mQl/4TV/pRoYmn+OXv5vlh8VDbblmropcfvaz5/b6mV6kT3LrKP1o4QHN
pojHgmkf4qaq7HImIsiQEdu/g7qf3oziyAAa8Y7cozN8VoRRKD3VCwjkQGjcB+qaaVPM+cryqLUF
hNKwQ9vOpC/d/2HJUqQkEvfgHgx5r2I++UM2Uo+iMMPVcI81FBleJhw6Nrnn1P/DH0IjYapnyPH6
09p2qITD8JDxUdq6EVtw2jM5MdKSjJDOC3Zy9ZYQOghaALzFeg4u2YfkucudGNmAqWynd+rM0c6B
K0uW7c94FdXn9RqMYt96q7cxh04nlnu9NxoOjvJnw9mO0k64ZiZVTCfT5VtziuC0Ae2vLgRid700
KrD1Qf4sI6HPcrqWc5nE/XNmBzFoyciKfKjOcXwH2dLW5pOe7CcfDyKJ+BjZVBZUDjADE6bJMEDo
61eMrVNH9gcCd/cigcJIcgZvz2tfnXTmFI2kAUQKnFgvXXZWmkNec06WKHIJ7n+QA5syqr7KdveS
j4Lx12/r9sDfkgOJ018Tmh98CwU6PdWu9RMTcHMcE7HdbqEE5JOpw9fy1qfSv/uIDrQL1285YSZg
T7MjNTrA7mDVZISWLwlo4yHwEuGgQBwxDrFfoJ2WuxmOZmpL6kCuu9jGYkPyuoM+NYinQc3NRv5Y
3+wi+GS85V488EX0Gb1OnQYInaxCNMu5G6UMUzxUgVJ+Yk2hkKky2A93w+yAiPN+lJ3ToczVZpZ4
8zxEG7RuQ0s0Sl9N2Mm7N0Haost1YR63/vgrplA4b+j3QdW6WVvV/Eh5hLVY9uyOSMLOffiIO00e
vfO45Lxu2vwNgvxcuEmx9DFyU82j9goYo/0X0YMj/L7AjFIaMmGL4vLR9OqErc4x0x8v7hQrqhWC
knu0hb9Ok3IrhYf2TZAW0H5yhgUkEdhuJTqEK8WmFbbdu5GpGO8Q/b+rtHkKEMZlq0nmItrfa4Z3
bLheATnEYNqFd7o0l8Fq9fTHmBahNE3P4AF7B0xe5gLXKyOU9bTUtbQR7L5j1ae/fkD8wXLTjLBF
jC9q5cUtcBqL0Xcet1RWhxa2ZWZ1xYbg3zs6gmrpMwnqkzFfEctuUhKX96EnBsgEGB2Y6s85/kMK
3kIBNESDZp7F71V+Yq555n6G5boFqbrwmz3reXShSs+YKU7F0II7rUKjXMHEbv7+CAfUWtwsETuv
fw7Cdm6WvhtForyhlX8mtQNP+EncLn1gx1PlrNz2tMVzqKnLB/EC+geXglZWXYNS0O60PXXpia98
4lVDixOFfYuqsvEr/gg1qDF9eFR80IjPo6IdzL3YwoCWU8/QlxW6hVPce0G5r2yw8LMf+JT/RjY2
aUJ5cZxTTfr1MlORYBqeOOA/AfmZhPANbdwySVlurNiGGzn4JfHAL4ZG28AYdP6M0dS3W8hBnZsv
jOj76rvQdo0XFI5gevzC5NiKJew2nNJBXtkBV50gCPcvltsJrCULUuKOYnrTFqySmqvMmqcBis8u
sT0LLILio0z6QE7ga4GFmwjb4kfa0U/D+depfE805BFjJxQZtBSHXs74f4nemhgcUIdup10iVGDs
mUxPd7hIuj3SVEWOhsWo6Vyiocx6jebHD6hxjs+A8iL0adZqb2qA37m9/uK8C5lXnio29GFwf2xO
BJEH/ZnjrGTd3WSau6lKLEaTX0Id6DRKRBzeFbTNEGIub4aXGVf1NBLbaavKqV6r71cVrGDMJQn1
GU85gMu63/uvI10j6h7F8P/se30WvL75O/C9u/JahvHsOkC1Hc3TBsvn04iszaW5J2LZ7Dbcd+VD
P2YQ3AKbilc8vK0xww0jl9G52MzucYEFFFNSMcB1bHboPP8RGAbIdh8lxV6/Byzk2dkPfu562Opy
ETVASBcA+QD+miY/Ji3+ih9zpeNTrsV6c7Rw+Qlaofi6RFGQ3Y9xIPgC+EX3VacqOmiva7iI00xd
qcI//H8O0JJOTQCWUpHBTUUr1FQxE8BdT9oMApU1qugU+vCHa4xDAzWqpXiqa6E7zHCJdddY4C3L
UYPJbfCkXNqAeRvmRB3LrhL7GZR/KFppFkzwElgriAqOg+OwsbJ2PWvqkyrLOk47z4JWbKfiDW6B
0VJOLUurWMBvIotfSaFkx+zIu8q5J6OX0zxwV1aGftCbM/SCPSJO7Ft9MG7A/omT/M5nlBzDkWf8
9zENkW4NIn5HOS1LzRa1ow7sNt7WggnvR9BF74W0tdjFW4Y5koiMbGfAkZ7bz5RoG6bTHrT50U0D
A0oP9QSPOw1CsDOki5ILp4mG282tXTbfq3uaQi4ml3TSJBAicIWkeRMcw1EnMCG4pgk52kTQ9fhO
/IwgtwpkG4QIppOit23jAeZHcSduWZO3gxZgcbLBR1pH1fGoprgAN2N97qKY02OonZFGpW1Z7PGe
mPooaKQpNet+/kbqOkp+A8Qv/ym7SRJ6IUMTLoji0RDMKZuMGLBrkpNv+sCBX1v8/a/CYnt8Xkdx
j23jQ/mbHUUkTMjHK1dDLEoBnMsrpe9pBRO6KvPaAFyBCU2ca6IqIvEg/trA4+miUKobx0gQ1cUI
BwIG3upn5fWgxbMH/oOOhhujjaOODY5L4S/7JLoF/57VlPkkJzrQQG0XDwKjsvCUww/iA/SsdUwN
mhPMPFYNX10xUAXQwgtGcFF+N6yCzx36XlY56w9HnbVfdEd0phqminFpDy8u0w5ijOW/F14R4k6/
WiPoIyILw1pSLzBTQdxdPrt9hM69BN1HYop08EivQed7LhsNVY6wIhnuOxwaZzr5bmR/qLbMaAMj
1x/uNM8H9NTdDATHPLSYrEothXjDpsW+yZDtw3R3VXBYTvFy6SQtdyeHdnKM1O7n2q78n1ttA4MI
NbgM3dnd6XCeblTjMsmLLq6MT0cwBMh3HXqF7hevf4wRl7jtIX1xfn34KE9F82va8a5/aOjvqCuG
lzngRzcTjdOoLWtNyJrbhXKVYIXZBgMINtQwvowYaUquZ8Ri2nQgzs4aLT7FIuD9tinTyQSkKgak
noxPcKpcH50R0vu50HpAJqRWpgkxvdwP7yudpU1h0iahdd1861XaAlqUcu/uEDworG0yn1ocGZLU
rYnrFxniNcYoQqLdDsaBHcDmioym0BgAJdu89Is4opoJDzYBlCb9eCNWsD0rMEh3GMRLcPGKrmTf
uqkEUHowAYV7cXodG1Pnp8qUxCMIvJAx7huHv06iqDZS/J46NMQXYuw7JI62071JISRHCQPiqIOI
0wHeo7tD/nQw3A7ZoTe7g4TRbLimBThyxGwC7eu9+c/Mn0Fhczq0/bFn9s40e7W8Dsg5kjd37TFD
hyDUnkczHKD63VMMAL1axa+gSpWfy3Pkbv37/cxvjrqdnJPJf1VLbZF/xEpQpqEe6RIqc9pXaIHy
9P+Q+9dxKI6khIPbRu4GNROTekiDZrARSM1bsOEwqVHuu6GBz0OZd454fs3wnTFuyMxL5L5fZyVS
5/reNnJs+eC2XRk02mIGI1oxbWN0jkRCOqb7lKU4fLQPqSf845QK9/u5LBlYFNdN7GgrIsoucZ31
NLNK47b1szUcJAvQP5JLyuOwKomWt3Et31YnOaLC6e/EYJM79dAGzvymAz+dh4UHUqJG/NjHS64Z
NEBHP7yQNV6bzpHbnAgqCNLOpg+AG4quDdDcBia9QIA8GqvecXbx+iEuw3u2zvNox7cw3edWwZYb
Cn/ubvoLyHkruV+dyFMmN86TinhTYo8q3s204rftz28tFoaibjE3hoib8MQwib0nF+stJF5YSGqR
pd7+83pKdRxcqy/eSUxDsYxMXL8UhMtDBlqPojlpreDCXe2vxgvJAGfOCtyeKvAdwPn6J0+502RN
rLNRz47i8mszddjdiMjSKeYkR3tMwx8/h4vklErgdd3mvhDEAsnTXBFAVDIcm4C82iG2aVxDBPEG
+VCt6c53g4Aqs/AGuW0e+3/LSs2Md8dXuR2s/hI8+NHNzC4T5K/ywh646Rb+HYJoRXyv0srMe6Ta
8ZqBTLG70Yx3lcV01rF/BhWNK1f4tNoZCW/+NNz80/u6bC/R9lERwi3DokLa/upJ0huuNXaZ+l2Q
HlYkLP32TqQ6HVSpwizfmk6yn1Je1907uWUZX3SwK4AWh2UjVPGmV6W4ohtj5BtBjqVe0tc+dsd0
GGcv4wLo4e0KJ0FJKnImgsozwij2D7W5Oh/zZCj/eXB2fvuFFi/haQaRd/9xdPkWYazm2RrekZ6k
KcvDXYzIe7UyDwP1bD5yYH/3inzzl72XseYNBVGVWRz2fS7+MO5mgWve68JenGFEmCdZY5IjoSOY
aa7ZiTlbcr1ZfemF+a8mKmenHrEUbNmvwuUSAcx8FgJmMGZx17O+B5bSxk4SJK0LfR2yFWYRGXGT
EcTpnE1lN1Nc2E/PfnZaaqtbdsK2Me7c5v2NIsWbXVcI7HdBcFDuKegUIWTsSt7tyo4WBdPYzkFL
fDqI2Ls0I7V0Bff1NUumOHNNaP+wtdeXoEG9sTUW1f9KTqkiTyE+pr11CKTjtEA0V/+v3lV7Cw9N
gWnG2r4++yeiJF0vSxtguN3GAnaSXbCYpt4JimfL5A1EmHCTOgX68U+ns/NHW9E6HQwJ+Q1/1Tbs
hw6En58f/T60iqpD46pcakE0oo1Y652F5s2cdflFQchV27QMajIfrnIR1t+7MJSAbnHbdzKpAHd7
Bdvo3OW7xhTjZQ65qF1Yae5MVak9sXMzXtQU/EqOKDKAM26BR01mt+0yjNhox1i4SsHrwzq4bmLD
zNHW86NP18OW01sdNzFAMR+/E80OaYbgxnfNmu9EDiFmPRHVID8qWYROqUEWZSW7DBRJYgDe1snD
xsitD6olykXC/k6Cb03sorleuEj9TSkaXfzcTVMYwwGcpfemF1DHBFQuG/ATBL72/F8ll63HLU7D
OPg0rwQXH5refZqIqOlAYPD/EbA/rPasfGjfgSSo5jRvovoJO/3jFx6u72KaUK7xfhgH/f1KP/e5
Ej6Ivsg7na4nRHOmMiUxXMcObwYDk4/qFhqF70H4uTEsCtdVDY7QlmHCsBJLQVCn8usUWDEfCfbe
hg1/Xzv0RYGeGfpbtTTUL9CGg/QOegXIiKq41vXjbEgXDW8fY7kDR6WhNH/330CT7rrbf7E4gOo/
zQRlBZRYzfTa8RTloJQoVSKzAMtxUSxhAcSmtT4CPAIPoo0ej7wHXvbiQ0dFSpq7Kp4MKrrmCE3G
Ffndzguri6Vndd1Zvxmu5kbsibeP7l7MSKehdSrOs5gDIBrLeW9xF4EbG0IRBWm/28rs55uhkgu6
r2NXZAIfEyuM2gKhHSbZPi9b/5EKm+YYSfLl+NSlunBdir0FYdl2HfFRsgCg7LT5oAhxT7RNWgBH
L4XB0aGCw2G7lYWeoUJrZZEOGvnBA2dj21j8LCxeNQMCwrFegvyxRP8EP58QldXmHi5SUydC+aj6
q38XkPhqjhmVx/ZOeZCmpBsBttI5gcwdT/KkBK5XyjxT/3Mpy0NqpeFFUPaLl+B+mmuSKzchwF0k
IlN6IRgq13E+f1u6r/pC/Ei+WG1W7C7tTLNvc+QTmaBLLu8YXfrg2LzRhSmYfVTJy3FGOqud2EML
jUMKY7jt3iJNLwywnAFKD5JjMyckRKmjZyeMC2Cz5rpvD3OgCHyn+zP2QzUy16xFdgRUcav0vFdd
iu6rasRkiAeF2lrYVECulwiFpxaBICPSMxNYlJSlXoww+9xtXWhi+OUHbhsYddQqPtHQoONN+NtQ
pjewJBIxy05v+164WkxsmC7hbYKlmhkkq4IqtGriN1ijWhsnVwc9s7txVfZtj9GrUp4Mj5DKYw3O
coBxAwMYPxFLAPuzc5KryGSxfZpq1IJonR52rYApWpMG9nh8ay6LAifjdkInnP9FjEJA6fxYq+yj
Ld4CBBz+SNp13tkY4zyQ9bK1u/1eSJtvUZK0/yTkaqK0xykGFbzk7pM+ilFd/7UMLFjYy3fYPFWy
/OJmDebGr5pmZPqThy+K3yZeaVzzmfpcNsAyXBcgI0QUGYjBz+Sc7dEmrjWRbBCuFnoL5HicmQ4v
3D6DJpvoJPuX1P0dRSgqTmdJ0LcL5L/wq5RnlwcvkDLBZOTkcPBxJeN1L5IgccH3VjKUkFKZyxei
fJ41FRstTsnhRJGoqkL05RaAqylTNJwqpzDiNMlZmqR+VHF3cO/7CUB5AmMQaNY0brmIVASEyFa5
G7IKLXotjPaR/HI7ljNcoonGGdcq4ITo3blZN2f7Kq5yZwdVS6xrYzu2yIQHSWYlWXtPqQzhlu27
HMcO8lFb6IB6QgRNG5r14i84cKDC0RUuxthDJZOCzuXWmSK25yyiGaH1V2qFp+nLkOF28QlR7A/y
wVTfl0FVrzsn++HVbkAa2f/zWMdzCOODKpA6iV1b+Qh/vYS5fHJL2uZHm2aOoQpEz13QGY2p1ItC
2p4A0EzJKyHYLhjvlNX1cydWLfI9WzWr9eOcUn7UFosGqNQMU35a51/axiV0heXi4N+CcM7y1IgT
nOf90uYv/8aY7+DavJxzwQPA8JknnKpv0kFLn84WXkFDRyAUpZ2AOOFD+0IszUtKM2jX8v0Req1t
l1F3GiEDMjp8A0Qc8kn46OA2vaSmfFgzpzQZNnQJZkQ7E4duUU30JFBdLX5vQLF/onKWFydwkoFD
Ro5oAq/nWzFsZ3OC/nszXWLcxs7+O7xRyPaPXBsau+3mcjbolXf85fWaSPwSWGEhPJ24NlgSesSx
y9U7NE/E0S/LMLNNVH8CYZOX8WTyOaZ8mEmvAWiGmmaESaaHOHWblNXX4vTt4WzXPm/opoXTWAEH
vsegmrztXYLekxFsj/Vr/x8SxwArAo3ZAJx9Sn+lZVndxFyoD1/LXeV9SlbJEK3TLs6khAPld8cW
pwZLPbCqXFne4XBlETRqDnpg6JCFDkKAWX5kkgP7cGSBFubt5dP7WaVjzXtY93vScywDpZEHtXUj
e7rZjSVxlPB98NKF6ibLRI9asyhAMJi/EGni6B1qhvqNCHFoDpRb5E1v6xxnLTNym8RY8CIxbwYS
RMO9FfM+DvIDLDcCblVFiXkFyzAaLs58miu9zZ1zz5Fb0UcbN94ygNyMMk0UsILnk0VHyMa51ocR
yU1UKti2eQTrSHZ+ttm2JpqrdAgCzLGCjf0qJT4Ot8OWRGLXlPMq52tcpdk2+FG/WSjpBU2DXZyz
zTM6PdZQ9dBVSSEkg2EKi6hIRmcYXii7SSKBg5tpcj/T7mfkKb7ZcCtmNPcBE6hX104uiVNcZLU5
HKSB5BJJt56sWuOYdbCRkHmtHohFxqw9S9pCdRGHtZCO0zT4VN6IuhJYPjr2FBw4nx9TxurerlVj
1Ub09krTKsuhvQ/t/KAs6nj/rLv8NFnhyOrO7UZE1IWGwS1CtM+Iwwh4Bxk3WbBB052lPlOg0u2n
+C3VWlg0LgIywDYlGVvLDBqnJfxSdXUZH9/lfAhPoEHA9ruW1Mj7xTSLmsC40yiDSZ6VeS7MqEfv
HIo+H4XGDyorkC61AE+TSU9veup5loVRagrqrRvd5lnYX5vt7Gz1z9Gqy9KsRfNAdFXjhIoR5Q4q
2GHErWovzHzn/3zUoDFWxPgmoouVPlDvS0LYTW61bYkaPozvRSJ7g78Qm9fkbMaeLAsavVwJoNHD
zzlcWhiEqyLpA7o1jHP2j3fvSLgPaIcrXOvKtLBumUyK2kDT1OsK62JXRbxM1RVbwfiKlx7DhOSn
xweTWK9+KIcoq885x4ezFO2qTo7tYhqqyNAdeCNiPv1o7u5lv5on48pedrta+yD4mf9tkS3WzEFP
ZatN3fUJfUEQxQgFqQnBfYBPBE3KLODuGwFX7kz06lukukcJpx37CcFmUwMA3PBzaUbYgTmIyJkC
s/prRvscI9sW3DdVtTNdUugHu8ONye7ouEHoOVy0tH95ODzA45VxLxpo8/mc4Nu5x3Go+4alfWWK
meAMzREClNx+j5T9ppgWrCvqNT3uCKc40s9b5QRDtdti7uchSKXNjIZiZfjbqnr23SOvtSuL+yT/
2lXGVd37Kl9SRuqw4XYO5QuvXwHgMG9cMmkggAEGQM/HOsvoNkICtqiTURUR7tlY9FjrqLyKm2Kg
NV2HWczgK19D+pYxn8+097uP1VRb4ULoSyM6LVeZfRYLS1SVU2UblTXIpkGTYMpaX1HF/VFZNs7G
NtJ3EA1oupjpE+n3dXmV+AubrRSpCmoZ29MlmdDCcMCu/ytZRXyBtLErewq1rjgdVMHRcUjuCwXV
85zkIFHt/RSb8dpn7HyS+7F9FwWLD4BjHTRYacPJqxDtjd7GmWvC2aZsl7Utv74zgD/2ZbS5zZKN
dbYpH3oE9mSNFTqxjvHF+B2DmnOmNdSJ7XjBipn1qo8K+rR/e+oTuLqQOiCBUTpMCRxNA3IPyOWP
n5peUXRzpcVQ7lrQO1ewvmY8YS4SkpzQmCtKSluiwjhctObxc792kgyzV39shkUm2jss4CW5oJux
qfBfOGs16FJZQ780aEKw7MklfzuodO5U/ZAiiGJHa1mjE9qmat+PRrBd0ps1ac2Ry+AOarrqR/gB
g2tur67nxQmWjQd2EO2lcPOtIdiW5fdhZk1ePbUfDwscAlekkXc1eOyEF84MQxOt5Nwajo1BXiXx
os647Hqs3PuTPSrCnNCKeRtJ3/25Kf38VhZ4t1YwrGNCxhd+doB01P7Xn1HbSBz/vdR1Dbb+a44J
MgXCuNgc4XYdbrsUcIzF2c3BcWLXgHa9G21GMcHre7r22m2G1ZU/HymcqKSZgi/rUm9+XbbNwAia
ZLs7z9AgHdFTQbIeN8I51UnkVx9o+tw92Pyq0PqcDoJ2aYaDfBigYzglX7F72hTKmqvsm/ypfi0a
9kEMyRGN0XDkKJ0A0f3nWjVy7A/HUENcWC03JxgWSb8tgUx8JYCY62rtTpctCPX4Xv9uvoSLWNkP
+K1WItyPChdssuOJEjcRTTVj1+qSUnUMRB4yGbwhh1yfsLUdcA4K3FTxFzwDYHH9MHNHtWAtqHpv
6JMXxRSXi7c2KMEGwZR7HUZDKQqJPt66UOVzExjCvjQSOjKFBPsf5Qg/rg4+KHOpviYBYwgNwYaY
nLH136YlwzODIJYdNxWyjO8AMmso/RPWcvHJwtZJArKuAZKhA6h0JUUfdVo4n60HU5TI/LoFg0me
qnFOm8PWY94bUfTIsLbHbFfpR7e82qcRmjFsQM6KkaOEEwyBmiqHBNTL0oygvAqJU1ui1EbQzGZM
dJOmvZ8YV0HwiSExsyMae4xg/K1oU2P4G4CiEQCM1wd7C0nsjs+Ibg944K0VDHI8hQeqd1Oo6aX+
wyNkQOVSo+uV1Qci5WbCOpxke3K6ycmReyeVniiu7y9a198gC/Rv0mUcePLct7oMKd8XbSvo4ZDg
jhHOzx5lW122dEn6K66uMO4lSG6RfpIP4vLUFuWvHV/FuFuQ3+AahxFXowAarBgjz95Rx8TYeeoh
/iHA4JGU28hZf+0ERzF1XSHyNnFSRJ2cdH7J7DF92vFwSYdGA/05RzsnMEDQnYVUF3uVuGv0aESS
Oy7cocCdzbpXi9KYc7jYX3pr+V0fkjoJSWzcALyENr+hdLc3D+AlVU0elJOrm3tT+1IhUucIlBTK
zodFkg8M/UDHKcl2wxUNjYUDcFAw3Rg8idH6QrlWvt7XJfmRdvCiM/Jpxxr5sk9YOLMHF6zpM7t8
pwhthsylxFNP/KNC1tXyynfQL+l6hOK2W+FnBEkvldRSRPf+v6J9PCWPMIiUtOX6E4Jb454LgYBt
1UrygWlykJQKBKNIYMSiKNuccUbKaC/Yei6/kncJDftgHnW1NsVIk0zBhS0CsZSWxU4eW1ptDXUK
h3XaqojXUMM/3T8iv+sGTW9OzQicIJDiHj+Z5r3/1rsxxLXEqJ8vsn+4oqSfnZGW7nr/WEc2lAwI
sw9377T7f8bWbeufhKBRfX0Yt4L6mzHdxay6cpy40heFc2XkrdAVmzIPyOGDCZDFQl5dZzmslrSB
4bTPsJn+AK2ia4Q5k02sBWB3iDoIwNSCtzfD5nppH1GtBsokK/MXTS2+JJdUPJQz3bBsRWqvtv6C
J2e1lrhZ+Nm5xbb0XX7O5/rPq3CYsCOkkl9aBLilWVCTjMl61oBSYI0nrB3yvdZBAmf3v3Pwhqqk
47w2N6hMu7FTg6PR/MZBEnYZ7VscP9Y+xdZmijqwSgJYM2f20X9LvSidKN38DygSQpRmR6rGB+YW
Zt7xCxw2DJLqfki3P3KILVLgByb442voLl9j51BF1pszukXNPJlCD+fxkmgzoNFnKOZU9qcX4pPV
+UJ4DMmaNh1iYxCY9Lxu/pvkQvAsGFfFoppxnBGYhWApCVo+O2AnBb7scNQleoRvsMzi3pJ+tz0/
mmu1dFrtPpNLg4QKhqWGLBCcnGzJ+iudGM/oHutLSz+Pv68s0UyFS2kzCuL9g2ftk1jYow5NEOHY
rEB90+14Hf+yywCZ1/hOMNN58C0ZBWkcodW4xZ29z6xsN88Qfb7nQv+ZOzWA3EmLc1VQf2fk5GG6
//2hvnUAQ4sH9bUhLDqAdMZ194gULTOzdz2Gcfn+PZIM2mJX7A5rtnmmGCVYPdDZDK2Nx6KG99F/
Ga4kID9M8VvJFGri9vQiyquD/69RWStQ/CuLSgpHjwMinGEYqq5qxaSXHokC3e5+/3DQoJQGzRcZ
Du+u7kVkxR/ZsBEmR3qjwfZ5zNC9MCJXHbPUyWTNhaWodEY0taJBc37bqQat5F1mvTZd3Ip1LP0z
9BEqWBHxh+6azL8yExuZ4i7/u+pLPk400Ju5AIhQ9nIPogRSjh91x4S3mmwM1Y2LpoyKQM6BFSlm
FXVF7+/PY6hyGGfe6pwYOQaotOtNY0QHbE6Qsu661yLbGrIWhsJbjIBr8SPFZa04Mk0OQbTZRkRp
V9FCqftii+WbgakOrKEM8W6PGMj7TMvoTKPG8UE0msyQ9Qw7KNI4asgmGrzFMSnKZFt1mmJ3RPq8
dWVNcURT7dZlRjWIVKn1HunTRPSyHI9bqx60/0Z3G45MHn64zJDQgLGi/581cMxweo/SlwNgpL1r
EYtH3/aCAAyGfRN1+Q23dITpf5Bi0TuB1TSwFyy737Mzc+GfoEA878p4/dOcyJTkbNDgTOuI5JDV
wqwzVCeBFa6EIEMNImbC5eQxeC3gcbkgzuk+DqxM7vwSl1ltct2uEnp6HAZF50A1k325iVZsUN3h
Ro1F7s7G7ICe9oTcPrKI3dnQ+JDvHYKRBvPc/sC3yHK1Q2rVYGshKe5LAlLe3rWUpSJqA1DCFCd4
4PLjPbmyFZlzaG8AFrh+gEKyfS26NuFYCYHv0RPzW8ZJlPJCKWdUwRaUtq1xq2+ayVxEHjKbqpOC
qhlO4TlJHHdrinBYfvTs7tCr4pP3tzssfFgzpiiI2EKe01Z4wD8nkPxe2ogqtswjnDgQBkT+p839
svxU2mcEQkhu37wzKeeqSnWpS7pFmxYKUzCIjUt91vZC/lROJQ6EiP4B958In00olW2v0R8QWVwb
zz1DpomyeEFWLdj7f+YJ3iW0QzAnt0bUL823X0EqYn850i+cq/Kyf9PfZXqPKwl87Re+EUfyZblV
UrU5PUQzHtELfBBpSavRUud2MfvkxUAIkp7ejubhyw3q+i2r13k+wALSa0xEmIHOwURn5k79POdO
v5iEAqIvOrPofHZg2//sGaOW1p1YusrJrXVAOXeNFfjdO+Gu7MsGTNa4OalQAf/lvyTZFbXNpecH
poOCcbUonn+sg/QWXgwxiclvhaHn3fsCvcSAJocn1nbxwbCv91HkF8vbZsHG2OXkqBX7F0kReN7B
Tb2zhoR7KHtqJWhJRfibIwU7+Ornlgmy6bm9tWZTY2Fa1WIJJzCxVgM9qUaM6qnCa/w7MAnv5ACS
kJizrr0DTbi9+S0MMWeISLgaodSAS3fkZqPha2Q96BbvZTS/zdGLe1c90ymuXFjaQC9Fc5aygSS0
ZmO5LLltQTul9eHBWmAL2zP1ikVgkIZZv/12OrTyll2pgCs5+TVsPIMaKQczZqNo0QBDzd9L/fOp
5J+SrNsV56UBhVKp7d/QTLuzPEZOor7Uxfil/e0LctcyOFRaHkw/QZjGxpDorUyNpYoH4CZ7iOTn
nn990wNa04L4GqM8RNJfE26cLCXw780vGA1YY9+N8G42C6NHj7WbzQe7TUIqufuR8A72dGJ1ZoEB
gCH0V/ZVooSOXUlIcMuqtLKImgCW3fah01vFeS2p7+o+pYagoQqV8b7pK7YtfPfSEvTmgZLtNVXu
5RvMSuPZfcZNBbO59AYjyXIv8NWA8jVm9820Lmu9qu8p6NMKF/n6YCSSDLsgQrGr7+4ROfCqHkOm
jtcM3uNb+FFPzDUmUKHjTIdj119DC226CED7HtYFYJjPJjhoe1zKSj5L0ZPvavQc9hCIyjcbdV4+
sdEDhq0GGiCfQgMjGBLQJAShtdGl0gd7TfsZiBXMIraSTWCD6XbgO4cEs+zXU7qmK+xO0DGocFwc
7ougzXjCXZg65beeXm+5iLl1QMhFJMqai7YQwOmgBwhzPwyyN1CMdWqG7nzP/AMxM9e0UgMAHFT6
Tx3gDw1Q5JpnZTKIdTef+79pZyPx9t2hxQ0eEaksLTQFZMdOY5vihUl4fj89kKe2L2He27h/hiyx
+vTzG23KA3xx6X/lPX3xp5loez+onMWz8k4LoWMOq84qTeBG6C+enGtwG0SWvBhcsSvIX6YdIKw4
YuNGk2Vfei8N3e7PjY7RNBj1UP4O+9t6PbFOrxX8nsLY7VK8lSApkhbOkx9oEQjVJcqV/crTyYtg
DKa0v/qiFkv90dZeOn0Phi5pMUvB0Dz/hNvJEtEBqBTjttihMzUvBa5b14KkZ0Fli4SbypCtY+cP
rBWkJDquUVzAWwwfHm79X64eJ+fEJD4Pb1OAbNWc9eOLTzXbju2yp2Y+8NlwEgEQvv3rnanCxttw
y2ixN6Oh6mx9FUMKqjibppczHt6YQMWXyijHZVIfLnGUj23wNqnsHJrKewUWtpl8A27wmoM2m1bO
Div6Ls1SugI5TwTUYmhbBDVOan9luZKzZLQJLhyGKD+GXvfKiJAhvMGHNoLOOxg/nAyoJb3aLaf4
kb3LHg6m/1VPXWcqkCxpHzHk+a5nZ0ftMVO2vI13nAsW7Rgf3nzDaNoj8J8qBCHE750yp1bYHO3f
6OogWzqRdRmAyn2u1poqN46FsOutkMu2+jzKTeR4LxlQ3YUZIuRsrDmBnZm7aKTm0ut74K/TIFQ+
dmUP+ChZ4IWEv9NpbXfhLa5nY9nwHrXBav5jlS+9Fy/FqObKZ2G2ngkOjqiafIkHMGtUpwvuHm0d
Q2iEItsEycgMkLkbGNcDPQS0PilVK3/6v1pGgMk+rQLz4NxCc970emtmiilstyHYAHMZSJqa/oCw
jCFeBmd8iHlRtsOZZ1w2goI1803r5CElnuomcGrQlZI3gNsvbQaH+N5qDBw7TdViys27eZAJNjA9
NzBxfcb8ux0/TNFmhknrEZ0XAm6lkvs0UFlZZsh42Xb5a/b3lKphlGM03ZSMhp0/bCaGRMEdIj7e
sczRvR32tNfwNqc5jguhmuCymKDMETqaNhA8R7pI6gHErk49xr5E8IpIxY0WrCU4nCWbiDuMYWOu
GOjR2I73GSd+s0yORZs32W0McuWPum6rFXkcztzFBkNboujZAeV6lE6pahDVQwD2bBMJzCVD/RZS
tlECmQcbfVzEKw0SMWXdjA0BXyyxj0mhgI9hqKW47HlfxLJgjacYPUEkJoOh0uaLEMFPTUJ+q5r4
5wS7KP/sHaOkDRGUcTfv6BZOsGoEKkzRj5bgsiFd+Mn9RgglW0YaQF/KBOnq+OK3ROLY1vq3DXvu
0BCAxQWbOcZHRcCHmmAwQrWNnTPHBboexLk+U/Zrf5rNyipqpg7Gtx5Z6eEXYmu05gKLhb5SWL9q
z/mvEUPdAZqr41ZtdLNCsHJWzJFLP3kplW/XsyRSzCR7Ki2Y2vPD0HcxW2dTvNA1MEI/8Oh190Of
MXUBoLda0tIHB9w1itEC7l2GHD0J/GFDNA8mLc45F361afKRYsbW/jWRjyBodt16D5pJiJ1oK3BW
fLNNLB8pkwA7OuCWLa4GMzmz22OR1KIfwVt3f96D4ZcvQ4HhOe2kGoTsPSzqRc2+GDALiyFG60Nh
bCUmtgKMGica+353ZEH/RhRNd/ey+TV0LIpoNM+D6DOhqtXfU/cF4D9+OUTU8SWJNfd5tv3xxzz7
iGcf7udfbrkckAjpe1m95hTaGl2fWXSzhxed1QVmHgP6mDjxwD1M1o3zI61itVH3uiQcRWwNqOOf
y2Y2S4WBT3PfcS6gjdNjy0PHOHiCGDy5BQjBmIfGfSth1+ONNpRXJJ/nQFvO3g2nabeWx+McsUu3
hDbS5u1N0SfU0wnWIWb+y+uzeyymscczai9XOlIMJZKW8pEOj7N5f2SpZZgA7htuNpTECTIkiAQA
NoCb/VJ7ee9a6dY6oMaUTyEdpILlnnLfP8UvtwOtV+dwxbSNspEAeY+H5qaya6bSZNP20kzSTO0r
+ig9ygK8YWUwNOBC6wV3BJeKCXy8ij1f5GGzQ04UKdj7CP2q2ff0hh+RVtvvnfQm6BvW11OuUSQx
K+FKcMamG7qO55ftbj3ILFFN+yz7ncFjra/oDPve4IQ2FZhUScb8JOzzjbAviFqlIcNJZwpU+9Zc
ybYHuQeff2HpA2MMe7YHxfd32nsFKvISW4FSOYBZ3xdWzhtfNCHcbvlKJfaOfDwYiWQt4CoROd2C
+YBv0/rb9FqTzSpARCI1rR6eIdAPHdQGeKEc+dhqbjzXhpNNX3+9+55wT0/kXaVJi9XFDfTI77m5
ixZub/Xk2I1hXaVwz8HPY+2G60W0oUdCE6zcTEHRo/0tsIUegNHUd4NCA2S5RvJo8l137Gl36N6M
PVMEK6eo0KsPr18ddVnjgQuQq3iQ9LHRTnHXwzK/FevGQfZNGoh+NzuGZLRnGLB4GQCA7psMe4/c
WXsv96bKkU+AD5up+gT4QKRykDzA8sHSoNMGgrVXzI3ux4OQ31BBgBeJuUQfMwtWH8qQWYvVLyFU
MC9887NYN7YdPCBhWbZwKPNpmeySAPtYwuST5dUAa84EkCY86z7GKcPFWkcWTmuqcW9jJYmN5Fae
SUVzyd56klcOPId2enMrJ4Mq/UTXzgGle9mC1cusJq40qgjmwg7htJePugFpFrk7HKfc0En2Yj6e
yT2Kd6QHDcTpOOpQzaD0V6EV3NV6787rbZrt4YGFUKTOZRZtCrs/pOGdEn6UxzGFPbvxKyTNR8YR
9Wny5cn+1CVC0HuH6S3a2kjBJGkMoDgsJKW0HeqF9PFhjQNPOCn7ufddEotAfdg9fqa1IXFeX09z
oeGR/R6fxJNPcp7gqc9dBuG1z2csWET0xf+UvU2jPBDR3m4Hfv2fV1ONHRl3UGaBofGt6M6HDR6f
t8zcM78N50b29o7IhZhSWqWH+GBivdHLiTYppQ9f2he+0FFEHcQ+v1bR0YUPAR6AeCDN5FdmeTWF
vxvDLQ6ICjRjUfr4RXgycLlc6Mpxdr1IfeMJrxIW69Df3/VncstWnGHnpwkZSM1FHv023yBPxK2d
AvHOpgtY1E9cp89EVI5hyPdTzM3jLoCg88IK+kSlssEZLjS5WaQp2ukKkqwANPaslUmaIqQFbXMD
R5SUT6ypNger2MvU1V1uPzcxb77MiEnirqCv1gRJ/WF1FNLSzfPYWzRY25ZxQrdqzDN1vKO7WVjy
/JwhjCuq6bZTUSetNwZGjjc4exI+v7BQ3ESKbNYe7CPf8n+6F0LRk5nugKHmQHm6LZVWXdhZNFln
vZwLozTC9L80laPlaQY9HQIwlVkmCyE9Nui1uctit1prenyRuZ5uyjj4C6aRJzJXTFvmGkVnC5Xe
hUvI/l9Huz8U+PuwUCWKlJYFvZbv7KnI2kc/iHMc0cgSI3sX79hjKzeTnU1cHJ+IygOgrwb7kmJK
LokUwMoFY7anEOUp+t0QsVCbVdnO1u1Xd7uXsqXXu9ZPDIxEkqFtqr7jxo+InniKL/cjxMrQTX0L
3UNF1W7vBxAaD/Ko5iecj+2xMrTILxc6aiTLzmM7+zrzLzVlM1yDYkeuoXyvX8DAAp/YR4Lo13rq
hodTgKnToYXw5OC/x+c+KoenK9IaaCl22NG6VwhgnRjTSxPd2etM+UCOohhDC6UKuioIWokoTCIf
BlJnsQ2UdAuAD/FhVxbV1P2wl/qhAGjWRXSYc/9avNTPi7u1itchIDbxcicmPqFI5VRAnPj+gL4B
i9GgJHK4QelFr/nlU0JGUBAukUBU9Co5tetdA255+2kewHvhwXiwInDHubtyvvAvbnGpqh9GVZdy
A/x2cfaEgGMpVUYt49c6x6lK3zjSzsWIwltR+Py/qCJ4AafrdW3ZvF0xqKGPkTvvMCY0CqfgV7cD
MM52b5VMpWMpked7notAtnV/dA5Glut09ZmkIVDXY4ty3qmpQ5xh83OnTOEbXsYfjie0tmRJQy7p
syfnyiCM+JFarlc/FBEaFbPxnX1hUTc29qRn7ZECza4c5T3iZJ/S8+7dTjVEimLGddjZyxozbtci
dY/lH3NeigoXcDBxImUDDZLqQjP2uZXtXx7GAOjPdGpg7zW5VnM0IPP5xbvLpgT3y7qLWRzYgHHC
S13QBef8Bwo2btHHWTGNUuREXpOotjRg6IWK/f6fS7lMlpoPT6qcx91PW7HcbOQPdwMMj19W0c8z
QOQV5S5wla/Uek+NaVHAklAlqOFr6BekLiej8NrMeB3XRTlUG4NfZyLhk09vwBmdjEZu1JJCYwiL
R0RsoEm9Qm6ICL1jJMmGdZaTGRsZauDC9lXsQLSsfD/YFXkJjjIVR+h2ytUu9uJ9jmd2Imz8sqjh
me1CAWVHNZjFgeWIBIO5vFpJjSDpCCK1NwINQZv0v9w+UzTSoby5oNmfGVgxDMXBRpKFv5W4mpj/
ih/U66XHZhPIT/wlI1a/TFHbfhUhe9fK+ChMKomeo5c9PkVKMSwMvTFbcBh82WK3XB/Da2TR0jR3
Mc2+V51M2pTxxVQZPxbcPB3ltWecSyZH4UBmwMVldDHF5Hrhe75fgiT6ozs/yJfS2pa8p1xYmV4k
tMb0vORjSSTpqtCNrNjcN5CfQLFu+wZ8/QJPbCw5k1mQbY1plXn3T9B52nNKHnry55CAGnPWvQUi
FSun7JW88jwWQmlEK9RBOLiWE1pVrYpTe9FxIi3bjpVeZx90un3CacXpJrfARqlbRRLLBZciXymS
QsNlzCdrQxQDEtCBTRZazcWtEahyiThKHc3piOlGVjByyfigzbocLOtUW1HaN+JQLnw32ZgtGZBd
IBNKl+Yh26s6PzBTsQZ4e1ZBVe4grmuNre/xk2paxndodKkfGzdMXMlbE+G1z+FawkWWhuXXQIlh
cw/BgZZlsSOL5Hq6WOmdvuzCmIqG8C9vVEdVktx+wCh3RYmLibbBLroDgi0EyHYhlCiJL8HrL9Kz
LnaMgphIGgPuhN4EBASNInzMh3en5ryiN5N18Yp++L2AE13O3Rq3A7WX5/ovaNFLPsyqzLufOezW
n83jqYH9ExOUY9v9CMjl/Wl/KaRL75g9Hix54jMGiYqh7UXTv0nyF7BPX+M/vHCCXQgxe5us+wL7
tHsA8VAu0IUd7WMQDtkLL2r4wyX7DuXJQuI7Bqj5pLBJ4zW+qA+xjQVSXz3Y68Ab8jb5aKEoThgl
+pCRJWEWsQ2GeCBimMoWncev+4f9C/fx+0w6lIB2O66xcuk6cnn6Fd5OZ61Gmwha/Tjlk1LObodP
isertjrKQiwduEY8sWIpvpbkmBc2mGz/sMaOuxiQhdbDyGNa7XIttgURZuKFI0Kc5rR9N9R4b0ZQ
qvEA/LwNRF0MOHSw9Yqzdj1LjNf1F5U/XdpjVXPMdfW2fQngurLXksDqJdSM4iYfnlvwdBvZVxM8
Ritjfdq2v05zx/JKnMz04lCG3pR7ZVIIa11fggIWbhMpk9EGc2OBk/ZxHRhVUrPhDbGzrPSqsUY+
p4xfr8QyKoTs6syxc3st5zJ8b6txmvaXrbd/wT5qDJilU2nZTYUwfeYBCL6F7RYre+xp/yU6KC6u
Y3HuFSwx/NFyIW/I+t/Wm10rhhZotZsFzrftOVW2VyfDWAKN1bVXs0Z83+tbWefmOX9oTHU43+H7
7t8fUumkhFze3l2m99vqkjS5+cejcMC03bg6rKI7cfGWamUVl+V6UFDM5vDe6nPolw5z72ReK0A0
VfHKEWEKJBdsaZPnzyJbp5nO9f9YHWOnWCJCNgCki6hJ734mZaCc4k2AnswZOVo/jOcUsAW8vVWe
1QWT4oC1tLtHcExRZaMS1CYTH8v+S7yTdjCKP7Ag0geW6Jubor2va3Ksvr6QZMrRHFQR4fMCi21U
nOKdfT1HuZLj9jjgh8uMUofU0FrrmTBVLZq8mGUhlEf/AA3ErQjG82kfaLGCTu068JbBsXoa03sM
IxLTXRyYObYkRn+Kfd+0RYIDBQ/RDlt/regsNHGNkIOmOG/f5RVauJCONn6Le44w0ZGahCbfI5rT
sK3Q/c6DVG1k1f2ArQd2QkMiWlXcUuAP2r68FhCDkJ1Jmlu+5DJX7/7bxDi/xsXPq9QEDPD2oxkX
WdYC1m5FbY/Joz7ZxUTBMU222AnW23S+VtXESIBTD6WiArpWAq0JrjgZetOJMHT/5BWVDhsE/gKu
j2nioWuDRbFt4LzdeVr+a35lP1xbdHNyqwdIXmbRwuRfC3juByHWGNABgdYJPzCloBMcPjuTZg7a
YUIS/BwnwAb6ZRxuDJBTIVOTineT+UicMNgqviitd0rFZZH/fttFXaGdl8Es/v347rZmsnyse50A
CsaYSJIQAEZfBSAhWF+Trnq3Ez7Ymh7XI1pHKoag9b9QjaIP71hXBwB2S3NqiqksZBFwfg6ztrVK
keYXOPeI6pOBnnRHRGVkRsB6SSeHuJoVw5kGAoVkbwzhpZt7Nofr6hSL9fO2PzecRDDQ6n6G+Oo0
FK3b5CWSaso7pMCjkDd6Ts7/lh9g7BIOClntkR2k+pr6QkndhD+tbKo00yl9r7X4uGk6Mrx15pBy
OSwLZcyc9za6Q2fjmdjRyeCUAOPyXstbrTkCrilQoUVGROZI6XQpQlpLyonXApWfnyALAGll47sf
vl9Hx9AAhtywsWgc4ghQJiVMUSrimwPetLALJk7JOEd25RzL2n/M0YEB3tM0Ao6fwYDZrbSMXWPF
K7loplD6TJq6s/FnFq6tYk0xYRoRc3Pkz5id2V4krPQFinLftgQw5JJzcQF+depp5WC10c6PZ8bi
lRHXI3tZr8YMrHjYxKNVP4z/fY1FJi2qcwkt0RYhymEifuIXJQBC+wQdXLUhOId6b9bGmHZGjl5F
xlXWjhlnUh8c6m7YJSdsTaWNZ3BnisoWxZdO4jPuHlJ84LYSVsV5YC+fXc5/wVJgvLWQ88b5hmJy
6+2MbFgsXWD1s1/sQ+tiZeFZBmdgCotvTaawaNcqcSCuRSYDT/z8Z8W65IOeAycKW7d/pvhiEo8+
ng0SyXgcQTKfjGAlQqfLSBpQDpBgfdIUOnAcCFRDgdtwJUgmYS38NcaafxV/1S+xJOJXOVznWuDJ
qgXPicDmFmoDD27cyCcIDyNweI77TmkvDHYcpAzVCsG6lSW2eKLP/6pzKTJFAfs5Qus4kaAsshSP
2F/1T8/5U5vECBxEFYrUwEHX0xcF7U64/U7PJ9oQsIHqXdqYmM7huxfLVKRIa/iyxhJOfpSs0yp0
SKlkZ3u3FAgxEq0Eh/C1l77KZmQcMqSYb/gI9c4gmrlS4NB61vEMkrHUZ1xyv3esp8hM1Gmq+ghI
YH43kngNQ5KEA5b16yG50qhZVSM8iD0feGdKOQZnAQeKyA7jK74ijlu+zeJgbnNNtxdhiGcEkpsy
iUSBCo+4mrsE/uVgrC7oKed9UbuuOkFCX10eXrUUAbHReYdGVxB07YCYsNvfn6FJH9woCsTwHTen
4yVrGnl0J7BOuKgbfalgijw8SGdO+ll99dXkU8CEFhsnZdR/MmjxzOQBe8UdmC+uFgXeMGwW878P
tUb/bGgtkfMFvI8aMbGyarmwYnCdF2b7NvsQ/3/4gMpdzN8Bl995LE1Mq9c1imVXTVdb8QsgePbv
LpPqYfyB0/3bjZsLd3g1e6ShTr2Q68lZUGNOagsMx4BRvgiv714G/7NodiGdRYA7p3z5/eAq8vin
pruNznoqSEp85XkY8tNongZfK43un4faeOGXzwwMxmuMBl3LE8UP4Xnk7sXgz+VJmNTxRecncDAQ
/g2MfOjQ/segoiTyjCDGpWhPJrGoLLIL6vvsQkXMLY1v+X9vr/d5f4bzOhqfg9+JUDNnP2eMovXY
CeLKoXfLu96L//L8fpWSP6Z6z1VaKmKHlNwZUHLIDfoFCMAxykpWORQ3eL0w2delbQkr15eGLN7F
J0viqqgsVARmL8i5DHdKJOWlehZR/89mwPG+oj0d4d1BEJ1oeNDlqRfDUKf6RMTSQ9P22CMjhI3u
kBqvSwr60tYOhQS7zGBCu+aYQbxZDY5bv6DtRL7uVhskIsGLlxixTNx/mABUu08YXCxz++RV9It2
PSqiQPLGxCcJ0DTpQ9CRbmaqSaO2UDInJmaqWsT/J0+cUkSwGIAAe8/loVM6BOS6XCsCUVg+HtU9
d4ipZnXWlwtZGhOn7UNBstc7S1lVGSnnTFkFa2EbXUHaogi4p5/1876uYavf2TsBzXFHqCsYBMT6
OLNmMxvVnm80nVof85HpLJ4lIyWLslpWwGWTBUnGxrkvEGO9gSAyA3afeb3Y02Kh+vOoRMRwaH7L
/BU5RhsT+tdbqqN3yh51DwcA6JViL2cC//WDW2yir+I2P3k9CRhg2BVnLDDHqmmQ1xJ9p7MIpQbO
RfmfHkRe2d5s/Z6IcmSxWzTz98a4rKVwiEXyZYjra/eEkXM8x2xUpnYb5VnlJJCkwQpTmnvm6f02
30vMHN4MK0fat1yxAeUAO5CoE5G4I2sQ5uQd1H6tURdip8qMcRkykqvLGzms0/e+G6/9qyovzrFL
ufN6l9Hn47ZtPkqRnXt9tn1rsNRkq3b7DO9MuPrgLdXkidT77ke5btNJ51XGl7hRsChay3aH1W7E
fLeTwifycN/msBdjQgvLN2QAomoanlEK2LgHVw+TxIRd1mz1sCqe0hKBo8pFdJz2e/3iV8Won/dY
Ybxn2i+43XvWxba4OGD5/waoBvtIn1XmfYUUmxqmfM7J1HF/O20RONuG0+mXJa1Uy9YgjosFzV/J
Fw+yVZy2N8l2WeunHgcQvJd7Z8ikAZ4bA4ZKaQ2Y/v3p6UGfzSFH52+vCV9v30bsZ9y52mS1vwwG
g2EdhmLNAPxyCchvBF/s04la1F7eHp15qTSqbcnHXr5KrC+ybGP64TZX9kWkeOU2lgBTwwKSfoFA
KX+mT3yEtBr3flh7n0Z+5uqLVb40ULVYi2CUAv8yczUQCn3I8AAbpbfeo/uNdHmlzxLOm5S8j7Tf
IVP0nGUTHrCi4mAhinpeYFmwnS8O3YgIwZYLlUkG7yFzJH4XBqpP1kN5Q6/Id02hagzfI0v1H0w4
xjvBSCVZEkD18UY20CFeeuTBzn5fqdXj2GpOO47SQLIhM45Wa+3eW3qSchhsm8FhUNWZWVCErazG
OJvvq+Vc6QLurO96zLiu3pGzvWRpWfaD/I7CQO2HrljdEdORx98suEFyWh4opZbjvqb/x8EaEPDe
s0l3DYmwSIcLV6/PkblHe82GxNJl56mN9pxdXlJVjMzt4EPhDYYpxjptxRIGSfnpdCsF50CNp3xY
dOVkeR+j+AOjwD3spZXqLZIjfvO65tFt+st5MWvbUapLcYpbHNv+yJpwCGPbYXQ48hWeL791FWOn
Q+iUO4F9CDRCPcshWxaBzTRsb+Y7PHPF3v1gNE1ca+wEwPVD9YuXw/gcuGyM4o7aEOVbDUANbDRl
hctngH/FEoG6e79iy2nZQ9S5MXxP5jNoMnwbopMKWp95Ep+BRwwhXiTYvbWI3RyeBOg6qCJCAD3q
pfYxW5VztmekJbaU+bAkH21rgIFawZGXBtQKJLbCoK8yWhRTa2QOrb7Tr5s7NidDwMLKTpHH2tuU
8bfMvxVIm0/tkuHEe1Wm5RF17S2Yyb33tCv3p+I1nqFTxRmozQBfFIkgD2WLy56e1qgVasbOEjk1
e4IiElGBJDT8iXR8vaEcOYrCLCtiLq2AmyXK9AvVgI/D6C+MngU//sF19jCaYoYMqNfhT0G3dzlP
Q5/Byt1JLBHXjnoDKgkeFWjndMti3NhZhZGjo7pcjGjoN2bIqVs61PcSNU3kJ1dirBFKmYz92+e9
2+DfB5Ulott6Yzy4TUgbQw4C4vMAzxLFkKhtTBy+hm7MQ5ujYa7FLpYGZ4TXTOIaX7cMKQT4/67s
+wEu6/5IpcavjKt+rwJasFnDoYuLPjwEgGIUw+30T6z0VlX4B8MjyvZeHCPoDIfmBYPRT8mC1bTm
sMomsNo9zVFj4JYZKvGyKzckghYYSGR5YctDH93NANruEJNDNYkLlGDyRKbuF0GZr70825fm5OSX
8dY8y6R/w6dVrg0cTeJqBuU27mBuzPReHd51q2Hp/p7m4GwJp+TnCvCMVc3QfqsHocv75nmV0+eg
+aXVaRZamBCO/02cOXyBdQBjbxHd+/RSsPf1/C4leukvbLlXK6wiRlppZ1LHfbVCsU0gPZY7PZrJ
CI7rvA75/8temkQjs3SnDrIBiz3O4Ko7laiyF9ckq0yUtBMvqefvEoxoLmy1dfipOlS6SgHDIwGH
HrUb1Mhq9nkv6Q077SxqyJ7s/+2x3V4/zvdAVpOR/wM8OpWmNSPodkD3KRzkUVwQP9TawcTSU8AN
uQHjNqXrW9zsq90YMPolUNcCAsxJFnqTVdb0mddyrc1yOVu4LSPTCWc+oOZPwIQDO5n13OJQp0MO
ped136wObjB+CXDuswZ9+RzWenMSAXlP2Lvhx9ZHvg8cQyGKlI+V073wblRWkkG8StCjgM8wbzgU
njix3S5PTrPKP8A+ZF5hB7qE0co14zbw2dV+pN7WZHNshyB9Kq77wBhEcNiBT+xQFYIr85inX6Su
dTGKRoFxvq6o6JTnlD7M58VBuOy/QY3SAH7MkdQbEyCeX9nzjBvCwdWCeDLX1Nc/fsURU7nTr1nd
KA4JnEartX1soB4eemctZ1kRNhrSyJLi2D264VSrVVBiwfXzzg8X0//bxhNmyHDDFi2E706kF51A
jXL5q7nDmpLNGvNbnNCkgoLriJwUSz8hpUXO3bDtdHCwK/AFoOnzsIZu1tRCaAtYqzueEkZ7mR3D
HU7Jz0bSv8ehj/RrIKASYzCtrblAwyFu56E2tEApIF0o+VC4p8vonx6/mjmhvXiPR9zzYYOsBXr8
HXNT1bObPE+RqEgD/Xx0VbJ0mg5aC81Pc4pKbmdlWWwp1IuUqgCrY4lyYWZpL0TVqIkCzS1Nq0jp
fECfCuxAXJhKbdbliddxKxJQltosEkRtbp7OVwbh9ePtQm63XF1BpiqPMvAiGgBUXnGhz2Oumc+U
Hec2YKLney+HINksoFF8X4e042P5hOleNkNIedUHQj5dp2W+iyVuG1+H1l7glrvFZB3SXipQ0Mta
3UsUCxY/7voQT6dunxXrftKORN4KjMwT00T/lqO40QeylJoqWv6l+cgoFxqRB0Uk+eoeuXixdQyP
0+1hIiRD6tfjrxC8wyFKMfGJBSQDKa01Rfyz2GSk1CfC+Qdb0baUY25ww9jnsTxqUcxOP9ZSWr/i
qqtKkzWuzPmWmYw3rYRe1Kop4UtAOktEMzQkEHVOy0Ly6UvEaQw+m0qsdVP7TnEeVueP9voZ8EoJ
rcKDSpEL3hxJD4gpIexfxbXCtc1mdvgQhpJiagMIucUyUFbC0rRVRF5lixoziggPDv0H9qJFlHbe
1iZ8Dn+zFUbGV7tjfgV2/nGHJhbSNgw5fmtTSXHAfSaPP08ursg6ecT1FiWkrRIfjDPufM3okTjs
ag51C1UzLKakmN4XUj3kZSeI13S3Y4ehTI01R5GOr0XLuAyNms2QPkgZm2FaZ/baMoBFpI2XvjCP
FQBSyOqyQmSp6SlZglOkuLE816sO5B5Vj2ZtByEjKve87jZ4d1GWe4waj1PUD1V/I9z7excpBP24
JcmPOJYvQlrD/6ii5YgQ+aUGQehoyis7jYl8+bj86nh66Doun1oCUJdfSgXnOWIFnJgCZBxjng+7
oCfDVKGnVqxbMGdDIv6cT1VAyTw98W4snHzzDL3dTM8EOsyzaswM9D7z8miFH6u9wtDHB/y4D7/k
Q8IRH984og6W/m8bo5/bqIFyqewgm9PiPJMvWSfCqfUnFJ/KYnUEfa7ejKtwLq8pn+tEPParMa+Q
AvieVUbvwTtIaXQ2jnwD9S3gabhVpL9gfd9f5qysMb/9YIl0TIrsFuof4qCAa301Ky3qJuAJhbtP
7ShClRwa1k24GZ2QVKb9HkIlld86JtLfUP62ZozVGCmbGL4iS6m15y4sMHyJO1nagNYthThrUs+h
WAPtm7NIcs+Ll0Rus4QUblgdyAsZtAUmerYi9oUHdsXTmbmhqGMZoylaj0sOtn2KMMENCP6rFjN9
ok2dIdD5f72NBojc4zEd8svw/qBR6ZN57kHi/QUQIIQ4UWQMVQ26NpO1Yd8tl+/MqAu+pBR+ntZx
4ByBA/HKZwFBPIapKB/Gc7/br2trSsLtT0mJd6Q+pNiuzbL2hRoNyRb7PoDdR76VXIS08XDeTWbh
QGeG2OwzVCzDPgRga83C9VGo5DYJZsTWCvBebloh6c6R/8ypZ0tEgVvxDeOk0BiRhiF4pyoA1TBt
GPL6TjNCueiy3Oa1Jo3eSgSs0NBB+SQlr9URIC26cJ/7HAbWL1jXKz65L81vQ+8Ns+c0cfJDthBx
vIdDZ3jQCJp3dUPulI35cQ9O1GRPg8ifFzYsBmbYLYNKFliQakwpmHYfmwpSKvr9jvNDBOP3EHji
TPzwPJKKt+lFhzWpWaS9KCGIWPpxmKe0anWb0/OVX5/K31S/obq/7CpZk88LQU/90pZZedYkcvDO
Vx2EjjcSmGp3SC/oM3GxTr0JkecRgSpFYf2ZVuX/aMjIu8R0v/Qd6QLiJrqRHdd40VsneTUEOtrH
V6O5Nx0fcMUw9XBQl61OXg/P70FOyEPNGccpEOp0A055looqaZbuaVG5zRjvnnM/pTeUHzscnB/i
F/sgX9ZOWDM4kPC3+Jqk0hi8DMHEfj4G97EQGLpV24ebsllnpuWDXU3VVb4ZDLi1Y9npQ+iBqsZx
RxzwvpHUKiufHv40803rpLCe7A7ZJOE9NcojbdYFNdmYBkm/l0jySUSqQBNhejOjVc+qqQBPFfyX
SOniGgZm4gt/3Adcya219u9iAgveikErPb80vG8I/G8VY382jNw57aSg+HkWOxUF8UFNajsu6o7j
HUq3ihzXJJIN31Urqu+zEOvLHV50Pa8Vc0cL9tgvBNnFEf7s3mCxXGkndEjPU39sIxDc8nxvPGsX
4xUA/oBaKQR8vaokKprQLhDbP3igwn1qAI+ON1C2r5ADz4OMHYhRCGQVSrZ4m7qaDh5pg+O/pp/1
eVZSlXc3OZHbFaxbJ5I5yRRZLj4eleD9DY62b4r62e6tk0vy4MpOH77g/HlXHNvD+aI2YReYmrvh
yyVSOtjUHHv37iDsso3iup5Er2R2fk6QBg+Wu9YSLMAa6v6tHYkSQXb/iiKo/QP/wucrSa0fl3bY
zDOhu+GjGaFVtKiiie25x4eM/YBVu3IesHtIt/Ql94Jc6ImxiuHiXnFKybor61u/vtydOYffWBd4
GPTAR+j29AtzotrkmkLxlDsE6F4beUAucFsA62lQwRfT9X+Qfuq1SQfCvo8AOBpEsXLM8sHcTv2D
9+oyKApQhxW5h5UluppJIn9/nDNQyRyBGzHg1VZUqxR028aGyGCIgdjgHV08EKtApftKVXLWN4qi
8DshuRPZopmE0XdnN4SSLr8VlaMjXJpoASb6CcBX9/WOL+dTbQLIZgl9lkuXuOkM8Fm5Pnsr0nPK
Hl2rfBcaPb3AYGVxjqAyWn1lKuZM+l4R2s6CYr5XiVJnw7F05LmEbDlnYoSguVSH6Xn1dkxXflil
ZYdRPJcW5OKFpRmVWJgwe7wtA17nSLmJW3z7ZlWnAEINlcs5EKzNehm8B0S65dfyhU3I3tWJwT8T
B8azPvkNS9SuLBsrNYUwEw4ir6Y7I044L+Ye7cwpGjBHE55lQvpu6hZm9f8bq0vtZnKVJKsiAFS2
cfDhQV5vAaHc4Odbp3x1MJ4yMrJx8Lk/R1szUpC8F2xgjvhjdHZvVN57XvaRThJznQFxt6Ea3d31
dKE2YmEA4UVOOY2sQ+O9Yx6heOkLsTDdQiSY287WhNkPCQajqny7JSe7LTFr/RZTPvbcgRhS+z/R
PujZaS7xsHPKN8iGsnATQs9wxstupenNqFJgg8qwhJmCEyVJWqZCMJWYiN6A1Yn1a5SItC1fwlKK
Ckrlu+pFIuuBYCWJAD81jeO10hoXjRNgyky3opklPfVCb6BQfmdLS39PjiPvU7wHB+xXE4VTtwNw
1A9EibbdJx8gOTMgX7SUB+h9ldE06oV6jOsRv3oGGAiCRGgEWgSYzvtVEIwYCZuzBPAshBpHsDWc
VBMb15IOyt6tuSImO4of3XvR4zxuXqm39BB1QsiaxsiljG7Mt4VCxVXsn67Qq1YygCNxJ5fF1dKW
tZBjh0efkn0Ohs/w3okTMjbWyE8y2YjvxnDltigSiPo+u7hNMYK2nhY1jCP7V+oRiWZaRi3jjBUM
TOfbEdXAssKKQ1VdPU7VnWm+R10FEFQhMJvfk10DBgB8kvteAoqitbk5sDIOd/PRIMoa1at0/yhc
PzlNLPO9h5Q5mrhmQkHf67pdTzI6StoBEt8mRAJthiaXazxHdl/SjeONxEzxvQ05c6A2tIKIWVm0
6sEC86hkZgDp7m0Dr95DJl3hhvkm7w+pqX16Iw+00y4vvaVQnBbXFy1+blYYjmwx5+TJo4LjuUMZ
LViZKR6ShOAyk9WYd6SYCwPZKILVHOApNmblgxsLkKmdKAZDXfnIGt654CvbNj2N6eb+KTWutRD5
7gFPVCFa6sRrV1L2jhylud/cvO67xCRRvEMki42tyqzVHJJr3aNqFfvhe6Fj6hsjBTNry4xs1pGy
XoML3YtToXI2DpeDk3ZQmYpB9/aPAKPHd3l0gaZDgcxZfBEEdsYjEGA/eFsqzedqqySRVqj3sLiF
6yMbSbQyQwvNII3IrSdGK51LAyyA26sL2HD5HYwe0VnX6On4/Ua53wYENKN9Fbh4jc/KS7ygCYwi
SOsGAR3JBd0djXujM0mfjjGB/41JdE+whciQqsb7+1PQcOEv9R97BJ4ReLODVkhqJXiPfAo8yN2q
JKfAFjFuuigui39icVxNvHNcdTJ0Xx1IsdPtb/RMd5jxkBv8YOzY/FFhVUe3Qut3CMspt+ZS8HMX
BwGVGfTzDzK8UQ1I5j6ybcCCvgnYRxyH98A8XsBBxL1yPpPdH0znuSNqKmIIsI92/7NcJFA/Iowu
wLrx3Cm1czjGi4+7uIRWVfDuTlQD6pHC81QmrmuCnuZUJXqhcx8NMvQSkZYyYUrRswMBh/pN/uL/
MfxJh3djt7UIJt08jRLUOEVSn+TbjhrS1zWA6BoWvnRR9v5wH0p/o/7bb0Uxu6up3zoiONS1ID1H
SHAw3ECMBP7CYwq5rXFT+/NCJ08NDcgieVYDkZDnPn3823Yr7OmPwt5907JMnjKtA2CYvwyfh+by
PgzZ8AoolaImNNkTymwgRkezo7bSrQuejU6pB1qQp0+GuC81zfLWKT69x2IBqDM15dRFO0S6hdC3
NlE12tYLt+WxbCQ7tCUPji1S2nwZ/dnPw95ktFIA8XLcfFF83NvLzku6xDg2C1VaDmznVrBhDP5b
rCWYXOR1YejCPeiP+0OUIKufFKVN9rF7TsaU/4J680hHrPdzzzYNUbH6ZlaZbEKgsCGYZQzGXTS2
FueJvjL62ckcOQJk0i22U0v+3HpdC9ttNgKW4HgsC/wMacsjy1u72Jcf6WTQyoCErYQPzA6nFgw0
pbE1UV9E73uSmGzO2a8zWgsoyzBWgG7796YMOkK8yWuieBiktLSpFQiiNlzJjmdz2ke63vv8lbSA
Cyt+MCxmhSdP/KMXtON2EhnwB2dPsI7GSdDn5q8bwGTzB8c3NGMl5legNXBFUxrX1egNQY2i277h
vmNoMP1B5SoNOJUz2t/+fCV0RT5JEAxGwmW/ym34tFKsv6Zim0WEn8bcC3y4lgqyv3gkv9xQNxnv
yelcdMQ2eF4UCO6NF3bgncsXcEXRGoM5OK3RbwuPgHQ/xJCSw8jx7+4QrXdQ5MBk4q9Vus+ORFkX
LTHFgWlzL+yWgc2handNqZtn8VscA3qlgG3bQPdKTIjO/bRm3Vb2Qyva1m7tS/ujsCD75T33AalZ
LkksAa5ZkuyfphGmfGIssSeYO9OnCX65CkTDTfV2pdhjgW8YLdLCMLvS6fNvLCAVGE+B8rNqGxfi
RZ2mqwd6/urZ7atX4ifaERzoPe5P/1lVRyeAT8R0+saSy7IKtSGBm7RTq78jgBWkWUuGyYH3et+Q
XXOGIjEW5jWYDg0TBZxEQ5osYfnZZORGfZRN2O9ThSVR17ZHyMNKaJPCPnDZ8KPRn7KsziYjPNcM
5VofXYgVaBaAEpIZ93nrVQJeoTTy740zEvuZT0Y48GejZsNL9YWAmvz0wo9vUMKN0rmIF0covjjf
p9bewNlOThNHaJFycuzhRw1n6M42fzCTSQ2wmWH24bKvPbrmZAcw9cQzGOFmG1c3GivdBhnJlOSx
eR+yH6nnPT4S8/6KbZAJDx3re000jsvt/w008Hrl96PefNcRtkrEXpTWdspJXkMhxyMoYj2FtO5c
D6uFOse+TFdVDJbnWqP8+XyNSKWh06EbD0NlIGWzuf8M2xsYFuCAVZG0DY0/s5MI/EwmVbvolLqj
sr4LgNAbviQfzWIqQJJZzCzsZlMl+d1ioeoje7cYYt6NL0PsJM+jYgUDkpC6SjGouvmU+JnUXddA
GAwajY61SpH5M70r8nB55VUZMXp4eVPlRuy/CzUzbyAWNMkV1ZZav59biZhpEPr0aX7SVOEltx6w
JGLrugEN7XElmKLiwUZ3kUqbLNuFD98CJisNiTGoys15xCMkmMPV1sINDZb9bfAdMNRHGUg+RzOK
SU6MOQweVlQKO0w4EyVa3X6N7TZyhiOl+ZGzjA5/9wehowIWYkPTTDCPQ9CoxP6olnEPA3TfCoT6
a5hD/nlETvTNJZ5TTZYldEELbR3JvYogj5N5tBy3kdXt0s1XMwSCjW5lQO5367hMWpNJ98iIbMjz
o6h/MbEnE0RCHCpTzHV5ow5922hMmUafvkZwebxHz+TAHNnnDX+1W5twQrR7OPBWQdoUPML1+tzL
7SPGZzJkKoBhZ6wahcHPolXhd4Uok2LC2BcC4B8HcpkW+arJgiXb2UfkC+zJ8ruIfVDnh+sNp4GT
nbviakJpktdNOR/EF/VPE+jqr+TmmTX7DXR5qgxvrENNmmBSXt6FoUTtwE2Bqs3Bn5OSODlHKN/k
a3mO3552AM/qmotlWjRkoD/zy8Xnt1vBRvdxsm4GWn8LlTwhUujVVBhXpPaT7ydEnsU/4Er0q9HD
7jcvu3GZkwVI2GPebtHPdjDnMIiaSx1K5j16svTg71Jw4HE3+TjUrwIIlOIaRSeBuFdDckMJyT3f
osOaxxcQN6hXVAOSqg1Ey+EzAmlUQzsOGlDe3ylQkGmkzoj01iQzKbOrYdTbmS46N/kF1ixuC4eE
drrLFWhwh+FctJqFMCsnQSHytAgQMzvvKZR8JYMy8EygZi3cKqdKrMWVJg4na1FCLbjYfOU6K5pF
kCj+CsuFyWwcQOBMP5253xJoU5unRiMfbIdyfO9kk3bTSjG9Z8XzCF+90nvELCmYQuAzIg8ppI0H
UTMEqbfAdsThRv75yHMzD9ZCHOuxD212An2cBqbkcEo4QLYmZ9KHtwQdczNo5Mlc1R0eVWVDBqcR
vV0H4oj2jX+1f7UokxCcBpET+A+5sbvXKZbqO9VEqtm4zAqwgFbc7zkuOMwxtbwFsUljahAzlypT
xIzRZFtKfKEOaKQLDy1zXvNofCWbeVafRWSc6AAg7j4QKclXrxhCMmXWupowXppR12BTj7VyLr1e
89NO/BLBELODa1m/MqbT56zOyRHPp3NDbaJ3OglGFiARkI8yLRAvF702gKcn63H5AjmdQ2tTn/5R
jDQmH5xgs78EAaZH6W6GsxNQYSDoRVXC67HHMczSHg/F1KG5EnvEN3v5oOmPgE8nCd2D487T8v/l
TeP+c4O5RnedEasyQvzo9DWiZkumCjymzYZ6bO8gotJMtWqJufgWj0guzKYVearpHNKkzH8ueWgW
pGOXGsXhRni27qJohX12pqqUUeLRIZfV6e8R7kUezWY8/BZ4OqOsmESmV2hjK3yfY/2oSgHLFL99
eoOav4Mz5kcvQcrIp+GFZS5oQrOFlioU4+L40u41tBYiNnLwbX1zwfxHgOXQM9P7bP9eneBa2MV4
0k8VNhbwyEC3MncJnTLo18AlbwT7TUQ72G4LoHP0LOSSiChtmOvvZzqBSQdj9EVhm9oz142+R4pU
H9jTiXqEnhDWSSkVkGSd/JT2GzxVqGK/K8gTPLypXzl/V+yVu6eDpKrKfNDB/kaMKD/jL1eJMt2d
7QO+31u4jMLKw7cfNsBgITSVtRFdvlie8z0jxWzIM5ZSu84elorbPkLTaYdCzkoxQGt0EvlZPUK3
O00AdZuHZ3cVdWWjII/KpBAKnu4/krnpWTnnqyCtXQXgEqrE8ObUBnPsO+gwSW/rP4ewO0Cr6xtz
XkJGoLq1gqCD8roqIfWcLFVeBwuzhGBfZezlRC4gzawOJPiZNhNCe2EhPncaLZQi1WScLYKFcpPG
7BHJf9Khv9HGOjdKqhVZa9cGWHRcoOBCFweWK8ZEXBBa8J0YcZS+IlA3xNQpSc4JH7g22S5dNVPL
S7vKSKtrIEOm43V/M5uMWTWVAQI40G2xzFVFa3NvRLkrTDIMLe3G+E1WaIx9oKk/E7VZDAjD086u
sbMhe/uky+z1brsQFOKXKfgNBq6KHWB6hNuHk/REtyRncVSyVZmAjG86YumkRZZChiVIL3WY9VQV
KvdNFZpPprkd1AvV6qHFL0KitvfYep3oe7SZoPW+dbOzt7nIazOjSpEt6u7y9ff6Te+eklQ/z8A0
kxtS0MvWQ/d/WVMbrpymmCzXWzALvvpEgcc4uF2ZFba3BFckfDQM9Nqc3PnPEXphOfzxbGlBolnv
wWEJ6rvGhBhlFviascwqNyjP9DhvYQac1qivHs0ygkIfIroHw3PJpIrBP59OrToWeTOdlOyDe28a
K95XZhsiatC7i3AGHSHzjTI1vDfYidHfcjJvmKVTBCFFR1bEnV4WVtpbAUelw1ShOMs6ANdr+rWu
OkQYH5S/u4pkjLa/BLbQq6xuO/Kz7j/b5NzlXE7W8C18yCHjO3C254h52pRL9z6E+RtjcepsY2tJ
S8WYBABS3zVpb/SWJ6xyCuwzkd+PqoPsh4sYVS8ZIfKvCn9DKcaUqMAJgoUzTjF5Fc0h2EBXHBOW
jXWaUeTzM2Ans5KAxvBPrAGPkvFgK1G+2JE3hBjUXvZOWede5PfSp1FK/1KldnmWYlSmopzPQJxg
KLT6rWYaAbv3hFm+rRUkVXNNzARaPlSOnEowl73z7alNuoVuAwzqm+GARalW5fDB5acz0qyWKFRv
Yo8BTjs8KTD71OH8KyJcY0nSTDQKrCbL6UAY/k3qElM+1Thz8/naLNBH8vonMjuNGA4mAORq/OFR
N7HtU23hOrz1ZK2X5AShdmbfrEqlDntpNGBi4xnL/VGPKIDG0o7++4U+uxkw2Fwz6OX9yQvYXUoE
mVyGohZN01v+Mkb4Xbt1lKw/3nBHSE6aa34vOYFg2kHtWHwvD/313NnQ+IM3q0D//++wgs/kOqN2
D5SRpXIUY1qkybxIQg95cODqfACFP0UgJQzeTek0NRgEExewiqXHYRDr2RbwlorisnBeh2ELCJ4l
GUtOrZH1l2l56GQHKHF8ehzpY14IB/m7gukzKLoCRfE7L+hpVFVk+33qcygFkihgmcmcEXX4Ddbo
uLfe7vTcid+i6mHdW5XQuTdtR+K9LGRqwt0S8LODE+PmWEvCxtHZ7bAJAXPZuNAdP9qoQkb/29Jy
jXb7ZikQFNQ/li5bmUDvwp25Qz3zCvoJ8qE15XTOHp9Jmv5L6TMgHMcyqtTDCLKETun1vox4uIGz
0wkgty96PlrownQbz5IwTTKwdSZES2wkCjiCFIJgpzBhwt15n8ydtg/ZehA0j2PR27BwWxLUlF28
D7sOH7uygvFDCLdQ5diwFfrx5j3vLF8e/LdTFTLY84nz4oNA60jNojr1+AROxlmPrwDzgam1qvHF
8glMuGodLtTJBgWyHoGKUqG33hM1DVrBsMHdR7IWU96VyyNZtKo2scJHDJixsp3kn1+u5VXcZ33z
XJKLRO1FpnK8h9kecFKJkWrCwbKYNapAPJD3gEhVqqqx/OxbVLWgZNJGshhLKlfDP2wssqfQpIof
1HVsSSnFBE6I2liAZ89Vf/haUUqVou6OD2N0D9hZ2EY0fR13SFO+VeNdTYGWqI4mdWDDFLwxQJGJ
wkAAd4LLLTaNgFYuZq/KFl041JA9HzSBwHRRcpIEHdixw61AmJPRD7e43qomRKPqCOns7DH1JsLO
lUy0t/9NyCj0LYKnsb3ovu4WHRTDZ9/VAyKFVeTeJDPFpYtXIX5IBVAXtTQIZECvCd71d3J6n7r0
bR3HtW2XLaJOdYFCtxMm+ITvzZTvCGB/fQ8o1qbXVKbtQd4qDEyRWZZT5lkoDK224kF9CcVhMfRG
XtASrCBxjSYsEBdUZD5FRcBx3qECP9TDzDBq46iytqLQ/GgtoEzHgXSy1T0UJCon3m3FCATy9lUw
oXt3jepNPrBNIMEeqH0TB8hZAscxc0MuclI7zNAThRl+SUOHrhtdXMmEw5kJ6s2qXs3IqjvEsWvs
vJW9VeeYjAsGy0onMubvc/Dvtt780UnAszicLQCmpfLMIikLtbVMv8xePm78WtGWiEa0Kf1v3awA
UrDWcOMaUH+qWwA1YMMXK8c26i4kQgz7rfIeIYlOtV2+lf2MyAIJRD/D3lV3MVG8Ze8Ol5JssdtW
Tpo2mXDVi38ZmdX8vtef+tXf6wGUBv8p2KUAPy5yTwijl928NZj+gQscQG4lCZcz8Ld0BHN1nKYY
CIL/oW3ewSNQOeCvaflw2aUdYIlvfRoc84TgI7qf44Vvsml1zbELVzn1lqvZf6Cj1b4w16ze2j6F
2A0mtRDG59wQMtAmMbLhM6QsyuL6dIvxfG8EOYoYMt6w1LrSTaPoCurzxiybJcVCwvD+Ex/9xjtG
Oi6+fHbIyOsksolxq0cK8ecB45koqKg4qh56s2LJXAMYmrdAENMXiWAFsDyQ9VpNBMTD8BsaevIq
vnDwguOP02g6IvlK0zou/77Ikdc9VqLGz3jqyXyHBLwkKmrBrKZvYJbaaLfIhNJ0I3ogzfLo6MCs
tWMGTXT+6P4LwbXEE7DKkqkfDY1uoHvB5wy6IkySzRp/FzqnZD9Sneg4f9OTO4cUv3h6WVM+X9+L
w26LGoiFAwlzR7OPJ8oew/eLNa1gLmvBivm3zRWmDxaviX1ypn/dFQdLulDjOIzRGrq6IdATpOel
OpDjEl2I4MT/oznt2eArFSn0TbrytZwQLOq47I51rSDH9XFCnKE6eaiJyK/yl2TXk1jCn61by5P7
ecSbRynMv76t7NZ56MD8LvA9BgcfKt61mea08QuwW3zK1Qgn1Drcv674K4ZPIvS9oDwkVSG+B9aA
zYVE29ZqrlJLIuuv/uIIFCaCS4ZOM8nCpD0mOAq3+PFjgUNpEVarbHISCHDI4pxjECuC/x2CmUBY
8O5/d+pAhGoixfOcCcZ36x6oU5w8rVKkq/MRLfTVgY6BksTHkRYHOh678O/FcosIwIpS+/pFGSoG
8demkxRA4ibFq8QhNA//tXY4uZw20BlFHg9uZG8FaxQwZ9yjFxB7m4IHu/6ubawIXxACAGKWymAo
jaec7kx5i4XxGXnr+32wyO0ao2YDXs3snAFeCenevLWZd644DsuP4uNEnrxXxJlJIfPov08GoXnK
OAlANzXJBUR/R4i1rOB7Yno3fvmyOlVycBW2t4A6MVXaZZMNOjGX1Q7lnp/VFQ8CLmLnHFwog/zv
uFvjeJbbz56UxmsDYHBFfIKNxWZiSiu+x0P/Hb/z8SQmT8fbg07W50+RyjVnv5S3GCdN+kyy+Iqa
Ki8HFUgGzTELcoF/ElQoJLL7j/L9i6JbXoqCQNFjHFwAgBMmTGo/+q91HeO8CUL+sPRzUzmvuIfB
YEAyfsnHxhLWLi0tlyThloY3cpnnvTkmbDiH9enyAZAIhr5Fsgei1CviYXDbJ5uNImfsJUn0SQbK
vb96xVHAYXdPHoinU+yntBWUDaYLgfFWiDsurLaTQHP908Bft1Yfa/lOLsb0r4L/oIoJelZdtgBA
FnrENbsr5UI1jCdfL4uW47OZMxfteWLaYlW+w30TiZIomuMZyWc2HQy7LzNI0mXr7rTyzKRO2Lfc
VDjuMbiAZZ9YDOalwgbTLylQKD4iqi0tO5jwNmWAbycVrPe7GtgSzIqNRp2FDEJqaMM6wFoqfjw+
P5M/d1ApblDrnkvnDgIWqDpMlrMTmVcWXrUAYL3u3OOlI7tDLnFV4u36SJFz1WnwE9/LDW8+/HTW
QkHlskM4Wfxk+5f1mwrS0DS4vlF1G2TC2zvLgLvFlfGSmDqSteM0iWWJky973Dr6iPBMgFcU13EL
7bo8qQ40Eams7ftu1O+OJPrD5Ib1YTZ1WVc1we7DMUsxSMUY+sjZjL0QMoO8PzFhU/Mk2bUmYeuB
YQ+6coSldxI7VTDDsdKF5qAkE9iqniZNClHxKhtVlF2/1sPgUY1f1HU1OpqM4S3AWhD+EL0Z7N3H
9FEoYfDPv0GDaChTKwRAH0PUAUnqCPyDpkRTw+07hDWKecxm+X1ygmS4rK3Ul1lijduURzeujvgt
SNNiB7zxzWRh4aF6vOl7YmnMuMm+ztjILKwX9FDGHbs2Ou/4Johalif3YtiBZxp2UDAedb1fUQG1
loMTpT9/2CWftxzx88O6lMDMOOLVwtySXlrTgWeE+U3EMW0pwWCkIAOYDXCcT4DlePvKvIVjmGVE
lFcDcI/FH2LlZFyDikn04EVsf7YzyXT4NNsUlxF+AgCPhb74mR4nWyux9rXnHjp+4jeJcO5xqCAI
XzdFnBQMPfq7cxKc12QKfAXEHROT95clgxGhsXkrUx4bsZqA77E5954iLxYu+o4PY/GZOzYPzBVZ
Il08V9FxsBW+xCZiym3FoWgGW8VhFG37HlWRZVT2ISqDSoxMZ7jZCQkuHJ4PMROl8pIexBL6x/dp
NZIP57qdKzRr+TLr+cz1ofGOjhsqoKi5AfQ2WQGF0u5xzWgKhNgxwlN/2FsHCYiOw3YnzSWpzvU5
PyWqVRB7R+3hH2ydS4nsM3r0X9qzuIYPdu+vIwh2aJx9TyOADohBFOMZXxNtB+5xFrjZR/wm2xy1
7C7US35SyBaEOdMAR3jNMMjiLfEvcg8zfo+6ggLaj23kd/EzHPmgGfQjyEV0gPKuZSw7A+7TzdCe
IBpv0Kvt1FDnd2HxS+zHwg4MkltKbKLTeEGR0peO3YBl98au3Z2iwX6s2v56UWZLQwBzEqGFTVET
JueDcSXdO5+kN6CAsBB4FXyom5FDaFuFQRB/vS7OLgd2LdhqnxAZAh6lITtFcosZZYjbx5n1mjHe
afjLZoCPJxhsjtDbGhliW53ZuewB3f/iLAgPXIQuuM8BDpaPwTycEZ7jpKFbVwuEpq8EOY3QCut5
9kF5SHYBiitBsrvCQ1GYMJVk0gQLAhFa0QwPEL9RMeoG/xbWjUAuOgoYm5NjXdtMXi/lA5Qs8GW9
zEdOCM4h+lS5Ey0xcyQIAgg5FKvuspAJBH16hdU68s4zWfGAXmQ9Dpo18uxXp9kkJPIHiPeIdbK4
tKZxvS0eeuwDTBNqsQVOa18WCJbwe/1s/22rm61hZoU934CMfz2pZsXsu+sH7SAZfL/cg5sp5gNK
R0UPP2BB51A6V9pZkOXs5ctgeFwuI59La/jPZvcwNHq6nx5ouMVzUpeBMiySlPR2Xkc1qbXVLpc7
so6d+717vxrau4upN4sc8KO5+bq48FWsNwI57WOY1PTRoW8dq/GpDP5DCPa/jWCj+tyOhKsD+GNS
BqU/l4gVrS0N5Sn/ET7Dvwnvil/HUadiPclgxbFh/3ymD4SSLS87gx9X1kxULmyhVf52BpyqQcDQ
GmRv8BGkSLq8cJ3Y0P1Om/5V3blmEvGm9AA9tNGO4qO03ROZQ++qXWInjottAFI82KBp/0GA6htj
GdAb5VkjrYiRHR/l1/5yymmunuIytmFcANNvHz9MemjLXJYKpbQvYAQ03YMvxGOPb9xuphXItgWg
uaA+Fa/h16HwAY8NJ1umDfbZr0HFCmYv/rq1RycRY/jqj2dypx6NoH+zXy4+522DwkmH42MAtnEn
jIBYYfjXMSs+bpjVD2QMXb+UgonIonZVpSrZs/2oGvFUqS2CrGOsueQbSumeGV40wQasPKHglOYs
tTxXgjsTCd8atmdcDm3EVTHWeN6zp5vwfNkmztXTCORrHSVZiSHQsNgN6N00lAWD6OKBH+q8PvBf
2IysDZEFzTrfCF69wAxBDVqYjhUKkF/GBzoHomxXxlSjNx54ODLEX4OU5b+aD+gbem0S6FNE5Mu+
PeaNHp7dUdJceN5yAtt8fVvq2FtPknhJV6JZZ04hy6F43uLRZbTb/Dxio7XAkP3ZygcxON82+HU9
VLH7aEwYvs/4icVyJ1J4aSQVDLuH8iRy4rMlSqZKhE09K9RYdKuWBehZKzsYd9qtpT655X2kxh6P
rwqr/lDv2xgUMKmwQRX2z41jiv4BUFncNY4KFYkvAxIdf+Xy8oR3HaWpslroj5TTUIodTB+lX8bi
FuP/TvbcyKvWppLIbrUTJ3TKMQsoH7LxmHR74nfBcEUETQXp44jLmMh4WeEW/wdnzGQSu0Lcx3/a
1ttAt6joDVJTWBMCy2qWi+gbhrJL0ezHOo7/mnMds1RXxt7cISw3fyfJhhgIpZKBJ2V8ERJU12ZK
iqqpKaD4ilt1Nw4OKqFH7JrpGvybUPkkUTlYD5NP06r/rIL5OJHhzmeW5+CgjSoTvV38xIQbaDe6
4F21TO+QX+er74RPuWloRtZK0kw4sdV5856rYVc2uud9cERtpeRkvaoXw0r8GSFu0iezuluPJHm2
zHE+0OIL3xefhiuGQ42qL36VBp2zCr6yp3HScUU8td4oqDhBErq42AiiVlAPSqBIINaWD1qVC+q/
lGkrlXljCFQjEq15sFGBv2R328CokQGfIuaUVCq6+FodJaUbN8cl6nAK77oe3GKv6QKnyebJ4lnx
8LC+BUEMiF71ZJG01001RIapVUgTcU1/wkPvPjTMHlGi+VWZWEl7nzaMUBE0Ko+0ahqQq90v/wf1
NJK+Z1AOrL7cXNmU1CZJAwIp9552NUGwa+bxdEjgxRXoxkqyzshqD3pRKPtImcwJ6cZaEMxFfaXq
A1zK3TIzfIOla4CV2GzcERHNfQs9iTtT3Bs3eFEZb3J0HN4RQ1+5FaN1CcEQ+TRa/ZR9YI6TKkk7
5Sz67fkg9nnU+ucfpvFrxVUbeAbYjoSgq71BGRekADTnZ312JGJs+IX558qT86Y9ZDtFM1hpQkFa
aSgjbzlLIt2UO4E9dDlIoz7ZeWnTnD7zh/meovoZNa28a6nAEHjq2YWXDHvg/RzKnTMxJ3SMHIEc
ZdMUIthIlGu/ZEl4GF/SBIr4sVN6732V9DYpCAOGRcxk2rnB/zqU+waYt2y7UmXwMpqMxrazvlf0
gaSKwzD3pHn8DQ3uVsKLtsn1e1IHiQNhxbRYYN9cfz5m1zVOMODMqwW9sEi9wTaJSmcG8jJGp9lV
TzPCBgvjwV0iJM1m8vO70Pu2EmYCaXBBKq6UP4QFt4nZev5kDY16l8EucgTLmF4bHIJ//6LLyC19
/sQ9+SpdbX4/AeLs73u7FhRWHSUSjITF8pUR0KXcZAWuorPRRUiUMP4fWI5mKJ2Z02eUcNMyFt+L
ZOQ8F7PxKD+2Hy5P1AODKm6Zz0BciP7P/N1SMwFISqCqM8xvjcwdNsbbrug7rlmDQXIX4JcUI7l2
Uillfmuet1abJnW+v4QtMMnYySgoCFQlr3xnn0VbRXV2mAozcRDilPv3KFMmKwHAfybQde0f1GJu
O3KrlWqshuYIcQiHUfMcuMFKL5N8ROCao35d6q81IEd892UwZViOAyNwxEMA+8hmVPKUJPHf1up0
m6vtD8xRnfGhKCS1bO1KtunX6HxnS38+cKfHMCHAr1LQ+qwR2rZpCAUDLR+8yDaLeVYeD0ylEmin
Idc6xmfrPRTDdHq97+rRMvyDmJzvSeQAThjcKlInMc6Nmo0aTpnTD+gjEBdXKP6jStCgUtihI7KN
VJ4fUjtvEFL6qksDOPg9//r73YtyW8Q6dAmfMkE9jJrWENqYM/6Vo8FNX+3RurK68Y9cOBdhB5Ps
oy7PyJql5KTrycd7sE/SrojqssrzvPO9m4waUC55KGNXZidw4nmzCBAzfHAEBYQxqulmfM9iYvhq
SS1Yoo2wtX2rbShkaN9eykD/bizGNIarA3Gz2UfF29zLiILL2vec22dYaPpjJNqX1Iog2IViF568
UWVB8xRdHVAvDzd0/CIt9DYvRjb7VI8RJ40VjW8eacO2tipMYTkimEW975Bioe5iIc1XhbKZfD2m
M9Gdbywlutp+O0iVFcGL4m6vt+tZRgC/N4WFKm8IceCuIxvJRdQajDz72hgJP/QRAw7pLd9tUcdt
A6kHjmTWKs+BDGT76rv7pBJpUAYTNXAWRamX1U5mehqOPQbNReP5WrJ/JEPsJGkiSxpuytzXPZkr
DeXyfRv9qPBNyflsMrrm4prVAAKGtQRpQGs4LSW9G6hOOkR/EvJRad/bE++2p3PjHNahkTzgCgg5
sVeIvP98SYxEtXMMNwLrLMIhCIb+l5TfgItAQTQRdDbnv/MuO5upuFMG2+Y3BrNzj3C06X9PmpiL
bOXVhWRDpwNDyDuxm6NqnQetsI7W4BVdMLX97/LeC6ZSeUsQM6XsnEmrX0WPZOV9vjGUq13XNMD8
s1XFcR/Uzd2OTogzKFgr6Gz0ID+4128jgL+qfQLbNzTlIphZf+tMRqjCYTLV+zcgRJuJ6QwKUDhC
eWoes0MxGKvIQnDZuTl5OGN7jux13TW+S1ZaLPjXV89YW/0gYbaxXp0h7vP3vO60FMdi3Nop1kcM
SvxG7Jw+l+3z7PzxuLnb/unKlgAl/iqFxTfmmUQd7Wfp018KiUR87S49YJgCmbx2sF1n32x/0Hov
Y8V2hmt8/OclSN45MhR0+Jh6mN4ENij7/C1+ULc9C3pOAiDT8Wu2PVqsSpDrMJYZLnIDu9kK6B88
pN5/qcsQYOf0HD4o3QQRe3A6CkeaMFSSwx/kG3X5NRHkPm4riRIO2r8NPFraco+nxBsHREGxyNPE
0ddm1ihBnr+H+BDAZToqHgFKUpCv/UD5+JoGMPXyQOFfWnKe+89dTC1yDmQsqFHueXinVXL7aC/M
SeXX/2k19WZg7CbpZ37/JHYLNSXXSuNgHRB9OJgfycPfYLUqNGtdIZfyC9Z5Qd1yFXR45xyUScg6
xQiQ3fn+uUyoZQILD3xffcydSZgCq2JSVUQeYj5qLPLN03iJGbqCqVWDq3PyOw1XIdVFWLUU9XPN
6Q1YH2wbUDa/nkwZWRlDWtEUhVU9+hTBXJ/pOXlTY/7/X+94waxet3o8t6wL3oL/mJEPfUWAvgEr
jDnxmpqY2UD5hRZn4ixScbPXfXPRyV5Bdp385Cc3MUkuqLMqn498nwbQgN6azstC04KAN/W9BnsX
LJR4v9g1hSmjk8UICVhZkUYRYFNDFJ7y0MjGtlaAspa50HjwG56V5JdKbf/v4R4B009QO3VrMdfr
19wGjOSrR589G8Ea2hRVyZFNzESo7Qs+i+VSlDfI9FUpU21d3cYmYfjf3TxAShF0ZHYsViY2Ozgo
p3ceEJx5KnMnUf011lAsSP66KlRbopMmARsBnB/2kFndqPj0Fd8bkg3HKp82ZIiHIiObINwaLZUo
05PIou91CFRNM3dFjwAKuJUPnJlUJLo1hN6OWGKOEb5g32BcGOpBtQS+OHlZkDDmF8uFxbIkrUZ2
9duHGdeXB8u6V/krEBNokN/K525byHbZh9EdUj544sQLgZrvxcz+3bIyUBjZX/C2ymycd2fB+x7K
mcTgXFbxf7iz8NTyatGrw4ZAWtCe2767+CXd8sO1kG1TkBloYnUoH+fARKP7mut6CIMRrloqmjMz
VBJMbUhLcobwO8ak9PdgCD4lwwZTTNVVcGr/plcd8aAnjGL1QGcm63xNYWvA/m9lUOd3oxju2skF
6pQ5lvzJMptJpdJny/jgXuW8tyDomXxZ3eyLhS8O9G6SedJFOnrF8TcHZYfzs1lo0yBSjZ+ojM0z
cSSAUS4w6jg+5a+kXz15hNEifZK5ufiiL3QlBbjuTyLAj9mzqeBa65XkkuHJLKf1Lxu2VVFEq0lc
JR6SIuZmNUOXU8TlrT+Qwf+dwHOTLfl6bhR5VnNP3R5LTQMDKrjlED9xQw3NnUwPbNdambl8tvnB
3XqNkPLqorykJkAftRb8xzCr8yALNMfDAx8kpKSWOvGaiMJPbGXEghzCqQMaWr+slyvBiR8VrkQE
IRf62mm6qKosAYnYqNkRCTFYw2zujON+FBvu0WEzLfmT2jKpQZ0MjKuEcOahOaNa4SMaEKfVJPRy
YaUvTvtQSCXL01AJAPeOUyjj2kJrrhat2NuV/KOfcb11+1vtqY4YDaeroLy8j3wLbbrtHDBkmwvI
9o8PGCt5Ov6JyUY8BxhAxVjKm7Cd8RjQlfTYfxqH3RVXAb+vduxKBr1nc8cyHrHvlOnJnQLBwUp5
msk2dPBiwU9vXjaN7CPizzPEJ7gz1A7V7vzVJ/vhiin2s114/FvsQk4XrJXgCKOmmO/Y7IgTOxQV
xoE3vOrlUBDwrpmgjSpFkhvLOaIRPYb37EidaHuKp/PJw5ReMqs5vdyxNu0GaxO6ByXfFUIFEa6s
o/mTpN67we7njIzFeNm9FxEYE2diLLsTrj0CL0J9fXf/c3MZZ6WER75behNXsIrLDqJ0ymPO4tvx
UZOEEdCzlgFDqrT+xU6ysHXCM8n8BMT6tsl9VArjkudqef04pLGAeEuwRVxmsRSTwXsLDjNlhDKH
wITndrYShk9NlXXAst73hA926zZC0N5JTDZNZqqBcB5DHCe9MWhND1aqzgeae6vy/N0k9d4yOuGU
+S0bDZITm932KtVL5QZKUCWlnMINK53bdeJQhvzjAj71ZsUrFGcQCGqayCReMw32AsD4x5kK+92T
1MjyARj1HZgdyIBfXKtEsVru6wreS7V/KtmQsvxvBTXZKnHFlXIWmLclCLIozgJzWDOv79Q8K4N5
CGmVD0Uc/gYAwQxhZkGhkZi8bmiU3q+QO/CE6UW8sZptPoG6uwskaRONW6hvRVFJRvKuVwjXQkDB
MBnLMIkG3jcNp6/YKWzsmfbZrr6KWmogrx193KZZh51j7KkHF3eCmrTAHSdGvK5ig1IYDr6SX1kV
VPmZMFN2yyKXw84sjGiASmubp9+6QqyzJbcRebcAmpivY7TNgfVAjE8pS6MFeRXX/uvkU4Q0ATYe
6QpLMC1ccX/ryibQLcPu0ArRikeC9WQ0/4STOiYJpbe0sn97VZx2qnkACMhHC8UlZW8QtAzK0N97
UfkWfTnpZFBxAaOQvhM76oJzhFrOnKIrWapethOdZq59269L+rTUo/DOwd8olJ6DunBkx77HpW2k
iywpgXlgJps1+aaEyP5cYlA9ua4ErabECS9Tf54k58Eh3olr/yr1wtF5rbenSMp7hylDYFqAXQI5
zFgxgb5dsSExf5K1PrR6l05lXRyiu2wmZPxwx5hYabl04/d1bZgTlLhH/2VYk0CGtxT9rdQqXD54
yrLasXPkBhWfVBxvC4guMYiTaCmgxKSSzzMSOZqRdFEYUkmcCONCvWcQiklfDFpzUGwaJYygR1yu
PimJXjOXHmwmMFPJ27jfu0r2JnmkNgYK/wh3Lp0FXvvBxV+UEaTmaAFT1gKN3KzK+zJTusrBK8ug
bO/QIbBo6EpCuuXREhZ5CwY4ZIJ4Uh2s92Ps43jR1HU1NqpEpwVh5aIofNyQ0SbZIGlfOqrJ/Vrh
tS4Kp1BBMr9CjOQE3RjotdxEkiYfBZqQ0a275viXtQGPMtymt18aWy/+4CXQYRhDTvkrJ+bxVf6h
CHM5IHspWQYUds8ZfWSJ/I6Xp+H0DYKflaKVPnPhwKsgIxYgOgz6YnMuekIHuhMZc4laWR8KqKDP
98UB3E0ojS6B8JY6aZoiKBJllDIvYuiMcJwZaWXw652uZRdklrZRUFBxbrU3eI3xsRKL8N7vXJsy
7hgu3r6b+0bjlHPbltECegzti12cqJNOp1uGFyq/oFkPf1XLT7rVBXIfkwiNhIuJBZK0jl79KaSu
oa88lnRoYALOdE0iFPLlAUfjbsxsbznegdcRSoHHdENBQWi9vY8VRxQsRewQirQTbSNrcqAsdZuN
3wmTKtkK5ZR83iFl2jAG5kjnjqwT1nhUZWZny+F8pzDQIIdDmXiWvoy0EkT+x7vOFdqKGEO4IcyV
4VpVQxHABfZTWhJLC9gzTk5EGhrVR3DDfmCYVdlAcPVD0sZLuAyO4NGUykUwNb41TGYCrDqkuZnV
OyqWUkqW+4xA814VUVGplxo3+9d0Gw+FjWWmfFbi7ZsZIFo/INoZmlEBkn+6qnRKN1qi4duEX1UW
dVNDZZyvvakLD4SCC7NBI8PcBzTWTk50uuUdtePGAcS8VgCq6tbqOg67qQ62aqSlpbbb7Fm56avq
WJ5vbxOZUBAJnkVZtQZO1fzlRS+ofrSwHV7k6kL6O6mR0hj3lTP9Sz461Mzgs8rrpm/3HFm5ikzn
6xHBR+AzxWY/TV/z5IDFgtcPmuOx6syJGqCAFqpb6qAK5S/JQscgUbY90vAr3PL56nqmI5amqjkJ
W8dzRNM52l6L5/AeiT8+IcO8rKD/QJCgwBR1H0zZx9Qr6TgpZISGm2KScHPZS5KyIi0VfN/5EJG3
JpvgjhWHUjULhG8wNdouvCEr9jI+WCFvGm1urQ02wNPhzsiD3ma7Y784RO9mxLoZ9pooqmGz466v
Exli+qXioIz7E0vjZjTarJaZCBTCx9QsZ9pVGZQKxYVFaVHa3tCsj7kEPb2sDHGF29HVnBRoFDQs
B/0Zmxu4Iio1+KwqSBifBgt8qj8WlYhtma65e97XrtNEJU7lESYHqGSWQN/mRbZk8t/cYPyfo0WI
DyTDaZVEoopOUQOwM3YJSrfYwTq8SY0VNgecjf3eLbQfEB05jkr3gHnSZrkbrBSXdthErWemB15W
6Zr3VF3Ar9V+pfSya9tCAaPqle4J2GQJAvF4LTXntCXq2nd/KdxeqsgLQW5/PQ9/DJoSyNEYOjkO
15qUKKxK2tA1dof9xtEXKGEP1L3PP7NvxrtaKPRBLvJ5p5J557KFjk6pjh4hupPUe6f3a1IQeALZ
IClPIhQ2pv31KdeimsexM9Fxi+LKEZCPA0PruaTJuCehbKOjkpw2VETHvzcs5Odn9keMRAuFy7Ej
wP8uCTATiJUV2eVK/qk3oQgLTwA++0I9cs9Uv6Au1WMbi08QsZxnRNSB+AyZgtDMCs9ANawJpTBB
mx2EhVoUevf2OIHLfDkJhMooLLktAaLknPxshAsY+8r6zKopZLhHJXmxd0X1anCXqsr1/kOEAFIg
LsnwGxIz0I2sUTcXEtAM9b4iFff7xLnT4J49DRkQcQw7FzmjjhQARCzmwi52VMZo4FT/fbh+Wah8
eTya881eAQni2EPkGC0T3wPI5IR1fNCz3hyWSZoXKtJZmnubSvVOCMz0FhVLM3Hk1nS8qEMpXZ++
52FWLQrwewPfm03OGRd++IvLDB4jow2NT2DfU2peWTIS7OS3DQYa5CD5F7tYWmjHDQ/T1xcoewiG
qCS5JlNA7oWNFXjQn9Z2Ig7aOBoE5UKHEALg7+9ARFW/TrIC5PNFcUL8876DbXmYeItyDtbFptkG
jZMVw0xxw1ECZzaqwY65iQsoj3whw54kM609ln9QVKLd5Dug5WKKvBTv4N8kKmU/Yf+8GcdxJ8nY
ldOszRPs5cSKY1mV8Z8Etzmt+phRFYOTa/JvJbunGDU9r2ysIWm3rrK5Vu9to0l5OppE7SfsBumN
T2Ly5HWb56jnCrTjmarkSAx8jV7lOlPgdBfC32J5g84Q5wXbzyNY3Z9RmHYFy5k8UWWqeG9J/0ai
Z/EXePTjikn7TK2p2ADT1nDywgM9YzU7NNf+2hgj7YDNiOHa9mLWYA+oWSpU1+SEPxWlk0/2HIde
GGLNSwBP5ofaNVpRv8IcpiqoSusncUohovYf8HH2xD5rGFLkydMgaP7mzhIPd7wFjhSuZXJbC+12
5vfepHOBp8pn/oMnnbZYwR3To6DYboFsHWM5nxHH9wW0Ujkd3w80Nb5k7HN8kJNwy5XwOG0Ktze0
EE2bHmPjeI5LpUj0d4h05d3+2KKqPeLo+0PsqmQmx0/yAv1APCXx6cIaSkKMWJSZ8brp/vkEpPSB
vr1n0VkV8+fzvFEXHTOOWyw2etIe5Qu8CQgLuYFvdbGz9unjYgNNRhuYJI1cwSnbnp1y0DKUo7OT
rqJHgN58ck4roFHoS4r0g9GMzkRbFcq25fODWGkTAlBplB4CbNj7enKZJRc7IpDmgRbDpEw/ZU9X
iDszXKrQwPQPQlwOye/MwZ2pOav3AIkLJHZoyquuyUDU9h+EKQlAFSIjjCQyE2NtiQadRFNSbF3O
6wQFKoXqpzL+MWYBBjaysysKB4UOYiapZCqL/pNTrjrpwa8mEhNAlx4hVcw0js5faZ+bkWiJ1hUQ
VFa9+fYkVBdMmfmKbNw67kj4kHud5t0wjixXqtcl6m9x4h9H6lJyfS/ovzGQrK67lcbidY3U1+O1
hAlsoaJGh5CnatsCjzSWhCbGJnIzA1+nvHt08RcOlqswsPLw6tbCXO4d8e+vmn7u9MkkkqQ53QRK
b9HAwa45zwHw4nsZry77Vi7P3nAog8JBeCxWcAcT1cmSAEN+dnWcQ0ESQN1XnbsPG+8I6gZoD5tb
0ZaEJjXV3bOEyg39iH/A1XY2Lra5lu+0kqKy9e7Mpg2ePoVlYbCcNcSXxntA/1U3swMOYz84Iw/v
zo1mBWrLCo1YS8OdxcE1ca0amuTuDEba3KSgCq6ylNhx+TosJ9zFpdtTFa24PqHAqlDDkLMNk9Su
2jwAVu8Ek87VmkpDBkcxfGGd2QtUSTxhjy+PqKp2yI9Ef8WWpNT/SKA381Eo7EGaqAScyQW/LaB2
Qy7OqZg3/8dO8X8N2XY1kmIeVcZfTrzg4EpIPce5f7UPh+cqBp+18TlNgFMpOQmATaTIkQKegsjo
mpLfoP6lQ4QSo6us6sNfLAiqwEBuEANxfXGxnQKixvHB301NemZ/EW7TvKZNM0PH9biuX4WjflZm
ALbpPovykKiNvAy+QUv3PiRB3MF5CFMnVBD3qdgSdAZb1GdMdjuSwxzBw9M3IK2MotCz1hZdKrai
mrMyhM3W7CTVehuOoErxm07vl5qMEbp6DmjQemFcPc1LCfb/MyBl1jTZWvYuD5jNVz8+QXMdnY5t
l7tj4bbc473PWpp6g7ScNJRPAfkYYDLbCkIoUDjl+rN6GRe/UR3JnFzJhlMoy84bgoIfwbPvj2nR
K/Xg66bTwHpzurDCrkmxD1EtRxeP1v5re1q6rHmqnlKk+HGU/WJ645z/w7NQ474I73m1sbNV7s0P
/9ecfLyvBc6z38W8JkoCbo44/EQe7qDfsS59FoRrU/juzX09iqBJ4cQytwu1tdpUXo8vceZ1+7w3
GCQHyHFIrmz8jE3ame21Nbt2nJYXqrPrBw1inSOkdQG3LCyYXqKn9ZEZ9HZYGXrmWazDcLRQn9n7
dMgC1hp3vwWj5yqhArOISPA2zH4/SXo9oizig1mjb0j9gsVsNPUK+CzYX9n9P42grl7dkxWt6Y00
6e6arKvBNMKdBxKT0DCR4/wkYj3xEJAsP/7+wxNbf/75ptHssYA534tMKKk4UW/5jAslklSEDuUM
cW14pvedT40INWbw9Oh/f5nTRqIdhS+pxwnVLaydQq73IX3tMdVn008VTiAW+Ji1O+O1d5J3kB+R
dcFh0CIhYyiP0abheHkiKS05PV0ANhGZCbt+jVjQX0+Lepn+v2tDOpNJM+KsG3+Avq2o1zBmcYQn
3rU470TGypWf3lsySV0U9pRLkpPveSFBUkpYs4TWHw3OZh9XtzKgZj/lBoI2KsghhRmsWqsiOmir
9WO1fHVDNS7gNTDJZdWNYRYIkDlB/NeFOd5VR1Wnzcx2uKX2sWnGA1MArkhyfGlCAagjgbMsQmAL
lRuIagfbrBB+cU0nEA6xVzV7U6LM3V5gaxQKiyFhWf2mQUyIZ3IOH5kBeRCrgEujFoEq1WOUzFtD
fbOk17oBhPLrZFglikShhsd+xCsy0Oy90fOWkltm4b/EthIZHaTwJnwpR4TN5pXq4QJVE9fTZ/ya
DYSNw4VzwhBkgD7UfrmmoNx2JXsy9Ug3cYK93tJNjIA68qP7HGC5NsOQLQe+3veb9uvYR24YblCi
OBi3Ckoh62tE7ZjRKNRpmeMS/pVyRcQPF9sELm5rlXoBMWPotoMGD5q8o01k08EFs78MzZDPNhOe
0KytiBNr86Iwisg1zFVANX/Tytw153nwoWNVb8GGbSBZaFbGN7XwKLczAFboyxa54dAnxMrNpyWn
pN8ag2MXJ/IZVGl6/KqhdoXlMY1tVfgDfYmfNAM5WFNodEmnPbh7UIUOgXPyPHmYywQkj6iOVWQa
X8MPsXbDdPBMtqBEU8AdJwUl/rLvTul/deHTFLxdnVxzCmJQ687LzQLMiVjT4huBfCNvK2LLK0VN
lLKm3WFHlb4PoHHKtRaQGAHslwnZLz69a1xhs1FM3HgRwMiT5g3V145uQwm3Bf34wk9a5Ss/rNES
7tQoiXIhRGF3K4EwYn02qq0mGAAgw7sJavIsG9qyQN7wHb9piNcQ0js58+FQdtmeVoRMLy7uasRd
f1x2I9UCtbTmHEG7BtWt1CbgoCqIF7WcpjyAfq2U6YFfhM9qrN/iAMDwVJOq7xqdCPVqb1YKTuS1
kh1cSuknWF2IQHkfwqNLFpFwqEIiqByX83lPtbvq4i15O3gPre6VkTHByhM4scmkk7r18OuzuM4z
p1H0HUOljgGXTHQOrSBGfB405xK4ycrPS7GZfkJIDJP8ZxW08G/U01sdhV57UxAJzXnD0QzCIKtV
Pgb+3UUbs6Yua+iiS+tAEz0W7GzbIIdofymq114dW5IcgWObnysLnpX37NbzNFlCuKmaXkudD9Ze
rCq3FuD5xERhYAIhKYDT7dgA8/+F89oCUJVgvTW4fIhTBRbaglq/Uf3VH+ij0mYGOT0SWypgs6gc
2D0u85xk7hEW5RPk81b2NJxOyMR9/vXu7AZReEazGm9XQazXSdHHU7Aj+M4JzY/f8wQpUBVvK5cX
0I3qIBJ5XwXkEsa6bPYBuROwquPEZhWGWO+26SWh2wMysTA6nrs+6tWIAEhtevAJ90nWLgMPCOGT
VlZQHZmN1rL8BzsRarP2vT/A/h4fFMp1Anewog6eNWlJX8mylIwcVCx7wGaxab84WrBE0+Wv3CRz
AHDWB6i1n6FBzDze8ux/emIg6VzXw2EBeJd1qutQiQGBgS8imyAMqAKBBQ3wkb9WLk/3KjINL+al
JS6soSWQFOP/Q20ExfI51rgXk9+DEHd17LaJaCNOs7Y77FfCOiNcu1hCUJlnOKhXclLVCK7bRrex
rP9OqEDCnIjjOxE/oaODVr+mfpH7e0xR0G37UoLogHK8ImWXxOkExYiV3bDIrKIMF7qveBHqEyS5
4idKXrUDSaC9uXimUQIUSjG6El6BShobHusfdq5n4eD+yTl2glWeteKcDomk8d1/lLWqN+7GmiFF
9JE3J7JG+JXORP5nL7PZHPoiN8cFMuJ7GFhtoKo0Unuj5UKUu311SCh16URhgwzMX7GNezcyY8yr
xocJBmF+ASYiJ3wQRCPcx48K5BN4+XnwpQntHwE0MXFto8Vrnb0bw8xVfmU+xtW0AjQlfrdZ5qCs
FUKyB/Rp8nb0j/HXGXVWjqxk8FMiRMGQKmqjdfz3Fk7YHa7fxhe/p+DUKBqiVL/Ii4JucUfeh0oL
nUCzHMqTLw9UYAv+apuEcPt8aw4fyN+AozrNFAabca8G+7EIHxILKLwKWvIhXAN7spwveA5P/JRZ
c9JExaYYqln+9HWL09AMmByt9VobQ8r/1Wbp53ok/8xWRmqI5TbbCNuO17ItbuU6DQPBf7WjiqFA
dxoAsvSCvgmldjVuHEz53h56UPROQOiRw3LmcOYBNY1EmXZ8BcFSVTBhvnmDCxVHGeQLXJv1CKvc
x/Kw2IJOu4YdbzF1jATwIjevedhjoMbIbqsETHS/cc9gUpYSs9DAaVaILaLi7kjqSQkWzFg/uWYq
ybSUFtV0jRDEwrbDNIzNUoVMHPqGupc1J5eGVCMoVmM1wjau/J/xD89lED2p0hLemQ1N2eNJ9/iK
ifmT5MNkYXIYJDTV+BTFdORluiarGmTikqK1j0+vE6IqB0R4bE+g6E/jrbYcl1jLhYBo9iBPR9RT
7FKAjbQ2gyhzOGk99YE7j7r0C9z8qMqUyVmvvm9ObopyMJZazpWREgve1JDshXADnP2/kXTzdm4d
VuKp5yUpA/VK+LaISNl+zghiMmPXzFBjfFVliVbpHKcIKozFAsp8LG6YPgHWPx62M2BsTkCxdk+C
zUPp8eJCBLZ4v5pUMotmbcn0uvRBlBxuY1rutWTWDzpGTE7IzrAVwBmbmGpNTbLy3K5m7nKQqKjv
hyjtSfenXlvSms0QDVTMOx80n4fwb6kBDnyid8kPKly1yMTt8sM6vCFxVZoILopK0y9CKxVgqdK/
BqHJT4Y1wupA8oVK5H5A9mubCGnAc8SG1UXxyF0AncdqeTk8Tos6ebQKKcPQjpoKqWyoSDgLyjXm
owHYpx1hG3bURVL2eufXGtZSq/1pBlomDKXrer8y2hJspneEO/+46EJpXWzIizIBT4plOBjhlt87
cd9vB70hxW71Fs6EKiC7wwVeB8/t2HciB9fKSqxBvChLvz1Tite0oYCSmx8mOZz4T6xP/aFuOr4a
hXlAsJeT6p2lNlLpEg6TuSh8kD/F30nI4eULKvUeU8XJwYQYYCldt6mj+dqw2kf2gEcy84YQC5dw
G85JgxVKp+CjmkQlGWsBvFCX+ym/IyqDPqblzyftR6qS2ayvb7h6e7ZoudDEgIablkCM0OpTrIs4
sEhXHiAHTCmpznK5XAwIeZHvoaR5FdA63qCVcGlVzBissJTfvQeWJ2C3q4LI1qw3eZAmCnJ53RF5
pJkvoQLZZB8o0hoRe0Iu8yF+D6UX+AVGUBcZz9R6IVRs70cNGefp3x6F9UQQ9vA4jN7gww7JuHZp
bLlPm7Xg8F8+EeA/sdQlvpWZRSXEf3zvkYmrengAx+N0UIGsbOqs3KNXpeVaCrEEfKorGGQ2f2CZ
5VTbZojIO0iPrmHtOT3oXWtF8tS/S9IsStEg3HnC8bNYt9uapJ6KHDzHNUNDVbqlXnF5WEBD/nt8
vo2aAnf5mZ+yqwGOq0E+SCUUrR4E3egbSq5KN74CETvCT6MozpJ3FLLNmzLdWy6vLc5zHvHr9MdE
17Lqk/3onnS+sV5nK3XW5RF+PNbk6K2J1BeLkkcwqwly3cd+uOvCK2XBfNH68b85M5CQVX8hc1GH
4HK+R+VcY7hM73LIXR7dCd6zxEXzoT3ueEbbJydTNMyGkxxJ1NHAlqbB0FLCpgBp6YA0z4mKdUIo
eLGIY8roSpAjsGZMstpZKtD6EGXkSJ1Rpfs1ZdaN+RujcxS6UsPa6+f3P/9Wa29H4UeGkFh8Tx70
/8SrV4zCvvJibOwnSIjxcO0fBBMLtAIAWc2XB5ttdxhVnfsaS5g5BEF9MHxbyp4U9vu6Liyo4FVi
YgCJRnDOf9nPtImBKnHHC3kjAYLqIWizTjuWatacgdDW3QDoD/6lOGNka1+5AdG7ADR3BNvy5mKT
SZCIFQdEIw7YazPdXYnOFQtrmter1T3s8tcAFWv3JvM8dOKn+XVUtphnl5p4A5Ar9ildo/AmrVps
PXzYB0J4+79XdC44W2CIcbPd5J4dI58L15KFbm67TLZGmqFJV1glIn0lgFjsdA6qh0hH4l1NrFDw
eOv9NRV9iMVjUHXicmVNSMKWSFrdwx9zUdBtCNEUlZaCBb639/JK6zH/RghtUlrQbmjc4bR0SW6g
8jlYo4XApN/qUUhnGUgzZz/pV3e7z5nKWAIMvP9iKifaYG03Yg8JiF4Qi3VmazgzRMEhHLNeZoqH
6eQmy1S8SP/Rngf19H6gIR1/SS1zc5fnMIP43GP0GP/IXYyUeFIg8ex6fi9wVjwoQ0QWa4uRxUkU
2d5/c12pTUx99W8YbrDe17EDvWr3uQRKO2fd1L4pGW+aizoN6n5/DIHgIiiN08vuciohLYZBIUFO
ZUD6hpJZd16buq83JZS8ASWkFDuTwcZQChq6PK0+hJTG1TcI2QGxKn+DKVHvl7d8wEIh+74b6lSB
AEd+LLCi0Ea+brjsuRmXpKgh5bhOqwtO+fX0/bkUOd/oWGDuhaTNG5v+Z5A7VjH7RavX3+THX19Q
R0ppS19BjioGzUx5ogEy6AdkPduO7E1r3MWV9mFhwyINbgN83b3GCOIsxdjompbBsmxtKFtZwdmm
WosuFSvdFcroDoWC8zUPzHrGojGegum5AEEthDUlNg67LUNqft/X7oTX5XMPmRgyhOw8waCDQw/a
wpiq91uVEb+m0fWnW3pbKfMXP4Gmc/wjHxgtdf4iMR9pzq2dSIR94XkweE0Med1/SFJe2F/GMKM+
pIvl30od7WqjEVNkYdu9Y99s5loy+kR1dBnuay9SBWsgFZRGTlZbocPFXW2H9Gs+l+L2YTQNa1Wm
S4ydQ/c6ep0idsCGwy1au321xcrRtbyXLb5WSXJc3Mw0+wG4kpLKAb/z/BCadSAjMrXuX/Y8dQCl
SafD6NfS0xZCskWVQx+OjlUIX7TDzDYb1PEijVKaIzd0Izw2T8NECiNwlOUJsatT50qhEo6grCF/
EpV2kl9ata7qYrcFBxnNtUykNQ3tWMzSLDYINEmjunVgoBxyXdPPw2TOELNO4CtcmZcwSZHPeSp/
tCOSj7vseWRITtkYbBCSJpdt3SfdQySjc5Pv9tRiU0UquM0T4dF7xmZyWkGSGeHzUSf+BPJd3du3
c7KB+5yTWjn6ZaTqhYk8OssZImEMY0RBtDfat2BWc72ItLNKP5jEWqFvWSPdntuVPtn1iWxlUxWi
wovk7WuZMSwvKJtcDZOfFg4u8qjqBKVfX3gJ1QQTdXChA6C6yDoscglKQBgMbjIyiqhWRL5Y/qwE
zjdmJptA5q40K0WW7m1SUacWFgfKyYtp2RD2pQnxQfR0eSYAeRs7lCTnc1m/+ICAYWz2yRkHELTC
UeXQOzwujGNQZMY14tc7TUlh0ChxYEuc1c0ZRx0JMYbx78lk6rdfIjQP2o5GJTYr92N4MAVbH3nA
cULWiEAPYgkDM0NQ85kxfHgnEOBYqDcNe/TnzEluVYS3gM5l76S8icW391abSyKToUFSzPOCIHzI
v/tpPYaSG9RrDwGqgU9IvJJbaEioDg16bSPORhW0YFH7qC8DrL8AWxZbfFyCRExhe2kI6j3D1Nj3
rlp5ZXWFtvdWi654ZRkTTsfZL9SetDnEhZJb9PcalY8a+haoXGN4IrXMzrqvvN1ilmcIEckCKBzm
lRQ244bvGFA1St/QfNZynPDnmf/Bnu15ifOfo9o+XfQL/w9p+jMwgn9/tjy+9ZSoQeMxOHJMc4vu
zn8nkxoPV4MP9yEIhzrBXJGKjHoMsIA5NwF00zjrD95Oiwh4XnSyldxYIN7lb7DNaKZZcPjOH6G9
reu2REIe/sMvEkbM2n6l6zcSesMxnZqxTI6BA/5nRpuHqwKCW+ck3YcfwV+n3kPyZKNZS7+yVSXs
9mgtxmPqSdSmSfuLYeni2/JxxhChTQJc6RFzBG7+ohAj9Uyw45YXebKbJS5WFoUQxUtW1ZGPvCZQ
qhLg1gsADD+39ZyxjbhMOiUXYqjZw/4euvbflv0Y7+ptOAhOzHUT/cl6gXJRDYdcx90lcevg7P2r
+YBtEEbXKcE1PpU+gUm1KybsgWLoLfCipoxFLF1wXqLKgf4ydPM/61nNfr9qZrfHpTif6PYavE4+
7+r3QP0dOV3kswGZ4LMs3yFKo7iVBy91TYnEVRFwEpz0m7YLjxZ0vySB1lRR3838AtUOwHv1YL4w
pZoWt2pRt9paCXL8mnnJo7DzDDIT0hE5sZTd+W2R3xVoGz67nHK1ESGB2eW/UAqwI+qHSNKRi7+l
3sX1hAwluvjAMWVVViNjoI+2MzRRzYPPtK4RnOsH+nhQyIqt9pLx5bzGfX9S+dx7jVvsy4ABNB4R
pt+IMYy75pfF0jDsDMdD+owVuPioSJ1AobAmiyUu41LMKinygccC3UX1QscqrEeM/yhsJ7NVgcor
cUxI+vzwd1XXWgXnodGXixYvvGhb6gPJ6oeIITYcEs+Zpe8Itgt7eijpyn0NuD7gPj5fibr4XyvN
BN5mvAErQ+9UWNadd57/1N73eFm60BK3FCza96Gjz6TQOIY0Jo2B9UYhk4TNvhkkV+OM7GDrwtAK
sHgKSlvJIp5SPT0vNmYTC6SvDAp+irAbFCnqaUNVLsI/waE1bFlSiwi6a/cGhwyosq7bsxYyQmMb
nbvkoOlXO5BTpcm1LFUPuQtBOiR8MwyAhtG0/Zb4pFeUTGAmYyxCQaNl4moz7R4g6FezkykgdmIn
K2ZW2Mm3/1RkTO1V9btJs4nrBM1zQtAqecc4GaG2r1Jc8htI4CAbsaaTL1WgnM4TOEkgld33+3Y9
lANLkUKI1pxqWrCQzRPkWXsDqLuKuMT9wm/w2bK0wd1iTWhctOB6Z5QzPjVehQvmMLMEp+U1Jmna
dTiXZVMFsVnCeGozG+Rp4eeMJ1Iu0ZiscN7+mZDkZrojMm7lrzI2fBLPrCaq2HGajtWEpumqiqQW
wDvIZ5EX+YLN+qBHOYwlESo4d1f6yOXF1m/UT3pi6n2y/rI5cxXfqTZwHniyOcxdFbpAc1dam2U8
lUGWgNiwbEwxl1Z0aAUXCaj5NycyoyEirCiXXENRe3azXH7mDX47t7REjxhBD4gJaQRTNf2wk0cg
fUcaW0u6j6D08U0y37hF000E5sDfAAe/NVd6bRocpXIJzpk1c8ej/FkrOT5/lsNzWcUKq1KVd4Qn
Z+ieTRh4jevq5aY/31d5fxFy307aZ0k90PevBENpkKaQ/x/hF+v1EVWGFPBdtBtz5vrnVpKEqHf4
us3zuT72/CZaHmgOJtRFaGY/hcF5iQqQRP4G4B5wPOgPPADBZw07aYdy5j0MmSlQFd2SvlxFDdc/
MauWFciEoPWl+zBywnvGE6acEEd/7KJ0xoVx3T/2CPzSOiwy+ogxF+Z8z9lbwJQ2XVWAMFQxYJRF
s5jDElksJDVs2DfniI37qY4M8XqPOvdbqdoaCNU+kyAXwTl7PZY7UtjWQKFDWhPFB+SiGL2TW42w
ABJr5PpsVr1S8wEeR3QyZ0cDyyXMRu4OVAX2z9c+MzWnJP4mUws3XiGsiaodIYqhJ4A6OvTIatr9
35YfncDH6vwido8b+gN35/zknQrQfUh5i9JooqdR18AF6cYszvKTrYqA1s7Qx+Sr0yvT0dexUvtk
dQUN4hOXTpWrB5T4ckpDoeghqoydmzVBbQzzsF+qJk5XdB2Iz2YA6FYWk85YwFwkMlfcVSGp+Csk
hdnTHw9bDihEiuCsIicQcX0R/0scGpyrUIvoqMV3nY2icXrCQeUrN998VBtx7j7eR6r8PNezq4DG
KUMO4Glbl2XCRBSiTeJ1zr6r+2/LKDHcZilohq7hhbZl+chBJRJ3AgQumaxn975l9jRo2iKXUc5/
kH4Km2bGWATbXFTMG3orrh6XiF33LEV4/mPDak07cMP3dPlaktF+bmDrNI93tBG/kDEhj7xWmNU8
lvE1Pu9F1zS1Bzyf6L2D0of1hUyLuy9bOLeiHhdOS89dHQnV3lF4RThhiFax+SjowevlUbPfdZwd
yIE5PBW/nQlO/iEPfmVjA99S3c+SGNYPR8oUCGbW+1uUs3NURJGVca/jcZ09VBeM4sONLpyNjUc2
7tlgXPI0FV3kKwBuRh66v2H04YPEtJ2z7d++xGLkj0BJ4lDalE0PVSgU7LYLasDusIiNWhtS0m7x
2v5kAZTT26rY6MQFlOMvFtTNds8OH/mOWG49QNapjjCY0FgyYhvyHgBpeMmZwIAhSkIuJfW0KSzC
PZ2JP3eJaDdRJT9APu+x18r2Q9YBxwaKUkMIkuX4KuvOdujRczi4p4vaGLdvYabKqEN4kXT51rxE
tcnaYKTuDib1odRfZj77lo6nefDbuikP+mXQhBLvK3a/bxrN9x5sefEmw8Jz9AoVY23vGv6k5lub
w/nl3Y9xhImD4fZbjflXRZkFivOLMyu/jYPJFhugBro00bJZnJ3lUzYI7JUPLxvaYq5nqAyCk4G+
VZL+lXR15hrtArU3xwVKwCAgfyxHobP1uSx3qtWeI9pj29sIPWBs5yenzYY/q8g5oF+WnWqZ1AFM
h7xFqKUpvxktZdBJ8bxK96gqYhPTdPRq1tKY9RwSvbJTsNkKNjLRlq4bv0FKUlTqMhyB/Ed7SwE4
MXNdqPIrsfueG3D+5/ryyz5UFtRuwC/noCdxcCnkpZifYU9xymwcYoEXJOh4tGqVoEvsq20lNn1M
VhlRpKcCkmrLWM1jh0F6XfdDM27OBpyBpBIXLXSNUUOflz/jgNQuSl/nRSrgHuUUYHrxhIrRc3Gx
cIfEppxRw6sfH7GMaNl2WaRrDMIlD/6tenKESxxq0aRGXbN2QnoFpigESIr3IdqAt2biokSxSb2C
QhIxN4SjOUuicW31FCMdDxUqAsdC3HrGsyJHX+OWJBs10jAU1twMQcOcxxn2dTNN+G9gOlXdlYrt
LhEA8d1SvNQcggO77H9T3B6wHrKSoDZ+6nfLaTAzu1Dv2KO7/xBR2Fpb5dxtinhYW8HlD+sSrYtq
kFmMKud2igbdjnwPrNFIfYlbBNAdb5F2PTfxOPwuIOPgzqHOcQUkALGDgB/JI8CgjREGW9g48K0k
bIWtCxMG9C10+uSCYdec4AvDudBmwh2rA93hNZHPYPm0Iai/CsJ4E9mqaRIA5NqKknkQqOkQSf9y
BVbYOnvME0gUaVQQQTfs6I0oBr3wQMifZoWg5uS3IgCtsWFloxj3dOIXiw8S2HUFf6OvkdWjqpZj
YNDOxWB/ZXSy7vEZrnu2V19X74nIWtZw7HgA4ZDKcqJZLlxB9dr2Bac65GaoWb4lRyGDVqYrpACB
2+Ev98UleSmIh5QW+zTB7SxEGBZ+ADO9NGjlKJP6b3zHL4sUZYNvNPboKIfBkXcXj3aKQ7B/6mNL
FDDu1YngQ3PXwwYKG7mjipV/1iZevLXKCLTVamQeQEA+q1Q06Hhz6WzfpIcO6E5ZSdNnyu1RDwLI
JiaC+zwWkTXqh1mkB5tRUdQVJT5EcE9pPMABnIiyuDKDSOiPzVFk0A+e676SAp1BfKyRLgUgDEm4
1KPta7F+q2HtaJwBdbXWgl3XItshIKSrHvUah3bHUbn4rHyxXxWE5qmmHv5rAkYaGaHU16cPMlrS
DVY2EjkOzUCfIyJ7HShUreUS6E5vjEbqtbRe8I89hvshyoT5nDB78/X1aFZdvSVBvmGxROCa8QOL
EuW/gmYhEyv0XO2uerrawf0qUWzUeO0q1kQbiOVyFCWdsqQzsRkHBOw4WNAUhsw0i6StHsGkWD1Q
pn4+dCvvP2b+58d3w4Rwv7xWGuMbGaI2bRjeUFZoiW6pXjg8uTfVv9jetzsoY3Cn8lpaRlXIaKi4
ek6BAZj2u+GAnF3nH4z7z1oHZyrcMWgeGSWUqt1COIx9PwtgwjOSLm3H3x70fKZGKvhbXCEJ7pD2
AYMyco8Ne3Ve/vlbjjGPwZeMtRz8pPagGxw9uT5G7KDF1kccgfrI3oqZbNiADzUDHaadht+/Pblb
HcFDCsosbOPbngLPnnmpF59h5iqmvIWHTTjki5Qyk3Lz+bd7xnsuzT8PSc/F6MyMJKVuGT01FFdA
PRiJyZBfgMI9es+fCAEY5o6unFOzs75NZNoGKpbjPfC5K/wnB92mWSYx0zegHd91+QV8INIQbd9s
3CB7A4ABiENKdg5yTfzgsWv8K0IAD96ppBzPDIW+X0P+U97OWmvGepP72v+yZio87Lo8BfiwuNR2
cB7luNqeo9G/kICk3rvF3SxYKe/nTVlIvSOpZVFb1tAlbI9N9eAoZybOJnNBV9oQyIk+m7d2icey
rA6BazDUusZIjN6xw7KkPodadle0HKEPD1ZTOGZ3NRNVF6CDdulgmCg/nwBkjzgQ5qlidLkCdINJ
2zlqkzYn3+qsBYvUWgnCDt5REkE8dvvHcUs+C8/njYH8jL5T3pKKgCzc5bXkWng6adgX5RT699uS
xGUK4Y3JnP0BIsdv3/5S7FQo3hWwujSwSo28GqLN0J6yJUBKhQf+EIxU7vfLVHbLZo7xRkFluA68
FISSM8/hrCSIBq1SwdHZhh/95PSRZjuqICeE1hDVh+vdkrq9HGur5HsTDMDlVFjxub73G0XB3L1G
g3KqW1yIYOcVEwo40JjG6partoWiZVArMIBQUHT5W1H+Hos5/kqwCtucYDJjUqpY71HRh+m5UKMN
vDH+YQ3nBL0Kmdc2Coyooeu6qppgNNw5qFsSTI8wt043eXtwAJdQaKOc2wPxGRAigV/4UMtbGm9P
IvstRrYzQlBwueY/2vU0ISpNkrsHY/qDhBntL+Y2RIYmCyb6iHtg3JDWqGOPE+5QOLxYFNkY9Z6y
NfDXtci8yQ85Jn5IilmlMSaJsxHUWYiKDwx6MXXYGBBkfJ0VAMwbfnX1G3L0XnMatHXdiIoXX0m2
4kFtZSfGvp/sNP2yVm5gigP1hOSjTDQV9pKJ1VB7ojdXvAN1tiM+kxppjWCI3eF6aDbQQhO0H6v1
hwHVngYVeDDc0whCGEUv+vGkqHvoZUJYxmkw5x+LvKkxZ0zYYOXdWRDdxqmc1RWcNTtf1ol7ffK6
DthNMv7bFW4moUPGwCSlr09SEpws4pIIVUcLOfATbxWijClxEKgJxVE1JobwNAf96g0L2i0vRO96
nbPp7l2hytCJ0OsnGkUk+FBe7lNaebaWopoFNACCh7SvgJh+5U3av6EvCRyzlWUF9kikfQCIWYQl
619lOSxZWp6CIIN1G8sT/GFzzlKlJhJ4KYXrKmK3Et344SmYgG6z446ZW8URhIsCcSM7MeT98KFh
gp4yymKm7X1HTjdnaxYNGJwyGnW3IHqKGI91nvGBBe47SbClVk8JCeb8Aa3il0AlH+OdX/LK+JhA
r8C2cxTmgPR2BbEQXcuHkz3N6qUHVSpkpTTSR3j1/dr/kcq5v+rD3dKKcHAQFxRs5768Qvf1lidl
0aowqJH1o3yvsZpt7LOysbGeRutD1+B/jidYiPouysfxxmw1YJt8GVayE1hIkHvkv+mQzBsj//oG
go3lcUlxK8kbpqAiUEMG5P+lCIZLOYNwiVo0g4km0w1wGTo9lIoAEgXSNfAhRN46pUgqCzp5yYHt
rtuium3FmhBQJtzJfHsOgyisZDSWW5C1qB1yKBtG0b9QNVIyoGuFLZy9cPOSmZHrYV8j9M5cwocb
7w8jAuNwX3Pel0LOv/S0zRTsjkIbnGybB8FziWqROh8NmyvSRpaQYQx/V1MrRWI51KfZSHPBbuB8
mfphGI+vz0NpqovFJ2hRK8qxnfDIJi3hvkpwYtlPsTXOd+zS9/ntYAKuPYD5q7IUFXT4UB0Kt3Qa
PgVpwYidcH6B/AOq+g/NpoJtsWFZ1x7funSiCofgsAJWPLbZR7qqvTv3LZDD+ErCsJPRTNakHl1m
OFhvQSRE9vQyvVSKLnTA10APcmXcgmN6lnxvHBLMi3/mbnZEkH3HAWpLNnV03jZ3bvsfWg0FsDz/
n3JsxNtBCszsa5Mf58W+IVu6mFQdZU4QuK+MZ88oFh+HjK405SanbHrHruyJDqg+C2P+htMoSg+E
nrxUI6Zhb4eMOkAE0dIahywaJNCx96skYL3zLpelULXU14fkP0UkWH1h7nvIRNOM8bNE5ZmCdvoe
rRnRMQv8ODIKZBYPxFJNIbXbphO2Z1mp6lT0P5HFxUvJ+QtYCdPilWjDGp8BcrS35hacCzL8mSBF
3Mfo6wV5fN9FYsjGwcWRhqV6SIKs8F92s3JVGQKkLiYHyy9u3Ch5zSR3rvnoJ+4eAwye4CS7h+h8
zq5HUci7O5jzYYUr7MOZEQcBbjIDYiryR3p5T9RlA1TWd8y4BQb6LZnVZFSQCDRmKbKVd7QplDU5
2jK4EkRNXLs+dvLD/FUe4M9ReJH1GayFHR8Jv/M8ooW+OPyndYfCJ0EiEtZ/92LhsLM1uyjPA5Xp
K3MUIWP7U2OyFWlznGaZgxKHwYLUtuVbmsvfQ3L9054rlrYLPwgnA5PA6LOY/ATGJLAjUmkf8Mr8
MjcV+92NejO+H59/DwTWwxRoqc4LS4AZ0pu1JSsonB7Wf7kgBu07rnt4+Rbf5VOwQq7Vvb2+jqrH
MyEs1rOSpczlA4eIA7bk/GHvcfQiN4wx0/FrMQzOZUIGRZVTe+0wgkbZK+wFZutx3ug4ALSrtlsR
aUU+LmV2vCBqgjmRj+dY2W6DsnMa3CVvNhP5Pccr743h4wdNP981hbkjnsImQourvVDqJSfp3vUi
8cDJ/fMvL8QF7PRsE0KGKMCiGyB3JiqEbi6mEz12E4vrRhVYc5yUNbVx0mGPHH/BuNUNIQ+7Ddjz
sVBAXyM+4ZtFA7h7jiF/kn9PY1ZDbfb+WPdseyucLOI4Qr8FHNeuvKUcbs/CeaYEa87Gc4zV6Alh
lhqFtOF6DFx77KNqlzET15l3eih+P/bCcekZAaw3DRHfXLn7b9RQWavIwA7cyFqIXuIBO4F3JEz0
WFwtQ9rqFoU9OevCHpTXc6aH3RGpHQGrFUEvcnr1oNMPzoolKVavGKLhOsJFPt5NDyAFNFouWwsT
hB7ameXGneWl3edHKpa03WeATKeeIBT/qIcJNUKiH0y3tYja2QOMXFosSPFHJLCnTwo1NDU+m5y6
4THSDqXkjhPAX1Yg3BIAkynN+3ISbe2Lc/fu3ve50M7wYKz6pAbkJ41duZcuAO9MJtJo+i4Df0oD
/1J2PNEtKhk+uV4ab4UouUL8wojN+K13sj+eHSaep3ixyv5q2/T24VwooiY3vK4s/XHtNvYlpCYi
cCqmaAOxmv95Cl/avdQojhSLNWSVsvFnoDM/mDJJhD58sWIJ0xhx85uu+glwYKzWWJfuTgSeaKc0
3Fi/Ze0sbcPiW083kQflOhkGPTepKi/Lio31Vhij2imEeLltXNQ7nSgybk9I4IxFRTCcVnYdKKyJ
cdMMaHXXqeApMJ4aAgxiBNEiiiFR+2hDgvFT38vHMFYmw6zAiL8kLEyXtLGbWLcgxRs6/+/m+YTi
SP9aAxQqiDAT1FeGYWYM2Aw9Zt/utDPPyfm75yQcGae4vZfqP2rRGv2AZgQhepvTfAfSbmAWryZ0
piATWdTka28PX7Q0CfgQIoqFuQE5PFnbZC5s7+nao9Knu/vwLUr6LVyvqzfYJ051lCprNoDm5WyT
IHyxtEkj1mM3W29RwQMdMpw7V3TZorE14NZiLlY1XAsNdjQ/2RcHHVoUtO8cY0SWfvzxluoz3MXY
/oXJjXHZDHYcdtZ/futTZHaxjfl24HBIwZxy/bBiWd8hvcLHRyghUl27xQmnp/mKVuX7vfNqVggk
CM3NG4Txz/Xz0PtmqO8azqN/PDdiRov+QPSJ+BGeytpGUxTZTHt5UyDObZhK8YfqhGZBwUKQ67UZ
KrOc+xrofafjQ4XDBZyDGiWaHifhb6Gt8+ab4Fu0ZhAmvqBP/Ku2ch6rqHpirdQ9HcFWDPm1mBqK
NNgNCLMkMnbc8UqjnwWPZnu93v+WgGAO2CEA3D7Qo3A/r53H7LVQ12afwUKoomAi0un62vlxmDAf
Lj9iZYCcqZoT8lrMgK0EPyL0UHeKCXRZfJYVoKIinbryZ1JrITVreK28XP0QmueUv+WxjsJ9YDWB
KzpqIDyVjvEi5DaBSbmGSY8WG5OAwuhXaUo/pirZJ1s6zyxV7zUhL+7lCKaE0LzBvgfZk3gFGe4W
Yh702JdOlcpvWus1WVbAWamKbLEdb6ekondh7CXP08aqIM+Hv/gF3rpJPffdxli8Gxk+4iO52hsv
+RWCv6IItvKgm5GrNpSg7ysFkUpUa5x+BeumK9K7p9v3c8UPbczWBBA1me80OOyoJezlJqO9qZHL
f0ocneWDq8/QNvUTqDC/WNiD6W/Z1Mq1RHcAu68+hkPj1K29aZTAO7iI5ECPQti25G3t1/RbTFCu
wK2XP14I0Vu6c8cUdpdeNOk23mghFYzoo74MqhI+SNZovXeU1LJc1tkwlDWZTWmhdxFdsFau11AZ
xedqNG+6gXju2DO0X/e9gahBpSTda+vQg5ysoy2HXX7myRF24cTp7H6dzkQoGekR5iMZ9SZjpkjB
Ic+lWEQuW8EkQlM8noPjWSt0Vx8l4t1CkEt3Ivr5TCITWSYSeFOz9ugnjef5J9KujCMv3cjtyNfr
Dt/Iver5E48HCJ1HigA5eM9XyIFfeEDEfdx/wtBZozeteJKG6SzzUDSJBSuV9pf0PMUxJb30H9q7
tq35Zv8hjm/S1gSLPLauvcI5Ral+NkgNw4rFJaYUGmJAIazEs70hPTmA+9k2sawyu5n5cColrE3Y
YrAhP8yB5Nvd+rT1PL0vUTDbXfFR++v99gasWfZGDeY4lUS2ZnTdCaCI+zIFClFAo4BjHfJUx5ZG
IadQh8tD/xqNIpRqwEm67soQxxdYzYpOSOdDTGqngaFAghc9pzfHNsQdezQaH93XO1U8QXmVNNhM
92mlyH9NYAoZtuDo1CKaEa3MeoUVtMNhgHOqOWaaUauMMmBJgyUQuyU8ALSjAqXqsVxXOlHcefZd
lAPdT77SzKQEFWdzqcEnPIoDwHuLSWKVuoiVUvG84XNum43mn66reOenbfIJXvWo7ekpQ4O/etWh
qWW/dfSjR/cp/VRHVqXzrnSd6ylyx5sZBJhFXgGGrRA1SWyv8YqVHGdo9BwsiXcEJuyattB64xsf
TXeOPfdRqXY9Esc4Jdh3Q50t098ltQmq1BiYpPPdAnuMsRhwKoNoZ/HRg2jm4lrLP+tHkk21aiUO
ygvyAqtWy9T1Ofaw2T88CmRhFQfysrcxWthfrAew5LkbHYlXsLnZgnVteGhP8af0/5BpLmoD/ON6
PBsw22vSh7HvN5pbDgZO0onP/zpaChgZFVD/Thk4Sx0WPMd1ci4SkBujWtMa8Pcxd6Pb/+mZcthL
vyEohm7achbc3gM8C8yD49XyNo+VQse3K843fXt519YGZCm4v23BlzX7zLiunxujnf2Kzy88wztb
RpsE3vV4r9xJiS4dED1bG2ARXbzr573ZfObcgAqQ+Eg0HMWK8hDUiB5VA6W04QBIestuOKU9RzRv
p+5zthahldnz/wzzHJDXqv5pMI1JZ5J2mhrWH0hehscIkC0Q02qDod2/36uiRvW+p8KbQbMywqNH
WoxXayhy8MNiEiLe4ojfQVVLHuo/jlxd9ev8yt/BDWrniyRSKXodOflF1fzabpXLcr8Ovt2lORxJ
doA1vuUhFFuBEY1oABmKLkgsun4trkOlw8v/uo+AfHgeISC4MPd/C31Q3QDzQIkuvbvr//iqUzBk
IAVAHZ9ebRBEM2TZ7xafZukyRO4WFdh3hSEMdYQ+9aNxvHLfxwsHuYwsiMNJtIM4ufhoS+vHNOzQ
Dz6KftEDckiWJQWwffmviKQE49wJzF5IpONVH5TuavI2UECRxEQ9VH1fH2QVLmSxF9sYbkZP8KHs
zE2nmpG7d4alqNuUUFzbH7x3opfIQr+MyluvwfWb2gFjHmb05KxozmbT9EeejVHxW27vH3bl3kLF
HleCwYI6VCv98wKGwFZ5aKlWqYnlEgtZLfQz+7DfsdZznVAlkcwbFLUI9pHJ6V+l7PEL6ZjmBQc4
Q3qR83pWG5crABrpsnJ5aCo0SsmjPSxDQ4j+jaT9X1MJr1cJdBiWRA8qa4eUrIwxWdRohMaDkdxl
P6JPxFSdyxXEfyTZhcsOSq6NkN3bulZKGPlpsnnYQbJHUSMdX5+sWo2VaDb8umPUiJiQ+Dtxy5ql
fOe3VRLg6yXognCInmOvzD9YhYhYfVPKdKxLgHONsMp6FPgts46pr4r/zeb+knRx66yq2V3OL3MJ
KUdEvwZQ0uyGLzS90CXZO1MM5bHBD2s/1XEwhEtUoSykQCVgEC2lz9zGS1A76NXWiJ5HmuXuF5vv
Z2vunGwZHbIa1b1NFdqaGsnyrgCIqW4dFxOSS0gM8Tn9zWxErQr1wosUyI+ro0kxhvVwgCmH+adV
8qutCLxfOaoDVPyZdrof+jiuEtR9g/mt3x7NYlSkuziXYlUpVdZsp/m+cdOGFymSuJZ9UZlShm3F
LLQcxmZoXP6XY3D+ZJDlVjpPNLPuuJ99+SRoUIX7awGqZLU71RMoiV1QZu2TzYCHJ8FGagTij5kz
Z1kAVdLDslYdcDdDMr11XaEZ3SiwN2H4g/ES/9Eb3dC15GH8YUyJFGBBUV50wrPqvJGNFS9bT4ZZ
lKa1lIKdlOBkzIimUfe38XXE3EqQO6nobDihYnQUgKQjZT2PWPkRFu0C25Fe/zJf5GgqRHr4WxLa
rt4ZbCE5u8IRxaH9pcFQzJrU5yCGpsFpkz2jAkGW2oS54magqDy/kEhTKHQW+SxR+e3O6jkz8HK0
cqh/4SuZgxwM1X0qVxCr8z6Nrerj06nutS8gpJmwWmxNOfr8o8HP7MZ52xJlvxAVUMdBeDgWLM0q
1amyAfePZC7peVx+59xownUKVdQ8HpA+QGK1UIHMh9ey7K5qNfi13w+flbf8osHwTo2motnIfXOw
HaTBfdt1nfTNuYWD5F6x7yB96+QwioL2a+syvMs0Q8Xf4FCRBDdq2gUbKCSSpegL1PmzOUZETHHZ
0TgxM5wW3tq1erUQXpazl43s2cd1+nNGgvOXZZYdM/BIMCjfC+91Wg4SuS3s/WlPEx/0UHJIOAH2
NBmXRxAuYz34XNHaIYJ8r+XjODEBdMpueF2buz8FSxBBz+L4unpwnwWbfgl8tx45JHqI84skFz0G
Fv37S2UqhLJsa+j2K1pxEe6BOXMd01AVYj7HFOU6heBYwQLEnNUiV87q2CtmaqiOzESiQNhnO88s
NOuT/InfjMhRUACbjm14YZ4eyaqpVNTGnVan1u3Y/CFbbqf6qPNet0xZph1onwkaKiTNKBua8Mty
qPEWG5VkfkBzIv9KJPcg2aZlhJplIyzJe1FLfihpW6Pfnk+FAu5+KKch03/2a8nD0qzqcXIHr+jo
CXUy0SJcsDgob6cKik4fTfaKHlZqsjsBKQUgRGDyxQBHLS1zz9DASRRTgXiEqIE+YEjz5XZQ/rQ1
R165laO/Ge6WjfR1p7gjbse0/+c8SJ46SbKAETlk5JiQrikWoeby758L3uPmxhPXWJrf4qipXInB
0S/HNTHfc9NQZno+WDwGlB3c9ierkzG8frX7O6UA8WGNndy1SLhIaCYqbvpgTW0XD0uDo1J0eDED
l+B6fn9Tk+9nf3ATu8+t9VAaqVBc3mPjm7SGbgqVuKNm1JePncQKLJJfCAW2YafDewAfg1vd9b4t
WGA5Z7RcQtYJf1Ss2xoPx8vSls7t4r0eOLOaECzoWWzGWhA6YRU+ql3iU2OhL8CqDintMSP2FGDb
/vc4BlpvkwJbSjQSNtFsWB6MJ3ec7QF3dQ6mSyL0NMweaDimLUCNdAPXsM+64LaIzE82s6Kcj2ft
o3noHPT3LFYUQt9OKDWWmkfw+sHSkA+lsKTTeaOL/apLQhpIrfTLHL3Axqy4NEIphiGKWWCcLHRc
NsSqhw+aDje6LEeMI9oYBlv7l4rTbVJiH5HASx8N3F1RYUu46lhlXQwIXHffxAWIcdNGYwh6ssEM
/cVuEv+9sg57PRx+aWTIAl3ZKbit/unExcYBXxNFL/UDCOUEdufIxLywuFfP92kiwfBfmBZ9JCRq
qkx32EJ/Q3zxiU5+3uiFYzwv5oJEgni7i+Jve7F7k5RlFXxDKiM1fDf8Gb4/cYW7OvgXpB/30zdi
oYKiZ5SHJ+zijRBxIRZKr+rPRSxQiU7gHnvMIDqmxipG7Oqq0jvRCbRO6YQHgl0jW4Vi/kzsTBRG
yVkVWJZFn5WMbDdSDUDvA3CaJuaMhHdxvmsjh0/QKM31akk5RMx/VzSD2KNlKJ8Z5I+DETXkvKL/
VDZsEnjqdcZezlmdZPnCNCp9eSuSh8gGqdmx7DDxu0PIka91kBtwNrVPo18OX9d0uSKntX1YsOnZ
7REoWAPKLFIEHwQ+06Lo+DiMNWaIceDllX8WSeRSTC9uhb0+ArGhy5+dkp9KY2dzXpzWtWwCiJap
9eFVb+hrkysG2TcXbHwBQc0nmS6TRKBQYEAfdPj+4DxkOU8pQXmHkHN7AgZMNX+AEfQevImleUeA
sYUE2pAfpzRFZu0phIykUgmqCeelRWKktYxMEWtdm8BdcCqX7yodD/9zIpNrQWEqRqyIh1gqdTeD
v1RtJ4WrHVoMXlkzx5OePPa7lrTW1p4EVZH2OnaxRl0qnYb/fP7ihslhTv2/AcLYVLlgCFiRtAAh
3uitAXCNxxb+TInspSu7xAIGIlU8AI3j+Yh102dQzc3T/7u5NZGMPPXV1XJKjc6UL71jYvrdDdCX
azmT/aEBwlGQBqFMML9CGZ7Ve/mtvXqxMeHMqnmhG+eJPcFB1CE011NwQAPiG9bQoYt4hCXgDbZD
CytUXGx6GDxaPfVWRiJQX1SbccqsRie7n7yVwyzuypRKC0G+ZgVaxETTMEwSMLD8HlFWWCCk5MJt
tqp4ZWzL1cua4/Bz1W3MA32/h7y9jQwT6YptgX2A2zV93xUnqQ5x37UnCgZmQJba5XzR4Y9QzFvs
UfQBVxaevVbkpQauu9TicAr2+UmwpERpbIEppKqfS4dwu4vsl/E7it1UBcUpMAUBnQ+yICX5EnCv
cj3eQXaSnwuwE7N8hokOI/yesUuXPYYtC4xLSMTyd4ycnXuZm4sH1HYxw83bwvKaMTEIUaD38Efi
B2PlSz5KKTReqBpOJigXn2M5pAvNrfO8zTStH63IG7bJ7gmFIibqcWfNbgLFrkFnMfTW4MgfV/lC
USw5ebw9UJ477Ibu1HxBKrw3z0Lk9K7VqGaBI0iC5EQKIAQAK0rJ+t6iENnKj2lC/7/MFCkujYei
hj7BQllR4MfXvKG7qpoLXji70Po3sKloURfhHpZnC2SI5SIfow3Wx4+eMl9Vem0UTV3pcW7Qw8jR
6X8yzzEDdpqCfThEfz7TjZr3hWlaFYuvNrgXSDtOKfGYtLO9vJKMpsYUXuGm+X6Usld2KX/WmZ4B
POUQ91f75GcK+NT4G8jvKBrZEFxz22XrbHuhfjjbaW8btglDNLoDgmxnIv8MVXiG8at+9S+p4zZP
XK0TqvVNo4QRpxOJUyCQ4FsGXsC6lkN+SWogK76JLVUyLBPcQ3OGZr9kVYWF7oLEuZ5RzqXt9dFA
H9WKQCmOlnHf6GWLEmBFrVTE1m/pNvhx9Bjg4PwbuQw0Y0GF818XEdpIOGIwhH+xHkgcr8bwexaF
Eb50zp7eFVE+lKVJcfqqFsmVgLH4lTYfBmzYFtMWyZM1aSGZHFaS9EPCGW6XKuenhKiIExbIlcUD
YY95AHa0I0TcHeQcZrkG9FZBaAzTiu5XQXucu0jSzeYGyrDZR7B7KHSVWy2rzYlpxDz2ale26dfq
SxfU7lxKXh+tvhqAAEqdM7vPpAVfJtz4qsO0itDQ9o7bkKbFm7+cVBhDPypmp7tO+pcBIRyvE9jr
v1BBV5ziNcweg91BShBR84iDZx1hL41eHk8HNvuXmHp6SWP7xI/qE2xurepHxaxwOrr2ohH46Owp
boe/QCXanf35S3p1F0I5WTCoKCuJzTy5gyAJqqkbFPrTjujfbwuODvly6W9xZ9aUUzbV38UAMSD2
jzw4O2gHCW+ul48F6PU6SKM/uxQypNP43X+sbeL4M11sjkgbJ4ILLobFCLgxCAGmAuAn5PZKahrd
HSrXLYxEXZUKgOHFmWQ/snzqb+IN1qZoJq/6GrqjdnQ7AbfB2u+sTPPVthb8W6YR1x3PVDyHCX18
7ga+mIH+PrkCyLgzZ4NeNLY6Pd6qvDH8x0pyWY8jUfGfsTGgbw5i8aYhBRS7qt4cLd1cIRLCfOFn
PopEYa6hUETf9w/N1vKnNqBXSBWDQwEwy7kAqk5QYtiW+T6fx1if+I+RslE0ladXoilRWGYQmr+Q
1JjpGH3+Z3HqxHrgDhox9DiJhEPIg4162NeqmTI8l4yFhiSYo1l16rn8XOPq5LeoU2+Xo2tS0CoH
zgwBxeUaMLMnH/YdHW8zNxMAPtfpAV/TXmE8XSRRudRbz+PMeySETIHe+S+6tFzAaHu6qFTdUAUt
ngA34VETV0L5W896vb8fafGcJBwq5yNbQjd4Khwz/D+klvVJpvEZdwr0J8Yn5YaJw6TcmfHhoR6j
MSKFgxBJ2EZ0LLfNI2Hl3ZP4tY8jCOBCOzFVyysDIbf578aHizC9bxXjde8Gu6hRcg18E/+JHWFw
AxmEKEn6aCgtTyVBNN8VuNE4MoX7FkPNYJ5vQxoMOfR/gRakdPUAL5WoQ+tCm4/zlIDUMfSXuUAL
YF2GLdXKxzf7dbK81YWknL8duwSneCxDaAzpWrnh1WE+qz1tH3bu7rtgbTuQHn05Tyn8jTgQOGxN
KsDzbPpIQlb+Kg/eYqo3rC1jGJkU5dxTnnjfoPHzVXBWL7EJdN8nGT9eKbny5Au4O7PCteufwDa7
43kFvFQsHsFsVMeiauRuspmrjoGHO4v3oFrXEo8n+B+UB8J5Ql/CGHPDn2GWFhYh5fC+MvboWlRt
e0+ooWXDdYgHCKJ8EeooTPcN2Zvg3YYGBmrI4OVBvucwlwR0JI5al/aiEUpupbJ86FCG9jG3j0KK
Zaz5TGGwV0Yao1L8BuXhW62ZOycZDwth51SGBCBq8JbNYS+Zjw4ihaPxl93cWQR5aJJLXR/lFaAp
5rg+Vp3/zjz+hARE7O+6ylPl+vC5h1zsdLmasH3TeArHxKuV7O8tBHlSTuMG4ASoTWWYJo5YcscL
+MZRS+kb7FyyTzm8zAZtPURPnfxtUvnTF2I9S1UkDdMGgTsODvQBiz2VxUZkvbd4u8Ob5TWMt/zf
0O655aR/PmgqM28JR8UccpMYgE+0xK31Kx3a4zFfRB38Kizj6R+lSFoqOLQtkC/2uwwuwWHLDtcH
nCwyVg9WylxqRdw8evU4NVr8hJYb0oPIJ0wBPdRqlr6h/JHRGRCxFKym8Ywk3+KARX8VyR/WTAp0
BwCyz84rM9vKt3dxP7x2y+MydF19p9m5sKY49l6lLK9fvT4EgrCvplk5M+2JdbOR6VehD63CZMRj
qgjMLYx8vpqBg8TDgcnwa2+dCkjslfhv/TxmWSAKeR/KNLqWUHOnoo2Cia+DCpGgy3EzmTuV73OA
4EXPPOYc36iowfOFSHB/pglU83PPrRV3S6P7d9mg77S4berTW7fZg7ZpGd8FlmL508H6xGV5HhQF
N6rFPXMqYAfJYtF9dHBRUIvA6RjJ1fcbXkUas6gAPqSjwRimG1o9LFTgRBQVge0HEV4R0VvgUuwx
y7Oq9bradnM36S0zLpjAyXHLvCWUeMvtTQrL9GfAOMV8bVUy8HHVlltFqf4NGM/co8O2q/oaezI5
+ITOVkq4lXPM6M4Waa+pXck25547wnCOFznabozj3lU8etolV9r/CC9e6MAZV4F4vhnKILHr9hZj
7g9tnq5EFh7+a+SVHLUVifPaNu8uNXZwc4CX+EY7cdYD6EERhzaeHgBZ7LFki/EYEScEMRtqLm/Q
SwZGir11oaEmR4nARnZH9SZJHW9GOOXllwe834CUsWe97Fsi9A+4qLxEnQj3+bxqfXegYT+hMUfP
V1O5aLiUx7fbaV0BwG5m1LED1egwP1TpnrXBCZROb37yS5NeJn7XLEUL5yLtF/3nBXG7+H0m0O9U
6QxvOyjci8Ppk51Xuf1y2DmNJuY1SUtDhu2UyK6ImmoWmF1kUwGl9p9wAQlfqdXPumFKtxRrPRY6
EO+CCj8pdHNG0UxRyph4rmyFxiqzRk8vHfEkGeyC1WLQDb1eum+jwawRozgEYvg9kbzb8CtxSn7q
0k8gDzqwRJgYoFnjKILG8/n03fsr65Vy90RD6p3VcrtFozaI0EV+/bxMsxgFoudgZd/87zws34or
9okE4TR2ZUgkWHHYmN6XewknGk50vp/Vg7nHsX6JNP75L0dUFsgCCZ0feJHldfgiizsjxWbIU8Pa
6rf7Pn8XP3kx1QWltQn3ZUlAqUostWzSljhhHk683Ubc1jtGNwge2JFpla3YHZvhtnENcOuwVat8
39DjA0Vr34O68bGcw/1Glr65H4+DcIaW87MA0hQBcsrYkMDC2c7NP1H6ecVt/j/1qHuHS4cIRHiN
2M2YUWVnwGG1PCmVMEDsRXZCmSRfREVKtzehFhrcjzGSJnU94TC3r+htGd8MMKa/g6qC8ibfA/Md
YfBMxrl5F8Mwk9KbDAYo5pDbxn/tqbTZdokzS5uHmKOjlawjAii+xJ0VjsXf9bN9YlDZswQURoWw
A9eht4MZhhE6an8KVMzxXe0hU9ltGEinzB4e8REJbgCTmFmsvvv6TG0gg1pTAsrTNUTcqdh6dIgy
Wdaj/fhh1gOdfXQxUEhzAcrVT6iOt2GXRGR016T8ee1KIlhRsRgM+2gyrngxnPRusazkc6LJEkI7
dXLx+39td2PO9Zk1ScBkOTuimO+kFOHHy5RmEa75U65jzWoW858/l2oK5pATSbzOfmKti7Amip/s
C8osGBcvdh0jK3zE0eZRZPIWD9bCnIQjccopliq8jsFalVggqW4nh839gTzLiXS6DELYC7DzbT4y
+C8r5AYddTpXlyXkIlOLqyTVrMmesI00TS4iRfMmdsgAptFoJdS1EnGN9drXPJGX3omozJ+dLeGm
gZ03FcC9hGwpiUV9293wnC4RF7uVsFFdsEDgiE/gYfRlw0CJIVKwgoBnNLprN5g+6jP7ppE5GttC
jMpHRmheTs7somKv7iq+8opeRTK67cqc1dFBbVxewDLoy1L0yzmTGZujKJwdllp5KbAWnpqajRl9
pHypiMMYs8/s8ENAz5pvZxW9flmuqjQeu31z3rg3YFKN3PcPCineYJ0S3J212oSoDTpGwXY8YwUn
BgD0Y8Ty9hQWPLtwwS/wiz+it8lrzs63rmkJv3WEhcz7QZIA7opY8NmSFdoRQrRvJGW4AT7vcRZi
YNaFj4SmGJ5nQiEiVh2e0qtG56TPFupONQVg/KOoYGv0qYdVLT7TSX7iRXd6CJ90UaJ59zJDjJfO
WgImpQKoGIffCDurq64humq4p1jC1TXKsD5cMlVIybfIEw7bGT7NgOup2UC4bJ8QSFw1PvHQ9ygi
FuVx7So80PsfIuPYxZcA1/LKSd/PZeXthBsr2CjhZFb4UioJwtE5ilgemsqXMP6FqfbpXOMnJ7ts
PE9bjgcUEhN9BjmvCruEWkp9I6e7jbtRPaszwx3Mpu6MupI8Jh2ehbEHbeYDGb6Z6fLseeP4ECCb
RfBKCpvYel3KaDt0Mxe6pNUsQZgJJt8KV7vJu6OaYCqTc6hnGi8zgJhrMFdNMc1nK1J7f80pL7r/
AYK9Q1wnc1T/qSYQ4oZ54vXXEA878BFJfh8fAkwrzxakhLBEs/FeZAkgjXDgZ4pD0FfcD599KZ1O
8FQAtBYpECW7TP6E73JPrvLOTTK5gU92dO/hfLcvmiXBrKawqgmNrmU3oC3SwAAQ6PBFJI4MVyOz
md7l0rdlSQ9cEGdii9lTj2/SzJtvHdAxBhR3K2JotAKZKmos5BIsta97MU7OCc5yvfiHU+dX/uj9
/sAV16uvbl8mhLMkGH5CbdlVY70fc8Be2w+2rJ64TsifNhjJyrwElxbrHTw5kTL0ta3vwwKvVvn/
3F9UreSASFr9KHHhhwIkx6c1qIMT11cst2CP8NWfXF4a+pbzroztiWO6Z44X5WHdgeT57HHXiTeA
5pqAuTyJIQUXkLOY0dt1rLtSEbXS3fVRz+jsP99gKbZNVBsKQtbS/Fml+nCxWJQJabKyNnCPr4Zv
CFl1MCmOyxx4rIDeG8wiolLH5fLCFIK+ARx16eQP+QguZUDzRxg3UEakakPImy9ShpAMeDtIBynC
X3ztoHH++qnSCKcgU/ACbC01aFRwG44hG48qg1wzYz6rDCYlPAvKuWlg9McxisUVNgI7F0T3zFXw
FtQZeGkFIqgJjRPHWEvjsaZcM3Tbs5PByg9mLG8gqovl7jNWXWRVQcsjpi2D4A8vC50gC0k0M7+2
B0+XQWFVafGhxoQYHTAzciZED/fcPAcz943es6lT5UVM+Gqj6oxP5fK4XKnrMvG2nzAn7SDrPVbY
9eKdGiOAycq+MM9QFnsFnkYUTR/FlnEsK88z9szqv7i0wcQgEy2Ej2+OLpL1GZ4VcbzfDeFYnW+7
QyX+4S/AzMVjkLj5TyKs0KnMX9gcnBlQoLtkguyKJu1rh15NxZtOvHl28YH2KU0QstEcypFUhFuM
yzjvIwZ7nGlarxevfSBkounO5XC35DIrEU05VKRQJY6wEB07J8KKwMs3xtCB0y0WJKjQnMdLVpr4
kjcdnKTOXt+L796vJK/b4fzbVCPqfkNaJQgpV6j8v6Mdo/cJrUbeBXvbFTd71PPy5sSgrShaAK4Y
Rtmu+JUWtavMsb3mzOYoW/gR2cRhal04XqapNCyZzutfVJ8NdL/KqO90HAVRPAsDl7df9Ec2LjSl
T+WBx1G2Ye2dnevtrhPJR/odL8IVTO3835F2rqXaoZ/nJdSpMmhbd9OXPgqfWN/O92dUDPWc5HF7
Y4GcpboD7EbJdliTops6ZWTv1DcdX4pYZ6ovPh3qbxMU1amw5D3Tto8Sb9Mtv1UWWfifM+ELxpKI
WSzqn+A6YvrUTyMyRQZOA12VPtEkC5lshBGzDR5IexQUgt+5j7q1GPtGlohZnDpv6jv8QFC7uDx2
yPu/pJriBRh8XXdDaBdaLI+JptiZOND4M1vax6C5IXVj4P3ZXkrnb5sE6HbJxlCduJW1ofGc8CbS
D8ikClBXI4wngqDkNGPggIG1rR+VstVrv2x6s7Crttl3U+GvczOcpmmLY0oBVc4SaEs+WYjHUewd
ilW4K1FAZn9Ja5viuZkLEaRWbMUGTLAbBJIJShqEelCl672LNxd9XfSS3wkyFAWJjYgMvNKiqBKa
SQfgGELjarUMvG/Qmn3JETA+/fAeE7Sa97MJulPPyF6luiT4WkKjOWTDyEQVn2wzYbBKdqMdkYDq
ComBA7wmMAXjKqXZEoDgiVbCYof5tEqgoBOpQfPIEKOKh0P6kWwCbb89wanHgVh8/Wi149otLqBE
NwoRAHdf7NNhoIOvX7MEUGO1L8zGqCvZrGC8U8dwXVNoCTJLGv7acIVQZvhIGmZtZWt+FFsDFF4C
x4oz+VrelSUapW0IgQL1jVn6Iktfv4Ogo4PvEYaUWqlS6bf0NHKo94Np9Lhj2jmlzIa5ZFjihcLw
nv7zMxqzZsWPWYYjyImaZDjTryf1vmCe3rgCEqEgybBWlJ4AtEKo0Y497aEgH8jFkRiTzI4rjNjU
Pi/qMjLWdv9T95xsdXEaG6UKiiIOp2fW6bYG5L8+rH39oufXkhEIlvenz91ILXgvOBrm6RYwaYNy
cPdjtHh0gAi8AGDZzK2+6dQ0p2J3QAzZBnp7JiC4v1FPC54DCyefV0QgHFnZAAEScpfKMZMkKxiG
PDtINwwgz4AUyVjSuWf98Gz2dRUI08tWXtvYfB2EHK6GdpY2GziJM/K1dwafy42GRld+dsyYuRI1
OI38qLrAPxV+OgL45pdmkmCKLY1lJv5s5DOJ2gSy1rfLTHk6hYDIUxdz3Cfa/MfVklMukDhZuio+
JHWnfujqv7toe7AaXFhuH9Fw0QBsP5dfZSSol+YzQcck/w6nyEam+pbxWOweMA14fvUEPsCBI9NS
762wTUml11d0CjawmlkLeu/EMKKriqfODKPSgwnByHVcxr3Rhlb3yCAztaFFw/u+0iUAooDMPbJS
PbIVXIT+cE1oE2ZqctPtbeexauRiVx2GC5sEGhQEQQ11FFKYyXiEIYdZIF8VByemk/R83noge0dF
yc4zLCgFGH7l7sShaJxxoiqqIkrz4X612HcbvdsPQtEDsZZvKb1c50lg0dLKB7nzo2WBC8/I8kuW
fKcA6kM2j7lqocO6v8KLIgpztFJF4Jiq40F3wMs+s0m2Hb1qRQYVRIBDWig366G9c8qXzsCATDAa
qvTW/kz6w7HQCuxLzZ2wl+7BmscB1Zw8NLOdoEItc4gb2Jv1AS60ymT9r/UjERjqcYe3cP9v9dJQ
gOQ7HJ055IQZjcqhhvguPNJjfCOPcE2wvUBcA9WsDt8dVr8mvipj5ulGfxMvESZfrOIVcO8NRD2E
sfr/PdM+NRPfnu7Qp2D1ws3NOSrBlnRn2vTiWvCisU6ivdsM/pGE62m2vNAsMdWYejXobaIThWeV
yPoq5mCAWg22rmMtPSky2c9gREDImpjdZZhxkAq52gGHoLolno6JZzOLEmL+NMmXodzHIuTK8SY3
I5zCCz7fJiHSPk742YTmcjlyape6rY+hxy3EGHaI7ewenAKZ4Y/kxllFBvE4qa7B5ZCLPm9gKMdk
/pI71YZ3zeUChm9jpJfUlJFJ+N7VOThSw1RT1/xgSg6NrHEB/4YRjFZGGk61AC/VUxzTycCWMofX
hH90AFmNpp5TCu8d1ycuB+hnaHKy23spLbYiz5bloNpxR1ILI0d59HkxK6gBKsC5vL5fTl+qP0p/
8AU40KRHmYKMxpyqEyANP+yo3R8L+n0GLe4A00a0GNqQyDtkpbbPYi+yLu/XKALNh8kDHZw5oN7o
5dm3n2Wnj3L2Kt21uBnpRA70OaGVhKBahd6HMV7iz0Du9wY+D8fj06IlatAE8uWsYeRxogFjYN4T
a9LX/ZDiW/8JWf9842TXMIqFpESaUKrqdn+c75gUvxhcQjWVXgzMNfOeTKCeAB7PfljZxwSs1hzU
a0EHRoSy5A38MvGVS8d/EH48XfQerkbuRDFzcn8BXjgjoTL8oXVpOvpr8M8vlc6Wq3CazF9wqVKQ
Bs2dgNnGbzQ8O+mgKE8gpqY5j4849/oxXuHyim41GvoKidzgx3B1vmVv3MpG9qP7uonDDdXPDWKW
F2RCxxOQV5ruiOY4avun7XDq1xgI/95r6YCtzyjeokfPanG8C76yOgFnlHC9wDd+708vtBdhCU31
DPVcbCX4C6L63OGw0gf6ldLcci8qAvEIiD8XxRk0GbIrqOe8MyZlywtDF+VSHg3dwyORNXs6zE2b
5mi4+sBGrBpf5HwUeKoDNdkjiPKTUjrbLUeNXS2w4bLZMLQUyA+WGqKT9SbrhXfrOZqgwv5DtGap
HY8gUnePg8q6z2tXQRVXfnCcMdhuiqmYI6ujc839xrYNYYpdHX0q8A1dBC+JH7J+6JyH0Fv/MdTd
w0mbu2rR3sBOK90YW6VNa82DhqA6WQPt9Soj9p3O5mhAByhRdApW4uLbQ1hypRXj3EuntZJuAKUD
vFaDRoFmHjt1quiH08NhUnxGfL1DrfLz5isciG32wbrN2tFaOZlf53EVaE8bMapoXnq5bjSsz1ES
i5teePnV+3VhiWJrQ7AdZ9xN0nsHOWgmoS3AfoXB3wCcAnRwJdQasCh6FYeRT6L/scjni093MCfV
OcVXhj//zfXynJxEsC1jJQqak3X6YRatUNAMxIQeZxwWGAK2aMv9pNqz0Zy7JImtJNP/2zUlNEy/
HukfOSIpJ3ItVZUrTf3J1gUBEMR18xaYozSTpcH6AYUADb6Tcg4vLPCekAtnrg9i2QeCBpgrZLu8
JNs/ELjPdZJKAKaUqpLqw4pA73iT/hgGNNgCChQFF1wR4V9Luf+KsbR4uqiDozFzOG4v5vwrUGJ0
trHRVvmeOA4HcqkaY24HYCB8AyDMLQtYvv2l2jX/HyEJ3FzcxR9VR+O7vaqXRJ5+5rqSTElwhVhu
p1LxPWuAMyuU5PbbJsloi9Bsleo4CwmLwEzHhXfYjmZdTgc/H/grOYwxcbwIfNWRKIoXLY5bNyS8
B1u8dyj60yHdBUVHfeJ2idanJb9jdhDq2IOKvKkHoLUqYQI5scV4Pxzi1O35MAVPg85ruBeSMx//
6bMVKkkG9VMc7IXB9pFNyQ2qUqyU4LJERmmcmqkFCnKg7oHMtwZzaSdXy5q6PdvSxrSqnfESDI2O
PIlQyK9hW2tEztZGIbMdl053CPlv0EeWp7ANQLQeOnAG+YLAnSG1mICBJmD5GDzxTL9A+siI08IX
1aJhZ9TuYLGmU1MX+XeWPVeZYnfEqvB6jUhCgmayZCvEnFuMCYrhbOR81f/pm72T3YlswaXZGeJW
Z5QA4ckAsdioJyC380k/NtWsVnolqFz2kvOS65XLoIh+Ci18ljUpIjy7BJtOWKj0fsMJkGW1qEVU
TTZ6OZiz2GiBSE8YSh1NaqfpGum02qLa3wx0j47TOfci+nKLpNfx949l4FHmQL20lV+Nu3C1cZ5x
SAl0smOGvysTE5ybPzFw9MHrOjUwgAVazxvK8Ss10yEuW4kICOj/jtZdqMkeg2jL/GFHR51YUVMZ
123uzzW/ZTuTTM6QNM8KzNfVVBM8hH+LMwLu1JVOzYGvcuyMFnEsr/poVbmR5nrWw9CgMTV5etKN
yLzAXsRGy1Ncc0J1BuKtmqEaJ6yD3W2aWamKH3LIgGCi/U8WQ0UYilqMUTWiNQf8u0IH3QuCiVPZ
qnRZMYOuh6Iwyoe1CurlR31DaYWKxoGAle4Y2uVesyDnqsOaDg0Jm3kMZzcaC97hHMZJoGV9kHti
EUcAWxpf/sWto4z7nq1qqpSLDagFl9lkZm/Zp69z1W8ZdShsCflMf5ZdOY5jJkiPC4VL0yvxeOnu
GFMWrrl8hj++NwqsP0K58rAuVE1Dwz7njM+6/vjlH16mH5oveixlZXte+WwsxmSj0/c6jnCvN628
THCcKFrD0SyihwcTLRS3aXmW/guSwHdMo/RQ3k/sGZomgjChCTi0ZGFtkU9DWh1CieC3d0sYYWlQ
jNI5LgMdTbiuEO3PGE9HKqXsVhHRtljroJKLGke7tu9pAvpovKTTHdr/L5//LsV6Q64pas1DPDwH
yudSLPHxIR+ffRfWlRLI2izej9T19efBsgA6W26Fa1MmqoxFLgglgt+yyk+LH6+J0KO6ic5h/V3w
KfSVTNtOS9HlEwHuFvaJWkAozKjrEBkJY4jn00Qs4BLm/PGNWyJUyYbNCjy/D1ayhqXtBWqXUlNr
AHVyATV/ys9VbQHORegPTNsxtDIXcFQKS7Kn+VIFy0qp+mNwDAIG60qEqOYVeuC1xEMsFf7pfLIA
XXi3ai6IEslaYRLTEKagjXYqHQ8/HN04nXR5UzyUdRPE3WYrR3P9jbGAhoHiU9BktSdhwTv+85J+
c49fNRzHyvjaQdtv7Mku8XnlGjFaHOORo6QMU898AwGL1jysYB24TNI8NXEo1Zts86TB/gqDxHkB
9bHp3B++B7718XDiQQKuc6XYsZIRtvGFMnUuIGGxCQVNL4Dntusl4KzxjeZr0N6yKT+FsJg5Lcvx
ZKyCkhv9mjyfTOvN+G0KoEE6/2k0CgDJrvQwry8gW0cGacCkyYWW0Q9+K/wWdTR7zCLzm46ReWAW
AjoqV3RQ4Pf24/upDkBwM4jAcgY5mPKrveYuynxDo5YmyBeyRZBQwXBC3EboDGPKsbs78/5PL4S3
bQU1Vfd9tInStJtY8WU8ZFpModEfEA4diyYqUd8k+ACRUwHOOw4qc9n6j0nFWCl9nddzy+8+p5RK
8/R2MTF4PXzb2r9XcDGxjzkyQZ61c80t6CVmq4Ivvz6hkcKFaQYSrbQch5+QwnBb01tIo1xEEr1w
ClfSq8dmPXLq6GgA1ZIVH2o8fFy7MKWzasRmJSgzRVmEi2eQFSUI9Cx16WEbaw8oxglYrY71VDm6
zsbH99Xg5T5fKHsIsGlTRDgfeJdzqpAm08QDDm8qM2TSo4EZWe4OX79a1ju/rx9zIRnVAmudopvD
oU+3024ep2Znehf8nDjEeiaX5YIVYFeedoA899Gc3M46Y5YJDPPfBmBQ+TV/Icif9DmckAdtqxmS
qnLR6nnWHrjAzY8gOey9iMvgYbAnDIk8hQDh/xoXtTEKnj5uw9K6m+sdOy4MignkgT+424T7RhUo
n7X7z+gVChH47KJywohbzAuqAKWB7w9+TquW9PfmZrGKAeggiRdaIcZM0JJtwsVPhRPTHxGccRR9
bidNOMjY8M2Q5BECd6TGkznEExeINHQPQ6lpC8AIF0bzcHynkq1pAM0PguD+xU5L2YiKfoRnYj4N
WXzqi3rPYFuuQJVReyw36AKXZ0UQjuPVfkx3xe4QX9gLY3Zq4GorpgGyAHixncdQSC6EeU95blGl
zfjn0Mru2sglgk0uHM6xQ9K/m1lRho5t98etMV5LV7enL99vIctvPTyg14C3KeT3Z20BjDJYeVqM
8VC6M2bJbTNozu0rY75mlvuNzx3Lsj1rKe6m+fGpaHijro7fMCpEAfYcjvw5xsUMVIQgeolE8lFW
EYphcbf5ZaO7vt5aI2key+3zDWFbWkdGh03kZpLaGo2z61KoFjzzJ755zR0LhITK8XGEBZkfSDIN
9tNWHbKiFjmga4ovQ2auAMfkweuFS0LyGVSOvRimAQ7DJmsA9Qm94CahpwNIVEDiiyYgcgyveKNm
OLelwqhBUJfrQdWF+RE4eiFo+3nqci6d7OnbKGg0qx9EMtw2t8BmzFefYwIAfeZKrvcLfpTShwjP
Z0dvHfB6lu0m/7x01J2PFdx9e9LcPZ1EqgY8fRQTcMBD4QSbwytMgi4wUXBI+M2b0jw8QYpvs7fC
06+4LQBGINLE+Nufjt2+2QWz8eCMEP2cQN0T+O8ebxmJVvgmwkTAR7F1Hl+OtlUQor+fl+Ly9kNL
Gj8DY4FNm9WkJh3AJUzgPDvXC3HgE+40nByygZhllEq1FyeIpPACsO25VW+gfEBnudVjfsniCuVD
w5yptigXAbAoNPAn34LXcGFJJtQO+l6T/ze7ttdg5pGwyUo1y4zS67ZiTcFfgwgA5p2GloYHIoxZ
xbl9+0Q6KPvmSjD/0Ha9guHP4g31KUa1Cn3OZmChX4lhnNDdtZmGHKXq5i/ZeCv2DZw2lmWxLDYq
aNrSSV54+WeuT7MtJiy0I/daCRzQt9hK58Z99QNWZp9jtBHfstAyMqSCzpy5Mh6yecGSu/z9WBwh
TdLfWhsqqj2POOmcllpIlHFuHNIVwaO9v1El4muSibZH0nrJr1kVeOF+Mjb4wmBEO3gimeFVmcet
XYCXGnhr+02wP1vw0x3TJxH45iJ835jzqOe4xbcTcwQjT04h9U+4UU9wtLzIE+zD2QbRiwPtRUvZ
TIcv5coWkresXrn2rkkeTilkpJcHt4msjm4q1sTgaNjzxbkZynWCFuydZdF4MoYk9XLoP3a95R/P
smHfT2HDDNKzh1Wigc+Tm1JpyQi/gw6Mky9hFU0/QE+2l5h7fYyql2Qt6ZONMWgKQTQNMTXLLz2L
GGRReSbfpdlmhR1qWIMU5wFC9HundqNndM6VaDjrCGrrIf7OlU/gGYssDMH5637dgyI8ccv8ZxC0
7Q1VzU0vzwxZGLxV8XNOzH+wO6+j7itKdaA+cblvaNkBOpESiV61fUe7PFIKKdztRYCEyUViU3CB
bRiKmq63RY6Wn5Yu5aI5lz5tBsLtkI8PlPnauaJu00/UTOm1TNHf09YOyQfOSsrbRn2Ldlv9/FLx
Hny4+nJJYf62QSZJlPCsFtfWWuoKm+U4RWBq4xFC9pxlnj7zlMUmxjrru1DjB7JNCkClqhHOtU6G
dScJtAidsrhngvxl+IY3dYlmJL3DlhfI0QV4LxjnueXEGTVTI7bKqd9VU0w5vPp6+OxtxeSNZCc5
rT1gOVOiHQ1QIz2na4UW39ghY8FFqwaH5szShGJ1yteIUAyWH+Zc4wWDO43vD5/Xf8kmjvZc5Pdq
Mu/IIUxoXr4jMne07bb3qA084KZ4b1m8JB3KOeR/x5cbk4xVcFyav5mP6gzbFz8zZDLm1EH7UL3N
aPZj+L3Y1Bw0jAopOrtfrIGseILgHfElv1Mpsp2JdvWehX3t+NPZ30Wrw8QhymgO6V5l6u4NHgMl
C3qi8F0Rd+HHyOdxzuYVQVf2QAGgoZESFeiLcIqN2KrblNDpmGZhoEarEBSZdEq2m6tUAxlTZtOu
Tp76pg9XcCVzuK1/Kg0VrESx2lBKxi+GDbKIIgJ0TNTn930jZC9k8Sl8QOg8ON8c65eKzDa4fIU9
Ehd2YxMw2FpbgmlQgxmM+EkemaNXh9HzzDgV4sIATytbSZnBVpBfMq0AJvak28fLnSOSga2aoJK2
zUd/BT9HrvYxrdBj//Db+BMjNRLCdxneYV0FXSTnw5FtE2IafiaVlZBUe2nZ0vNDG2PZ5W3oerwB
yGGhIFLxHC6NqlCCYV77dbKim1HTI10vpzjd4y3ozarRao6fH7wckFkgSjf/LbOiF67fiF5xVC46
Qjod/8HxcD8rkq7Is+iWV7rKLsinBxvml4tY3+MumIko/5u7jZFnTW1VqSphtMUgKGETlTm/lIWD
LKx5a2YM5V8glO3Sgq5Y5JnC7TOxIEX8kMHzwugpPIBK7L2yDjBxnE9q4vvufWuYXRcymIhfNITK
Wu040+io/INbSlj6nQDB/WFd0qQQw3r3wwulAJMWn+vzip1HJUxqFRsX6s75605dCVypqAsSfJ3j
0A0kg+lfvTRmvpJnDEGOexnbvWi/yAUmIUai/zgihG4HBMrY7bJqreficcGS4ey/HASVbhwikAov
veqC5xlQ0quRhrU3+n3wDjCeZyBozre41j0TLg6pfMnB5R8F7h6cOxVqk+Qm8COt8mlU07cdzQvJ
FGKJ4zfo+lFQWLDu4PNr6ZODgwLxo4tOHp7hcpeqRTjbMUNF4M3xtcEFVePsF2gTl3o00opBF79a
cMQD+QnWhzXzTudM+JvGwg77keevtOgTfy62MRtv+a9wPATLaiwxE13zYvzMYiAuOB0sVuQG1tJ0
jIIr3+Fs0e+MP1HwF6ofYct0+FXeislFRH/jwqJtuvhqoSPRCROm10hVqBJonXlep2A+YYknpfgv
zRSSLYGqhH06tzz3R0yb1dTK02v/MXsqzWAewd+nfQHCqHKBc/7py3YfVMPiIyqAENKuX+plwd4y
b69qiA7l0Hf451eI3rTh+54BvdAh/GEYPdQjOZwlnz4ly3Reml1C6Q1AFQZPtbixCbvV0Za0ZwLf
KMFLvhzYXgdOk+rntaZP/kGk1/OluyCogwuqegjs7/cx9ymnJRgBl553fKo7VYyZo8dZzGmt+7qZ
YHm06TrQklXFzolg3BVwPJuwdfW77kx8OEz9qA+VKsIrmaHCJ7hDc6laZsoDpASXo1j1IzYEtFSm
kk95BAv4obDOWqo8V1sUxdMe26uWpuuqP7MBl44iWkqw4H/SDrSXJykKmBWDM0EyjYbAM6y2tKg6
Tu4NgZHMlKmYFPdkwXNrYJoU4nsOGGKLb58CTmgNYBfhck47UtDGCUiK907JnH0DgD5/bcdn5mx+
8jrqjoYUH7EdcfNx1a0B0G+eEITbupNiATBSUyP7cytXVj6q8ayA6uMzItX75AO5ycgWSAp4RPjr
tIm8FptpHAg9k3q5XCp2EUgOD0k1JxvYXoPZLRZyD1kQn9JtCs38EXydiYd0RV3UiJMP3dLfjRbG
dikvyzuRFPfE+E0n+GZwJVYIN0RQUaLaDi2+SlVCswTfbpkYk4KqPMhmroVrdaLQqh5/xWhNtLr1
5zbmeFxxs4Z1hnnhgzQ8zGteXE+tjiLe+gaYNg7GjYpH7BFzOVTY3xGHp6b5bcm3FKBbA0Qe2HRx
YhZqmKXlL5WA2udmmpo8zt6b/r+Ut9M94yZjg6bOLxgOegdr3hJ4GY1vW403ZpG7pvb2wJtw6AJX
br2uBHrRK9H+CvmQmodRt0cBHYxW36U4l/OIaJ8ZloJtDqPd4gimILquZ8Ore9kRXj/vFTkWSPaB
cGHUfzQFBK7XqON6QYjcyPRwrDNLQLSJ6NjkK1BS50SrVNhe9SwXBDYUNcc6ff/fA8qWT69qALqg
prHdiNjEACBjEz9KB+8hucD83PhV1OJxA5CGETz9S4FhYpS2oFebWZUaAu7kgfyVoSqnNn6bCL1K
ZQHgbNQhPWNKF2RS1eYQdecrqlucg+Wgu+KK3NzUirnxj98mtJHLS4rT59uJ5t5/CenLFJFUneuA
T4WIcMElo2yYcF+JzuAZ0e8hJaq3G8l4KJZdE64h8XlyhykAM61Yx2sWww3ZETVIGYwHxioY4vmK
1KYV9GbRRb9Zwu2zSNpPDr0/+HhLqaKMrZDUXWrhOAjABMXkVSlne2cQcRidkCcWqL2U5xj0J8jQ
pLGSbqj3QAYk5vARRyPMLUIWg/lgwoO/vPlCv/gE7DE1bPNzuplxy+xHe4SfALazjMdRmXwjZKP5
udB5hdiRyo/iu27xoq0kg4iBEYm3kD3C0njEitQwk4SwMpV7yRLAt5aVpj9RTgx408qAi5/hGHqL
DHqmAOWDKJwgO6HVZJvyU9tSz2tYdsuOwJqFArl20IJqInGwr1A6CRulxarv3Q6x86UKiXAiVyY/
a2Jnbl3ydpGhJ1bYX3dol4rmAfEIWd/KPEZx56kFr5/65EhB7lPxL2nUqOMlkABnlGNG/gZZydUh
XVqqU4iVaDoAx6RTTNPSn5HsFztgou2b7W6ZuoGjuxg8Tis5yElY4asEyEkXhkQT6cjYmWRyg5s9
Jqb4t9F4/IlPGTrGwU0WQzKwmfXyO8kSwX7Fok0all4L/PRRGUEPDxf9xADD4MNTN1WFUTRNBwRk
Jx/uPrU7IYoTCbw27RuKCk1LTSeSwpb99efI2LpVFmqzrA9qk6xIUQw342+qhE2WUP1eR3fGQ18Z
z7BNSuvA3afyPyKnnoThjsAaehqegJ4N17jPT+9HSSp71Veipq/cRrRseJd97j3mE8LDg0wAJ37J
0u5XlC/l3cg5OojmR2cdBZHmWAYtTusvRX4zjzr/+bifsW25ebWr4aodT4gLp5Q04ZqbcxcqOVrO
Dsvk5dQIjqU06Ajs5CQrGVvQ8mN+3/DnrAuADySAyfzpqF4SAapTzmZsmxebwXKQoIwshwoGkTPy
YOrzU73KZMfu2YnyIjaOOw2o8NV9vRMTXFcwIqZ61Age7s/SYZiOols/zrFLEoCF5qJBi3iy9n4+
TvgRpH2hkLDVzGxKovDzmgYDqrezL9WyiS+mm6mjHWT6Gq3oc+DJn+OJG6JYU/5hGfI+N4lEv3vW
pVrnYnfRpYNJZrD3urWOg7lsPcSZEYMQ4T4FYIEQ/CP9YSpW4agghwga1JDqrM03UxGneaR8s6Y/
Y9ccAt/Niv9HPUJKwseGwIvr/XFevqcUOj4p1oJcLPLMTSm1fg0AmuU/AOfW6TZ8kLo3CvPMUQ2B
3c5t+cUCC1leoy9JsW69SAb88tnEE5j2414Ud93Nfq8GYrzYo0KKSm1HqqEhQOEmej0hpSUH6POm
SceEJmoDEbTl3Xyl8Tf/oNpA+6iF2pMLjCRbC/QTA93NUHmoydywvzysd1qJjXrWn40nfIY2gVjP
told1bzOU0VOwK5gTxC6ff3RFOeqJReDpSTr8j6d2yZilpwJlcFNEQUMl+H5P8jO+NEVApW8/wVL
jTt2CwuOfv3tpiW7IEtykGOkgYKy0Of3yTLo/COe12kPwreRXbu+l/esLE+xg2ewHkwycfZYXrfY
KS/E4mcc9ywerudFHXEuFxWET9H6/e4thQd2ecVMPZ0P4ccjvSNhwKpBcLsjBkSSLiQ8W1NKKIGO
1ZcM4F4ybBaezpgqmmjQcYWeLNs2RerRaqqlUupHtaYfyFVH82aqWqmYbf6j7VLIyjdiz3fdk6Sb
AX2lSWU7FAOo2wTb6c7uaX4ExQzR8gc8mv/kZjpVfw1kblAX/i/4HKKm5FJkhq54Ki/N+5+hqSFN
UYjFyvlxEzkMUP8YAxNp7GtEEAxMUB4uThE8TgTHr97gcnJrpScCH09PCMKXOs3N4VRUbqBrumdX
wE785stkSdvxTG8sLl4eDduA/ttFgAZiNnFldba27ZrzxH+vBB9RA0fWeddw1JbTqje9ZGAC+v3/
XIFOm9zTqkjN5sZnVRg/FJUdGss3M0Ba2rHvTTLrp8lZWO54E+o3f+xiqY5YMS8g8okkr+QsMR4/
2WaVDKXccV0bh+YTBgk6B+P7PB9ahrrxD2wnZ3J2Gsjh1EzuAQJjL8+kbMrYM9pRMaP+xPV1X9Xh
4cJzw0qO9Uj0FYix1ZmV59IgX3y/hNz7ABKFVAGQqzAMWLwXuXUaDiDFuzhrJsKHWe+XvK/Y59df
LUAJoEmNOJXlogcNK+FF0S1Fxd312f32stBhRFceR+EXnwQpH9+MYm81N8dqfJ6Wx0cb39GSpnQL
yI3Xfe9ozi+eMCuXiN7DWXVj5zJTmmDRw+RQcPvjPb2Pmzu0zRU7Q/qb0zDUSgAfGAPh8pPKnIqe
WznGxcnlF+F6LxYnerqXXdN7xBkkcau4ZHUOf8JEH1Kx9a4m8SUaXrxIA67ByKQBEH6NmtI8bxfy
K7IXNKVJZVsZyX5a+yYbXov2HTzzIOfayXtGgKBTrL6Qx7lxGvcP4yYPLDpneSXbgs6XWX2IfIH3
Oc2RoLbLfQ4eql5UqzkUUJeitgu+9xHzs79QbVB4NIVJYz5MbZm6s6eLGyhVqBCfd6Jk2xEMwmLP
Pudd0UvpTDARsZ6JT7+HwMrlf0doTuoCR8cF7Bekq6bTKBtDro94smRkrK7/1n/7L6Fh0B4Vl411
7u9elbIos/1FyyE5nbB8R7ynJK1lEdz0OwBH6TYmWjTjN2kttjbjE4TMPwD0DI1//UNx4Lsq71Y5
LWx5EkhTCo/GFi0Dga8dxMMVEGLiRqBYNx5BC+hoZjklGGhyjpyZ1JjkX3rTLSvYe2Yh+4v1+ne0
69OFIYusvStAe9EaoV+ggdGEmaoTx4PdVuZZcW8oHYSpSPgVAyvlrTJQLio71rjkJukWudIqUFvR
CEPwnuWqPG896PZZR2tmaxgwgarG5BgkbIJ7y0h/i52nFYve6ifethTznoVHE6aTbOHfkyU1oCXo
IF4ox2TWDiFyOvPapppL/o0gRpO3dHl4M64nhj1EHT+TFovamQeKs5T/XxH9hnq9uVf8WuqegPtI
AyxgewuBO5Lps7ly2gnTNQfyQ6wz8a09ZRJLn7jXbXNAT0xzn8A/GYsC+pquU5lNCn4wk79EwQQx
ktco0rdomxGrSjIJjN6eitdGoahwgaDbgh5UjpDyo/zB78wVKHZ9qXjM0AuoxUbauXHc35GRapNa
W/HAjemiavrP/OkAvlinkwyBEtNYsqsOcu1v0u6WkY12e5KeA9eNvb7d0nxU1+Hb2/XnDdaxOJsn
mpzTvLr187uA8QgDv4hu6dumsld+9EF5/hV27nufzl5W4jNwICBls769n9m8UiSc31JDXgsryR67
HCqix+spvEvYYoLps9RYbEmj1UaYhpF4qLREkfWOMWjMlTAJPhFRNmKV60C1mwqmn56sl7X0osOC
b2cLcAm6Xo7MQ4bz81vktR5vfTIE3P3EiCyhXkcgW+h0kLEVF9YFwi7TW3ETs7yUuiJfcQAKVdRy
GEk//VpyMQOOpPNdwPKj2PlXTsrlVOfOXdOSE0KzPJhR7PH0KXHYWVhtSiRXVOV33zAMPU1Tg1fC
iKs6OI99i/xm3n/t/6B6cbgVftmpRZKGV+ax0FOSqar3bZgncWBiH3B8ch9Vy0ZqvblfWweePqT+
AZQzkiHpb9toHXkJP5JFDZ6tuZigmbu0gOmfJorH4WR3LO7fqgUgBMca8jjm5jDJnx5R6AEWAEnc
ipgJw+YrqCE1QltbJac7xUiki8UhnoSThRWXrzmytcZWSj3G9InthHBPYzxt6fpKotToHcHUY9Dn
VqwxPMB9xS6IDcVRovfE/6MzIgjgs6UdN7I+eWDPw78937j21hTWmPKEt+THWQovOBB0XMLmScI8
ngar+I2teYUjcXSMtV0tY17gSG1emWNwu9OUMxytjoBaYNS13RlCuqfDa7/0wZTlaeZFK1DN3sgx
crmE7nmS4X6aGSY0PIAXTnCzc8F0MI6YKD5UezC5+Ts7/bILW0igg7vz8WMUt4XynQtem6BYBWei
AzntuYepm19VKqAi4YLRZ4LIytEUaQkSwkPoaHd9N6gfM2dUBxH+WdxHUcDhLQSaxVUGRTEOlmUv
adwlxIyMxDYH+PTbmy36TEtQMcmV7RypqwMN7yjbEdk3ZQqO/l8AsgHxuuPDztCaG07YY+CUfbxI
LYv50OWYQV8Fc+wsAQShKC5togDb0LMa2651YFtHaWd1ewJ3UmYJ79qM9oyCsVDp30R+kD4GkD1L
OMu8qzmixieOCdyhIh97hWajAtWFWoOlAJ/+6FHnRSk5fFb+INeK4KAXv0Ph6szblgYy9upMrkz8
mK7FmjOQpepOklRGh1uYLDGEYC7wANywEG0L0dF5gZlgBbDt+kKq/wCiTCcVmvu9z5Tig2ReyeYs
K7nXwSZws7cS4cab3n36MxpDqHF2Ls8a5w7WaU/PuLuAIQ8OgGzl/jTswOmktcQ+x34AFObSj9nF
hJgqg3emxu4wz4BrdaUKzcWAlxpRXrFcXemd7JxlikFp8uVCct1uFb3txNrJSWN1DLpNIa6tOzDD
L3zGSCSNy8epL3IR5mEMQRAc5jGEInD1xThubwJD1zMsAzKFOtGELDtMbg826YJs1nQBZ3EhB2Ri
xrrL02hFVRoTVNLeRxzMy82kFkNNImE22CBM8yjRKaDYwQkdhd94ZUo45YFFAsGTECCVRXJCTmdJ
UgM1m+UZ8a9srkwRYWHwXVyRnTxhb4qeg2rn7Cp1uNKMSX5g8VQtai9z6rXvg28kDRqomXPnSVps
mj/TSxifg0tx4cPhGcCNWWBVwOeb3gMeSU2xHimuG72OxVd2YN5UbDGXv0gUtD8R+mVes95tjXCE
7mpxES82NZ1ITu+h4g4bUlXH/chUK/MMgXiBhICkG4b6qNx5BK3Dg7pt3ys8iIAfZySKZlTMGpre
qu1DzzAug2fcFlEzQLVjd+SkH4kd+ETdAr7LD/8RC2PA6OF54jwNJTUKgeI/GhNNZ+BCu76kRd96
3vOV27UzH99BgLdEazddBRgfiigRdVIji9rWJKdsKSOmuLHpUJb7pm/BX1ZCk6QMlwRPVUVG5ZaB
Dj5YU3I/HcUiF0+AXsaEAifRoOI2PRqBVvt7321P6eSNLyTCaxc96p4+4AHLM4tJ+ipnuKGSOncV
leQ2kJu65/mXBx1BYeLwdCDTd+4FObDiAeA0CT3yvHuC+yP2iDzFWuZonwsY+fuvBFb8UiXpopZU
h7QSBPtAOAyD6eScT7vAYGXYEzQiEBsHM7MZVEebHtTQmnAOzjnXvfOD/ELiWQ5Hry/csug1D6a4
6jZg1pKGKQU1lGUa2HK464kIdcn7bdqBLxTGOIL0MaYK4H0Z+zgO3KBQeKUrPWD2FBFT7h2WRoEN
sReBF52gOuUz829Vr30a8gprKkgPjJ3DZIwYjhzI6GMB/i2jgmX3hhBAo/SyHfH0z2uVp+2J8o3q
MNQOwXy9X/Vkiyv18jZ37qYfbOlfG/jSsi7RITx+eHNf+M9gZP1rYTl/QuD7mYoDlBD2GtGiquc1
GemL66iW6VZ4hMu0sHPv5CiYzrh+vdA+BZ1rMxEKD9wPQEibv2YTjezh33qeZK4mNt4IHmt2nQD7
MxB8j30zFg15eSP1cgnkBYdFsZgRYjnpJ+xQOtCPuiQlZPHHYORKNnv/YqpP1X02uxdE+MbfcErm
/QQyiCjV2lAcJMUD9taNYzw++DIjEvFXNyoifh8x4Cjtop5oXxk4oDnrTaMwLv7sTmHNxDRWx4Jz
EAxuQyd5gZ3/dHPcbm0lXtG1sr7zgkLft/1Kx5l8BEzkgZEppTSda6vJtoWTptGsceL4A+Plf7Dg
EYa5TEmEryVE5xDJLms+LzqaJ088ZFJ1C4wAw4RooEuib7/9sykIkoTZqIJFeAvwFVozvDQH2aDM
T1xXfrrZaEaCCO+WUWQMIH2C0X8h8642A9pkW3gYNty4PFzKCDLhZlAvyNKbnJnkS3eL7zjGNFpo
S7Jh02WjkfOeSc1R5DslJuOHxMIqXgZKwCAy+CdrvT6WukJ0Z8ko4hAqCnB2JhLCs+ElaoCqOyMw
Wp3KnhfER/SXqRxnlLIw5xe5p7KnibvwCDvmZCm6Uh/r54fAgNPnOBN+Tf6sUG+W5xp6kGOvTXvI
8aAhBoLSDu/nFV5N2gkkqLnypdlpanPqEFtHJ3Cjh5uHKDstBqKYEd2MyHhy+UA/WWz/NIEup1yr
mIlvPHiIWCqbrCq+q8EtfNI0SPUPX/cpb1E/C2SgM5vkXISEVpRzwdvtntZNzYHkX0T8K50Z8X/V
wgRuS4ykiAP6brVPkmZuA9LCf3qTvHZxHXWy7w6eUWRaVVCi2o8EUdfuNuZOfwn8LD0RFKwzashl
DIT4DDPYa++Mkve7zQOUiLSS48VDwhVyP/frKJjji66mJibwj8GgX9cyPtTcEd0DHq9D4V2LNWgO
g3mUehXCLhZP1DBr3ytxeHSNy4WG1VttAn62g5Aexl75DiHzbkkbOGzi0MrtYehm9bzf/axFJyre
1DGDfPmSQo3jo7wiT3DmfCU/tRCZXSw/2IEPcGkZfySWz0YdqZHDyJFeXOlj4EkXi/s+n2U/3aOt
Eq9dyxX9yM/jzbgRvmlKMQbAqO4jZHWQwLKZr/ECKET4Bbdczmre0S1/9T1w/us26hyTrr5b3LN5
IijDE0mKL50URUSNpenBHhHoMZ+t9k7HUys84z+vVyRiRVLQJNKPSyTFNfz59cVE7Ik2ZeDgvpi7
AJY9LM2DJk0/PIBKi8UrNzD9jDJDo8nFlqh76dfLfCPJAeeZaVu1IxQnTOplXcgwimPDutlFXjtD
xhB//kGCO+uwrZbGPv2WFeVu8yWtSxUneS5163SXmtvXZ+yMSU50TB5mkr2UueZwr0Lqnr0tZ73R
kSLFJviyu+uWZFJK4f9+Nz2gqiwieFNDckjuSMWQcdC4L6O61qcPGz9OpbV7Pcn+px3eIQJZZsPj
wlWt6PSzXLbaOMBnO32ltUZ/1BIAMbwkdBn2tD0zgxstQN3WzmoRn9Sk7DEylGkQ8yqeaovyTiUe
ersG0Ch44gDz8+0+Q+BXvEBkxNIpimjmQC0Ac+JdoHhrAuZi1c5Kg1gbm3MFokdVtc6JITH7rxGR
ROla0daGhgovIt5iPzc+dzgtdtnE+7UIjFNHJkmT7ENTEfboKJThI3RsF6cfaWv7aTkXRanx69La
/LQ7fPz/ODM6iWqo+1fe4f6QXnEeoYftbSveR/pvxnKSFeRzUybXolfNplN55DP88fM4ncpCADuC
UN6o1o3/EsLoa/ASHfW9dGtq8sFUCOg870HLSB5+SH4wcCYvtx1eIF03olO3UP6RjYxYOTIvzHwr
vWbNa3CFABp+v/+3zKyzd8/AHYMQ3QyH34QqnjVsls1XxCcqJQ4X5IjGs8FIzLK4umC9GWP1/Y7y
siYhoq4t6ht8jTkYkxnOF4jwubSL8JaNRjAUP8rQgmMPzIlP/JfZ7AkhQHAjE7AUX8YH1z7q48K/
eNTpHVi/hSLcYZrNnC7Dy0DbBM7IXg3JE1zn60YdGsN1dui4hqcnuZU6A6I+NQgxBzHU1ucv0yhF
4lNHRaeEB4AJJSZfzc/X3AOtRKHZEqLoEvRSAFqGUcobSRqYvdrV8dB6Hz+hsAaDU3P3SW56PrpS
5zViJzQOpCaOQushIdZZcgHTC0Mwgj8GU2HOQ1/0uAHywiNDHiv8T5i4FJKAmFay6L96rvowBr6+
B2AbBVqzl7sshNB3Mupvgy96dit2komyrNhfI76RGKQXaIuHSjTM7bOMEv5c8OgdXmNkuVMFNzv0
KGc7RPa3XGNWgq3WU5uoo2hnI4pxnVKMArP16yXtGUf4Mu4cOuCI/jr42DoZf3nxRJ9w2sroEF9r
7FYsNIvCozrw65TFkG5LdM6qphZnxpIZ6UXCQsYlUCpZQgafCIdyI7baoa8n95yqV8LeGBsgOQli
TbP8cBn2LNzFp+xjHEzFG2SRhZDKEwEqqFq6tteRH+gN02y6qZuLhCS81z47Gbt6fYs+8Tiy8nad
63QbyoZ/ZmBBEVGufEvYpu5lfDgsrrT4DAVLI4ywo9bkA4RvOYpp4Kp2dwDa7NXMWtGSbk1b4ssE
GraN0vR2E7zAln8t3pj6rbnNfQbBcZ1VPSDgfo3UkZ3DgR83NWXS2WVqPPg56cUOG+e+fDGc6mKj
Eyogrc/ZlqrYJrWYPMwSdvOFGv8rZt8YYELl1/8NTtODXIsgn7jRwLga10nkuXVpegBEj2h3JYVX
3N3q0xuhUFlQfJpVrCE340k3ww1K5IXs9kcKdeeMzJlj+rh9SuO3aZjwh6VdSJMtM1rtSmd06lFN
JeIWcWFS0eIlcnPdloWg+O0+yihHnkbo+SqhV+8zCptj8VRLE8iz2OsfJQEga+jlNazCEm43SdNn
AvptjNCGj9wdlJnj8cfjoCcYJI2P5ErUHZVTSVW2PuXneY/sNtj209HyTnEyj2Rp7otSKSxb2J42
2qoY+EinUapIkRJ/Z5rAX7BU2D33Cb0tqSkufP6ftqds6qY7tqA2cCEawsSkIExUsF/4qOMvmLMC
wIyF29w+wnOdX2qbzY29JG/faErOXvTXAqOZOrCIscf30g2i9qnibOaGTFKl1oQA48hjCOyeGsLW
mEwj52H1nTU2K0jEH/pQ66heDvNkdKxdtDWFSRSdn61GF+9SWK/slDvqkNxxso137BO9VCucsKNK
VsIYCxEQP8ECxgJhEMWt1t2MOEq1coaSRCAMkzLG8KN9TYL/C8ONbo1/IkxyZ8ggMdZg5zQsRiwm
5hx6e6U/zRhj7W0f8MqGyc/mweAuBFGYIPsQXDkV88TYz+/R4fUP97nWRP1wyc2pg7J1wvvsNdX1
QP5wDKv556StqvoS3g6oCjPniRgeKRAyBn+h0zVIfDcIUW6XNCJuNib/V5X9bYFzwIccNdzEHOwF
oERyYbvo4Xr8LKmgtlLJeyKN5RUTbH3QuZPF0k5sCBcZFs2k9/FriaAQYpm5IHXRzF1Hgd4MuY+1
IGKMRah5gYK+ZOdJDCshiHyeGhysoFepgpZdTgVrtDLmG/5rAfuDj0RniJqL/3m5ycIb0DIkN1Ha
wJAmOBpdV0RawO7gCWdcQrJM7TdqKdn4Zsy3ALb3QorkDmttnHAq+RmRnuhfXurZhF73jBrFoy9m
B0HtomEX5TwjI0mGIgHKFAiMx+Gy5TXXAMnOY6bz/BEpvUdrUOG1aaTGkBwzfywMLwY7OSzxuRJt
xFsdeM6CZv9F/zvuxtGTtTjOdU8lU4Jdo3wk415lXrQBjLXho4EopnZp4NMgLsyurZkMjN4wjwSe
7Udrs7VcHIEKmQVatE9OGMgI3SpPfDOIrhGZq5em5cFkIJR33b9uZsSLQl1Bgx2OGSd+QCWji8GF
PCb018pZX/IMMftN0r16wprCudiXRe7XnL5zk7OzKwOMdS/P+k+ZpHH+sle8Epit3hW8PgHs/IkG
Ri+VGWwxjCh53OLgodqw9wvNbDXFGtQ+NSChZsgWZddmn+MaqHDVcRhL6N4d8qF8l/Hc9bf5b9GT
rHXwvsYeb7lceMFpk4t/x+SBKkDWTkhLmHyI7+EfE1hFAXk7Me0EktEkSHjdfPuENoULPLsCQRQy
ntBCPg41DxdoiUH0eCa7nPmqeCqTv5/XD4kraP41lJ/RkA1m41sb8jvm+/yzibammV0WEPZTyzT3
ZbI7bPbLZOHiYh3uxBIBkmEC9LRC+uPpYplR1wpA64fruNTSPauWDqJ6igt9XOYJRvLqYo5zywIQ
0vXsxCDWk71cJnhcfF2Eb9T2RN9IGxa7MDqpc/xinEUC0EYs1rWJv0q4a+RCnTL3Zl2xqeQIUofP
I0XO7R/XKKOzRYnX5pQHUSQ27kl5O+EsJlpHRe/4BbwC96N2+21XMwkraJubHrAJjWT1FhU9Vko5
8V1MWNf7K4obwTd7zHWUuqqBA9gwQ2QxnQlz/w9Le4HK32ZF5A6wBh+aK1VOW2lizwRPhRT3G6dQ
jJR8oI6SRbRx8ZfpEvw0LDPv0l1Uh7pBi8yS0s7+58d9QbfA7gh9XvzZF7VXWq+wIpoB9eM76wxW
+fhmsnzYhitS+Qa5ihNR4PRSGHaXW5z3dpvRnh4uFULLilwMkOdgADI/1L64MdYBjlizWa0qbc6i
qPAHz2pp+K1rUh5/7fuB7zGc/xZQI3DNXiL0TLcM0xlltN2k4xRtQBHH7aJJR8wGXhksw4Befgav
sysonIk4Q0IjIaybw8h1XirpH+kvSlw2cOiAmejXA+ZJXau58DZCEQYfJQww0jTMbQ58p9C+86FG
aQZMNMS95ykVN3yeduW9G6HXosxk1+AR58wINlJCEspwVHyPTbu/Kh1LvfOI2vnhtucU8npBx8s6
b/ZwEqeZ3twxSzMiwbp+6t4q9UPFDN6s5N8NDPIuX7RygW6nQ6mlxUkdCJO06rrWIiNZoYCVBTqX
X8w0omznAQhaBpolKKRo79CcT/bbohATxhVRqK6gIYRZ/irn3tYvI3YA+vDIOKssVqLsp7QNA/Th
I4sh2TK6L5aecadLqsec6jZ6XcsMV9pa+TzeANoloAPz66UcYs9/8YATYCAwTTsscb7rBCbDh0RN
YkOcgsOAj+DuD1BMtqhHnY1qOefcgpwVYqHbSq4eOwiWEL0/JRNzyMVvaGfKRJVCdRz5FEsBLT/V
TDWlfFugWL+dG1OWR3plLbgCTYqrVBsSr7+Q1Aa/wdp+Wm3bPhCbop3kmr7lytOHc2naIVgzMYCa
CZ7g6PCuKPBxg4InIbGFqDt4IdFDmsYgnCxnux76o4nKj7d2oUJEa/F4SFBTJogeXVe5uVCf/moX
cBAvSYTJPFicPWkplwjg/3Crhm9cKgDm+GeSF5H9LujPWFWkFfF4COrY586jhRK+wcLXBMEp/Km8
avv0Da2jvcnbS9AWkLVz6kWNgyLaOPc6niVxMVkB8OX3kEqr5UiW7NXlUF5SGw6XToqgLlGrsKOe
LGwVchVVo2GqlAC04xsq1pU8/qLHberseFzeioEOzkC921Kh4HbrCcAWkcKD8uD8ID220yU1Dl1u
ih+j7EhYddzEouHZOy4iMKiHChMKlaNlTiKO40a96o9dTHQ8lzosc8NAmUU0R4b0cV+0ZOQL3Y3V
unZ8vKPd4s67xH+Rrjq2cS7Fpd3YxLssFpF1EFe9tv8B//cDrrfvGW643SKpxCMfNkqqysmwC13b
8o5AO+ujLIjpFpsHLf6Dms79OlI5oTy90KV2yM/TtGEcFn/AxqjecawmvIGceyE7gYvKV7UwbTW4
mHORZstfVwzhIzAKiSsTSmwTtA5p6BAKMAE2NHWDd3dh+dXrIkXOkZKXDdf/AnoQTG++5qsngUc1
wgCZbqNI2E9HcCmNSEnmClsPCXSxMmTIXeEf0WMMhAkIRXCGCfxqO3TAq6vQa+YFSMxXKue0X/x6
1KYZtK5vVTrpGM17iUI6mFLlZjiGyefh/08ysQ8vuhovk7Nw2EAIsMXX2pzo0Ttw/EjC8V+AU4CX
6P2h3fdqr6UMXVejGXsTgywqq5kloECL+cS958xPgm72FY3Q1YrEDQ0hwFShK+Jzhmzcu8S6SJ7g
rJFFEce2XR3CqmyeF+EkDflnmH4buoflKStWrVDJbhoAW6K7jrZ+L/qXgCQZZsGZ4uHqAaUPy6oU
xAsL632ZPwUe9orXPh/CeK30/7OC3FgHyeK58gmrnWykGv10eUYgVFgaWp0tcc/Ru8Sgd52Y826B
s06ebYE1dPngnoPKICf4qy0E0aHDLn9sPeutBwqbTLFPohbQ3ZTkzxZgJ20+UA9dXHjKsjObJr/7
pxzmfXxy5dmO+nPbTFHbRCrAR1dTRUyJT2vJQ2GL4xjPLkDQd/J34wIZHLR7peUmtTBTOsAG0zZ8
N7ZqvrMjNoT/z+0TbSshsvvdr+p+V6AV+JmkdFZXoMYV3Vs+ATzuv1Yc1Qq/WSgnQt9lv4dC6wsf
n691TbRhe74DoqcWUzPRBfRcHSuXs1Gzkndk8g+fIZhtuOl52N3wDnSphLrhVcm0k9mHY7sQNjUy
yhpkw6cT5nLtXKRP4q47xirWiC/ZbHXS2MHXz6qUKqkkEvcBCjQuwy67YHqJBhCRTzSiXxhL6BrU
cIjdKqjRuRuXynTDhULLFmEO9AgNvJw91A89kP2J3FxhGRV4B0YXlhQ7Mf39YXomf6TiB1fTG3z+
L3/0OjdH53k5TfqGrWtCNe0FuuZQ/3BSmPGIksIu2b4WwZ2VuxbnnQPxiZzQpmYiqE2rsSGaYOCu
oSQl4OxZ0/bQpwfkMBo7Ez0H04J/T0O4vSCvaJuQO0KsfrkJC7KUph/9oR8Sz0L4EDZNLwnCsr8g
Cx36SIe9t6uJrspXcpmPJLmz8qc/ygiJ32nTrMDRoiYVmE/MAVR/KEY/KsniK/6x7GaI5A768ruY
ozkT8rGCX4a6egTt+dz1VP+ptYaL8obixj9HlwGElwe2RfY+n/6AMVii90cohh8fsrXtrlC2wNss
WYB531HUKL/gRN0k0ExKfh4XysRLLyvpphOuDu9GXgwckIdqV8ILmjGW8Doh7Tb8X86PZCWJ36z4
p2sp2qv4H7BI5SiBGvzKI5E0/qPtTWm7lc6qpmJsdylAuvha+d023IVJUryU9w9Sbk/NkSs7/8I1
bNNIIET9QRVGSW4+eijC4OfQofyzXGSmWEVOrC2bsKj1e+YZ2Aavmip1aWGCoiLAGu0NTudPiWSY
kl+6nGjsDWXN8r+sNpNlFnZ9vYN5F5Ceb53yG7jxCXXHUlLzUv1FGNoF+jLSpAjH8LzpQ4Fi6QX5
31ewazRUFK+yliKmp7u/ePNwViLuCMRPYhtNjZTWoCWmL8DqZhtm/te3j6ekSkghJeS8f/c5mg9j
3MgZOBZoGjhi0Pddy0GyUqzekR2IOJhBV5npKxos3R9aynzbujNc5zNnwX4gO8LLO6TaRyon0NzB
pvQkWiEgZyfvOhxPPJt7Jamk/n7Z4k+Gt/b6Isn9crfmCbJ3h2LEWNe4y/sJ90u5g/Hfh0UooUJT
xkiySJa7gpjZZFG69EtzgmwCns/nEFiqZFlJvpZOWEhnbn28AKGIF9yHKdiH11w6uNovkgI6Ka4f
RmwABgR6Cv7GaeVDqiKWQgYA6uK73HrvkrNsxb/pzif7uJdneAuiafyaUN+seLDIgEqVrkwmiw/l
lXLeSaHEyH758RDiTaDVe4sYU2kG+W61G/5Rm/kFk0/+vj3+1MGIB/Aw7Ky5Q6LHSepBubC3/XMT
FmkbOgqjwWY8vScr6EkEnqlu810Nwqb7kUUYamY2422WRGnXhrvscqEXfVAPKVYjSwgj37jXmKLs
00qteRe2WN6w/S19n9I8FxruAtjyBbSxL2PlCk1RtqJVzC9J9Zaad9FZJ+Pq12XZPwaDzPqNue6R
yjd12OuU+tbeiEYVprD9TzoqfCMw7reh1gxqVg78IZBP4fJIaWTbNqVOrZ4K8UeaRRsV7ZkksjZU
FKJxI9d1T+WY2tTvQmwdc8vx+8nmutuWbgdMwiveftAXXcbwdlcvC6ZXfSXoiqAsZCBl43ATfddR
b5sAsSeICrhmP+sXAd93qPxFykLgdPYFbef7mraR3mKhvczbQGpw7JU65TuXNsfbElmze8GEu0eK
IZTnVMnDxeWULgNKRQSZOfAKaKpkNfrrSPCv19tSBVJt8/cwEUIXJ7lc0F7AgOQyDA6xEZIkxzS+
K6Ezz5zXggdgy6fvoKnzptx3NOclamelvZ3iHM24IKWf00c9aIpImL4Mzg5Oi9UZcABZCXDkh9yn
MWiCblNluBmoGC5oJaSygMW2yE/T5aHX2QZpYTZsrYRXiwSCaWD/XMF0Vg7yUqFRoaSVQaNkD07X
NRPTHTpDEQW5usdTciR35+EBJguvTLrSLlincZIke9phNMAp7MMl8EXUeubmiwzN1429vaywBmaR
LdQ/R4fjVKwn8VCbH182qH2qXI5GlI2W5GnTHjCwQJo8FFlfcnH/jsaP2nhO12fuJFyNiaY7Fvei
UU0D4zaCh9SELFjWf04dOwApJoX7GbMJkVlf5eze7EWWFvM/9mkYHD2Ex3HCtO/0cmIVzWxNykqM
sOYdwUQeHnG3J03H3ELvTkPf340TjXVJ9Fvwr6sGfkbSBv2uWUdqKgL1iKzENtKSgs/G44b01Brx
koNfeyVdupUjkC7m9XE4WtBLFNMpIprgMuq9Ce7mIQpSifA05a7S6UO0Tar4WvWZ+EyUCv4gpfJA
CRgVzyw4zqdJp0D4LXjjQ8ueTaZu//RwHRkxn5ODStL2+UBGTBRBxZXT+MqQPypK8wiXuu8l6zZm
+2cT1YlQC91biAXX5QWKxUktJqZIFrAekWDOz4PLKTrsdwJ2IrsfAEa0U8AagtMVJ8Qkzaco+BFw
kxvSjRSNJOhXrvcudapNXsmSvAqtnhN8ACLOdS1Dh+eZYxhJ8vXhL3zNLKTSxNYoxSmID+ufLdv/
Lyd0ZKSroIJoi95GQV2t0E0oZwliDFrO8TAEc0ea3k7x+H9aaw43cDhUuNuyTsa6DROc/bM3TBgd
hGnIEIdgO72vsKuHW6oL41x3N7sWo5N5YCm3Jl6nPCoG9GN+AZspmdj0NrrUDTCwEp8EAgm+8S6l
6Ain9uwGY4z1qoiKLFc8m1zGYd/UdEb+ioawvXAy4/OFP1l1sNT0PG6vsI+LeOY3kAasyW3hrFCj
1/J5ltm3bRTCOjrkBQE0apTVveQpIoKvtMhUIFR+OQQg8svp8grcfIIDG8zn+n8IoeC31guBHtgf
VmZgPZfXYjCxoh+W/NCpFzu8K2puX0lex+b3zBUN2ZUOwMImplFlZRXOr1FK/Dx0NOuhnmwWrOyq
+bWs/YPSRmkJ1XoCHq00ZxSp4U2XBZqyAnguke1KgM0upR/FdMzgSbNXh0PiV9gtbUzoecH0JkSD
V06u2FGfW7QLfxNDV9NT7sc0uPNgloFf9WsBRG1OGH9fFiGnej5amYiMXZCkuGen+7Jbl7Hs6O1z
3MP3LJb47+GRlg1f7uNEh1GAGufdL/tDgE6cRYBzrdPpzGW4T7jDkvQJkrl555NlWdrdyJExT63s
SPgtQ450R6WXs17VaJYgH7Ln+datgpk0kSQGT4vvFbYBAtyypAgDzR8RKLb2jRLlWyOOR1rc3QFc
LloRB9pd2YrpdbtxJB80fiz2gPb+EIsGZYhGG+agCcoYQMNX58oUKtRguMQAdU1bo60sTDOoIyxW
N3yD7/v+ftGz4LhiH6xTRf+nvEv8nUXNgNyBWLgRWRHynhweK8ZMMMiIsf88QQY31qsiMXQ7XsGA
bEk5sC1YfqnOyNeQWCJ+6TUHpPYGuQcW3qRMrVCqe7pB9amK58ZteWQ5vEoyVYoToEpskrPo9EXu
UUEO5Y3hGWCGCq40Mx+yeDCo3Pa3RTXUL5K84N4cQcvE7h/9bOiEFWMCi9rtfNBLmAeGNx7CJr6c
/4MNi2kZXzjn5UgpM6n8X1UG2dtuD+CaNc7sacEkEVIY0jbNsqwpMhrkRT5VP0zRZyd9nqYfillp
nhAMlN/f0M6bnFBtS07/pphbeFVg/0O8kesnmOL7VD/060baUWylCJZTFJVpG5dkbLfRXsc2RSHV
NSi2BiKrqJwaazGumMVVaJOZmLQAeGvlRW/Il3FHs5UojTj1yETUaMDwUsLdgvUR/Gy3q+n5GAsM
0tt+cs+sBt4IMJLrsozpLrAYoj9dVKqiZ0RlwDjJ0KsyiHQ96KsJX1U8PE8XK8leBPQTgDmMcnyh
t16vTXHFMzqvihZQZohOHLPZ8N79uMdcx+x0q5yCNUf2G/ANgveLWw6LB7Oad++t3Bf6m0vyX73+
3BFv3mZ8c8Hnc89GQi20wRtKQHWDZ8AnHKYndR1k8sRVHDxr39MH70GsXLAlZFibvZdlsUlcgAcJ
Y6OjAO+XII0APhvWOvsg8AT5tu9X8jWYegGdJ2FlSAIHeCF8B7hXW6IMM/SLfm1wogbImUtBlPpd
t2+pGzhU2178jZb3JWM46cIb0+XDtymXuyPMLcYLAA+EZJ6yl7UlB0dJN9dM5OANsYC3MbQ9q/nF
iRRSP+t75DnFbtBdCuPnqIxVBXWlCrCnQkkzYy0AQ7OHuigK0qVXnmgluODibGrPyp4Xl6SNb/x/
Lm9oKb5K8ghy0vsaXCSGgpYnKKQGmjHG2+guLoZDEeE9M7iwC9zV6ytfInfcDeVYTA81daAbnjQ7
fCgdtm/1xAMdna6U3ji5jiqdOs0Bnk5i7tAGmI8HbcRkpQC5s3hQkgFjYM/f3vvOYJZLzAZOKCRB
0RBhNk4OhspUQ2MApYIPVAau66rp1mLuKNpWHl1XFh3XqURV9JFpW25SUXbP7CXghQmX9H1gfMxR
xBsDN0DqHdyjCzfqvrEUOJt3xeDACG1wuKm8wiYuousb9NB5qvhZCKDHIn5mPb6E9kuU7/j7Q3se
Wvy1xyaGjSMxYoOnURgo8FH16TW5GKBU8IeYuIa3uCQCSLDwioE8rUjShi+Or3pTMzWco8H6Kve4
UXOix5aI9zKmkS9YWZzemtMVFYSvSwPFP3h0Z5+RyWDe/zp8GULdmyneqaPsB9sK00K5L3lAPfIS
omZeAErChimYytwbUqtaw6hmQIlr1vj5AgUBJ7nCRGBeJKs/sAQHmjZ+jV+i/wSdmwSCV43BHeSU
ZmXzXh04bRykW6UKL/sQnuPtukof3rk30X75+LuB2FXGsdomQT5JIJLyBn2iMULMmmuLvMRqDxIx
b4EdSJlKdC65ALWAro770N4mj/KYZSsk8zlE3e5jf9kGgSE3BsZ71tIM42luOM7UNNaaQR97mN6R
+Vh22DH/CL7YOMxSOF6gbGMoAY7FXhu+fvGRCjEYdfRajMjT93O3Zgsr3tpJZyZF5aRkfBNWW5FY
6McVRujevPpg9FVJdvlsNSiKqV9hIvN/VhEER3fvoRW+zMUbE42youtY5eIW5k3DnH5UOgyrwIa9
+dywUu5YZVGQnRpq8hGmsC6V8YK7yx6IE3WLGlPSHcgM1eJdRRS8IGuydQlJUMXsKe0fOA2aq+PA
a8p8l5l8yRaUAYZpVKWOpGqTM5rN1N7yQcN8d/9EsQTm11uXOkfwX5LJrkWVZEzqIBjM0Nbkd2GK
eU8PHD/AOVb9uQU/Fj6VAr1QSE1u6xjOH6UJiz+V0RjmKlV59sxYv9yaJWpgSGlFpSx0aJ5xtIcN
ATMBj1QF2LS2PKimmuL8h3TxVMsqawXJfzudocqjcutlJqrVxSBRm4FPVC6bx7GAK7gCkg6ouc7d
ZPPp+xGk0IljMhmuBAJgcniQ9wPoEArRTB1MyxKW/IZtrBg6217+mWWx7UAiXPaS8/Qsk3Cnc6uy
90FX7c2cOthkHIvu13YEUylbtGnpWdGLkHmLP5/bSfPtFGenYVH5EYHAykZ9TufLrxI/KCQEgtqQ
+X91in3K6ve3gkpO3dlrLFd4AJw4QjEijDaFYHEGyuyBNb9Gaj17/LZzInS5HQJq+IgnPNnrMc2F
f5hs/n3UV7uI/unXqsE518MNAXkHe4EAd0UcYgqx8BpO3RL1LCA/6p2BERTPnLuooTWHzWexTiB1
59hDmjxnUFNUf5IYAD7uUiSBk3ozFlfYggImfnSYxXGsQMjxARLmOyk0HN3wnsWERtOgA8ImZHhW
9G5vmOjn5w8ScemKpQbMxkDaMFFd5+NgWrcSKs/NXIZ3i48zE2xyBy+5MhkKt3W7b1lYm9dS2p2r
YxWDiLPHfcpp055p3SKaJgIQYMeGnMG8Tm8HMOpudO1/P4R/WPYW8wL7GbINHaxV5nGwpqMx+HaU
Lj1dYfGHEFrXTF6iSoIPSN4LWX5M/tVtdUKZRoudDuLstW2/aTOp1eeO/P/zJl9DIAIyXmkmvtPs
gR4yOy+3zt8WO6T4mMCsiYp0O/wa/uLjq1zmeA5RJJN1RNHaLF9L7oO7ropqFKcXzMTyKuweFkda
bRiqN3yciVV/3BvQcwrwVbVLkeudeKk4yGgTNIv0ekYgNlYuMw6NrYsVAp+jZF+lcpieBW/2A6gj
r/bQls9X9dXA8UAg085aFFS5cMHBzJvPGBGNFHp00KdLMIlhwIHsLtYa3F9KuQgNadr+dRchACeU
exfYCqbGlVKRMheLpGGK25RwyvgpbAE/6PRSudR4hVA8LHuCwj5MsbZXPNHYdtICCll4FrOL/gOe
up7/a+Ph87VbDrvBFztOz3iVjoF+SbIS9OgtimlYyYRd7+u9j1+PAIUuvZl7OP0nRPUvKzUv8j+U
iF0jX7ngXNhZM5UhyAcmsUSPpQOgsNq8dZSx94gtY2fGwZr8vfmekAbOMBsYZYvzEahIMibbQMCX
pLLjvzTGwgW5d9SgoNUeumAETIl+h+uWKUHrZofmCe7ZWg9DFlw7R4mW3465+JGni5QozDJtFQbS
Qe5n0n3o0aAXSq5PMGyRDMyWk8Xo6Bo4he5tbPCu1AtRSJsNEtP1Lg5nLSLdr/orl8soOxEM8Gdg
WjC1z21parGJL7uhsmb75i6NwWoIwkN+VE1uBo+QMv3neZtl/yEvzQ/9unQAuQPyrEH2tYS/c6JH
KdDt0Ay9tgUazXNPjt5s8Phach+bUcpMPb+ASKhA+Lh7CfS/p4JLH/b8jmXIm1uOjQEDZUQbzOdX
hkppV6qVKDV+dNnOsdxqyLTqQ4EnLvxQSaIkWLE5XKC+mkGU+x8S4/gbU3+pDym/7oBsS9r4NVxo
KvgS8ErcguPRngkRRnBtrzQ1HGqGYkZMHrQA2Exe0G2iM/fZTI6p0OvbDMvc/XpwThNEhkkWWbbe
orgnf5P4r93YKWxz4lzYg1z6GSTEdx8kKZXqFaclP6CxQj/GZoMc3tse1ioUtzLvsw0/zAN8o3/u
TBS+bbEIAdggwEo4CQvXeNiKtcTktV+kPfcxQW64VCUFHbtH8NRG36zftoKAByuw3ECZv2UC3GH6
Dl2AT36q9HZcxTBtG+QhiF+OmJy3Ce5i/dT4CBmIDOu42MehR7RUugadcKYBkUkxg35E3P0j5Oh+
s+AkgfN0PTKdYqONHRjQ83fplaI0P/NBl9bSiMYF6/7oISZLwLsYl4gLjdJoPLk0v8KG/0MmloPC
4DydX3PqTk3QsLWZE5vr5yaukdzWbcvRebhQuM4sUFcVzQMXPPYQXHgKdWov2Ihuzp3Zou+oUa8+
x3zsyY2CJlTtqJ4IYpFcH0wVCe6bi/Tn4iLXvFejp0JUcwtcusgU9sQ8x7wJmkKN+9xbue7vEqdX
Wixf9eYMLc3fN5vTLrN1KBwz9dxHdnkSf32Y3zJpj8lUP0Z5uyYS3xmdw5A4XW8k6W65v1RAXsIC
qiZyhnrI90jugIi5TlUZr/ld6eDWWQbaIboSTttLSBr8l8xdZsHORFMp3/dq7JP2nAal8kElseUr
0n1VEzmdsgBik0Py+mHOpbOKQluBmeCswX9z0OZAV5/3e6iiJ+CTqe2kcie9v5NVB4XQXMUw5/nf
Ho1wNoZAx6jXxGx8JG1mTQb91x/kIvenuPv/BBFceaCQDGu+DtEA5GJgy+yhDvDtzX8YifnjhN8d
DzIEVBe68DoyRZ7ScDs+rnvRTJCBpKPQdK7FqkXs190PxDYbPbzPebhHnuAM1pgNWHMll0dz9beB
kgjf3GHKbosjnOvY2YevQqAUODZy2lQE2svFAcPbEUESecD9GB2aDWVhvUNCcP+3lqM7zfBJtlQt
P5drfAZF7+ITrfjNEzX0nZW9rHDvKck1NNcf5fJsleuJDNLBXDbzMitbeUf3OQKnCSGh0Qf4B95K
XafrPQsxnC+aMtWQT5Wyu3Yi0qmy5B/qS1jyz0BJidmuSkWbIywH/efQ6Et/kUcGgqOh/qVkDBx9
eEks4JQ7N4f5qcJdF/U5c4CUC88vYQyNwqHJ4A+7y/ly6TY+tOPzG+1t1YGM2mRL3Bcuy1BEf+aY
xH92zs0ZTK/WIa2rpHafAndzSuQLgfdFO+XbtcncLYTrujNyqLJRjstdaKuEppYl7ep0ve585EEz
MiZH9gHXDJ76Z7iPMhKB/Dwg+HfckrXIMTMc/VBo++qVw+fRBM2Cj/bWOdEzoTiCfnQc10fBbM5/
jo2k/FQIqiyTugsTAloVDXFsFnsaiqrI/rJwwQd6mfL11SHyRFcg8T1q610X982EZEbPuQpI7HHo
5uL+qQG4S9fBcdhAOCsV/lPAZFOXHoTT7dvT8ST0Fghy+i7jNlQQ2gnEf8R03X/5skpKmahfn43F
XfqolWlAWIzMPWegoMxdiLYuraGpautzttl4UeOUN9Me1I0vDVUPCqkk3x/oqsXdsZeP207FuLs0
IMbNpgHX9Bitgqb8Ixq/vb1CaRvOJP94owr64RimJPhDPG26/rZ0UTfsO8suJf8BwUsp6eyJ1Cvb
4bnFBQdAjoVQR+23M9PjYTPDDOuxLHIweIdkcLQ+RBiCoyaBiJHO0g8DFXNC1CzkEcVI64AkFjRF
heCwlrBlJiRlyaMDEvf5iZmoG1rVTI6TTrpNMxCZh87CJyXypoTS5MN5T5N/8mn5M4GKkdwkVeD6
2rps4OtZom8zEK0DYewJLgDkMLj/uiyXsyIG9FhBtkkheN7JcIkRyUK2uDJHxsp324EPJXWU278B
B32vwTT+D44dKH4E+ZgGy+VEGNHsOKZc0Y25ZqNxd6wFbjYrUooRBFbeBngx702UyvnwdDzJxkiD
xzeU9gbqg3fs7FhA0XtGwr1THYUMC7Oc56Ewh/FrdY0JCGW6Gp4PGaPlU4GkSfVGLH3oBXrZnr2N
vk4KI2UNeTVimHnUApf6XuoVkk3pBikmXDDi8O3GL0czKvVaOSQHQtzBJhmZ2f10nto7gUl8Pqmi
qkjuCWPWWHpPQA1BgOe87gCH1WB4aOBHyNWe0jhdP2g10IZ5OFB0IsC4Gwe0sV6fklEPTAcNXaYU
i0686nRqvbuilT7CjbL+OiRxyN17o9kaSrd0PaDY6qyFilWUIX35VyL99qKF/93rkIskX9DKGJWg
MGbJzKWWbfsUlyeGluRZrHS+9X+O6zmGNIosvlcxhWJ+BHWgZm/2s3P20fWFcfdCc0npgqa0U8ja
F0EDy6acc2JH5oBYlu3ml0eg66IEZqwjTYTj7/LeBhMZuh/4d3EE9NbXjjnppVDYdD4/n3j8mDsJ
mzrTxc0LxIhVUyD6ih9/x6Dxv/ZE3wmcsfYga6yyqyxVXdsVIfE6bmQnWis8J7Ea0E2xlO9F4gka
EPk8PKdf4yyFUs570UccFf1OQTiLqHIqTGMtvlejzB3yIuERua4DW+n8MH4wa3W7NOs9nI8R6T7B
Lw4HG81ulf/P6LgBJ2iPXs3XiVcrigOtjbP4KBRFMexIRPMsoBT/MuTLFZxyfdixALgvVD3K0YbX
O8mXSzbBfhgHP4RSAhfq9ZhEGIuP9rvCAlvWs1YjFXv7ugq8w4RtUzEXrShBcDxWHjWUYI5KSIAH
qPtJpAKOqpgMCV8NOxeDvo3xz/gQnOON+FBED5ylXVV1u7IZjxCwWwF9tnr8jSAXQVJQUzhGRniB
ad4ectu9zzMeMmGw9Wkg0fKUA7ApeTpowxOVMl1VnNDlHpRC3p24VhrZFFr+3YN8I/P3CeHIDKW2
qsPnP1EO8t4qxt2F/Oh0C0Uboz3EC3nEVysv93Enq6GEhnJSTWoQWeQcoWC3MBsP8jUwMGK1Pkqz
APK5QS4kkdLHlNXNbhT4b8RGXBP9FCMmWtbXaljrQosF9hvfew72LGPWm0zwd9mXzJuQZ7pCome6
/+Nnkkmh8Nrs7Tf9b5wqENgspZBGKhWjY02KfCNaNB48UPGUNV+LLr6Lqo0JjnvEM/SyPecPy69m
dSxUTfjswKT/nFRX+47sqDWfUqjkM2ejQpuJWs1NUTQ9AWIk8lP/t2RqT9mf9zkf6ldeh/lhtyuP
Qr7yLE/5NGumR7is7NHkPz+CBUlA+DFW/1IWzxpyryJgq7pKcuPn27hhBEkI/lXGnOgyOSq97nsi
fucGcRa4ksKnzXr7YR0z78iKRfENC/ghCz0XfEcjgP3e2UKqEvXPR9vHX0uXOfRNCsrjOu/ihlro
L5XFt9nlQvfupu5DgDUiO9h5yPSFmMdkFu5jYqHMNBi6eZ6HvK2F9qpFEtvIRfnN3ti0BpQBI8ZO
1aFjU3tZ/Xqj2nmdCRAaP6VjEs33ss6L4TWxob2B7DfszQ99kOPdHoVbURvTuDSzccGqlXz7dd3E
z2i6lAQtfuUPQ5VZm3hYEjr7aPu3XC4mLS8A3R2hwa2jrtBs3qH9boe749zhFCYOrJzqIRUd4M57
H2323eO77ro1HS93WIIgGGthe22EYzmyyIebS4sN6pHFoJhPUlx7Ihuw5AFae8kfqvI27gvbVk+X
sZYs3p8M1PGupBK0jmmdVNzsB5ndVErIu1EHlvSp6XjpmblLDFSxVeeoHg29fhKVjTsImvpaI4ct
0y2ASc9wRIEbniSqyu2eLfCUQGLD833Y0HLYXc/mDBAanYNS6RbZGQaJVm97l3ZfizNmmIbUjCaU
puRyVM7enMLldq6IOxNjVm84hmlsIRZZZ6ebNIdcfCmt6gLDpQ+EsxSjpDbSH3YPu8FCfyqE1kuR
jjn/Ab27ST8YYesG9V9vNkJYfvgThSAFpSxPfcvfNm+5AVGQ1pzPpIO+uhA4qrQsp/ieqT9vd39Q
fp6KUi56U/thPf4H6yVfKHoz4MV7vSzvocg7jm1GUlqKZ6YEYyGuXatzqkD6g40xm4Z0PGMYV0F2
x9sxfxd3ot1+gAsYMTBbJzgtRMWUS7VC84QkW4HAmIXRdx6JGR7jKTKnfRUs6egnuctugDqZWKGF
+ZkpLbLKoVUx3wrGE1UjuiIM5LEwBsEJJ69w/SJtjmtswvDQ/Xm/GcRfXrxSGUq29W9P7C7MmQnk
2Jh3zFQQlSt79aAwQ5i6RoZF+G9WjTpbOyFJs6q5HUAaN3X8zmCBIkZg/2WpfUK8zqgu5/i4+0yl
0waNFB/f3mEq+4E4kzvbOF3SipznxV5jpIuA06gq7Vq2gX8vwrVo1Hd1l/46FrUQuClrU8V6xDcr
4nG9NLtBi/FcsPpv5AeejZnRkpXjVsG2DRl5ym3LPem3nmNr/qIDpnt5ZkKwW96EK3086faaDjgo
K/ays/PMTVDG96N8meCaIpWL9CFXMW/2gF15rJS7lyL07hFCP4i7MyQO9cjDSoPwMMlU9Jv4MUth
5otWxpN4W2CF4vmIJJ6VzQa+fKs9HLxf8zhm5ZHW7urOe5q2uYrsi0W71f8U+VrGbQw5GyaRpmm4
05aiaNywygI4Jx8pHEL0uUtc8CDIEqs+ldWbnOCHZywZz1Zkj/Xbvh6kTKAjG72QkLcwj5mc7U53
uI8cyZHlNtXN0ahRH/nB0ejUV58ABvlnPew4UtSr3GduiJJecybo58DvXVHzrbV1QcB/J1ICyBXY
jsb1mzbWkZB5PKfMuNohpO4TI4m9y1JEEaw4K8lu5rhwFDmxpfO66vLBt+IwQzgIXzmtv+3yMEEP
tZUwKht8KZ1oatOvATHpXsMXD1vnXqDlZk675rMLq367gobJScZ91piwwLXwu/BTDtvMUGzydc7I
Kt8qGj1j5WzJe90ejEbGHs4Qpwdl/Rjlgw2QtyMAQRXZ69V1ftESz+DQCR+endSwUeP/4odxZklj
jXhVZIQj74cASud6LP/KtDAJWMbOsP4VA6WqrWCnFzFEaq05HB0kEgjLcQjAgv2DiWQqE+a870bJ
/K3o1smwIWTm0I693XOOLazbQp7+2MSkRp5yVP4OQ8Yz1l5+H3+7ykQk2U1K4Yck188CBv5iIOFW
r6ayr6tMBETDVRxOJhiucVJw7IfYKUK2HdrnLekvkdMbwt7MXuTV3VCTxK07VvM27sY/Z9Tg4Ugf
NHPmXRcq+C2wEJMAGInWQUx2SdAudrkj8alunPSlY82f+0SrOXYcUHYwRPgIvM9IKIVq164ASkz7
ToI1ErkjhiAm+JvnCpLBP+FcwodY6VmPRQr8Py0Sqna+WCGSPUFB1zYYmcYaeS21wzcPooBFLuh7
YgEuYqJYR8rI0ZLKjrn6DrTyljGmSNtjU40lthYPnybtxWjR9KMFOqpU75VrFjkurZzVHvQUPH57
LE4qsWYV4RjgeptB/KA+8y7G0EqpnieCfQWorybxkbp0NYQZeDc3jvjNOTJv0wFz5ozHE9FYvMdF
HTyMD/M75HTUKfPZlJLWcoNQVFYBmbuqhMenBscSGBXFRUQAEpfyF0FkDs1Qml/nPAU2dudyI20V
lyHKz0UewlRXqUtMG1+hfklczAPw8BgHsR4iqc3jas8PbWsEWDHMWxj4EXGsxQl9O/pxTBLnNreQ
5kUC+1bwe7T2LTkmorVJwjkSck1ENqSBySw3YuPui5BpE7FW4/LiYg8I47S3h79EaUl0zQn4kTh7
XqUI+kV4RjjpW+AD67inSdx3r9wf8vF/f5L0q0F3VGQIvbCXi9MClrZKCbxOjmB8RtXNh6iaiGYJ
NNb4l87uUPlmCNj6PABsFMdAuoMaroGF9zdzz3zBycLmx1UrmoqIcdU/yKrr14dOdte6RX8EwFsZ
rodNYjddBMztCL+iG2gLtzwqD7z+2mpwi+fNS96fefY/apwI4mBQhIusySh5/K+/KTMDlbIp8TPB
EdDQyQyCebUzDzQAOrOH/EvEGJ6mjZ8xG7h22k4Yt6piLmsHDsF1LQFprbuu90r/0NKbofFkampL
U66tz/15LIR/qhsfWYQDXyffjS19rdOMOPxMzemfsF99hmOsNLsJZd/SGkib0ff3kg2W9Dm/s57M
NTRte3EdLNaHHqYKFa2vWXD2y3kv6XVDtfcYrX1Ak01k2MfxxAAzHtFvsgeL3zNtqTnNvpn5Dxpr
OQ/C/ajlWkze705793/KKks2QWRlUZNwfc/g9L9a3FF2/MN0sy+vKLzoOMOiiWY/b30zJhBcgcFE
IHkXJAAzU92iFuW3GcPSFhLt+blnNnXpeXOqXKwkBXlWwYGfXq4dLXKY6QGnnNYIKwtRVGA7zzNC
hZD2mNsRewYCywFR+K9e5Aem7BIBls4QLOBynAbtgLkcsksZ8GZlNTTqauo4ybkqqBq5GmF2iJiz
kBMhXc+Dq7bnN7bem0qNe+7yc47+Mz9jRYpDfG5Rf6ElGpr86rCH01H6qttfxA++WQ29SDuOHy8B
f5Qxqg2kzeQmDIa1vylDR/5E2QwSLXmCGxxvppB0SIDHz4hXMz7ViM/zUHOgLZ7hPAlkKiGFjziz
xzJcDCLa3YKeuENWXjQBz3iZw4jmGuQTM8LzR9eJ2JHCMxYZ0MkhEh4A1+w4UBhH+gM+BFz2vW9s
VzLPFzomTpp88GnTFY0PQJSmiQiTuEWf8BoVDZ5Osnbn27ANXvs87OK25Te8YM759ix2mE1qrbuy
obMEOOlZnEQ4HKZEm0V28LxV2FqaTOTp0V6ATRJBJInChqXMtyC9y6iNqG/8uhczPOHqlgRBs8G+
KAw6QQMSrTAmLKtyNGZmP4Ta3bU3/10uGWTrVpSiLTDC+kR42yuoBzJRRrk1RTbmB5eTVNGpvRmW
JV7aRLano6lGgNbBiB5Yg1OBZZO+Otkk+DWOLkmjKDOA41hxEazgb+iM2VI6UXADs7ooITsCy2yH
finX6GrKeNVTMZOLOZGqZx5fF53S9jXaQLH2W2DwhGelPhkon6+Wq2GwA//9u4P3vXSCzNHEekEz
YsMSNxXIj8DFvMLkBj8Mz88RuyFZ38ua2jQlSYdQwDidlOj/KfT79hC0LVUBoQ3UmfIqFQj68Z4T
E57Y0TvqeNB2FGXOhN8AhAgwSlzinyMt/YTM/3/CpWQ/+NC42+qjOB7hObwV5kHlj3rL7TaGzUFR
Y32Lx39LPXYCs8ZQaPg7vbUjLwILzPMiObahIn/rjLK6pgj4kg5piHeGrThm8XA11g757lqpdfMf
CydOyl/TdM3xXwpmXxzeyu3njREETmpAJqw9CqJM+j1ZjvDEFqaqaFF0CmNL6N3rvy8tEE6gfFiE
BvKqhVzegrHxW/zjISKSjRzNZkh7LSz43bXUC+NYni2eYTWBJTso8SUMYxR/JSkOt3t48HmjqP+O
cCQDKn2e/H4zEae1snQ1MhhHpP9CuHLNhWsoUvtXpvgqfVu3TXyEonD9LJnV1lcrXOEZW/WIg3Q5
CkkCe7VeBshbWD4fJ2dmDZnamOLZFKBRsz+C2KP3bc/Bn0Ce6aMv3VorXo6QCYXXOIhe4Ngi+8BI
KLNkRsF2pvm+u9opJuLZZvWmUjMZg9sgokBNtT3FA9+bTyw2Kn04gEtwaI5ORU+RjNEDczYiFb+8
CH7BzufesjdRL4fct1E2PhtSwC21fi8DuV+1siZdW9UTa6RaHjOCVPmvX84GxN6e5/HbgcLBJqA1
7T0b8z3nPD2v0pldSi+eKzTZvDCOvBUfunCedZmxjoNkGinB7sg0/hYjq1cxuGwqlu6Ul+jEUwto
pxjVSgle0ce7Cw8T3n3AOmRwjyD1yZfni7d32gvGU+Vnx+EVGoIrzAh+UtjeB/PEUwLi0WO/KKhf
qaZEr+rUpGHe8rQfAfYs3rvTo0WmrdrHLL7KuHPd7ZzR7ujrCf38RDuJltJIMoLtFBqfRNLVHYiP
O20kGIIPEJWPmJdt2Qo/QPFaRKOcJ89533zZ6pAnlV/uQ8YuxzzAI+E9ZOCoKGXAjTNM8BQWTu9p
JYcyqMjuu7v08nw5tK3uqavP1CS3L1u4TFELtPIIZJtEOLSgxXhMMDyQgl3WFoUiz5nCjpErGEtR
BBWDzSA8xU0vlkBQovSt/Gpssh80OmtOwVRAbJmdvrjnHkcksBeb3tlXs3gV4dFmPY1UcdICceL1
/jpBNXSv5kwGWsfgBmRI4o7zJ8W5/+0XXGXgrjXwSSSrpfmZFQsdD1R0S5QSqS0DgAFhvcrhT5IW
9SMJOfbvGZhJOaHCsBsUIbDNX6RQjPQNdaMrSB91O8z05ThT/z7qa7tmTkdCijb56Xz+RQGKkZxv
DZghhxLGwXbS2pwP7Y6HNUKDd77crsmiPpuZmGqIgGWBaNbf//Sl1I2HAOTNVeV1XX/heKc/DXrt
YZ2v9BBSk/QE6MkcTZDJbPCBa4r687hHSF/73twlHUXmrSC+p7/U2BOv/AqHncAwsArnWChl7UjY
C8CX6DjnvPkRPukMnky0MY+XyJX4dhTtaKAc4q6Y1sWQerU3Pt9mYZpcT+ycOWA0VP5JpLXVilDS
IL9OIH85jBzsjjlwK29uFSTBbcEz5Q0pZEfVwYLD2gvfcCn4IOGnXrwRKBfjfk7ie379893HrUqM
EaMgrzqLAB16E5ugRjJF5cePjbJSD06krUhCe9i70j5zQfFJ9VuKoQFEVp7kXKuPEF+Vca0uPxzB
eGy3RxcQhLdB1Fq9KpKhi3LBIlOx02wq1nGQknAPJEY5ofvNwF0wj/8drikWLjVxLmOkPslUpEm/
hfDm+tU2eCAfAvgtRe0axNgLctKah89ifKSY6HueTJTXkhepjxISk4Eqt1fKoteca+HKbnvR6C4O
D1/frGF4wwUvLsVu1VksgtKmpAVspr3+krR8/PUg3iR6gOnach9G3Hz4ShNeV42D1gJETK6ltMSK
tX1hXkXZD9tIQqGmv5RCQsrZw556h+GVsruTqPTl6FjX33/hgUjAnVcIvUYK3o1sj73Rew8j6+fT
pX7wgRdnNhPVbcQ1SGuSOvK88W52VCrS9nJHpL6WelHwpQ6p7tJNy3UBzZ93COncnrRAu98XjeqF
wYwF/gp08fsvVimT4kXU0ABQuNjAIWz4Qa5Job29jfikqg0NIeXqW3TMHpAVKLj7TqUor9MRgS+7
vKhcahNEEnBauUOkzeFDwEPjsqT7d8WyFrs8xQbdDLWJx0yWMuQ+K1Iukx8kerBuOb5cTYjiTF2a
DCPXPWO3yNm/aUAmOOrsd/HTBE7SZpUnfLHHZbnlYralFSBwN8j24OPxb3n3lRifCYS1a4T4uack
x1AQju4szb/1hk9zqYbRSVsEctgIV++pAsfz5qN4D2MOE94r+h5zFb3I164GM+EAQJ/3kAORxVeG
diqih97ksV8VBG1OdMUCEb9AUB4E+zF7+Ed6IyVlF5heVPSQ/8WAkBlIm5R91XP9RnTyE2VGlxe/
SBX4AKTQ4/4bJUBQuvfLZzrxNa+PSCo6zOHwHigJEW0s2fwe58sh8nXvZResHR5K3vw8bwHzGtzS
Gbg5As25BVqNpKo82RxjS8YjAg1+aMT7hgafHgdGS+MWuThd7vZc6uNxKslxpZ7frMS262vIiqQS
uiw/x8COmI7s/4NoqvkU63oqeGgaNCd6BO+8WWEb5eoBR4SEdEugNr5sDJ+Cg7UeszacdJNS/h5w
r41dx1wxfP3Xy5agalM4mXbcK4OwYuCKZwUYmcBGjtoW38BnmQicfCqJgwxY0PBFG2Tr9mIm1gW3
n6Z3r/ueph/TUsQ3ifNfR4Is2SkfgQc3JhEha8427E8RBZwLezs6PuKHfiZ3GtjhxVfOPmUNn7jQ
ojp3aLCQ/plaax9BQ9gmiXKA40kku20n0kawQnsemqLZ8pnbywnA8p0qNrJ657yc7R3rl/7bC22n
cILZbXNMHgaNxGp9tuzPUG8sJRJhfVuc2S/2PqFqgGt5mGVOdfto6F01iv0nLX4pfLppf5vbjqhw
hVls3FRmFSrpckoYOMmQ1M2/YZQOPm7Kc4PP+bydLGDM0Whmwj72yNQbcCyqojrYh/Q9B5N/+skQ
D1XqwpkA3EEk62ZC+W6Um939mEGrdMf4Idy2UImrFZCnXdQQXk7ArPGitTzE6tJ8XlEqd0N4YsfP
W2WiUHW0K1hmiNvVplsoQQ/sLle3ozXFTAagsQu6wZthx2yR6p8w2DeBbHD3pDel6o3z1274Tcr8
nTWryHjIY9DJVtxjG6L5eRDFCUigcEKEmh3NzX3qq49ce17y8nvQhnNMgUvNk22VkR8pmcAXvNUb
7C178P7GgQNsIaop1Ub1S6Orio0bddRWQwqVfHeFHcksjpEWNqiFDIxG8LLZ9p7NdHMIlbooWEX+
A9jfmKDWn3ZnbXOUE44h0d+Q+X6gvR2SBo2QrGO0MLgUGWWVT7wl/IpeSnKfvCrArTHJitUInzwY
iB3ziJuCNFEAbLEoXG9RDjmzy2eK3tMrveh8J5Kc3fPCAmwOzu5XnkFof1QZiOzogvTwMg0z5w7N
KE2daw3jiRqJ/WR0iR/slPziKcywiwdGmobAGzk9paX6JOaWmIwnYeuXkSDM/uB0AwuQDQa84VC8
uzFrZtLcJnkC2NjbR/opUlwYSVVyB6zK/1IdcnV95GDulfFCy++WT7TxrWvXbkbkIcuv+roHjZwg
mmxZUAfoot5CnaqpF4huvzzhFda6qNTyKDdTj3vi14eLilVt0q5/aCcu3l0ahhKpt3n52oeo7CEK
44J8SuQrhAfHqjiF7OSirqJy7wl6+B72mmVxxXU5R5hLnXKuen6j/IUersE2kb5tvWrxBaST5nzR
rXbOKzDjFfnKsnNzvA7RPoYi5nuRpLbrGBpBJkrtB503mbGu7DGXtsvjF5VrR3oQOHS/skmjMVWd
wgQfUKBRScbBrYKaYjBusENVj5NbXQhQxPdoR2wOdPJqvw5J1Z8FDuwnUhra9vDagpEgMxfZX0he
nAVb0otuSFAuAZbtKUrE0qzh0fxHuR1jsJUCctSZzjYf3VNJl3zvVn6/WLSMUmETJnwVK/P5Cg/m
+D2lj3mHT/Mlyehko38qs7UAq8huLri2/T3INHuOwwg3MOhyusyy6xL5cz78r9k0O6hJdUdAhsLJ
c+2G7o66x/oLNvBHqGaqMvHeRQuhJIGwstZJjVJkih+wKqW08UgEfmJbuKYrjjBVG/Ppdpvw0fYL
rfU9/Zk00Xsv9VhqhxqhmI9S5ZVEPaqPzFBpOtLnlhXRV8iHRzfabXIq+1J3BT+AuWhri4Ehp0lf
94ruP6RGPuZTHItjdnFL8As6WXIQUGUJ6KeD330pivCD/jJ+/w01lyNiC6xTRNYEX2gfDCe31k1i
nqwwsEaWpzxtIefAJ4xl9+zJT4XQ2zsbBTzoqxKsnO3ZLMHBdFh52s5MoJGq+nfwlkrMY1xQXiK7
2dhiIv6tbBCXduD4b9pHuOn38gOJKcGI6pJ2P5NU/26CC2VN4wqPHRv/of2vH2DSl5fHhHWBc98H
ajOTbmiDWxCnHVYRghY1t6z37XEnMuVx36BRambx0oIVACbCitPtYk07YPymJEGFUAQmn4vFDHn5
v7B0Gnq4jfvcrAUqMnbDMicGKz8uyeBf2AS2QtEpbvXyj6C8XyS69DkctgIXk9GatrpiZtJ4LN7w
uqc9X2feTfX+9Rzs+xHY+ebvlOK7AHczvAsHz8IM8p7+RvwRxRCIKuq1QhQ4EuSzPQvCuP5ZRF9+
JPmhzW14hPL5mZrxB1HEKU9FpWR36c8M7fcGKbubL8dv6iyVnnGlSw5e9wJ8G2t9bTVhBco3YyMk
fSjNobRlJ/Z/nOdS3PJU4f3zBJUfRRvc3TpdAIIBoxklQDHYo4wjTFcbVHDKA3gPRE9BL6nh96w4
5x2KdEiB6/6YKjBdwwAqc7Hee2kvE2bxuC94KE6m8/fy1/yNENtjGfKqlzcBSTj3cw3C9P6i2j1H
TewLv9aCdOwZpYY17z9bIwp4GhBtqHOabNlh/QMBnR0mlWEknWKfSYO6kp4lMrryiwpr+mIHxR9J
BEDqiKgtN2hl60z0Y5swVj2cHBGcRi+K0utRftXiT9qg+IVuFv4OVqSx1e5lNJ53IHRN9XlouyIa
FWDVLTI65q/8czmENrFvc4cBI9yJi9fq4a7iHuvJ66PSwkWxmf7vDw+Ubh67zDvqKk4fa70loPQe
WwhgVdjCrbMsTL0uyi+7NAstkM+42KV6Q0CxZAYLMCzhwDNks0PNTOpbvbwfPuFwNJiZc+QDv4ag
ecl1yKM1Il+E1KAf5QM3U8jGrytBpX/JFv262oQgqDAGWpWbUm97FewLXs4EvyOxwNgVvkJKc1rd
QhNp8GDwxCG7BX7Xf4bH/dBYtOEbhwS/LpPFu3oByJ6lmWn+1nXlyPblQXnL8cmGC6l4lVe28WS4
dY2stCyrxB4x3v3RBJMw2mT2cKSxKSTD3vqCJIV/iLJF2uYf0DRLbGLoQoylEMIp5+5l16wKjCAl
lTsBoh6omb3ndVkdKVMfK+AgUrNfgj29P7ZOKGv+QtoM5uS7lgFFWhMZbD3ntenyhLuQXFinVfRa
HSYbVfzYDftPsy0qc1jYsACg2fWkvDXkmTwOzp1EDmGEE40+p4wpSBSjyqisAZnyE1CttnYl8jAY
x6H6DzhIbZq0428uEoHfENUbH1FPs7F7Sth6SF3Wxpx0hcgFE9vFDWQGxKX+MHjDFd82s9mYlk/V
tLLatAuX75SbbMoE4DX2mlJVRKNPlDajzUIdXcVpuj7Pkl75wkgjIwyVERndjNs2PQRiJaq0gs5c
N+W+XEqKu1F/eQatF1zcv4tPZM5uDwXrmlrkE9bD/gZ+3gzcqz52TOC0OSMy8HEi/T1Wawia2Pok
yLGX9m2LouJSwI4Ie7y5A0Cs2n0tfF8Ea8IKHCwDrrmkWa2NmqHl0O0jUIMoe/q4+cfpSOJZCyh4
dXQ0SrI92SE0y+vfqvuBz1MCCDelHltTuONiSPWrKON+p56/L72yTnf8KvvSkrGaiAFVMs544l+h
nInbKSkIB+XWqafvGpnsxFk1yGNafrxFnQiEfEFe90O8slO7BgNhdS+V1DaNoOqV1jA/UwyrR+3y
XI2GZ77xZlcvRUObx7e4eyHrtZE/b+UFII1dcpHCUSlS0oGEOjn8xICxlXyeBtmZ/DL9fpJskF84
sRRhNb8hyw018buJPkWGZ+ld5rlg2B9nfT/nVsd38lHxhROyKheNf6xuN3hfYEhoupssEZ1SV5XK
8QPaeYhwJipLNNi/a1do99YGnobJPb7nCkYoub9PQRV52YLnoBxM67z8NKzuKjaQxFAyxCp5hyBk
Qle7UlJRPamvuSo2ry6SsY5U7FkAmf52QPC1DAtKF33rGol3fArIwEdU1cx6/La9PLEmPhQPPZbP
CmYLt9YZQ/WsTmPRIyh9wrrJWT09pb03PB5OdABkdVfhC1EW8rhKjCQaTtnqBdZsuFXquP3gEDKU
BsRT8h/se6B/paJ7+mm0ExmQcW4TPV4Ska4V4grp+w/GIUrf4YS4p6lDEB3qw6d9OTNLyDMjxkgg
7vQAz8XJPV3/uk9cN6ke0GBPOq8J9P322y5IsmvZRENu7N6cgcY9Q0D01yNcFSjdwzh7CDTbLVsP
8HDwPeIShHR5i3/9rnvvkl1UoVpys6tGiloNy17V4SCVgcvkKtm1JZjAGb87fY8NHMR8XcEBkLnl
EtJEDZMmHdWqYcuwLaCu97ii5Z3gVwnqYNf/J3tP4Bty0UerMwvNhH50qtHyMMHjN+4umJtFvsly
K798Gq/u+UFtap8dxecXdsYzDYS2lc6fowzLPaPe66TsdB99QT9nOChFHoKEYBJOuFDjnuCDFqWz
kaI3MfgrW/WWVTzY8DQ3y6jc5YoNW1L3RNH5Lq5GSWysA6q/yQueYcLWN+ZxKLFdmThul6Y7laMC
DSXJF2qigvRA+9JpwH09cEZ5BV9ybHLqkyS0yMgF1bS//tTgT0yp9LDe7A1TP5tuHLyRPIZHbYkA
eTsva8Q5M32jHT59Y2Sh0E4VnXb6n8M+/WoHBsIUrAyhDayEj4W1wzbS9+zA881XVnD601ynHJWr
dQQry9agGDczWh8bPaLh4tVGfjQHfElFNleK/GYxq8Dd1aIs+sbeUwD7NlApDiye6Ai6pexa7rmW
8fzq0pQZ82A8tVdSJMrdm4zsAgoU3NSskeUjd0P7htavJ8bgScmlzuzrFh4NYUZgDhyuFSj3gDHS
ld5aXDMdJCbMwpZ5NorTdoknftif/pKEg+V5ICxkdpYcARQO9vewUNIjufM75Q2udZ4k36mKa/ts
fFgDRJcHHYcekwiVixuI8g/MZx1Rp923Yc+T0XKGlcutmA9ovmX2R9SvYGLkhgA64zpo7Lpncs4J
f3FQwe0fAH3U6L0r0k3DvLbLXj8kdgkScdzs0fQ4KTGTc7bCw8IJxU4VgZSYF9S387ypaQMvKMVH
dvHd/qcjDCNho2lil8hFMq6b2jCwXSEPHnfaGhKQvXMtnd8KkP51zs/S8uUSjimxuUphh1jX6cYj
JM92tBQMVzXZHTpHi3JlkV40rSDLTEPskqudYc2Mjh8nyNpr/jBTPu1cfQ2c8UVaQnhS91gb4R7x
HUh0m2aTd/r3O+VY8wW8JCUGXAU2n/pJwc6dPrx4oJN4MVCp4kanPR5dIKLTDOX+zPILOW3nFJI6
A37ZsALYHpHvRQDK+JZTII4a5yiHrNE3aZRFiK9M1wWphf1QdDp5t0u+Aoe3UXuuLZEDFw/0sg4N
CoUo3wic7FOmw6fZAuAF8p2WPP9ZUfvs8DRaqRFbFopy3S5or8geeAfQrLk/53pGOxv8qgstrjy8
L/eemrnX5lJ0uDtrnE3rkZ9ZVcYW0ISC11qXrR6rC+bHcuL6iGQEVK4v1aPueuPMGPLpYALk8A8+
hOPJYoiRodbOM6kokbdSo1JGSgLZZORa6eQIZyjSBnLc8JI6/exx18KytbhllFOEgRAi8nLLY0/i
ckvuUpDxl1zDEkKO1KPCn5C6FD2rHqca300IAtOe1aowKmoMQoVK3OCSFGivIGplYKgqlHFxFaR/
762HXSEYTog1LeZgEIh7jXHKXq5qqHyfSNdDwrVf+mumKxwcR2DBwt2+dk7fX5EgCSvFXl8Tw4qz
Qev26zhc66MmTVDk4KerT7bEZYQh5OgEEyWRisVXHHZ4fzOcuUuPVodgTo1apgGvCKWtHrWm4eP8
iuQruPEbhgxMSxjq1gYKQd2AI4DbXN5C7eESo9KVFbu9XQtlArM1NnqHiJhzv/OR9w5XKid9kuBK
rXZ4PuW1P1POm3+KVNRbyWfNvJOKXmE4KrFrzz0H8YsIDctqBkVg8VDZJQl3vKQnwZDZnmnfkzud
BsKcYULCK2bio7bNQ9fZok8dK2I1yEBkGedZock/8xUwDqiu7hmQD0U+N0Z7LcawPJAlK1r8mA1f
fbWagPoricdb8WNetex3jwHNui78fPZEFmTTpHd/z8QyArHrbmuRj1KQSe504va6pIcC0/OgEprv
EQbhVDwGj42w8AbtAotOhd06t6INbu/A/G1TuiXwBuaXw/0lnpGgDQ7Cjeew7245DcyjGB6S5puN
Ryxjv0c5DBOtMPzJNANVHIUiNYKdwOwOXKvJvPgB//quRiC4T52ZBQCgI4PYOeYeM/q8r+13oee3
rjzG94n5816unpGmG8s3qWL5xIi+Sf59ApzR08Wxn8FyJ1kU9fSkbtuUqNGwTS8EcQEwKX3FcDCw
T9BxafpQ4sMi1CN3do8A36ciBrKTfuaXleh23ydrl0wBkbeAIcO7Ez8ZUFia1E4+ZamrrwxaYx9C
miIznq3IEX08REGbr29Hufnl2OJ1/8YrHWDlgFogpqWKblFof96TmQm4D1TiJKaaP0cvZeg5LGEW
U7bCdjcrvaITPGVeJF8rGvnGdbKmcL9sT9AI0rgnnXuLBn6HPT3y8PSoQFaKe6ZdcTht32Pk5ORc
gQKqkWP0xRMfUcgbMHabp23Dvi92Ijp5nStRa/co4XQdyNtptaBLWVKu6+sADwW4ZfTosj291BqF
zMXdYMoqNT/2s6T8OBdtMSBv7WGvccceRIMgJ3h3yCjgkvAZhq0SeLAv36RZt+v/YejDG6CiLkjz
raBllBEScn4Z6TjojchdmhguvlZS+ZBpGMMYJ+sFHHB2PQE94rlfTk92dZFmE/xkVrHvQqxMHrx1
38ap0/R7beFlb8imlwQnWpoLjEq80fJJn209nUoIqvAYGEVQN/W2vUMVcny0Le9z+5h8X1pRQ3LC
H9yOOeYW4h9Umuq3DsvA6YPj/NLyEeSMBJ2p3iBae7RAUq8FSsJMmVbe0O3G0VkdFFqFQUvKIgLS
MiBEsM8ot7s4XSuRe4ONecOaOXqP2kCaANbvwY2Gz4Y1B/s5MA6oCmOi0oJ7b5NcVerm/x8I4stz
EvmCuGBWXkTLN8kMqhBRprWg3HaJAScOAPg9I4u4xWUbG9We/jlPzIqndegY3ucmes8pst1c5cYW
SjwVD9J7hYHxzzDrpi69+ow1q+pMMNih1H5699UMgmRf89p1c+IowH76dlsyAcmgjKaur7QgPFU3
axh9GsQy9LOMUSOBCwSpV6p5UvHNbcUu3Fts/o1ZsLkmtAxrZbL/YwPpjaK0/pEfb3iNbN1sjtlP
/SjnXxyuFctvv/0PrcncjpYtu+Y3kYJd/duYC/6T8xgnqpKtHeH1VHDnnh+hXoCzPaP25bDOfieE
3B+HhpNlhQHLo8zVy8zldnBbeEU6RV4oVopIO3iW91RKwphq9Or2bAVXrhzz2tqMxFBm8BTm2NsD
Ks9afYHAN2YvkCUNmUOCZOEl8O8q30aa7qB0LcGSm08hv/NBkhcSl6K8tMRMbm/T2PS1hJ2ilT06
oaDQlQBDpEwyTaHvL5o519+0YHCMwdYQ//ApbFmZi6TNRFTlpxWs9DmHMERnvZ5nA/jwztj08iRh
jWLMwpl85rWGH1ej8uBKUz4+dnXv31cDXDj1j/7PMO6IUcEDDtT+S2rFEXCKwdKL90R5C+faiI9h
q1wVU+IiqwHB9R4VuINHvVTaiirtXoesD1kT9eYKlz7P8VDWZDIBnPXq7xa9pMgQG0yenprlcRIn
EFD9Fd07nz1Ot46JO1+iUIsnKYRQWcfX8UFVvmlSfdzMUIGgpWUyHGKHpibLPTETdVUK0x3oinjv
X+ZdIYHTg08AcZ8Ycji6Egv81+tvwno+hqWB8qnOoy4UDo8K4BWQztnSrsFgQv5e26zA7rLI+LuV
gSf0+dsPi3VLyd0hd/siWKsC7BnOudtEoPVqAh25hHnrFvEMu9jTsLEW6dA3hYUMNiUBpLw1kEcU
viDYk7T5pZiXUn4tXvTEJorV0pgutruSLUYmgdE584Dm/sfSvtndBogOInWAD3zAfak0r3EM+SWU
WIrqMT5kw6oRwW0Qd/ayM6fgi+Ek5wi4XpLuw3FRMvdH/AAvo5KCz5gY3YjPMWOmdCLmbvFU17PD
2GFPEg3uXy8p8Qg2om/Bh3KKHy/KKyz/RdqkGKeVQx5iakQcj5K9nbaP9dMfmri/CHiMvSZliI2H
PltlHsnIhYKQ9jX7JnhJo3RfQYui6ntYKUHOwO+/NeOHivTMKeuqpugrPcn5IATM5uWWPm0bPB/B
TyHu8xnYM4RKIAwtvNenv70CUqxdQsarsuk6IuD4d8Du25QuMfeppJTe4XsZqlBlF58HUmK8dl1k
4pNOSszHP+QmmxVwRY2lRHCVbXe0N8RQvnpvW/tlp/L5OV8cGAvNMcFctVDg1ZQI2nxL7Vvw8Yrl
6zkiareLeiXUP0wU1a98XEMmD6wP7KU1293IWT/iJqUUqJasj9dfGig8r4mcYh2AE55+fG3VEX4V
R2zDZ55XDuPudH1Sobz2RdvDS7Gdcu29Jq0v/KtECaVrBcSB6zxKXc8ZwOyJLmrjywDZ5YaS8qqx
XvGOso1HhbLKU6AR5AlzoYqdNSV8NxvAorh5FHaV6E2zlvz7PCiXW2N44hMc0V0minVtouc3PQaf
yriLva4Xtfyc+9dCXN/OLqepaQLwAaH2Y36I/bULWaoSiFoLXLdWias/G5OADQOCdddyyh+V+B9H
Rh3U/U1tSuYSt4XJQ56lL6syI4tbeOqrJTYK4oJmO2TVji2eHihc+MZurDOyDfXPcH/i3pmU2i6S
J4710Q2YWP0YB3qF8lFB/vvTERM1tHEB4XJuhHNQMWQaMQM3z3C/HI/6fMHW1xQfG6/w1r+Aal/L
T+zaHxEoGwMoKgPIFr9kgi35Wpdu4l/oYMVaFNG6Mazn7MUkKdUazCmzgaP59VbZ7WYa/I+Hf0LS
vMmGbAMwcEIwn+tRxxjceublfwhEBuaT84C5P3QbMwU0kC+0E2zxX2dBUDmAvSJvGPKqUQHGTiJM
A+pgI+q8+DCJGWfAQNBkrTlHrZ7iI7sq42c4LhiC35ntf5DmoxjVxkQgPfb6o1qkdwQy+o+0hTEV
7P81sX2gP4gzWe/B7hPRCa4meh3v8E4+Ifrx1wOXk/QEFzpOcnZNIBHjyF3XoQ9MApJyQFsdkcjp
kv8wYlR1R78XxaGe9K+UWpjQanmjDe8hWV6ryQX5xNpBD393naw6I+/a/0W/ZG7JuSMlJXBt87yQ
5c//d4Pb9WIzk3nQpVICKQ5bx3iY7+EXyrOxbtZ9IEhAC/XID1jGLvfEOgygo/V2gWxYBiE47mZL
jOK9N155kFpShaDmYeqT5zrUqbmDFTAp0Xy9s5JgMHxdlnC/ICzmrm4casg+Kbyn90FTBaBxmsL9
IQ2K/5UuYmQGO7kPblkH/DuEBnVhHosa7gFhcEZ+se9UC7KordodvUyH+uuqXdafMwOgydzY71wH
p3nrhv84ixwSS7K95CKcB/vhvdTrlNLIWminT9akejTdd7BI4mlHwRWD0olY1RsIxaTVs8+YUwF0
kTuI5HUjHp/wmcns7E6awnskjCb3ELivUkvI8LAZyVcq614mOMOiEqQTk2sDeHItR0f1XAXPjxER
WGUR7Qb1kXCXC86wnoFtlFY3iGvaK8CfEt2W95MpM4yP5phwD4fzG02HHXIavEoSvNSLXTdwSU+N
qeaq1Wc4jKwSkAsLHmsm4oCHJuUuscjRLRFQ5q7oSGsLYKzFFTJxatyniHXsI7kSXd2PhokxP7Y/
xrwwwTqF1ookMvjYVfx5bdfTCpM+CG5co2Myj7bHiV8e+Ebk/sXUSdSAcV7DM6HaPNkGkKKGVUNc
qr0jCOnXmPfZbfHAR6qnD6Yw74V34ccmRbuXUXc71fFg6pcBM+zCqUdbNl81BS/vnqAMYo9SfhbD
IuWeDzCyMj3IybA/+OcY9INNrhsgaZID7GkswI5mqtOvRY4s/0fcDL7FjJwCppa3rOQ8Cl0Jgcdi
IOJorS4ShJ9OPKtqxQKlOBb4uP9Gj6kVH44SWz1d/w4fOMx8dpakGq/+0uAKxgPl7Rluvh+1cn8S
RlEamD4IO64l9gvtfI+3GlVkrctoHCOkWF0GmkBDv+kaLq11xDwswfdZJxRD2ZZSb4VrfBjksUPG
EEgtWg1G9nL3vp2essKjqiddB4FuOiMtcq8wgTboO+onL2PnpQifVbeN7Ihz0L7Cb8QjlNqGgSOZ
/u4qgggsogyBeryjz5iwg9GiGKz4I0MXr+JOm49zTlzaZPlkcAie9p4NU+5kOInuYnqA0dhH+37R
U0aY95UwzmTKu4XwsWQ2hcdUXbwaLu3S3MOtii2ONAzPZNEgZQJfUgy85Y56++BW4labsGhKWLvG
kDFt/lYyBGyNKKdJEiwKWbaYHt53OYjmm1peKJQ0p8BQMzkMOfedJ0sqenUneHopiDmYWP0yr7BW
jTKbryHjZcfySIrZff1AHolMVtwZ+TchiJkC+waLAMWJ0OhtmXY0Jx/15FyWWO6nf2reeQlFBdYv
8bHxc9WVnGMkgpJMenciiIhZUEpdLl+NVoc2qVDZB9WuKOuE71yHv+KzbhWfg7APzlwIvg/bQCIG
BH1dvAI7cE6lUe9s37YdXmC8XbMyr/8SiR10AMUXCOzFPAcAEpx2WtPH631RjqiU/h2AONjHQi+q
NWntcydu3uocphTRFi2ZybGVYqikwn8oytdQf9isjWfJUySa2cyx2zlK+BHQL5e5qjDwstn+RRqh
GIoinCKWcRJS0YkNYDv8dMW/RKIKdx7K332v/176fc3JJfRiM8wumDhAXkegcTvlJI0KjadWiy/f
JUq9QvsfhZjaWPWbHDs5+s42ipkrP/HB7zfAEpd7PjWAHw0N0HCaZ9CFHfsI2GDc5VdSmZPKH255
8cittFxwmX2iNUebsRQv3WFCY99CbJClTtxMUzMZLM1SadvvtHeE8Luz/q/nBko1MKFK4tfiRR15
dWJLoQwGwM4bRmbbtVpzw18Bfh7/qzaO6nKQTfG1QSG/pAlz2j6WZ9T6rESsOkMyuFLpdWUzriyZ
LsU9bnwH8FrORP7CQvVf1qwOMiq00l1WlVaNMfO+Ia+UvGUWoCF4VXf41HGOBWLKviFwRIF4lpk6
mpn9+9CatP6X6ZBB06B61VUe46b9Hi3gv5fmjZM1Tdz2QD3y9aaqg55+QwTKML6nJlbufYln8Of0
nSscUyvHiOUaHkR5yeFTN4/k5jFNhpcprmCKApoQX+OFpSPimAKGV5j5vKEzc5zhez/PEZ3vJnP8
cfSmlCjyIpMpD618G0965hobwmBBftHN8+zYuzJXRbTtiJNO7rq+0Zxzl5JK4dHNlzRSsMtqZ3al
GrKNwUSyweIWELwLFmM2ToIvdLhgNSLyClhWIq/FaNeAxZMeAj34sYAmnuysIy1I560uX3ko+sRh
c/GDJsbEohfup1hJznyWGXFinRGYVdDCpS80HVfH8nQOO7sgh/hWZlSLmaw02CTKEhBjPq5ujL1j
C5db6LD67M5BX1HmhFZSeZuWdpU6SqD+x1VQiL47sgqhhHwJtZou4afOUnnFkhWbJBGStf0LET5N
6yuNWyX9vQAbQcl+11xfm1YRWwmP3gJluFuLtTO/uobU9A8ObOdQJcLGDdFk7gtsa3cXAqGgr8Wp
nJZ4I20RWQI1Kmto/5zxdGk/u91c0d+154ar0pl5jDvhB0wz0Vfwd4h0c2XD0FtDGOjkDjTmUPRb
JhKq+KMJs5lOCLTYZQ787hkyAWiItuA8VorCUGQ+3HMEfWYJWvzxNirlpHgwziFSNjvSLxgB/m90
Wm4uRm0FzZsdvLkF/1cGDj3+vlm86DRYL2h1BA/AGwDfMy366ycfb7cE0SQxI+zd3HURDlYL/DMA
T/yaTV+zFlwK2Wd+7slQYe4rxccln/ldTFv2dOIolwiu1xG84YJxatkKUYG36l4oqC4BcK7N3Vqy
+wfDSCpl78NvfUdwciu7V10wMoaQtioTVD9wf4d5bGMrq0W4f2H48kSxT80/1jGIrCAkT+SyI7SK
xi223mrrnArerbne2IJIQdggO1/165SGYivlwRXX5/zW/nZYKs9yxWlCZRUfhKhelcjA8Gn6jede
b/Yll/VhIvqGYbKA5nS4zYVpPn2S1xO/0UvPjfFAJ98a0c7tybss0q0DzHk2XyBmjiwjM6JGTkUM
8tQxPEAxcMsHEQUjem/wYy9c96e0/6Yp/yuJI3lpS+weofhZ8sibWLeRyf9CPHJPqsaJXFtzKcYv
nM0D2AsPbLsD7cICyWcuzUth01gOwKlg4hHcfYfWIfcw1lIQ9QBmrM8Tp9Gj4tDI+FuICIZmpjID
Lz/PMhCvqiZ/EnuKEw6vpLDrhvN2oHElp080FCzlgwIAEYkksoft42rMX3XBz9vL6jiUQ19nsGku
H74KwHa+61ugvfsu4hHkK6xhtXuQIABfsseNk9+rWC651M0jR61YEywKBD01IBZrS3S2DHwfXLjR
bMrehdldsS505kqUkUxbX7XMBh/tAoUtnA9a1TjG+ySiDA76py6bQdIDtCdAKMUryLWYHy1chKRq
3JfA3gW3+Wc8UPT4tZdlO5+oF8Esw6VdW83zKsL3OazW9Im8wDdKpfZdNiITO6wxRkJT7wxtHKsm
2ADlJYGWI001oKG+oA1QPpxxhyHRiedDnt+hh+MT2+l28W8iJYuB/BKx7BILp1cIK3HDNVa0Vlo2
dyt/w+R4Ltmbk8LCyJ1R8B50DAqYhIMJ19GDJ5pglCTq80VChnX5MvWJM7Kp5YLrxIcMlKHHdp7F
LuKGQgfoQH8inqLXitrgWckRCDJZ5GH9FRyYo9FQrPKhppCC+o+WLBzmewSp5j++RHVUrrhcf6T7
V5lTX+sLPfQk4wf2T915EKLZWmixevRJhA8YpkfMiMMcRpaB21PVmDUPzjXUnGFvbFB/uBCOoBhD
7oiedv57+FanSHOGkFAU9lEtgmADFmI/RVbIR6EigkWZl6x01SSn1ULbYtYi4VpJb++LtU8+4fpQ
EKzs2HKEWTh009YrFl1yLlFJFdVt9GnxRWI5fx7D35TlLuR3LUzYBl00DGRRNikx2DQPqWtAflEK
5omA3c/iipWC/iLAqNoSxJG8cabV5On/DBhIvdL+KErczuqtsbrbaWMac9FVLzPZLgp0Z1hpHudz
RnJWQ/BvLEkyBE9GELV8V9ovQCnIYh9iHqTMJ4Xsp1nyKWYGprbMDO6M8/miot+jOF6S1OypdQll
B+08htcNK2R3lAhV+zehZDDQVmTee0firX9cJrcZRSd+QOJf0EhBBaDJKA5oYlyMvz58JzFYwSYS
VNA4KDlr/5p85UZi6VbLAmsIe8WfuxxZd90E7znIFL+LnKGJM6rb+IL0oqrC0IJ1pW4gt4rMThuC
B1CE5jwDxK6OA0v+8kr+vcvp2J1TTK1YyEIAtRGTiS9dKy0aLEAWfW9X0/urOU3eAwm+E55PpWQr
XT7ztsRpWLu74H5gfs6CFhyTaB8kPf4gjzU2hkuznzs4t3PV0IUNWz3qRQrFHF+RyDXwnBvyKdMX
pT+4joUl6zfGk78K7HkR+fUu6QMFZkSP6NRmcu9aB4hlmL6+LI548aFLHqizNHnKR82h6J9JUvEe
MFpLtCIAQvbmY6ZWkHjV7JDzrLYEVnsdhou77MPUC3+x/SU+M1bmRRZyJio7C0VBh4dQdlblMerG
LGiyMKtwmrYZaWvEp4jqEFfMbyeUz8s7y5rlHZsJZMRRrfN0O7MCOFFJHNlpUv9gJavtqB/x7cfx
7ruJcXXjh0aDBgP0MmtgUrkRUwuNjV9pQjRvDxn8PNwjmEJZW1+Ql+w4w2JC+rtLcIMdcVzHS6sz
DPNqaIx1RAspqhozskwhguZgB93pS6u7slBDmmtd5V0UYsaSZI9QjyuduVzZmvBNt+6CxHXfrscP
K2x+Nm2SSmIltvZTocTpoEEFs2g3hVatWBSFfKnMdBjjvvyvJc4yrlKHKsLYe8oik/GCK6M2noAF
DjT9O1aa177hqP1OND6YYk3AZme1Cgwmze+2u5sYU9Wp8ibWp42xhgviPCq2p6cFutHZv2L4tsa7
cbwMvj7IT1LUkIHQFqRac+miGk6HrLNAj30YfeNeH5D4PGGH2oxz1XB9QNPFWzfgishaBVyNjPAS
oeZh3sC+VO73MzAyZ+8itxywXA5qjIA5lkLocSMpOK0e8YdsFxm1FJE2ci4VhbbtB5gCDvI3mxdS
AD5uzkxZPgY/NqwubncxgOxmAJ6iZepRMRYYoyBbY6YXA0HuVRgeCdXuMUggwENNahELCp965JnN
IGI1pCMbSet50oUO8au7g7J1oNt+FmkWXifPTDEuleU7XYPD5Jikd2MaG7Io+v5y4llud+5XWxQh
7CnioRd4MBsFskQeqpXAT5OaWcE0qnu6Eghg+pbq1LtzhZlkEWlNfbNGu+iqYUgd/kZ2rNySgKwk
M00RnYRm5lQbyOwMljACi12CAVB/PnWeKM2epILC7rtvX/tYoraqPr8buZevw0Z5x2VnQ3F3PgbI
zL1ZMSux9T49y5V7WzEzu8Cg2A0EeDhXjp+wLoMGt2p7EgdC8FKv71eIxvzuBnjtV3o3Vpy0NjS4
o6o30G0Px+vQRKHBIsJD8bdIJLUymXO/vLMBU5JyuTpspvr06JSmDTmL8/8gt9NV/ALnG9EDdLhd
UoqSLgEdkfuYBe5WSZyEZvVzScOIvR38s0OVoNwsYEGuQt99u6n1yYDS2oNkBYvCpZpdcSGqVtc9
0nil88/CuJ/ggw7OXzBQFkx/Z4ANymEVlKfmSHbuXDlwCIxahm0UJeLL9Cv2Ck58LfGB83Kgsmx+
VVkRAsg0wDAAspdzo6kjx4SXbH9taoflg2h2UhTcewruuIMOrp2KPzZZT/mJ5aAR1TqMreoQvoH1
X8mgywbWCY2xKG+5LkUfB4feJawDMjaffloO5G4n4RDHkSnvuEtJ1GAfhsurAcV1hBDVBp/Kq8RM
evPHNAY0QwK5EW02U7W6byl2l7HKbos4xaFxChwQDX6cFIfonNpDjl4QM2HRp0xNTCXmq+zEgwlz
FgwUbXBIJq7Ad3WCWuUNF3/DhUB8qidEtFZfN14LGbbipv9DwgXK6aaSEG8gyg5Rjm9V57bMViol
QXWFE0sAwFd3OQx8ZniF+ySdc+okYxPH/mHlmxnCmBBgSbQfsYiRCoPH/zI9aKC3F7DXRiGgc7Zm
tKcpobq+UyJE6CO60YiJs4QEvJq+25zEGTPQBsOWdR4tQvQ+5waec9SmoDNZcaLL+ke2XJpt/Zd/
mGb2eciI6C3YZjPYEe2HlnKM8DB5538Nu+7+GH4erd7Ie4MccSP+Z/JWTMN2lHhu7fbEwLJSKm8H
XopUjnNcdJ5nXGIiAVK9lEMmWuqq3t0nsttjwBpU2B7rFaXbzJrudSqRnFOS9uMugT1qmJaWQ80g
DE4u4/3wIdZf9sMxeIUxBxn0PsqauJAaHFn3ywbvuMiAVNFcR82fKRcbkGaJbTdw+/myXs0HYUyt
8Z8ta8ObXtmMhetaQUDNnTDJJCCdNJv4m8iyLfUPqPUiUdD1ZPxAbvn/T5vEQY4Nped+K9UM0H6X
pV73EiSChOSewOTO/aW9TtcbP8J2vFC5FPIK5T4CaAs3jdfETWQFUObk99gipjYqCLNriaf2l7o5
Shw399zlS+Sti5V/SkJHNvbc6MFUrbbsb9m0CrYMCouyC2l92EpEBS87rje37k3Spny+YWjq6D4P
/5/JdYYL6ej7sjY20lJ0je8gRgFJf9gOgqg2Rc6CQgO3yoicIijQL4NES3pHh40yL/vsfRi0gMfh
ybHQPUHMGNlEcrE1GQGW6UxYztealJwbJ+zelBY8Rum1WYBc9qkxZILYYrMnU282mEONRLgLCnDC
U4nG8T/cCC591LQe0YZBc/DUXrx09G+jOba1flC+07EnRhDWnP/FQ0thU/zQOoYLEDljobagLO5s
hd5JE3BBXtmR6ESr2busc4U8RBzXFDVC9obnxdbSpSWG9faH9HfcS+icuAvGvnuLnDg+2WLwRwdu
4/toQ8zp0rxT88yrV4RuAQmi9B0aT4x/7ZntVJw2azSA9rReY1IAV+/1VW6YhfHDt7VA9sV8WBOH
UqhyQruPjcQ385kpD7fHplPen3AkYw2Uv/lwn7YfAo/hVyFZ4VN3EVqv0HGD1uhCOhqEZEUE5Qko
xE9alf4kYjduwPL528C85FYTuzzVb7ebL+iTSvWcceArUWukW0r4lHBDlmKSexBX8Xq/+3XoIz8l
20sLYf0y51SOCcBLYCVH8SIveKeMkfys/uwTgc07/hK8FSxGSvCMwp6lmSDMASwkgL7KLrnok2Rl
A7rgzavv7OVuJjvyBCS93mLlo7qIcMPoqELY6KxdGfGXQIRclSox4jMrAitNfuyGjaWh72/wAWks
itsO1UHjxC3pW88cNgh7PcxUlnkZg1tAaf+RiEnuFdPUJ1uo7EGtQw4PdC4NtULegs6o28FNp/d7
v9VXWcbzNIicGd/5YAYARgBCQz7ODmYS/MYKDm42iPWmLkPue1qMgE/VIJSKNtoJcFMcYQg/myCt
LQPC/q2TRhboDjhygWX407CKaQ1HvT30w0vUDFKRxkh4UVAnDCt9ZQRarfg95f+8KfKuj3j4twYc
5b9nK+nJZ/0f4g9xsGulvXDrLdbrv2j274aMvvkoFFZFVQVAHqkTia7ZJYhwP9k5Aw4XVh3Xxinx
Nzl4vBDm9FoB3jheqY8CM959YFq3xVjyhh4MSnY4iPc7yD8P+SJf/WNUiXCoiFv7cZ+6/hnjLAlN
oR/rNugnhsuH8DzqZluqQq4NpvBmb/gXXsVNO9uzTu6WNRayhAmSMKs/w97Iupta09Ajk/1bRYA0
4kF8nzDibK56oHA8pkBg2le/fge+geEOEIaGDldl3i+DOibrvETI7lwsxMna5qymPtnxT7Rulg1e
JtLGfwM9uuyifyZ+vFHfA0/b08AsHffcvMAY9Lc6fbBbF8LJ9DnEmBNjLEkbz8pB61L4K3iCQXiN
LZbn0aKKFYrfu2UiABFmUP1FJrewCUc1FGR0A+pduIYlh6okqj+Hzw+4Spms/pF62LMzOx02YuSb
GA13xdVUYlp7Kj26UJUe+AErxC3cp1M2TvPYVvdAcO20ZbjMKCO9qCTZZp2KyKjeoaLsRBgttyFE
cE6kVyUE3WqOjXYk6mhr0WT+uA5tj7DnV28Kp3vcZgCttZQrYV3s2/b4tuTmRWnk70xkQxfuKTru
r/9k0Rja2tO8vp5IFRURTu7HJZYtGljNeOKrGbs8gszvGeyE2xkQG4MF9L+kIZIiqbNvgtPbC1eu
WD/muM52ZMeO927iHclegrFC3Z94aDyLQuBuYD67nFpcmdQWlyrXQrvO7as4nIHCy8O/BuZ2vJh4
AwMHIvniFy0Tjcb1t0Nd807Z9Mb5dtLai5Mwqw2md+5AmqVhHcHVeJ1Nctp3JECQthZaKT9Ew9tT
PdRKN0I4GUPlHi+mGEz5c9sbtEYLV53m86tTzskSPXaG9HMmNYZ6BNm34wpfwhtXrNxi9vmOHnT3
3kkIUhAcs6t5Ls55/tmMDU7wXpyExnjvkM4meg+Xgu0j2gNnH9xb2T/P5WNH4RBYNaPhE1wkGfij
RV/5j8FULkdx0KipjZdoykM8HpECnasYLZ0/Rq6SgYhFT/O/38lXKcs+XfbwKaCiVyKFf10PPbvW
OMYztfR4co1tXraqcRe6ppuV/dpZxOuIvmrhlT8GA82wamf0Q419Q1aounu2ImnATVASsSmtVXmR
OI6CX9KG81r88Y35U9quJyRmzlpP0OBuC/+OxbcBjfJi9QFfQyOhxbn/C9PYMHfYyRFef04DQUPM
/KMTKBMf1uPFN6B2xeqFe7gLKEu2eeYSExydl9f6NGTUfDe3JDpZRYVu3MIp6uTfic858hsx8F5L
x0jef3sOfCeqELiRfjJS5kEa9VS5/hKqWQio2yBZ93zwooPWdh54MWLcaMHIEs89mFSDH801bpmq
c/UfTZx1SbCZwflvLlBT66WYE6MFhnym35I2pvo4VoL2SE6fNo+NndJO60vRHJSdCQdU17Nk1jcs
db1B4rq6vpHR/9wZJ6I9KYLtnUDaWoeQuBTxDcyuCTWmS9+YQNATzR5k24vn+TdsSwH/+di2k9ix
wdqrr1X0QogeKZPRfV37dUX4HgQZ66PTa1S3TWSJq5F//WkY4cyPyL5cr4MGhNu+DHgFFO+56ftb
o074tgkGpxFzDiXVLFeb6lkhm6iegoshpiWPNFEReYAlGxkHhcD4yQ/ipgCfcJC06ybnWkJ7Vtdl
ZG8VDVrpqqZZWKlImx1P1ROGuVBpqw9B3OYluMr4rCyVrcIAc1YKA8NQubcb0vhFkR1XVLt862UE
NdTuBISUEfR+HY0I6pCFGLK0yKwPY5PZMVRUghz72WkPCZ3CtACvUcfNGYzG7oIr2p/+OnlDg1zj
GSrWcLPWAkvhJxAZjGd7Q8grIMaWFAcoaMbz+dbq8/1oft0LJ+PlNPV8h1tWOwDuuzoTgRMTP6N+
O5WJGfsXOKrWnt/9+fz86tjJrXFPXfhUPuu+iO37Ha1fAtkLm+6RJWTcooCfrkI9StmsUVkh1mUO
D0NoiNwmI0NF9kHCh021axVOySM0PCLwK22sJI4syVv2gbobdpTk3K7MteDZqrFlfTyN7zlOR0ZU
A9J8hpKHPSTX9qDX80/fO67kjj/B8fR9p9UzZArcQG80AWp1LirwwyDv7bdd/gz2B4lnUMTRjX87
powBeXcHabIQQ8a7an1MnDWEO9tDI7qQSWD2cp6r7xWfnacdYyxPyG1HdMyad9RR5pKUwHQ9KzPd
uaFTtORlhzdT1+0oB4sfVPoG4oX3os+O5Wk/qgHuoZymYOeQwhJIi/Vnzhfdh6zdVc30Iu6LZdAP
PRdPmF9JXkPO6dVUyFNZmSowJsq8GopwhFtEQZTfAnIrjbo2hNCmGlM/duKsGMTPenfmrtdzNHj3
Hip4Ql0nuB6m+e2TTNBsKj1ZbH7UDr9R2ZOjRLwxPArDbOG4S3dCwhXpQLjNtsK2yzRQmr63gvjA
YfkXgomuemzoiFmierPeMOBr/7DObnZKxiJh7G59wfhxdvROF8hhf5wc5kiodqFN6RCpIrT0tN1H
hVXQi0t1c51C1rHLrqalE+HEh8sJi8LY6+V6XTvOCa3cEBQRwPdPoS+z6b/mLHTDnXf+7Vkh8VaD
Rf2h76aHAElrP3lywXYKk8QbFsFGX9Dpi7ZZqpyjxWWWe59yRZaB7MVtkUMMydM365xFsoOZ1JQL
tqoU2pheeEIzF+2KXjvzUntx/xIZwP4f7jlTN+AmCkgeVc/agbpK1ssxqICeS+AV6boojALwJ+30
4and2dyhFkVUSTnMdLCm3yiCsRjE5tJ7kXyO7lz0WCYEYoTJAQUIG7r0Bi5arh4fGlnt7dbw5ty8
XDIzH7p/FCjZmEPgQakzWsse29pD/8VIwwnOydLvW5fV65XfiTTMNdUFDpfdgNf1xQaMhmmRh6SP
IOB5QmtkMkmwXqSNTcKkcQGNI7tuFz/4o3CzwzyvJ7oCq+H8dhzAkoA2qda+KM265BNE8kAlRJuf
qxXOiwd0JRcsjfu+3Ci7s0ROtLC990B7NqdobPViOzb3N0euhGEF8M1O514tABoLVDZjWDaokIT3
XanJK7l9by1ZjGggPdGpi/U10emOCs0KH828fYtMjEKr0QASG1Ph0w26qExrGDo6YotkXLOQA9wk
Clf8wfHwwNSThKqP7TFEaL9t86laGvHyf6cuRPsK3HmEz09PuR2of9M2vxre7mmJW5MED+vZgWRv
oP+Xxtq8IennjjrFjPhKp6R/1dHHw2yOropqqPIT5B/p8OCaTTtPwzHiRKOSWXSL0xZNEViw5PyJ
iOWAD2BksM9DHTX0s4sAUUXeW1ygmGM9lWJe3FUDMRi19R1/Yi8fN3GVt3Luj4ET7mPsSDWOhqMU
VdpDrWZPO1xYyEdfwD3L03CAzljnkPkOo79fbxGuuyPHmMoolXFORYygzTKfLCvXZA3m2kdutccG
nyogt+Jl+HPvW/Y6091KQryM78BASCQUoVh2yF0PduC6L0B9q/OWBYpTbO6qqBManD7+X7L5C6sk
IJWMxk4h+bJzkmhzu+BhokfdBU2hy1gbs5ObdkZLfpuZNBJlq9ssl3EydeX+3bCFSnuO2KLDrHRQ
v/dv+lxJyGJ0YoPeo1p2ND8VmAhvy3fH7hbvae7cQQ/wgftIIU/S/bVrsepvvnVGIU3PcUXIMQbM
GYMPqu0JnHnmeYteEXe+cNe7KQ1YacEvMO01Rcc9qKbLyFzn0nP80TOJVSqSCmB5eaIKJBf9+dmb
6SDWU8wdWyRIWpNVQdvCXxSQSRdpOTV1UD4jssLE7brLnHLIkSfjQAVGfQgc9xS+wytla8gxtfCa
MVkASXT2inc02VfaAe0QiGzKZJb/fgFDJDINYj9mzph7VexFOvEyvmaW5j+iA+CATJu5FvIwu+QG
jhh2K11gHSf4xcd3AMHrQ6NSw2HgDjSsQ7J9oh0bKKN2hV1c1r1VrEYn30eIeh5eimI42VAXWu+c
1pAnib1tBRSwsDxnCmEBMA9MpD74rFefoTtjfcIeEwqkRIpWPPXGsLiHWL6rDggyLAfJE7zjp0Ez
B50ll2OkrCxa+HMJg89werLdhHLWf7ORG4Et814SVmq0iAmkeK7D2vL4iakz9Xce19De76uwkBCf
MgTs83eOjezej+r7D9o/IN6N4tKSem2wr65j8hUmEmjTIrXeNgsPKsTESQw+sQNCiEFc/ZvsXx/N
KJz1wL7hZNw108JYP/QxV6uKt6cSHTg8Ceo5f0aD3jJf8P37z/cgzd5SlXNxi9FJaeQlMDShBVVB
jsxc2p7gIcNKC8SCh/RaVdivjXfqd7b+GVYaUNEJCaRGQ2RgPUYBgnEUXixSu9tbDYGcxJfKewIv
7aIba8mhsPMwUTWLxweMmt1CrHqBfz5FpyHddqg/YGsrQZkK1RlLcRx4Bg61Y2P0yz3qNu7JxIi3
w55CkbkYUff5pl6KJVtKkel04pEZYewXFJ/muooCcphMH/vZSnWQy7/agXu7pflN5pGDPjGkWj6T
nv0amlvOBiLsp2hlsmGmCOmc/QF2tECqWxvu6sIovWiDrLTuoQl10VKlTAd1lLIbWlOI34O5oKTE
3DWr+3pbnPu0WK6kZ2HXosVF+mjmQrg3vCwVJQ+fG7Gzc93rSJwAdVKrHBdB2BAuIfWlF+sHRX+x
wlScxlpx1XKef0cdvbPoI+EMAJx+irV/jP4VkYeTl+QSB2DMj54e5XLH+TvW9Pzt1KyJmUan7Dxa
48sL8MiU+I7vYVKBFwLNVTuJLFxQ+XOwnqZql6wVJcaF4BWmJdqCj6x0rAk/ootU4QarXigVHBqT
OIzeP0vtw7j8EgIteTHa1VXn1HDTod/yEaZA/bQ1sHBnpvgacecUhOrWd0csi4MBGLPodwHFaob5
5QD9CEiqBOdJtqgaCFelxfKg3Li63ywiGTUYC+pXJj+7G7ALKXYHRHEzVAcle4kJvF7U4gc2cDAg
q7DV+yMOMUCMHGe0qOIomIxYIpS1t2EAl3sfQUS3WcnFaSRsAm4SUJhVLn+JwO/ilBnRXgZ/dQDo
y9N45/2HbbAoYEt9rY2Q4pQvgxckfKtUpuMOV8x3Mr0ew+Zq2nDlXlGaxLiKaTQNL2K9E3Cb3zne
OHRAJqQON5X5er2irZJZk0QLlEqxEWwLynmv0MkUnHUVFEbnaM04drFqfATnT6iqI+rQS9/KOcqX
nixrqNz+b/ySfMPmw22gIA80Tpo8dVKmtNoMs9bhUlp9Co20xyE1T/gAgbDOwVENGFn8e1pAaXtR
+IYvay8KqjiKDkAysjCC20Qra9rG2Pk/pYnW0A2Mu2zCQ9mnakLlQnViO7s8zVQeoPgMipDP+fLd
IPk4CxN6/MJeQ4Z+VEz//q6qVad+CqBZHroclRIHzLeEbfX8G8rQQCdsLDDF/lZBqWmTPCzV6dus
36en1gHJk6tAMe8Ah854NMgpLaBXd556pCpZO++tZxv6gfLfNoA+/hx6MkTELLHwAEhhSA8xXr8x
xhMtCfa+BGWklDs5li25qkFgF5fVdp+Y+wFJUTFhRcNvjZp/y5T3NPcnxpB3acsns/M5XepO2d4l
5vv6m3Xp5/CuI6li3bcQ186jjgOlLqK1SwogpDJNMdjddu7bthuA6x5+I8oVWpeQbt7JbCF0eiqL
pdvJP6CqpZHAAtgKqagXOSA093R0kE8iIjeBhuKzpyRnp/IL9EFgSBhlucxSLTTZKxnd5sxBgpLv
kckWXHwW/wbQ5eIF8kedrcU7zJprZuszTF7vrorRrCmy0RW1wEpNZcUo5JGEQXe5uj/ibpBj2H/x
KXzMw5T98sMlvFjFfZDn3azsutILeusPXhi8vUB3gV7JbcKUYll3jNc5aHpXQ4fvrGKkQvdPBM+d
8FticKPis5/Qt6XxGUpa9DnboQSryuFHg3rEzR2iNyHI7cjYwMRVfR5M3gdNf29dTRZXTKbWAHh6
0ixQqTwxXhn6d6SNcN/S9OzqujdTWr4PXV3SYu9eVKwRr+FEGvUwQFO5y0+D0Kp6wh/Qh7Loxsd8
G3N0Ly0MkmtLL67gH46B0sR1iqhupu3nG3iSJspY1l5YOO4W+mcCC8/HhGOJqZ1LM6BnPI1q6FhA
MUx1pIzxgMlPb/79MVGissUP5izDFXl57BXPIkQaUgtdYu0JXsDlYAIKADJHoPIMIUM7Mo+GDB6e
rKC2XB7omA3B9fkaIiLIFifUpWARsVIeXoR8OpOcFQBlq9U8KJPaGoM/k702vgXOXJo5u5kmM6/U
4pzz+ZEX/7p9lCpa4UGsodCeiKmd4W7IYBltqkGSU7oCql+S1i3qqQN59ySXyZZJj9j+/W07fSl5
tXMD0qJv16EZK87H8FB9OPj7eRd7HiXBLAlROYof4D9idBivgfzky6uLu747oT8DjGPSN0WgMCxF
VD++j407YLHXRhyVWyDb7JC3FibfnizFTZG/0AInieclkKnPdbDbaUQiGtR40HvPMdHDHSZanGHb
8UG4lkMk5U0cTarL6hDAA7attzudPf6nVJRjtXEn8P90AMrTGZyoyVsCYzJQ4MOoeLI/I/wiDNlT
Bp3mag5imhIGeeTHH29vwskK2kAFGYW+3ONioJyEIyxDUGL13kd/Ih/auh0uV1VAAVXA7xOV4MYW
5O18IKmIIFjfuo1klcnKmOVNcAjw3dmK3FDVfCcfM5pT07j7BCqCifd7Swlzjm8GdD9rbNoAEMoW
AHT30tjQ4xt90Vh+GgeiZEi5ETTibGCjH72FvY8vPBTaRxcNi91lT8mjnlp89JnddAF5ETzhGwBW
mUSFOM3GCPTtD/z/7esWM+FghOJOUegDNylAE+ab0sunY4e8c+1YtbTCIGgC1PUXDvXgDaH+g5Ff
uH8zT+mhCvzKmItlG+B/RgHo3MwVy9aCv9O2BiycJDdccC3Qo5VJgQjKwjiEquSAvysV7by7uzFT
G4Gv+/FYONYa0sSQFYGjwvxwjDagTpR72kq93P8uhi82bMVJAYN9tyzf1dPOGsh6AcYTLtRjyFKQ
Y08U9phfMDj1FmqN1HDiYbrNQkaTrhLisnx/HH0LfjjdkbleHR75DxjsExB6AeNTSwrPOTInzXki
LQCt0zO3L0h5TtXyNO0u3WnY0bD85QdZ+XhmWNDlZ+4uuTNjmIo43UFDc2Z66pgxxDnL1MAwsWp/
aTQiitN5PxJr4fwQbBxBruYwYGWJUo6SRca04P0yhSHUP/poDsUEecm7qcJqbFUJeHljWlNjKZDn
uZyGqLqENSwMtPHzwIozSUx3KGioDVP/ntNn0JsVjWc4hVMMEYVVDgyjbP095Yj5UV1lvcze4Jys
DBz+0sKjy29UnD03MEbZEfCE80AhPXZs1tXZ8hg8mqH5j4aWlQ+laHnzafH1iiQcBPucIYPNtjvQ
jiK7ZADpsD8ZIrtcgb9swLLWPnfLo0Co8VPeiEOXxHezwwp+p1GEc5UuVZ3UoM1+OcP9rBdK7De6
JNLrhXp2TR5pa9dKk/QvUdgnKP/6IeWs+GgfesqcW01q8Xqmucy9SnalL5gczwjtYvcmHQXhNFHa
qQ/8hLJ1Vp0JWiw8VQPky91D6bvY2heftZ19gF0PWwdxiJmZkrXFtyYBHreWeO0itLYMHQ6FF2K3
3a95u3EquwKy63aowLxPj9DPhmG4qwfelh8k8WQS4NBneqP2Q4AVR/lk/Kybf8sKuKlJ+nd284Sa
/yN4FcZFgmnSmzEv3Vy4LaxWEccbnEKrXLIxOepR2292WpcfsgTCgNDAXL1Kn5YTNP5gJM9gW2gW
oo4ccE82om2z6sAE59pnw9SAgqAD7LZivA6eOElnFXA1TYDYW+dhnIcYaO640H/hiquHDAKLTswz
H5Y5v6lOWB/zNhc02TZJi6k2URPOCDXlqAfs3Z5Oh/hUeIpJ10lbcMJEt+ZVPqryvaSehhfcFfMo
QqZw4ToB8THSlB2hLcdAT8CIZosvDerOeBfLSQBzAYH1TfJVLB2opIyQqHPrfOMBtdV8tlDrs2z/
aoRttkyw/eNO5S65ZXFI1HGwKI8VTUQcg0Be7WqOr25TacPdy8XEkdMsJW0ECuxgoCo+FrKDCaeu
zJe4ZcNU2Y9T/wnGHwsQVQA5aITk9TnyQeSveHkPF7DauN2wTE7Uor0tOKL3iRCV0/RbspTGZHub
4CAaP6A+m/tEKe7R60RJa/f50wvrdNzKkjQ5V6X+on0GJN0y7nzjFeP8HJu5XUbKxmvy+90owFZi
q3K4Pua9olGPmLarEQ7MCNtjY9X0h0V7Q8pj1hRoUTy9Iz5GcxInZgDDhZqWemMWuzOyFSa6p1xD
ilv+S+eR8x+/hcDQXFCbai/p3Jw7b77sknq3yOkz3tCX1zShWdjMx2r8hTCEFTlkG1y8DnfjCmt/
U3T3VB2tCdpZbVP5AJu3i7D4CmTLvNJ+lNOfTT/45TZukDGuYEhRWb0OvR6BubqQSJf3lxpfki7S
eEXuEaafWHaPPAJY/IVeyaZRz8YfF+2oNkpf1moV8gjBeRh8Gkm0DdoRPXbQtV4/TQzu/DVrApRG
Wk47/tXoDHhI1UwQ/SxrprHqX/wsN8CLK86dD8LaP0yZWFCnX1vqtB88DGSbx2eoffGkBmcUsafJ
YLI148ggnLRPDbXaO7Lw/VFxiUEQfE27SbnYGMXiIdw6aINzDQEdW/S+t/El3TnwfOePRrnWfVjy
5SnDQ+hGyNobXg6oFUiGKBomc1+6gibgm809NeKzPa16f1pREFSFXxMp0vxmekH6/S+TVrrzDAdO
ZZYpzTuLt8ILCmepVidp+eShAbWMhUESGtzlNPMP4FN707oG4l0ka2WmBKGjavVfSP1CIBuLBbXd
fj7Q/xIQPwKHvhgQ0K3HWaoLZbKWzz37wHLI3qQ4aIqEbd/apBF9vQrPfUszoIvL5YP1uo2wg3v/
FdS7srB9w4rtpSRVYsZ8fexRMmUEfuIAUQoCcrC+Fq7CVWKeiVNfSGF89qUxbW3K8SY1rpeSou2x
pkBIDZ9gTObDClnK5T7KLR7BVWQmpIAczGpXiUqn9ZrjS0rQtCLRXeYH1jKfKuZ4g8LZ3wecoEoZ
73otN6FpjMW2+hcmMYeKPKCv+zMeAwJuqmMPraPZdLEPbFJNH0E6Bqns7oiBnokbKZfOswoozGtY
XsDE2ZBB+sweCVmrs3J5GngAcvB48jvuHemvrHp0aRp6QHnGFlyPWnHPZlOrmMTiww7NoDJExRmf
RMQLygC4R87JCafbsJiPsVWzfXyMZiz0IJ9x+b8jTRRqNpwKazXqdqwsjMGcOneRf6q5Bz9L3m9m
Iv1PjZIZROZgTSkSxYtWF77SNIkwNaaYDMKSq06urOBOMQ06uNvSRJOYqIdMhHqNB4zwtHqt7Te4
d1rMZ4yBmsUzNrvFniQGjOKKdpst3FMiggxVItaynZgM46CWqy5hHQlJ8Rk0Be9SzDVO68mgMm7/
NHLUxj4i9k0CGQWZIxtWnkuFnITKRzLkshmbzwHCRWPxTd5rPa2jvoVburxhEhS43f+XtGtiQhbx
GjilfehR1fCz8rSabevBYMimK/g/j1pMYru64Pan0Q41LM+T2gU6rpdbf2pJH/5QdkDJBS2z1TqK
7FQ8rxYbo2NK0KG2ypz7iEvCD6Yi3IaWdK9wnN4yoCwfHpWwGgAmYDZJd91huf11Dn9vLAnO1asw
HcvdGaQyUvilccnT67cKqfTVsZEuXkSCEJ9yXWoxHyYzMkC7k1DAXLdTVzJCQj2kJQYma+eohVHx
cDeO1ONc7ytTtOAu8FEhYWq+0n4RQAmHNWLBQFseJhXrSiPsFJm0KbToH3CqUoGOhi4p2ijJdbUv
jjaz8HF3zlejWtTRZGPXe50Dvljjef7f9hEBVm3mlg01s0BU8KU7Lwuarwh6fp3thDD5g99z7WPL
rJzKEwTAcZYWbCxnRzAzzx7BPscg1Edn4S9xYApYDJySi4AVjmKofMs3paUPj8TCW/Cr+Sg9s4h2
P5Oa91+34pKeBW2Er9rSii3CPFoyl60RfNt1o2KWMrNE9xvlZAkyNpCX3Q3ivDdCv3KEvk72hXfj
MdVq9K08y7RMfc2UlIMEuD4vEVZldU0pkYxnM+XyTK9nl1UAsWkURDt1qZCouIRN3a/q5E9t02xu
W7vGZKK5DBbRFmcHezwQ7y54HjnNa/sUmDNcV6bpxCKbMQ3hlM/LEOrPAnWIxwseyMcF4G6XXPXc
/1WjeDUkXUDB47HThznPXzq3eKhuK8I0KrBGDEc5ixOMwJpB2F/skNOZOXkFP9ipRYTb7n9QxsV6
rkZPqhcVTH8ziFDLgMfE6h5dMS2UCbflOcmJjS8E41ior7OHEeWQcnpDYG2dwwUYLVyDLNAcsxU3
JpC5NXFWrm9FIXPZ9+ZUTJBOrmu4CfYuDY9swfRvlp/WbRwQ/HnyNyY/iwYnm6rMXaJnvnckh2Zd
SAjKsQMuJ37ZQM12cyW7/Czml2h7PbTy/2MRt0bRL77yRU+yKtp8fpkHbudKjUPHPxYXZXiQ+hy/
kI8tpY7GXOHA2Ognn3kpOK7z8jPdom5/TBhKfnnEcyXncVtWkKB1YzDkuH44FPhiFua3X9EwKy5O
II/GS134mfyazXU0azYlMZ9D0aAVzeiMI1+JbNIvXSP8vOAJfk9IjdxEWRTqVnXYUwOUzMiFVZPY
dvHhvuMXFUtKV1no106xDl12+jn1MJVL4GJNVRtI4xk4knn5pBPw4qNAXXoMI9+NJ2YRxT8Q/e/s
R0GsGTVvvOzf3vcUpYmcoOkIaHAQSTyArOlJ/r9XxFOi4egnf/uajO0t4fSMCFaNIIAP9VkFnXmb
PWykSCkO/ABymARxgZwTNxYH3trNgLI5al85rCjcXhrNP1ZrVFj2b0VBX348UW3VoMfBw4MS8VM5
9q2s2bekiO6bgHmKclRCQZmEs1yz1QNrJYyTW4jg/bIZBfgIocbVnUYWiYLzR0bAPTCdS8sjIw83
r4DLDAjmzX7YmhGcKEFJ+cSqw8vtVo/FvPfhdvF9yk3/RRRrEvXys+nT/FNeH/IWqtKKVUFynoAt
jD17Y1a52dORhFr+w6IrHFPClIJMvu1hD0DVka17cO6u3Qb3KKEC24WNyolv3o5H/dQULVLlW6ni
VELPwlFlmXEk4ejPTsaQJgguG95OxuW2Jf8KfbPigGa6Ir4EiA6AUjOTOT6IqV5lPQtbHUFZS2SZ
WZXsvO9NWzcK121JfSPyBs+DibyVNMB05HsiosDrAhaZEb7iimXUKbInO1Td1zfZ9YdcJbJzo2EO
3SzjaBA81Z9MF5kbQqfsstDc/VitFgIYyZVt+9bmkA+ABu4STCOETatoGvwlwdarYINLkotekT49
DZThi3Qymr1H76x/uHC7xtjnnxhmC31PNnMp6ZKXcMHyird/YCWRQ5M7UEHZhzK/VpvJN7EJWz26
V9Un1FgW4ZNXHWndiKr0GU9oxPnJsF057HOT3TT+xUbjefD7TO1lJp3pFILnK39DX5NIZSiWgQRp
6yUSOYhdnzOOMOUv6SC40d9lWPIf4yYZtt2CoOyZGr4g5sxPejisQHZ+WiFepavkIr5AySdAFfTo
/loUZtP2wabZJKqTiKKj0zzscUIhSvnS8gzWPf1xxYq0H5sWTHtikkKHJZFVlEOrRbsqzx+8Hupe
BP+cYeF339DZITo6JwXYyBM1mt9C43CaqutJYbBB5NhBea5hVHdrJAyjo/p2vgwqiqIcJTwTrhkM
sNY/3t83xHUCZk0G22O7bmJFeXIXXSRDFWaCI8c3DgkjPJ59yhSskNoP/HRszlYncLyUloM23JoV
DyL1DBUE7MTRNni1lqq+31rCgiKkeSS5Vf6Azvk8Yjo8AII5EN0nREVEQn3OLbc07EK4U8BNWNC0
6AT7PK9PdngK+YGFVY6rgNjy+4pHnMhXrxq1rydbB8is5S9ZDiuqdc63codfEpisoCs1qwi3tmla
wCBUfbNRAQ+thJOABxcYooBLVJA/2sEyctYhSr3xJCSGMzt88Z9ZcLoZ54wl5gFKVnAQp6Xgv68v
vvuxBbC/MqcwdoRu1NVzxa1p+icv3mk4uY64rN17ccfJKvZZ0ynDeaTvYX3cFAjpz6n+z54XSZ8O
wlXG7y/Z43UQVMCgQ8ILZf0v80IneX9f+J/WVfpzUClMP510tJqL8JSMPpSKQnj1sA+JqPMrlY9S
6WGTCM62bc0qJBAZdiQbv67E2wduK+y+uEC36/4zjgE+nzMUlPeVAqy8QHV4izbPP2j/vpuUil1e
YMZn2UTMS0VTGdf1O+jYStzAzQCweYea+tmid7nqlIDBsq740OqHV9iO54ZRfQvHyPQKmN8d2Cwt
3SS/7U/3VjiA1MKfywR5fUYX7qK3UoCJBDPeLDCMnn/rVw5LUg0pJR+8uoRMRb3AciGcU4HB+Zj7
i4yWR+AwuU/Zd6vn51ZHitoLWBxTToOg2kspCS9uU+8tcKHMsbM0+F+xZO4dYfpnnV+3sn2zpZIW
dH2UeAdxtEsKVu6P9F7PK1qotXmEik9EbWuRNpvOQORI+eJGipwohD0StuwMV/tGkogXNqOp0mJc
dX5cLhtY9CYPURC/cDbp9U/4WYtrIdESjnNJZnz6WzVBHu82jvSrJtEytANIKy22l37PmLzJFuWY
PrcbDM9ONZ4hWAumQ2dH9MXxO73Ha/zDP9wWIK1scx3gvUuRbNw2omZiLB5WFJcsBPaNbInAFn7/
kBOGUMxBxFBgx5y1n6F4rL0JnDR8+7llFuEEkcXAGJS+RnDZkEu+adz1DeVqji49stLxbp9QB7Yi
eKod8FeIb6v4woEYKGSUZy1FToEAqZ+/H9DTdCTogrfldzQOE98pi8gUN+JIfm/o6dGfI1SUU2b1
0886iv6YNSRSbcd9l22eeOE8ls4OxbjAGbSulZ8fJv6ZcRhOHpgM06GpH7Kly15LRzTYKTWCPN/e
WZUMgUdeNMlNqZghIR647CcDitqh1jjXidB1iiIwa0DKbo6ZoMpMwNfhZ6NU3ZYRF9gew/vwHwn3
H5USvTS+xq2ElxojNCFR1jRzEl7syA2uEIW6eS/jJbiVbcGLtq6S2jyb5sAXjRdB+Mzvw0SVeIm2
18mEXmzw3FZuioWVn6Ak5n9bmK/T3en4I7MNFBQOmEHRybfUMp1SQc0GEKjPXVcPSYthDY6LHSYf
Kj01T/AlYLSwF/rv2B9DXnYw94UqRuxTUi/aDqGoeHpdB2fRyGxxn9kj2cqN6uUrI2MlJ3qs90bd
KvcWst+eMifXVvnJbwQN4pshQojWZ6v52kzM/LubHJUDH1qf++YVMZ/F5LdH63tKHKitTMDBfWE6
0W/LVbHX4Vhr1hQd2aeOUFForOuaTd7KPVZCPEYMaydKAfatktxhxB5fgeTsVXXD+xTm8UkJqt05
j1IMjd4gDmAlgMddESf8za0feidTxl2f0aiwnZwo+XrVwCU/APjEmZ43/gSz3/x1PLM9iz4TlBCr
d2+/5DAWQyuSpgP4tnuTy9CZR58s8aFgLFJTIfG6rab0hCGqnK8p6P5mYkbFdz1yzPDC7gXVATBe
Wz0xR8SeSOxD+1Z7LlBkzc5wgNAtQztFMkDQu06GEU/yb/wwjHhunmcwaL8XBbkOHvWz0HVwwRLJ
IC8mlET3ICWnLz7f6seK14XBae99aV139I/N1pQZsIUjIRP3BUEn3zuGCIlZbvOEShofwXpOZs2g
3jKFso5AnQQ+546ovpa1DMqE9TSNBfXso7UDv0hxtskZNw5vQxbPLH1iQcz5kNhhe2uGXBlTCo+V
NFn2JXvjxeOUF8Nes/3zt6qDG8EqDpX2ZUqX0HJBFNsA9SzOCLVTPlKMjhSgyr9vVIj9Ez90xpLs
Jq/eoHA0a3UTulLKQV18Z4NrptyA0T5HhXyP8qF9kuTKLuYCMY/3CBzlWSANVS1HElyFcfdnH3Qd
kNzzSykpHsQL5s85u88JTDT2ltpepq/2Y4C+b2yB/YfLkofvlCWwKUNdnIXGq0pIQ1iqFov0CwTW
2zOtXQNnCfzgfOobjY3aGfVpNbjW3kzCesew0Rr4a0nicfwnHIShB5KyowluZfujso/z0HW4XgYP
PpllIdL/UPn1BLsxp21MY99dHBmmYTpoi+tM7LPA2nYtAGeF/l0OF7GztI/feSic4jN2T8EH6zZM
tFc11eXDUn9NgeJ1YmgkTi5VkU6CbKrM+9+1pBtJDQE3vefrTM3/9oYKfbhE8JnFz6+jb1rHNHh8
rTH+7H8U0um28FHYfkD7hZVIOWwTho2ugNmzDt08BjQlmL5bjqfQ2F/9rLLNOEMbzL68h3asdVb0
pW0hPmIryqjq4uM/xlc8t+FCIUf2Tl0v98Vf+4Zxmnrenhf2lwYMfCUAwm+9gZD7HyYGyE90/lPU
zniO7bCuQ8AMrXsv9TiRtEEFq05sgnWWgHeX8QV7jTvgIxK+F5y61t4RwYzLXixwpAmNR1yV/pNT
9RfzPc0mXvYLNxsQfRu1iGPU3glPZgj032xTJkmwErzU30MIbj1WneGBSGqk5G4c+Ijr9mtkI1O0
AnGbQCTNbJYV2xZTOVa3M8nnFAsOX50RRxwXp++/+0w7yPmS62zUus5y03dM3/jhGb1T+8NLHK1w
GTSaWzPyU/ty1UrrHTD9/oNJZYVgOcxuzzPo0ddNqqL6eWHSRxjB+7TBnOolQ55OMXKQlN1uRQ5N
Wbnsq/cwyKKkeMceQSllFdmsEiMSCiJrMSIjFnE/DdEOZJGeH9P/eUtRHpNlkLwt/msRqbPiQkJa
r9u9NV0g5LnRzQfPJxENlp/CPs7lFwS4wV9uM7uS3iwX5W579t6maXoBaEU3JMNSbcNHs6rbKABG
Vii7OeIhB3vgd65xeKc1Kr0peWc/YaXpVJV/tzTDjygKIfoSktNFoyF9GNk6996Drl4d703ltJXM
JFB0myTK6uTRkfPMUh4qI93P7tcLf1JLGuzPZx8UpFLfypWqhXBFDfgjbICpvPhWfPwCfCR4hEvy
PNMRpdLcQLpruD5q4IGa6nwV6V827fe6gY+Y4jUWjmC5IlqQIgLVc3IoSLskiVxF15/EqCew37tA
SqvZFheN5Jhq7cGs32sBevCqT56YbrZmOkOudtX/cPVuQJ+Ps6EhGBh+9nHrgBoBRvyQ/Bw0jja2
d3xIhYwbwRqjEkmZMSUHZjSuybbsn8fIpsjzzCLHOvq9XFgN3etu/buqWfucXuIu851FS2rsxn8l
zDC0qdGOJI8L6ZaqYRrrFR8vLZ6TngGdgnXqak339sglvGeGpnAjmy6buvBTWs/YBoRpzs3gEVGA
lzBAX4liIdmqkswPDWno5jG5cIq+YsyIdrAtOB3OIRNgVh5nNhzfDBi1cDJKk4pP767Y3TIDuG8s
XDC3yc74XLK9y4vm3U7TjM1zQ2JZUPIf2AyjLZ5oi7jFhOod9MHiiZLAZJuRql0gt8PKrSwFrGse
HE+OxrqWr58Si1Tgo5Ne+NYWyQ8zrwvTJYzIsC1BmRcAZQ7omTKdA3sllPK6+d1umnc/cblF6Dvy
zULBsiydqinevOhhBVU/8fuKdUwQCa2IQ9KDKKJoqB+gjeBkk9/2mLPz7yDdkWjA31JwRTsx1YHC
cN4TnOqP6+qKNrZBU6rpdRFT0oS90G+3xOjiGCPQGjsn7OZuxwH+N+blkWLf6u8wy7PA0F3BJxxK
Z2siAOmlqBmBrcyMJb2vh8qJNAF4YtoXCjb7MrCaZbUxbi/crmk4Ze3mk1lk/SdD1XPAnxnRuPP0
zP2V/IPtPHuOPSPARfsM/vTR5Z8gU1tqfJD3N5eLF/ELl9BI0ipO8u3TiakF1B78yDsMCW6XoHGH
e4Oq2aIu5S/2kw9aY1uqS7jYAIs9679TkswSNDUlekwXoe0BRaNXeC49CI0DKDBlJ/7iyrO9vxzG
T1uG1pczj7AKinPNUUjtH7O6IynLBkXkb7xsTTsqTtOuRyLP/HAOZ6bGkmu/uPt1JvvmDxJSG3qJ
DJ+HjKowSen+Oy5jxVXlFbb58+LOBtmcXH9/3bodwca/luN21/kwYAw8kVAYpCAwEILAxMKIGNN3
8Ne51ukafcv6V9cwJzzPwZwICZEDEmDpA3Jjg6fdOLEyKWBFMf4PDIQMVBazjLbtHpmQ74DalPov
v/wOVjLVUNtnyxEyfBuFVBBO+ZzHb/ksTAQFBay/19iqrVSdXLsnEFpjSKdY+XWx6MKhCLuasQKs
vw1aPZpvSyTOuWizSznmhuRZOK2jLXPDzuS0Y46P5PpLqsOA6bKc92udbiqec+/q1sFbFf1C9UDE
CHalKvJCF7eX3KYUILWEeI+9sDlB2MInTznYvoJ/DgWTWOEjsbK6MM5+ecHmlWILDKAxWVCWgOXO
XluobFGD5yevFbudTBhZx7q64DOwRaiRXMXY1r0H9h7I55ZXt29+eyZnNe3Pc6LMcCDbovp7cZAO
IEhd0N3HxoGAdcnILySD7gl7RkrqOWVQ2hibUp22o/OeEzUphghVkZsuH2vTLCXku3sSbnSugPlG
JqjyDx2bHnsun1fw8q0yVAimoWBm0sk8mfUBZgG2f0Xh72MM0/dNWZt9EirDG99lr+dhtQCCtD/H
QdxzJW017Ybggi9uFJH8UmooGvkE55HdMToGlYR4QoCJLIXTvc3yDPjznOzjql4tj5rEXgPhTTio
UOB9TO7KGo74bK2QP1Agq1xXK28rNwJCpAZtnZ7UaRw88XN9oCBdsa7psKzIQxbslYE4aJnErVAg
sa386bcMuDrkiVdtDlrhbF0GH7x+bRbMMLetqufk8rvJxwXEGRmjVq7IJM6QjOASxiZull14xugb
BkvJBgx0tPhnvr57sfVTkadtzjlHWFJvTPW993EjOoKKnGsHlX8nKoiP18LtfMm9U59JK0GKzDnL
O70zS1Xd5YY9g9tS2BfHHdtxX3JQOcDp9c2N6lvpvlmODNI9wakQNsoX6XEtV6ZOtMtmd+/WT8kx
GEnpL7V0T6iTM7mm9ECjSQB/xSsLtfT8OCPasgsfN8B4sImLCAG9GpPWlP0y6wVmFiAlzr9shAQv
Ytq7lJ7QZfjaCkhmMnwlFgom2q0VePw02SdXTmTI7/WnPcx7xJp6pToyz/nBRZNURQ/thcspEv5H
Jwi1LLCnPhhecQuhmKmvCMJ/oITiPe+MKWNal23e7T//j2bmG44+waVdh82L2FjUu9+pHK9nkWve
Vl9VGFT0TvCVWlxd/FwZEBjMoiyK+kstgfH7jEnKVO4f6JuKKWbUOoRdeQ/+OOq0HP3xNXGkN8TQ
KTwQ+0jK2XhxLCebyWfl0uIFy+vxRi9Ty7jrNuEN7Q2WKQCCeeKSn9yG5idqjDftU9eBjgZhZ1CO
+50OFawPMht7mYzSLxFWejGIedsIMDnbHN1ExftGH0ULyz7sCsZY81ePBCVW67Z8rXD6ijAm1Sa4
zKyNiADH1gThuMBa3jkWvYADyxF2mIvUG+hJHGs+odC/yPihoTZotPuXxPxbc4SY5gC45u/jYZlP
konJ3MyHT1EtiZnl87Z7oW17CUKHzCP1A745KsERE9hffTnvru6oaFmHTijL/0j0S1pyqJxT/CM8
/pJwNxgKslfLxc+5KkQAje0lXA5v9hqbkNvVnDqjZW6JwlaCpOeFqFbQncxNw3PA5PhyBrLrMlVo
jYj3BiPTe7rS1HpC+Cy10Dd/oUXr+NbOY9RFVkZhh9U+8ji5YxE8EeBnHWkhgKShg5GGuLAiZJq/
dZ/TUJMuySmygdIkgrEPSLzAtDxR93DuECUVF5pM1Z8c8o9aRyK6P6ChL6w8VIsnD8UpC2px35TQ
hBvjbSLGB+7T5iP7IbnTPK2SHn/J3dxuuCe5tnOpIdSj86LKo3SzgGbrxAilRK7gSxwFphv54dwG
mOMya4WGwnYzk+H4iQpCMdxinf4Grm7TIrTnx7XCoeIMtEgSHkcNHJ6kEEDtoB4nuvO+7UZsqfNc
nQP5LX9eRqb5XjohwqzgDcT2uCdqjSeQh7R6//d1tWetTcmQEK2WRl9X1Ot1cJjNx1bItefpPOIB
QXid+0vKXxG5B1l3HoK0Rt1j3OYo7XC/SBKiDQb2jCC6CgFLJM5gM7fC1RL5AyeoqbCv782zCNsI
1T8wOH+aGCl8NJ5d4rKkYfxcXUpTZUdUT2tLgdR9Oy4ixDQCamVQaElf5XCvLt28W6j0HgKX3Ipb
/FH5WPvUK30sncFxfEwGSW4dOUP9pk9R0njlgfI3vKd3RvEnnFkwSIm9MJp6fcNP+s6QMNEI/36v
B1Y//zgldPmsaejB8ZXKwondttaUG/M8U81FUKWCt1H6YBeCSawRUkSfxA2Q4V09UPL7ApK2JLyk
gshntoC+K02m+jzbd2vuiQNPKQ+y1QFFdPHvvRoxNs5lhA5pOPwFGUcphZbIEvv3OpAhXxmU0B5r
F5SaO3C5ukCaq67Pf22DkqdqqhFU4g+S1q3lsr7FXUglLNqdYd0Po73RPXUuftPBoSvUmK5pOtG9
ztSTV2qXY9fp3jDAa8ZG+LYOoGsZOEiMAY7kea5Pu3pE+D/o/nNNq5AOuS5bL87EBFy1Pp4e2DLv
qo6Da2hERBMPIESClPD7Lcu7HmVGYzegnPXOGtNbGgkYa8cc84moowwXeihCpCgKmfPznTIA3qSk
qWafZP4ZU82RoY8ij59YhUQ3WFG34INU78gJjY4Nj4E5ya2SeL0tWTOn0qFEaZURTvR/Hayk7ev5
Vpn4r+cjL0PZw6RQZyDMgehmWvzO7WwtR9h4rgHdYmiXcEgWMpPqz5nTP1O8CTiKINY+0U2UdnJ1
2sjH2Kkkz6Gapc9RyWxypHqdgQLcKeC1nDMTqm863HKagQ6r/WU2g+O42G1TtJpFYH0BHv5/T3kX
ACwG4uj1zNXjAgWBmqiK8KrXMtK1xJbJVEOx195bkV5ZSbgjdZ83aQxvpjXM1GRgXX7GKh4CjKk9
ivL8f+Vt2Y/GBkDDe2Rh2uepvWhSwCusy5Sop0PVX8qet9/uvFte2vnUUSpyVgICKoZPiNYJPSzn
LOCY2Bdzz8h/i25tCw/MxaPtdhqmAk3uchTcCoaMqVuqDLa3V6AsVEr4KDzL56TKywZpe8dCZfYM
bl5LkfZbngv0vwohfV+5I7kN6ieaSDLflZh/FLg7f3GfnJ1E7+lrrw8YqMlpuFPiRKyxjgEnr53m
cQqMtjNhWzUQ6HbGkwWZ98U0V1immCHtKM0aD0wUrkvLFn4+N+//MsK6O2FE3r21ZFlpph3PlDuu
+k5w3M8hoUlEQxI5ZFAEX2NYDxBOfHv8qVWcI0VgKDTuzXr/6nHcbqclkJle1VA85NOqHVowqZ2D
Q2iFdctcSGIxzUsBJ5HSTItogBpYp/b98xqAWkger3ca6Mix8q459SEXO/S2TAVCypIR3crZ3pwh
BDRUNZglRHDRtmJNPtu0ncYcSQqCc/wNJQu5Hho8iZs0gn33fmbWLW3ONB+xE42gzSuAXuE1x+rT
lJb875lC6vMVFvrl7A+gbxD7lxlCSMDWyrCe371vZgOwh/57XH1N8IxeavfLfS1lsBT9B+pyhva7
b5fVYa7KoKRLSZzWHd4jlRyN20EHFSzxqo9gouKsdifeEJUbGRab+0ID+ai0kyaI5w+RD4FxnNqL
GH/gqzCf8FH/F8vx4g7m0R8QWKLBYH7rIdsnSv8vbw0RagbxhnfLjbsUpPM+ZPE/j99HjZ0fY/GK
ZqDUdg8jBYLXdHRwfcf+hylPNNXQtkwl+xIQpNTAWtHv3XFsLE4BrO1t/Zha28pcCyAfPZo97hOC
MNGNOzXbTQsdNg1cTTxgASah4/ImGiRrtsDgBbTLKYPoVAyVMIKgyB7T5Bceu5mVmRDZRGgwGUBB
4alLy2pM8KVs68If1K5JEDndEz/cIzr28haRR2k/gsM7FQr74Vbxe2HIa6sym8wSfahpNRmSZFW7
HJk+74wQN8FQVtpcle7zskIxMYJULETcdC5NdtgidYm4LgdQhGRndQj3EyQ4TAWAapkVGTmz5k2x
bGe4TBKRX6DUgj5DtmobpoYjjYJjw5ACutg5D3/EJ88z/0o5VyFoV9jbGBN7jFjQX0e4ftlUFc3R
h3XkxaqJG9arv1xOHWMukXSYxOQwMNaQk0yJQjZw4DSlNtCi+wnOQZwO2Xxrqutlrym/vj5hRxAl
hkDswCVnE4d2Lt2syA7SnzOaZZq4tm4faUcyj3CUkafM+H0vNbxOX4lkbPMSD2FlnKeBegG7j22q
s4epQmnFAatsLq3AEPxImmV7dBf8OUkCcZSAwA17InJpP9CsBF7M3lGOfEBKa2QvtNN3XWhXxl2q
9zgWId+3cfeWMEf3jCrwOeMLP15MRBXQjVppXh9ptIPEwnJ43aPIMmTmDQn0xuKUZrB1lYEx8oJY
DBn2W2j17o54TzJ2SnsUE8CtzfHGqZHxNVSqJeayihxXlDwhYKSKButeGBSKl9/BObbABE6kO2jr
pkHqAMYtME0XGBYgpgmlCVHy/qOiLyYFC+wff6hQjYDrWodvocp8USakYzSXW1FWAKTiX910DI8P
kxvi1kVlMJFQA7Le1R1x3pM4l+VbWJfvepjJodE97oBK8P14nb3dxl+VmEf6FyWARif/ebCbgoRW
V4swuTYyVvriaF0W+g8J8pBZoUj/5rxcxoMdkZGFy3nJk+54ntyOLNv9Xr0HR88l5knSf6BUFB5J
x3IEAaXSglpNAXHNnG8CbyZpe4QhpU0ezcJqMhkgpxHPku5Rd3/QHYVEHUj5WgI6Bd33LKxcO26z
3C4jO1md9sWJGOjPbFciz+7+nJ4UxYDb4Jl6nv9wEuBNThoXcff7OGNGMpCNpIq6xAGqUGDGqVM2
aB0Eoz4+/9KUUBzJJQy7sGGzYJhkwgalPxe8aQCT0WaIKTYmDPAI4v8g2H8NTHXfgXzHHcN205KC
aaYKNpsZu8gi/n+1kOTpX88e482G7vp93Wn/8hNXwgoaYXA3f38SjF3XiLeWsZpkItSHrayVJjQd
iKibShS8O68mx2KN4bzqzjj2ZNxU9zfPrZzPtuW3h3qujbB3o/ZvYfbY7uiEt+lq0YwtU8kntf+t
7P+e1zbhxGTBtn8D0ajjNg9b9hDj+NnUhWXRADq+InG9g1sW+7/r0HkqSe52hnTF7lCH0SzJdASp
zgw4QTn2gmnTdULsNShl6yU/yeMyAKpS05eJOqQup/MCvkiSZH2XF1ycZq+btXfP+B5ASe1dZybQ
pD8xe26qgVQxYeUn4C57kyu+cf1jlGbVRrusv8MOIqW6HRGfYUEmfsI5brN7UsOTE/4F9wnBaGS2
ef+0VkhLd6/ieVvI19Gwb6cy68ZA5ud/9Iim5K3ev9eDwBjUeXIJze1edHvM9N1Q5DFKUiv1dtb2
GOqNAOiMX2V2NqQVpBVHQZODonlT0ebT0w/VcJyTy+0eZBp7vweJ7nl1a82/UYnQbpfrsgYgJY65
NW4KucNimpPx1tRdYXU7raLpIYdWBPDPyPc6CxZQqlo0IqZ8q2kvFHnSgQqe2jb5JFWaeVfJZTVQ
9wt4Ko6D/W2D8Lc1T/8D1pii58tneep7OVCydNhpFAbM7G/3cW9X4j5CzI1pmhF+oQiEmFEFy9AU
OOG+y+4KGPX02kNgjfW/5RMcRwaFrjk83EtvXRCpjjTEUFZlWaRMWYaeKIB+6uNvCV4rCMVb+gB9
uhae57UKZeh+l7Vi13kqCqvGuBevm/aL1tAzcqAHqbuJU8q/SK1f5gziEZE1JNzeQXV930a8wox8
1EjKUIidzZnFw9VNMwqw/wxzyFYWuFRe5sROQdDKaIGPPT+hYFgZzo8qQb9vFR76HawowQYz0fDq
vOJkjaipKoinj2CWc0jRctDvFInjh+PkO5lX71leRmMEj9OuucvSZDsWwxMAsliwFs+/2LHtPEld
TfwZis1+U3HTk8zr4DIgjBPniDoxsOL6PbUrqhFRWin5iKOEzkzJFUzddnQacT/xWSFIcix2DB4e
h8nTAEcYOmxPFLSzK9h2po6IvqtJe8KQfqgXRkmtv3QkP7rMcq1SuSXxjmCOhA9XwbUMRzayuwUu
nM9wliwRIgg/b5jgIwtX4LMnRbaIW4SKsaQdVTWkii8LznW0AKPQRkTKNLrrwimvQ1oop1QOdPTF
YjHbjACCKSnh2QrDsqVe8xwzBokG1HqrJlzUSon20bb0fdfWbX3wiBHFOmJdubRELSUvPl+RTbZh
vDEIa039RiomFTpXiI0ZCKNS05VOfb+NjK1oE1iPb8vONHVsF5UK2KL6E1vBwMoHiCoDdLbsRGN6
hzDVCBX5RcHhyUuxQll8gIOqeXpovmnOewQtjwZJ1xw4Gf3D7DKwlus7YbC5+v0hsxUlM9UycljP
IfRUX1cyutWzv8b/QnNxtB3uiRkNWAj86eNBumWYqZR0bEDZhklxc7PQw3AxzGd0TwVbQMp18q7z
EPbzLVI1Rr1LasnNe9gsHS65F94blxV2PfPny/mc42e/pVgXMN+Pi4r6to+Jak2hHsOtC2wL+5tt
thikmTXwFtzujVUuDvz+HWV/Fzu34zatxBKI6xfjGD3L+Y46vVf48AN5HCsVxAaJztG1wfbN4I5B
HYMqhyQmx555D2aH8X3yM+Yb+BX3vILnivnZmMkd8BYBeMALUPw0M+0RZdXWFNLiZa/W5wbH0v2v
E4BRlzWG4oQ3ybBURxrpIkg+hNpy9gyZbM6odijinr64OtrphwTgHNLrjrG19vVwn9CUpcE6+zeZ
cad7PZ+jVD/mzWQRe+IJHC8vKaWafLSN30NpSMB7x3IBgBEmx1Ga9Q67jINRlkKkoHu+wItZ0kcN
ag7So34DCotC1McdSHdvUVGkqXYRpYDiuXSRaWk7SO1nhntp06BJwvZPXPFgmDcqpY3HtJJJt1kI
s3bTHr6no92t+tMdu3HXgT31aKF4XX/MR64Sep6iX4oQ8FPDrT1YCvZvYyNgQqCWKh8SxqABAiAi
5MqqM8lpVyuhBsUv62SAE1kFDgtRKjroCaJ8YtGXwmCT4nbLfudK90aivbRPgTDiM8VuvfMFsnBq
91sKovyyZGSsBHUjcTo1OAlGQP0fegmFleUUuUG/w7Hn9qHY0oVmvU0zfIq9qhiApxChfM2nUIj2
OXqoB6OiOzodltXX3VV/AriRYBJvuNVI/0KhkpFk33oclQaM4JeIkJXzrBpZNx50pGgkVMcFv797
j+A4C4VWK/RkfpK55ko7379drT3ddtPrZyXB4R9RwUiv9XmwNZVWUYOaPomb6M0glkv8DAIzr2cw
9RrFyxD/ETY7jeSVWDx8CrwI5BdYCAqD/CsFIe/hnrjvScbme6dOZrr9p6SIl/kTJaw5ox4eifbX
C5UIbGDYQR4/upEiPgeQw4WW33xLuXdFYqtbKcNXEnDuXiBzMtEGW++LJtz8BDesiSrN5jp/2hPn
j5YCDDQwP98iOZduHj4wRdpad5vVVZasdVX50+hFI+lSp0OmLoxOoa0s/E2hwo6pJ+5eN6oPutSx
mpk6KG7EioYWYNHFVJIWoZOIFZ7XeTSvxt5n4lPp2vDxmtuotySNVF2fsQOC8Smq/bX2pmNqatzn
T55uu/cL5R7iZLge6JA1hd9IKNTFegMNEEVlF9YP+g+A8g5OyIkayyFN9JMmgb2sxt8fFQV5DFXD
2mtfewV/wDOrNi9onnZbChpB/J8Aq1PGd/S856H3o9v6iNMWMiqOqmuJsWvvQ8lu2kUWCC94aPtV
I3Qve/NJWwvRJKYOEdHkpA7y/JddS+QtJqoE0V/WsyuJcXPUSpCqyLv7KSCOgJnv/dTLYKALkivk
8qpUy4A3yVPkXSAPnhonKpCApMXf+lvnHpneo0lulihph28Du5ifkppgnuixW1x5A8A2Wfa2hQnY
6s4+WCkTLrGAkdVseOxCwLgJ5Z8vV2wpOK1oOj1ES/otjZUTwUXR0gnsXshvLLd55OV3XNbCpBQn
vMDcXQ2aZXyTdLba1iByEOl07I7RRJe22QEUkFOb6nqkA0r4RZL5QaxZn/b6g3LkQJip49MAB1Da
puTiLeTrFzFzkJ8oYwWqO2yTgnGWvBcqjlG4CiJMvF7ZdamC7zdRvtCw99GqVlx6ocB5g+BQA6Nk
DbWrFt9g7XA2v1hReuIff40Rwdrtj3QABpYfWVLutkHiO8b1IMOqS2iU176GG0obSPGmAMrAEgHR
RvnnPaCpCSUcfAQGVBUbamo/r7gzx/ghY40LYSLBGrVVUdBz/diQjM75O6bmvMaweTVbTA0x2ZqI
ZJrzW3dAsVq1Qqh1SovtnVNYILW8SIFiP5B42zVH0+bPV+DcarC9q73fXup7CHtxgaDU249fPJk5
nedfAABrD20PiI1yNgPS4s/1WPZgaM1JWt5KjkitlbHAKUjb6h9bwmz4yJz83At2x4hFL9pqGYV5
chY5JgCLiXZXZ/6ZnT3sNpFCi0jehA3K5+8WiqOmGS1xGSCahx71EzZRilzwwzlZq26R0O746+36
0ETxFTjqAITNcJ2Zepaj26RKJDFagqpM8+H340JsQoyosznrnc8sMKOV6PK1s7+RKb46PXWboGVl
yKfwDremrVyF58GqaR+pdlbBdmtoK7HgPNmcRBaxctyxEzKN4SXI6y3OKKmNgGjBnPmwEzmzUMsC
0y4ecbkHQS7zIn1bS03Tbr+bCkP3/lDZV45JO0WQ29EYcxs0Vs8JdLayaCDi3Fpxok9MKcNu0YUS
69hri4zq6oq5l8n3puz3YO4BgjQHsfnTp9aJt31J7GWkmEaVmurT9bumPzqgUtHHdbKap46pl/bM
rp3BocDFhQy1TvcLKxMt3wbJszziZYZ8r4WNwUR7YIQpPnZYnanVPibhTb3JIUE1Pyk+dVr/O7hu
obGNkBtJDGB78TWa0qOFyrcm69Lty2t2oUYtVQ0dz5xfsF4hl76yYXNdync5e7/+/IlHKiftCs5+
Zbm/2ujlbxfGdN4QApShfYigu7ZaAdV4SguyB2DvaUvvtTEvsbRSdMXxz9mbPFXkkypPJkKjEreb
UHWW7YKzaHwJnPd9QoRHbodeLFThSs32YRf6xoqE4RHk+osShf23FdDT4LuLJRjzGypGgz/OABNT
Hmq4VMkn+fE9f4QRhCt8jMcpm0FWMFqtvvpYfgJdC/TeMw3S74ShIDZpVgfmS9Am4VsZ2LfVcM1Y
dLxANzEY4onHxjdKavusbznb4wWRJqmd8tC2ExOuylWhqi/8nvyt5UNr+A3hRbHMDBXcCPbN7cuE
QoF+8C9A+QgJuTOu8BPYcuUIh66OObEpCCSvL/GdV+QpOlDDFh1rfNsm3UJetO36t5GK1iL8dbjF
KxilIsqs5BEgWL38vuLCoiRBtZT0M7H/Ziyn/aCwHxUjLVRELowazuuqFXyaRcYuSYiZVQ9jFZt6
gnoEdouYzCe0XwZgDfexcrS8GS6au8lBdwulcaRaYns/8Oft1os2ZQLK0QtXOyvaf+lpv+0GpaKE
ixHM//+MMK8n/uiTnYHMb2x0kKcYQ2BjlBs2dGWlVcPL9T1QbK9o9/bi1ooPu2yA2MnGLKA70UJd
W7meL+y/xH2vIzlb5gCmpIiUu/PN6ka0rev3crgXW2zmj/nAp0+r36iwg7ffd1DJ+B6dP4dpRpIp
3NC/Ee3JSFY/PFEsbuNImCgbCF/Cch6SWN+SHW89R9107WrpPXC6wVNAaZbewc2cuLEIvUBhibhT
+qOn4bxY4wVXjGwNtWSDsE3nikbhmoA2NFZ8qwmDipLbXD9v8FoJKrhKjJnW/DIkRBXZKcyB6ey8
MdQGGW8eV+p3vlbPG4GEQrFyE9maA8PTwFrDyzve52RNRcfSwzqlX4T44a8DjFPzeNFGlmD+G6qZ
+wRtgJ3qfMCmTWhRhTdaEgIVZ2fiC0IimQF3GGNAdv4YmoXE07QwGGXTtUzC3geJDqEBXAQtsblg
w3nLZh+J4e8RGBtRKs3/056iYh3/CenQt0lRd3XndCAnnSq8hqiYLBo0VlqPEnZzwSzqB+lPH65d
qLhVSpzD/fx+zhveffGHXTDYp344Suz76kOdXCMn9BqVYVQCVrffU70ZPUcvrDKbl2MNtW1ZA5Dl
gAOobygsgNbxFtwdlhrTw+Yj1PgJe12b5M0pvw9BmHxHpfHml4b5oVFeC01EDJXNXJwd2tqqV2cw
Q4aXMbcHnfv1IkH+t9tuIIPCquX0Yd4Qc0M8ncqWLihUMvKOXQd5QSXpvs1RUJgytnqI3/aGpzBB
FmaanZWsKqRpQjXYH+E1jJFI3GplbcVYY89m87wWv9XjvIvMZ8cZxCJWp0Rv2D+Kc4iiayDcPtCe
SAdcletIt+W6ELCWSeKaySqWtgEIHlvyTJUa7yrDr18O4pNhyeb2fJVaaq5mxNQ1y0Sj6665VQPA
j5xHJWk1GekhuyUs+ccYvL9axTMfY+ktkJBQSTABL0kxpjXJzrg7sT5ukQ8M+SagdGKj5CRuUkmk
UsYb72an+gJJ4+oNagR7Khv1bBaGqkPPBW7DGldeSWOqPQlO22OS0RhGF4w41at5zykwNldjKm/m
a9kaDfACgMkuayRxnMB1o1pyBp1cLTD+v4aoZYu7FGnK3DQswpVPtPceQW4Kq1kVqPWKsp4QrGk9
srSxLd0O0OcS+V8SzCWZOPhkSoVjHRMcNp9czYieTCx53Y25dWl5Gd9t4B7TzvfRe8Pyc9RqIDT3
NOXHGshCIEFyhIE3j4AWlA/A3LlDBSJPq7BQ3EHUjdtbKV3kmZJyt/dMfcGoFYFVXsqBQxCEiy5C
uEefcTc6lPJT0o27gYm9I7vxdYaAPAwmmjpv/46tnoRgE5qtI6oaf8oQ5NMPioTGS+nyGQkMMUmS
dw/eDfdThrWSuB3fIw6k4QKyp55ea7Clf3Jsmw/18JWk1gUjc/EvLntMnOyYSG072/QLrtcmFtmO
weUeI4Qdg7MlKpGj65ctYrO02EjT4R1H24UapajvdHCIzYUkonjF5wWKfUm2NezXQY/+DAik+qTE
bukiqHaKqqGjwZIT8AvzKbNUHjxtkuFoVzzND5tk38IGtsMSPbcout8YUISInEGKzpJoYuLe52Ua
HJPgGEOL8biKAWEax5L0W607kgHND9sippLJqC8idpedbfT1tMkS+I7C4qJ8v0dtooAO54VPCAuW
XZhmJH6Dz/LFq3epdCfiPmTVzzIbn9t+MYCSsTi4ftGhKiDeoP3+MyJ8AhYDS2Ci+whwgWCcMhAk
PJF/LTphd2DCVoaczzOaquhccwllvSg3nLwvPOQjXqzzCRqjDijhVqRiWigklS2cB5VhBlbTRcQT
METUhvUPkv8l3E01fu2rYQc/VJ2/AnDN/Liq5Q+pSL1dFihZy37S4ovqvfRkw0gjisKijYI5rzU/
O8JyFdWu36gx6S7cWay1jGzZ/rmkk91e/glLqNSduMj/Hr9+C7rtaL3RDbo6+S4oTtFrp5qhmbT6
SMCEM2H24JnLNe8Y+BeSL+rrA3xIVm9nlbPg9QVA4TWisP9ycil0YHAbwPKcDDvBE3wMt17q8ECL
oGghvDb/e3JZYWJOs3GsAr029GwXTSyf36XHWTaKbznE/Mfd0tEavsCKWJtn2c9S1SYaTv+FjxMR
dlK5WrqXKjejaKzSEpDGArh6dgcpqhvMq01VmOkMdE9JiVPLS5g5hUqxqcr7zYNZLD8zrYZAfuPl
dPD2Ekh6PdUBJ+5HV42k3EOCt+ZD9l0Go0bpMBFBtCOUTa6jpPB5H5kTUDuvWV4ebm7ZSxc845ZX
45y63hThdsNeP2QWnssH2//s3/4tGVSgGHQYYYMwnDxerH/2KphuYNFiAGGJuZ65PyIikaaG4p3P
BXkRgFBHctPe5c9WkPXDMB+c8x3P7Nb04nGYosPXLdDTMDq65nZGRPVAwtQC7e5BdiGNgNVS67RK
Nn24vezJIqVEFgmEqkDA3ZJU1KYoBryETv4VOG/BWgHx/TnVDMI1GBWeAcgv3DhfB0gYgRSgMLCH
H4MzAtOCPswCkXcbbhgVt2v2cX/Zki17ke5bP/QlwhYQtUQ6q8BOXQPgdUH2c9/YUPmFRJ6k9I0W
FvHwLdPt3tqbNrIpuvFgtDoMBMZFuuj0+j06b7dGpCInAKyYqampJl800o7h/hRnkWeskhoGU8G/
ZYVMEGKZzNDX9t6pXLHhoO13zPpA0IC6uBTcOVhaYVT+Q5cAQBY7/nyubwGtOWkHuux6/Xs+Z+XY
ypjq3xE9Xe19Yyxw3BhjafwuB7LymU/iNJK1hS7P9YbNMpWoHdaqZvKa4qW75dBt5761eSZo34ZU
GzKWOFPnMWOt20kqH37DNWDIsfGvU/Pxh4Wk9wCyhbP4m7yftvty3QTCZsdkHYlDUnaPt8ea+X+h
b//YHYRh785PwJWTBiX9iMV8nwRXX9zJ+WAGSU0p4gwkD2NhxMfD/gqkIwpwe/oQZZU2hpY+kcas
kkODirKnAW5kCjWV03JgyXp2AVfMHXiCvwNmX+bnuQv75y93CxaYMLhhfDCz5YNY18UfrdXmoIgq
43YTVK3P58SQY/FWcLfmttyjq6kFmXBY/6vq90RqG9wdKiVNc6VIAXS+fjkKwo8G0I2TmXVyLQDF
tu5MIa2jX4x+9m1haIBedb3Zt48GOcQg1sLgv0rjni+sN+6FCRAnMp5wgxQuZcS53Rgdyup1tkbv
83Wu4edUuSkA1yQWBPJT71DVGBBMbY8M3anockw6IDTbcY+MfbmQfRcGntviEnN/l8RT04kXpP1F
3TGXCHJG4J+2aaYmdMVzbWsY+6Ehl/Nkda7knUp/pTXPnjaOtiYXJphgDsv/2D0RHiHCYEFmj6tu
AYiP/nssLk0/pcH7wNbwGWSVwpE+PPjonMfqpUNtHoFKajHzOyapu/SgE7/G2pkS/np29kTeTe6X
cejoGJkQ1PNRRS4R9Oji5Wh0HwGFvcmK3xp4+xYUL8IjrdcTBZqfubNTGi1qezdeAC38FQ/IHHDm
TJiHxdWpJWTElekKtdlXGQs0ZKZXGtX4lDgViLH7Yf4ARZg8PeFthnDtY/WY37Tdj4P3E7hx0AXL
zQZIuTi1nLwidzTDdV987ETXxydCtyqkbtMQdnD/8zuU0ChDxTaHh5Q9qmQSjpxJWvNnfheQyFkO
vBp9a7EL0nZa52aac2s3xg5mfE0f+634my9pI+0ZmgIj92irklcvR5psOnu0bTZSdCDMBb2Dsi88
bSLckTmz5rcKUv3ifMmGa+EYD8a1cbGcC5aWPT+fDvjSNA1LdcHPfTtM+DzyX6B3r2pgXvWMdKP0
aGkavG6t8MtNduL1vAvlU3G1Gp2NXuWTDQFMDRUAN/pgciFeEtDKq84cFe4jFNpBVZIiklNYBNOH
KmHfKZbdt+Dkyve7vI6SGL3HXlRmmBc0XB+fAIYd2H1RmHv07uVvrpuyv8a7E618XHHm5pWy9ilx
WJ7nCF8VFbxTBJLHHKuuorKeobmvWbC2xNPcanWTG2mS9UdKiFF3RF0JXs+2YxNsUWEGAYJpzkKR
pyREibNdU3pDId4SDbG5b5yZ7XB5iHeMWB+wqWtRAanbOv6iIV/PPGi9+VC6P4oz3/e7Es1c5nDs
/sKEtJh/o81hlrU1BhLH7CMwXTQqa7fkZ1Nhkgq/JK7kJ6NIfOtZhvDlpADPiigYAYmqjqTyF3zG
6vsUV+QceTAcuCQ9JBsIP9v76FA/xWWOuGlfXFRhMl4Zm3njUCUV0NVTVinu6ACp0Mg6o+Qwl+sv
hoW5LNA+DcpuUU7E0XMjFvJKxiIjanQJ1jVfb1H/WpeKLZbNYW4N2Xcf/lrKGN3Jo0Vj78Gce9ap
26cEoNdn5Up8zXO3nc1ftmpreEixlUAWQ6kmpMEGUczoZaHyxmQKJqtPjKFBaFwM/917BwA3SkJ5
3PuYs27Lw6EaawFCVJh8ue36P9Am2S+zxCLMOmN0oMdYwFC7d5pS2NIU5uDUfu9ybPAZLc1/1nUv
UD6FvPgq1SZWKt0E1O3Drc7fDiXE56x4ODkTVO6FyVH5zHlaC00nUz/M5VE2m0z4+mwJCrIEpA5l
sXLldvsmbv5m6pPrlDRkEAUeCyS6OxdQrO9OSWVBzLEyHuOqyDoViZj+Z9DedMgHh+a85Ey13yhs
u5Jh291n2SmYaQN6HIOI5SP4Yz2YOunWHbFP2tpSPXRnoDaK9ZOc8y5YUae3jo3Jd0XgLPIq3691
eOkNtQgZh8hi6ox8MFJfRF55GzTRhaBGhc+kFxto2jMI58DJffBplKD/CjYZhcPJG02BAm9977OO
9OyBqP+wFBK3dt1A/tGg0FgjLkd48mSyUIIB0UetPcfosP8o4vKbnNAGIvdUJEu+viM+AjGAGVS5
4yVDyaHHEfzewjh6wXU0ZHGqL+Spxr7mfXzEWQsSvXgmP9uLJ8zzi1IeRsOLnCNfOLGt37RKeex2
+SMwZWwjEnwF6pw6aJ1/HmPJbhVI2NCBzf1YMbc2lpAdSvVTMBtAsknZNjKqUogIpsnHeCGgLAKQ
aXFaYNC5C1B4shWoyVLvof8clwGyxiMN8a/595O5tzzUJMxusjFoq9stHDR4DVuMFFxdKQaMx7xX
StTmZesw8KFgPTxIGl+6qeOl18nRJQisS8ceWpsAeO/z0IWAK1F1jI4PBBkq7Y1l9115nuPWbh8D
JZhZMxD4U0sWG+NykgJVZssiF9bzOXA0O+f0y4FQgxFNGyBKi3NcWbfSPri0PnKW/P/l0UmRBOEy
FHKnOGhiPAsvrf+m6fLyefxH2k6XQI9mL/gZwkbBTa0CEmfK0xFNAOqJV8F9gM8hpGlZbNd4JA0S
Y5Bjf0jDQkwf5K3jIavRf9a9cymZhoi2Kks65GllBS7CFtOp795t3G+DHMKRayTiweGW8bFR38it
fVJGc/Y6s7UP0lMCeNM8Wcu6+tggYjX/zDIHoVXYub0s6j4gBejUmAG2Oe5SjskdIdX0L+xDnbYY
17F1ksOZTGkpVlQjNdfhJrCAnICgqspWXZkDGKK3zgKGwlN4oHjVzvPbFwsXs1vWEkNugBDGFCO4
1RnHfKNIoNykbZ7HPVjLF4OHbTnJy/r37k+YXzYnozdPSSi/nopnLZa3HPG1hNAL2NQfHnhtnBwK
EzBN3X/KzWm9bbwIv6GM/Vbb4iMjhLEmjww9niTDdDaF+TGrrN17Nys+sApmEfjejrp4l3qoyyuF
uTXYOh8V3twvrULJNlxF/Pz4bbRQRDLmljzQvPoxJWXQtfpfrPBeYnRRuLddR/pnAM4u41VLECEn
o+NsuiNj0Od6qmMnUWjEhKtWXiPSt2L/XxaVqMJG5IR63JHDkOGFx4/F3Jzjqt5Xx4oBBEv1a8m4
e7jVhPFJzwz5Ao4oSv/a0tsxPYA9aThc7Cg9iTlWec4JpOqj6txDQdHZp3HPRK2yWS7O29GaLPXd
1tcMsqsyUmG7NObHJEuFsj79Bdp2MCRPXEbgwXtdR1CmsnFztdnuDS2u9L6jrM1Q4qe6GfJLDJZg
1W7kIFtzBurRXAx+q0PfB/2Fn9Z2HocM+bZXjKdKQe9WEc2kNQKv2ieBSMjASNS/dW5X2NHb5FuN
JIyMKDdOM2svgs8Lv6wXTfuINDqbOZEeDw5+fsAdOwj7tJXiUrorog5On4ERlB6B9q+HCGHlOyjj
IqvIQkdyG0fg7epG7XoEnPDKt7vb9WzkJNGG7n55G0gn14GX+K8yjihwIed1yissxhkOQx7GxEI/
Mrjr+aIiB3pZEGea/hDAwiwA5pdnBGhmV8KmNOUdfCtT/9i5EV4PuMSIG5PeWm5Em1JKN+mxR8AO
WCsNG/ywunAlITHj+FeqBHhhe8GmoNtbqHotefRQuEgLIPnVkSOeOLQrG8giH6p7WhZ7YW+TXc1g
SLRfK2qE08R8swLVCL3QAsgW/hob8mgeucffAvQrjE8r8icnX3Eyh70f6wCm1i+dWeiLdGInJUBY
aeV1ol8SeFMsXo/pxo4iXkG3DyMk8ltn5gDwSP6Fj6r0hvORSYT3wkcw+g+OCKFtscgV6xmFTS+W
YSBb2w9FfEjYyVlDpaeu21zbtnvT9TEgJjAQHq+RalAOgqzvfrfg74FcK68T0c/o/zpP97VqvIdR
NxsT5OYVvetFWWx1Akm64ZTtw5BMkUt7h6ECgI7iucKJZDcajhtTxibk25pfLv6f6abvNsG9Xc7G
7rGSDaH5/EerV5JQy9rrGxnSG4gf7LXCpScNoOWSjLRHFY3q+qDmyC6FMBusLVgBuE0aL+g3CYUL
NGOE6Z/Z0NaP5LvOUzpQHTtFGndsmyLsM09+gbcxk7qro1HgjFZGzC0PDS/KYKbXUohlMWxcmkLZ
lLCFuMN/EjdyvNPy24/vl/N6dD069Eaps7jbLEPE1P1BzIcxIa9k6VGLXl/2hzenB1UhxgG2VZuH
D6u9QpRX7OczNzjNrRXj9zS4P1wqNICbtaZTpBrpnas3kazaDSadSdLMm9M48q/6M8fUY4yZFjfo
9SRmuNerblBP4wDLBwmysjcl/Fjku5OklUB5ilBqcap+ITUJaIlKsRPbNiQabXCBwX3drG57GVB4
jGyhSwXcroKrw33OPis4khecMVdQ+d2rOARd1xwCj0U7C4f5+H5QFRbB1tC/4qYsaZe2kvVIFv4n
KGo7kCa67Z9bqV7YoEiYqzT91qwxJtT3vhaqiyf4wyt6b+NnSbE6VVyr51bqvdk3+XjX+0MGCKN9
wa5E+3JJHPq2URe8V6bucNSF5CgN4hg/LAZgkZ/Td/kBi8/7lObbzHche8MYr+FQQKmSZNONbfqH
0ZY7ANQf0vYJ0Klj4UhDk1G9ayUicJja6kAsDjhlk1gFfQ7RI+R3MECVsBWKzpqm/a51eYsPwH5i
GR90w8+/DTgzSJ7uiQcbDVDMxqWIW5HHVhc+8bGi2OFxqcPnGpLfENmRhazfaGrGzKCuARvssLOl
OQ/mLTzSO5IafP4qghRv6F9LYxAnZeHmoPVLsF6wbKZGvwYjqNJGThjhgjWQ2RzicKXpHL3qxDmA
ZK+FfTela7kKMW7cQtfYfyYqtzJnIvVACJNlgdtPIOehZbtEq3w3HGYWNeGydYFGVh4gmu8+IkQc
Mpp5ojAPxXhD1wtz23a8cS2jCDD+OxjJZW06GPYsj5H48FXy5APPrSnh1WN7ZImtTw14jx/0SdTs
p8FmtZhP9IOgiy/cFPsnOBKiYncu+bc72gxnkWkIMVUvjjVZvYX2XYkw0MJdawe4hStAcnpjaEFS
q36kaZV1Uwxa3UiYElLoJ8q6u+GLPxronh3oRsYDuZxySHCL42xzuZxHcPIQiGnlGBi3dmrH609a
S+160TACJmTbq8beMcJswyBEtCjC03Yz5SSkqVpi1QlSC3FJ9+eHYhBTeoIlyi7EvIqCWCYo0J0X
lFu1wM8HyYt2tyNSgT8bcV9ZPJ86utND2gY+SupjKsQLXeKqWQXamviVoVSpE/f+d8SB3yLfn92z
H573HEnQZD+FJQgKKRik+raKRtfGVr75/LTVjL6TnYmtGxaXjprBL+G6qmONE59TCt/7Um+LXXZ1
PN96v1kafKRig3KJUxyxUPBN1CE0HZTZJzG6Pq+QUGBEV4ryGB72ahwYilR/Ssxa3jVYp2iI1JzJ
r/B/edWk538955oD3yLtD8mkDD/1pwgf20qS/QBFoFhSvpQNKujVxmofE6K40iCy4P6Aangbj+Rd
1hyRS6kZrtm1vFU+MpRdCSfYglVCew/YSKUDYq7FThDPQkmWVytN9+b+KuBc8OWKW75rAzLInXul
r9iAbFjVGJtZiP9vkouKuUTpHe2ab1t/CzLEDkEwtiCxjP5SEyY9ddW4pDhV1HOJR7XYpJFBvBow
tWR3R9Nsvrd7N5pUAwhyxaM7gBH/x11fFHeEoT7VvC9vJCX70Fd3rJOObvqWYD7VU7JH1XkvP15R
NcaEpXveMUSVg6aVWEOEMSJfC9yxV/IlxT5szwIJR221/3qjZmdIRM9r40z6hlr7rNXOQWXfzIr/
WlBUXmS5IYqlPtHOg0FRExcZFISeSQiSe2F8eomHjB7LPgzVGj94GwP1NotWsbwCyUILC4epFJMw
5Q1ulNhKGsENeFPpkr6qMEX4Uef4pwxgiE8ZUxsTCAaL0rDjr17EnvWC3R1BpbofDWQ9Ak1txl1J
TjQ9JFJbL4Rk6SvnKmxM040/aqeTai4zmqPlZu8leIRfr8325vh6bdKaNe5cPkKMg5ilgy17iHs8
G8iPAMFIIjIHT7CwRghfWLqwCB4SSnj1pBfhRciNQCYu2oIQJdeF5vM9L8tzN5QKmxEVv8q3Umm+
WhWtgzRqJMGIQJEtzlOUj6I0EiAMTWLio+KuR77X8Bq8S97//rq2yhDTOlf+GpaOwuFsA1pN0pRU
w3HVuW4vLSawd0KLs/liPfC8pXbGJ3EkbqMjiY2Yoe8+EDK1AwR5mzRDWuSeezxsoSlPAryLI+b1
ka5VrbT1RKBdFg9Db6r9sCbO7pFymccuXN7MXcIHYIVYAZHSctod8EW256285Zso1Bc7pb++hxNx
ThBL6WkbpSxH1NWtmwk7b3Tu/4SkiWtOpkh0Z7nAGnsv0SXEbDcoeS/YH3SMsN91M/QrnGZopiDt
DFwZwp9NV2sARo8TdpGHcL+JVzDN//nusVrky6su2XL4jiUkQqWXziZQIO7dj7SQ8AWM516PVhKw
SmjZXoTQ0TozHk3DjXy2LISNZ78z5dvMtjmAvUBRLlQ2QJUsjE3KOrTl6okCNGnSoJPICVViKleU
WN+l5sc0VVD12lXsSnrcSd6RiRBbvSiqAIiWbBYgh+RzG3xqRRr4yD1eM7yx3JqVyqt5LIzBlWUo
nYekuiAg97+XvUYsDDXWlon9pABkpWqN9UgARgVXgLfPsZQmErHzIJCpWVzk9nb/wHqZm7zvCOnQ
gfl+ADkmBpGC6IpzMCiHrtTDRrPngAxfT3L3yYmEi/rDXnJoHlSem/A56wUbeO4XJXVnh6paEKcB
sQv0uZMzjFVUE5hW3mkN76QDBUWuCq5x2m9SznVE/kmuq9Lwc+kMO3BuGRSmWp/qxhvwSXsLJC7j
GlClSP6CD9Iw9Zo/ZTXDfQ91N2OttSjLODCfMeSaD81TGj7TTLccY1A4VewMDcuzMV+X8twHkC2M
rFyD8B3y9xgL+8cYTuC1nJMB1UA+iQffp8Pd1Z8NVUahUqbAskOcm+QiEnTVyFI62S0oXJEL80JY
2+Mm3vTGWFnxr4IquaU13aBXQZ9TJ4c+y+dIGpvMrw8Y74vfvhPYaUx/uxXjiwMrruSVIPMU4fI5
AAcGKnOfrD39v8k2Aw5iY4BWMQkhWpvAIoA3Ll6lbpWbHiiM9EEf4yl4Te4FtqKfgD9l7ybCF4NJ
c477WV+wO97miy2Xar2/t641ga0B5N3S8GazlrdUoFKcOXe1sF7pi+RtIln6PjVHGuaUgcpYUPdC
erM3jf6uLNo/vs0jRVSc0Ss2L1dQjI2pT9J/DWLXpWEd1wRZbx5rEhp+opIgrPONJMGEvQLyptFf
CKvesksgfHzW8h/vbMF19H3mx1HpwwlVL+WhHMjjtYZx12/4PmtYNECUPxfVFILbA2zMvn6sa1QQ
lnIwVbLaCa2RsDO1eNJTqdNQM4soSSUjhyHqRx3PUWg+AxUJRdI/e1YTvKA/ipmFCMlUpHu7PEhV
tFLsBPf5d1NuDa66pWu9317cVSd4Jpm+ppmmXTQBVdWK1J/k7KsmJbieGab91rXOg4hROv2zGmAX
MlukcZCOJRL5vK2wMsYIG/1rEc+XkhC5Vt3fpDxds5bCnMwWN2ZPPG2SNe+DUfNjO6JTnvErJaVL
bUPzEyDxuUtrUqhRxLktHXDiEBr7+oUtrFNP+A8Vrnxy2rE8qYQDfghnydr94iJTVtDs6gdzGtRf
gONJkYKvXXB69Mz0sIoI2yd04bT8M/yFRprTMCXabla7gGbknf+aaA99KTFJuisIufSlLbNL+7ZL
Cgab7wVSzbhj20QtrGYnPxgk7Dp1EKvGPNS45p8PZKLHRJeefscFCejVDEfHuhjrqplcStjDxNSs
FWvaoAmKpXiXbrD/8N+RvXuuG4T6isPWdjIAkfxqMkNsy4GNqLLlSmmz8yWllQsTi3Mtuh9uesVF
LBlUbX5dGhHoqZQdLw0xw3LKnJwQwi2YEmt/aBiDhIvKAc+wBqAiO7fUf8Z1gg3M3DzHbecv9i9x
zu6eoTf8mdcYiP35EtRZWh99+pR6P6bIJPAdcdcEZqB5qpTbpZ6ZBTqebQpKVRdmUlLBHhhjLNFk
zQ0fhA0Ng17yaDz07sR31CrZA1RxbP8kcbodrz9A+klPA//aYnORAj7JBRke8ZrMBuMg8LITS8St
Fcxu+PYLkYk+xyZhu1ZSPY7o/uBTU87ZWN4eUXJr+f/kyBNsrT7UAlM0goOKnGTpFnzwgfwm64VC
DK8MietEa7mdtihHwOEAZh6LTBVf6z32SlsgD15lCeMEuy35EjMSBIuaBEWcrC9C5sANZutIldwE
yTgmVzLKcimVeTV4epPjliz6+RxyuZswNv7lfily+KFHQltqw6ynkrwoUnUpAcfWfqxamuPZC7GE
rPt7aSJcjZJQe+p6ebg8LN8TjlqbZggksmFXSCNqtw6lIhoOIVQgUKjWxFU7Ckz8NFA3NOmKy6Gf
ho2SUHucmsNZJdSnAVHQHh3YjMYZYzIVweq/0tK3H54oc92Fb7KnvyMReCUAX8FTbs4L/XGzEksi
HBfJvSrtUjLCcdd7E+3ceGgcDbsxKg80OVfa+JlKs3pB9dJCB1N1uNN26oIwrG0Byjvnqmc6OuM6
BwjQfPVBsnt6u22DZZ48dLAF4if+AwONMeAH+vmZqNzlb5JfDWXKeEIcDfctVrboMw/8Iu6xg8i8
B7W/q/1FgjEYjBS5DjKPYwQtsCnDc5cbs+OurJh7UzDk/G63TZwv/LKiJxbp52OEUuDmmPfIZgdv
PMpeYRYU2DBwyoveOs7mrjjfedo/wi0qaJC5Xl1fB5iuN6czCbAePAR6Nca/RQkf/4UaEsV5Crk3
IgTmwFf3UOe21oup+y2DXuxfgztY98NqOTXHbwfG4U93hL8aHBQP5C43tRqj8Qg9r1Yqi+Fu8Qm6
9WermpSyu8A0rv+zncIV7iUCjhFQ6ZdUFbcqdW/BDK0jZPIW5czxZjXUqFsHY7vdOY6hdcsUGelJ
cdQAAgl+9rbNGmKebScRGUtc2YwdoPZD8Cn7cmdxOm7qkn30CuINOGAP1jOLQr7EsUq+77Uq3Ih4
6ULGuZTQDo0nK34dBUyu0TgRkP5CkKFuC3tP2GU2mZKwh4Dup5kglWV7FzLvUzf23LcqSFgbtolg
LGpaXA36VmsyTYzVLR4yx/BM9U5YU/gGCPOe2nKec8ZmY2BJi+D8YfNFS72YpxK4JpRMMdT3aFjc
PYsZFE0R+b1KZ7fhBl8OW/d9XXMGhYrx/mQ2vANeGlxoFi7piLYVn+eB9f83UsmIYfuhe2DfiJya
vJ8gWqQfuJHCXQ9RmMWtxewDL0GuMqfbeVIP+sGo8W59+aI43lOFYZegOYslaL2w/o1nCfPhL4AJ
KYfyx6tHmjNtjCfFKU5YoBP+34j5MsQuuCB3wxOYsqK5+ucpSQ/MSh6eKY3y7UWFHHXcMqQ2b6hY
zP18NAm6D4P55X2b2Jii8/JkhtRZNfCahqe3DEE5okPTQJLuJyvyUkntYaamiYrcOdF7fteMnwFw
Z/S189bJoYKo+HQ16XSdnxnii9qJfpUP/5BhX4VbEGXtwWcEgmirAqZl5u81O4xZE4+h1xVKK7jO
YlN2afv5GPGcG++sRzzxhsoohLnI8l+4knO+jsealprI9T03p7XE6PwopI7dEGDr29aVUGwPlw4P
sOTAYp71dgSjrLUfcvi4CsDtTuYUYnv6wP5ewAp36W52OIc88dEv0ws+1n4bjDGE+eSCSRemcyFr
JIAprG1Zdz1qn3k9mRqjxxoVMrpiNtUZrV1KpFq0kTxxuzYZKxR4VatHpr2DjnBlwUIS3YcQP+vk
hc+vrAfE0cZPyqryeEmUNiclQ2Bhtn4EdwSztkPYWqI9oBfCKRZrZ3SbFxNcwPqQ35VvEDvaFNBY
hTD5L22uZEI866Y+UqCXHThJ7EY+s5LX9GrRIb5S/WILa0+/l8u4vhHRGi2u+Ftn2ObGzVRcHSmo
pskFGTLEKX0QuMiGxQVvARGItQVssA8r1Z0YTIElpPi+mkFp/3AjCvK6C5YlBPZwZgn7/p1VnYv5
yPMHE7muDmAP472JT3vfbWKmf0TuTAxPlWahKzGfs6Jc1iqoV5oAzZGfTcqCZg/pMqMhRUOBSy5s
X9T8u0Kvo6VgLDQTZyAFDg8MENr5wNtvSWNcYQrKniDHM9ru6Pgi1+o7aKdI60GJO3Mr5QKnRkYI
upBKhQ4gp2zYO34UNZstnAIH+kHQ1VqMsEWs51h1GmUNCr1/S6qzKTmM1eNeNZ/ta7KYs/BRbQPr
HuD8MUW47nHUFp2wjIPuzsIdqV2XjgpMXiH6K1qp3BQvDU1El5ZXR5Q6o7hQM6jeBEE6O0gWBOwp
+eCVG9/DqS1/T69sRx6+kNsZROMS58hMK+gDsjuK+voAYmFwPsQWwjrYOVz2OJI8rENb6yD/gTJX
FZAsMoF3UMj39YXaRJ+tngCHo1ekZJeAkyb7kBbYmVqLyOobpwDQFpHdZsuI6b88Yf+xSpW74k7H
aakykWqitNyU8iyZMup5oSoSjjxA8Q40gS/6HBhCMiEaPrBJ9aq9Qw7D+A5TEAfiDcBbBucHQ7zp
cf0GRET2ZQAKmJoUjU2A1ALBmyKyQFlRlojnK8y9pcGFqRMXnKoufnHONjNt/7FNq3vWkLDKyqwW
40ggMPKMgza7dSJwYRgM87b6nlNP6hoBwzuN9aEMpiLsE1YwHwR2Lfz8znYeS64mDYASTVe05Cgm
SiTAzW/BPcDwcGOhWpgOdc8ns71QZnE7hTMLcjin1T6v0uaXi2sD/gAlwL5QpZRuIuhuaACxQ4Kj
p+GGihJvI8BraXZJax1+um3ajrjSn1QsRI+5mpBoPy2hrSlB/rSdsTinWVQqGKkK5QPcVWuNRpDR
tXKyrzZ/qAT/cYUoRHpW4OyaWtgONowwjFSn2KdfV9pZZVo+vMyQyGVoefTeRN6qmGtoS41txth6
XPXAlBTRYFHpbgXS13SVtPsShK5NAMh/TSCMsCJ41tPzWqqbO5h8O/CAHAsY+aEH7uWa3zDqZGVM
BgsJRkno8v/1fWXBTNAVivDs4Ts0nZIRDrrWrmeT78yL/Q4//C/pcEDI5kfWficuY1xKtLek7tiM
EftJz/EKozuUVK4mOlB/PaLsDtY2oHmjoDnQFzXOpk7qdjUJR4Rp/uJWAppdwtbeMdCr2lsFSs+M
cwy/SVvtOhk8CzWl7I2kUO/pea/j6C6E7VIx5ALrKMsEMU10uEP2u9TFlNoV+23g9j6wqMW/erSX
oawJ9bLcuIUYbRphBqkS74hh+FP1i1d87NinNNS49YsVVPcZ9suU8Z/rg1/bSjkAGJKvM+weU1d0
Vrz9lXavhCTu2UMMC0kZth6n+Ks3x8WS2Lm5+sXBtB6R6vkDOJ9l9EJ6i4sfjChm7beMmvJNRPOX
gXVgfcRWbqq8nF+we3Ua6mjmFSM23LrDzQDMeHUR0xNCIxyFCLOsGPbl3lb8SHf+qjJlVB61UTPd
CNutMabGyNHgmQpjUP7QdO5BQbi2yrHdf82ItKVQS6raMiQyscToDyNzavrhB3PIXtAtqHUUV+lU
G6MA+r9JdOSg4GOeL3o86NWPpAoRFGg/KkO01k9eM6W0VPfSYRTcn/vASKbiQwtTw8P0gn3lTpFn
2MJZ0kunCEJ8rGsZYYRqGXdkPK7jwjpII9sDdTF/bI//XRMZlQbM3unCIt1gnunY+dMBEP0TtpXr
+e8KIzSJSbEmvx/UCdODH1liUD9vVX5IqupuBMVhk2GASiQChrcMsGE+85JhImS4uO/B/NOJLxpm
hlXC8YXFJv3MEkTpJLmtnDkU7sgNIct5HBO8A9sOU76Vloir/9zYFoSQDQZFnbjOfl0Vn2UoQ5+/
0ROnxFL0xO5VNcxELEmv/j6IcdLY1aA3phf21KTjJMz2hPkT7ussNOq08huXGZU5W6+AvbYsCiA3
Z1ye2oRY62T06xeYSUMF0pIIvvFmg1IM4Ke0RY7iGjq71R9CY0lxOT8uii4gagBz2Jxr9UMHNXUp
/wly1X1veEBvKPp0kYAajQA1mf+NcoheJRsuyuYHi5zXDgvupoI5YPZcKfvGTFRVHAy/bjOTs7sZ
UCvCVmLRsqGUM8Li0GjGu2XhnmxtBPU66SI2rc0aIfqFU5QfFJweufXeEdkB7NzDOyPMxyF9Xx08
lWTSlyNwNWkE5Fd0kp8Jl9sbz7SFN8p7q2871gv5TXmW6Oje9RotcHx9D1LRd6EWsSzarseAjP1M
+TlPGJEukIB5Ap5r/jQFLkdnW6WS3I6jOoZ3SoedbBNqCb1HzvUSGTYc48aVyD5dJR1zDM3iywHL
aEzqZBV/7XUGRKatVrF38L/Kw2IHLqsQG1hhm1GB8zuJ6urLSRFhamWX49H0K1lhb8PpNfG4qoqz
rBh0BLp+Uun5JNot74GXvNKDZhqDw6us8Mb+tm9zYdzMrWfl+ZD+vPZ+T0UqlQYVaUuJPmyyzgXS
vayAKblqpCMon3nyQSDHFCi11LjJs/mnfYM3giCCUplwG+rZlI3FTmsalmITOcWsx1LU4eQJLbpy
V+VjSElbWA6J5wfeuH+JV25ff2p5IcbiIlRAOZljFD3O7W5F6Cf+gBYIwuH8OVkH3yiki3/0tErm
UshFLFMq3m/60U8WZAcdZcQjmo8zf0PfZjjDQvES8XkVZBWQG5cB7qYuGLfQTyJ75eSsdbCf49kh
KGl12f8035Q/rgu6IcRf16iJKLKYLNjaRd3DLW7NT2ZzSsfCu2bm/ViKG3nSh+rgQR8OFHGojSTV
cmOKq0RKkVoRTJtNzoy7Aoa9217UyqNoL9yifp7y0JkAnvWkMk+u8D18wugtBoVe0E3V67NvQ0NS
IlVwRLmF7NQjZc1kSpVBS5HVs2Bj7ufB20YsGL9LJvvbMcThNW6lmZHiFFL7UkfxivbqRVlW1+dD
ACd42ARtWmLkSNBoq/LLYNR/HDetLb88PLdJl1VGseo354GpPHaz0AmaHAlwA/EQEfCS+9Zzec4s
LR3hRfWlVvQaqCigLB+1jCOy803ssxWxuJpSe96f+qPJhVGZYTlR0nQR+fr53Uo81V2liXxv05ow
bavIMQ27wqwluMgeenmBVrr+09Z7XKIsLc7K45AsU7mDAJ8ci4Iw9i7zfo8/NsHQ0igeEGW9tFDM
YAysNwjCXbZAPkfUC20bhxpjcZM4ET2VHtURKyJifHNAssBOkkc8mkNGRpMTX090KRvUsHVoUvJB
CV3id3P4+jqzdqzSY4Iln6Yyi9zwl3BUEkV2C4Tz1RK+Hq/M8sB8KyKcnXOzMC8dtC1x8nABLaDB
SU00QXreP0+vQMcT/5Pz/MFitwtn1sdNahSDfEeex9ZTI25mL0SHrsHQWgltfQh3T200dVsGu1Dq
JTKkhemdHCZHdGN6W9EdibX5VGYJcc8oz/nM54Q9KV2rK5EGgEm4D788N7KDyPaHvBXfnHd6OyhO
yixMMFUb1Y9owCSRELm/W2fHFu2UOLDQIhT2VRo2V7Ku/VPt07esqKEqS5Z3mq6EFVlUVX5oAkSn
3zCqNGBnGPwTYPHZAX3Enb0KoA4uOR7lliq2oDhktLmNZO0HIITUc48u5v6BWTuwH2KlmtRcQ/Tz
65CmvNX+h/+UcRk6gmj/ggvgePOZ3Zgbyrug4LGJ7q9JlkA/VmxE8RaJp8+FCkHgq2BTs8G8HDtn
y4psGIQKlfeiEwnCVznLO/9VbXD+OWLgMsCNn+CISyJxuCVQNFcTBbtqEnef3JtHIONvLySQhRgh
hkFWkjdJueTBpBs9FARiTF/AQQ+ta7MX2iL/X2p0dyHQWo5bLrkWN5O70086ZmzBVl+IGjQUDV9z
BnwPuSz3uzpW/7blWGx9HGNCZPPeJiaCc+d6aEdFQpGjlCNREUMGhGFPO52Op6LkhHC6Nx4cy0Kw
9ezMXwEuO4bqEs7nH+DNdzCXeZxTtS2qgkkceVo9NXJhbkQsx4IL8kXRu6lE5UUSu88tCyb/FdRs
2401RvFflCF3unlNImtUNLpg5XRUBSFApsqBxV5wVV62bFfz86uQWmx1Wmt6v7P9f8042w+4RY/t
FWNO0+XIoeOXiyfbTeMwvyB//y9inLr6sFWP12YduOAC37fgyAaOvriDuTTLu69siIh9NVX7TwPE
pc5Q5MT96p/diBIf84+jXWZE4cvrcGiej+8vvif6Rtz6hL4SS/B3SKJ2Uqvwx/ltQdZQ5Qu9k+1f
zs0J35XXyCQJus7JlOkJXNBwHhuz6LMHBcqSgcjN0ZEFobk1xyq+tJ3rMwLxJQkV1KiwRDZhpAMc
L2m0KvCGjODErGdHUbFwYv/pXg3ifs5ts8/ZAJ+qxocNJWE3eAWQPA5NCM6zgFUnk4xS/L+M7ahC
hUfB7lr8MmugVfyMgpatkqBeB9fHoY+sh03KHQarejo79s9v3auO8OylVjt/GpWYYEn46WEKp5gW
UL612ECnxeoX3nTa4+KFglb6Ic84MPxC7UFIElqbw5GxFsWXmB4oRsaNNPauZPNnb/JTqLCV8GYw
Iar4lwUUdne1bOuqXKcq8pGOjNZy0V0sZPPt6d1+3XJ8l2jeuDjiouA+7a3I6Bsnk5JLxcwO04cc
Zo7si0Wzc4RqfQ3vUo7SD3PHBv2wcagnV/01FsG3zfs6AWlHVc6+q+nWZNcMjsW7EW5xHxHnDARj
lxpVLvZQdlJgPVaD3KDbR8OXJvM82tSoWKSoNbrYQF0zIWb9zQnrDAaICH9G632DL5qF+PKUvQKT
nHw8MTng+LuLR2/ZqzA42FP3gzw23c0RT8gd4b7UgZ9lSy86QNO5URnpk9DmiPqwqp4TG2+Gt2BU
f1T4YitE4av+PcRo+mma2Hht76JMHLUDOWE6B7omi1o49G00NtDxo2SpSKPpk4V2eLKszUaBQecq
7xywpNbHlLYuhqxvmfGgN8ARettJhrkbIQRjpTEnrzbIw6rNzfTl0valjllFwC3QOUnd72lbBAVr
ZFF9l6+4GkayJX1Qmi5i1fp8tNiPyrFFVmXAlV0+v4tNULPibi+csEpFuSXv3bZSYbjw8dLVICPR
oVWIDeMhKTVx6J1AoXhtQv2AoTl0sPhXrM8XsCNLQpfjGjMjdg5szm/vP1PTqaJutJP3JQuN0x5k
5B/oTLkoopf8CbkCF8Eq51EJLCZhh90s6seX0i9mNBXwPS8SwvhE687/gTWSPYFhx8bCwt+CNU1i
wVFkXQy/uyHlfdCBnuyOYLl0J6bc6OZpqnSpOimRL96NwtOyCFQ/iLjxrLCFuHKXw98PcNZsTPb5
WuKTcjD6Il/WA8XEqkAHG+/URV1aYvY1D36jZg7n8ar6ma45FeyTgkeEs3H+jTuWGUstkEVtOLsW
YjxWAChfMM2Jo5idjeGjFBacO9W2QrNDtA44XAo83h1nWWnMZpKhUClsPvOfwIFAGI8gov3AanSw
hCSt2RIB4+wL9Vw03uo+fs2nITV45QjBkX0t4gkXfmEHmcfW3h0ATxFMJWgNfnJnEH9l4io9HiUf
YxU63aZpljcshwYQSzVmmRrQs7hkvA1ulAt82S144OPf31jicHMSYsSUcW6cIw+vgkydH7+aCZ8F
vO+GmChNbskdHYtbblS+2wSgfF9oO1pSA/fPvz52QhPKW16SKfvcb5VnX2AQ/PHkuFraijyKu5FV
Lezp7+jhsDf6Njqn9bCNAbpUK12bnc3LFj18/f1a8gSTiWEyWB8Y+TuQkj3Cn1P2No5Ahd/8ZZyk
uYBBmwGw3YOs503Svfdm/FLXRPhYHE54kZ+79lWmKsSRFQgPaaNRNo3hlZGXkVpE7gxbdj9josil
AgkdTh6JFy7+99iUOc4IOYrM6muflTpFsaymb4+6vM28nDfRRyVKmcV5vdIkfaB+Iud5jeBGzhj/
XxDc/sEeszUm+honCRnBrDUvuJ96fkycSW3dxTCsYKI/KJIL0aNUEDXNgzHxYJMYPmhfCh+gNB5M
MnaXVMveDVx9j3hBHeyEGAigA4EHNZ8i7UBUPEM4UnIuIJdQVonKdCq8Mp6K8oKwbNiBOSBKvfd4
LLg5YBeTgbcajYxt4KlZns7gXBp9KsRlNDl8ngtJX2z9DvQTlBiYEh5JMK4alL8v3Olhv98Q3ZR1
ts/sj6HJgkP0Xz4gV6TrxUf3mEK4d61gzBp5FsC/QT+9CEdX0RqQ/1h3B0oCjtTboTZU9v5OD/dW
r7tgMmfhuoDsmLOJgf8Kh2sDCPLO9ECAKoytWrHfFoYTI9GhT8HecECQQjGbqgZVstf5On7nW4kG
796EHQ/UmKYP1imcPt895vUDtFzegs1qsz6JSpAaRWt7dlAUOsiGQND0BCjOD1Nbpl2gCP8Syc9U
SCon+80uTNYfiKBEkJebszgWXbCxMGsrkb1c18ld9pkBxsbz6iI84vBnCViV0On/7Boylm7L3mis
v4R9h1bF8vSA9R1zWibHL98eyBGasWhbRlNadHU6g7tlt1mEQTsfUeI6QKNmwQibgXzpTRlbsr4M
jTQNCvam31Q1MSEm+lTwagixT4Y7S/4orR0sfvccbuIkwKVZTy6jHBcRMzqG4tfTf1kqrOOto55M
q6Uf93+FaFH0RCDPzBGXeX+Uo0LPRcZWMxr8FgyzbUAh5qPpcBm0e4oQxye/CSbI4I5YddNcDP9e
BjAX64yrxRf3wMDma3nX8iSzI3BRErrBVz/KAsaTyxoE1oEk+J5q2Mw2nBsd7AX32bAdHlAsf+sp
IRK8MDm6HzKMYTSwgh/Mw5u9jwaGLUGGo14tvAuJhUW7pHm8lXxNnIZiOIG7o88vx6hTAQd7bcyg
3/AU3Y7fG5HkPMjSiNpvRu0Nj7fqB7BmCKhyauBBO2jolw19R+L/DUg4ycyHkIYe4SPTqiPuRG+q
BL/TlM7lCkOivNn6sFXhtdkyoRg7oTB46eyPDPQriEBKc1fYMTiiDE50Hh9hd3avGpUWLqs/T9jd
9+Bcv9iMQ/qu00q1UcjQ5AW09dK6b8T8byOnnNccEw9KviBSeuGPHElUcIzmtyrEo8MAEthgaXT2
BDXBEmH9QBFZo0r7JCjrSwsGCVwCcKnz+lwzzysdHNqycbXhDIo/q3s/p6J3xtvGYQk1ipMF8PKi
NSni2iW9qWjp9c3RzJ1iF3VR+TLgotc77BT3QcssJrRBXtudieyziN3fdwZLqUJH4g2ffGSzp4UW
nB9ARKXGrmOrMiq8YRVMkiPYCJdPLkkmVBdgwxIt1bgvMIJWgnqlCXxdxccSwtpnlZA2VX5zBmIZ
xvoi0UoZlxmI3QHjsFINe4P7lFylm+8kc2V2odcenW42NlQsqQgAa5q2I6EuYo89wfoJ1smc/hJN
w2Nwa2zpSukH2ilVXkGJ/hsczTwBM2TJ5caQNqsjzSBb2JG/YH2HxZ6+3YHgYSjTHhvW8ISD/0L+
u6dD4KEluFsIeZQbk2bIObsINjvEHynDQTn/TBfprxg6SIkrrbw5J/ZCXqI4AJbmn+K9igTpgp1m
XAblqCiracugSEmkXqYg/CfVROYQnAbwj+eFNjebGxccHCwwMlPjVG3Mp9eon8MspylC7IpVwYaj
lqc3IV/csGjoNPXeEJlJfXBQOeV6PrJjo9ISIJR6U/4ZTnV2ZBDtR9OvsYf/KecZ5rF6QzoThepF
aGkIsVbNa5Zv64mYCKs2M382rtZbTiUI6/bSGEIAlXp3m6BSmg6MzGc1NL/RUZyWHfNNZDvITvDB
96ya/jMQSu3cFQhVYJEkPwnjMjORlGoDdar2vlownkCeFplj85lJbVqqCGLbiTCyVC/lnjg2jhfY
AMTVS0tb57XzNjyFS+j4X+mtFvbB/Jm0EcYzUeLpa5514r5HPIdXscrDek8XZw992XE/eP1RVL4m
ZtskM0Q/491P1SfTfP06ilEJlZ77o7JgOUm1mx6MAZy/7OyVOj+YH0+7Fennu/OsFY2IENcNpDhg
2OtyftB0n/Pb+T/iuE+JUjuv1wynAnpi9etwa8/roV1SqR+tWBmvbSCbicCmx7sqagOQ2jReUVTr
5e0L+3Naake96bi5r96nQYnrEBsTytgp3ozU0U9lOif8oQHhQdaXDLWhKPgxOZbWDdahEYFYV2Yc
uJejjT7tVpRnPaR7m6PV6u/UJZmt8FVK6GRO6cFpTnfZTEf788aAbyDevG0GDYqm8xU9LntUUZ/R
7yQ/V/m0X2DHHoMcN4npmkQ27+Z9tBp572DShfTHnKtAZcXnnlDLrLEbyTqiMsxaYnHEguTFHS4k
r7FjrrGxswOpAOzb1MeZvJBK6/pDeOUwgztuM0KMjn/xZzwk13iWhVCCX9NKmYmZKC2qrckMqgSb
NSr9q2dAPU8IyC98Zs0sPP3LYp0oBTXCoNoQKtTyezvUz+ZAfVRBHTEzhfAkLo/zgnuLYvXwdQvk
wtk2mecmmfYHmNGkBbb/WXmxscK8HH2OK0mPahsxDOek2hAzhfuK8pc7i30Xdyst7RJlR5bpFCcj
GFq0OSooyquOXhOnXIj22u7ZVoG7ULLRl0A0HiGUpRXucGk6Qg1eMYw1dj4TKH3k50dXljNV6ANB
JD25LIn4AR5mXXQ8rKSqCzUbJ2aG33udqNB9RJz2i+upBNCmKHPMZELiZDIm3tDck2newnxBYh10
Lkya1xzzroJDGTmiMTnLD4VJ0wnabVmh67/4Lt54nUF3jf8fWVuUkGnirXJJQ2P2Sj5LrdecUXjk
0FWr5LaSBSCKgZ8zVabzJNevn2BT/J3YHOTnXiqt1gNCluck5TV2V/9T2xfuz3YIOFcRFwFTuRIx
MKEXsFkM7KPrD25Lm/yNdxZDb3E7Oy+MbZslvgxSfq+KNwvpvyhH3XuKsm47q+bmNO9NhRLAVisT
mY5OzwuD3cCfJcPHJEDilcStb9quCXkMzm5PFtOGBsANnRXO5DGzEG/IKcmhDbs5E1udlePEwWF/
tLaNeaZs0Ull1CPokwSLpTVkoMZWgOAIKtN2Dhip9avl9Kpc1vT5Rq2mhqo5B8UfMR70VTGa4pYs
20NOokKGr5cBaPeObd7sbSyWVuWP+lsgpfrZfk6e7d6OyZiE8w4UlctohJxwg+NhaLBUgC16wP/q
/8qMmkwNUBd6IysRpJ1q6++814LFIxPXq2eyd1pWbrN9hEOfAFwmO7+Goc/kznhFXpR7MR3kHSJP
QE9/62+B5MoYDYspR6s2r8uwLEvnvCXf2GwKM0C1yXg8iqFgIiiwoa+zZwwGvsxiQupO5qzHVekg
iJppbFGumKpUfy05j278xXSCHFTmXB6OwKhhuEgwyvVUVKvDIiSfM008YHHBZg3OJHaxyVxzN+s9
txtbOR2VfhLCLY5fBkMrAs5oRyFJqGwOKR2jrdq5H+FZt5E86pXHa8LS3DPbjJTnVyE5vrmJUlIH
l3geopOpud4AkDq7Ed1p85BGpHo4R/eHThyGhfMVWaoTjknpzv/6nA1/W4qdOzjyG96OZZud8wcK
tMOeLSYkuwH8KjNb1zORghEXgqgF0Sow5RhsTY4fKEOsSKdhosruVJMdAqCB0oyY0OFOHXcy67ba
ScX2Mt96n3N0mfUf+4NhQGnpQdiBJdTGD7uxlvZBuEYzDxkx0lNa6SIMhP2P3+4tm9yiKTf95kOx
LJ+MKHv96xSaYMe1J0mzW8m23plkSup9ph7a36BfTQDeDIRe4OQZR1LqVlArexocoxzcnbmaVXnm
f8zR1vk2aOnBtDfdzIZOWwRAhOi11PVOAGd+cOsVYDzKFfIprDuvZw52TCUa2hTrwuaE8ujFfhm5
zawsbB+nSWbbn1ClQNjNPsvq18IR1GD2N5iiy94A915itAHnUk/dfy0lWWe8mo0ICYkIm/tMtK9j
xc25ahou+BG3HmmP5Wx+diqcGZ4ghhvTk3Pkg8+SweQM91vhrpV6SNJLjcMA+2I5ryeE3QlLR9Zv
i/lKa8iX/Tlis96BuxUsyJl3dK+mDcC8LYS4FLPAFcVJe9Fb/t1aAZf5UmqLc7fuIIifXySUveBW
cVj075BABPzuqHHkdpeyJ3anCDFPhIc8uv5ksOFgRSKNb6W0YnBBdswZ4LFxwjxl2Yoe7svJEnFH
oIXyU0GeQ2xHmueetAruaOlS5v/20yPZjvgtOUF1Y6MOC1LHK+eAMyaeEOkcgiiuh9ZB/6wwJug4
NjRSluQpE22R8ZJMmWFGAQM8pOyPR/Ykv8HreWEV2vKT8uHTrej+5ZZTlXw3cb98KqPFBAGZVG99
0IxYp1KrkCIehCE9eOVZkqgLLut6NWfEYpEeLCbLNkb6i548AVZNb++45kFstmAW7URT4ScTrvS8
HzOk3YsadpURq4n3Hi9X14pHhG78FDTd8fITnaHlihG1y/urX77RQJWcewmPL8v+qQRahIBhVwy6
g64meesjh3zDnP/MhrxGCF07Ct3dsQDJI3VC8TQ5HhS9WJrTPlLmuMQNTyCN3NwbMaQeGE+Yl5t4
l6p8mtC1RymUcDB3MVrc3l+Mbwp0u6Vnx25kGQmgKN27Xfqb5sLuIBUgIC1KbxTEh1z5HeyUDV1w
UNWS9CkQc2/U7T90z01l+Xj2ZF+oxrwDBlgDzHJrVRZ6+di7bDazZ4oUK+Sd2FubuEEt5FD6l9Pb
OraNXvfhR7yYTse/pV13ZyHtrD/pW3EWogMeDV6bWr+KuMG9Ro1lIkJNOXOPfXmdIbETj9NgM2sf
617Yfp53RuRcjwy6+ozDpaSkKZ16yZAnCZmT5x2MbgZ9s+NZNIXGyWPfhfIUGrGHWCx5lj3OC6Rw
q12sZ9La0L4SvKJht1DuTJon/AbAkIRMTGn8rngUnE3MFo+qMu+eXH4F/lod6SmCPyUgO/echEV8
cEpSD8/b2vicg1assEzr+Mowk610eY8lxACWPVD6iO+FKlROCup3lS02noZ1gNEM6PlWVZ9TouZi
srS4FDdal1r2fDmcpDj8bA5yDhj80NC9Y3Y2SNlsOh2na07IZQsNdzqKMUJ3L7JxOh1Vvg3GfkPh
ClppP+XTqNwDBV1UvcgvrBTPHLRz0vzYs+PBLcTCXpmEd/NNLKq9eFDkqfigId/3edc79s8yHhR1
oGhGXP4tH9spijlLnNGrnFahYg5sLwCap5fMsl2EMsRP+N1u9hwuOEQ2PkQ0P5ngPsdNh6r5SKx+
SLEQ1/WcPDGj/R0AmJ5rs4taB2b4zC9GYQ4kVWKXKcon2atx+eSuJtobhxOllakfadZc3LXHFKWK
xXtLUIW8VnN3rsyYsWXlys99l5REQwkESA61eVzHyMqU326olBgALqsrXSb2xTP913C5U580Ml9U
AgNZJIqZMRYCjTlIGzgxTue/ShnXzfl53cO7kzZrAKcKzaBngukifIkuCo2rTmloGH3pZuoPVo2r
2iAm8iYuuluLxkvfP50wpnD0pOSL/wvSFpoPHX2347YI0yUPi6L47uyrYH3b02+7S0ydxJdOvdG0
Cqmww1YvCJ1F1EZQv1IHkFSHYGrh+aWufVdcVHPSNx30RbWDjI+SXN77saDmgZizgpUMM3BE0FjE
qUYz+3Fzdom4OL3J4RqUnCuJGpoFncPSshliYiZs52UGOWyvRRappDAL1OJ2DTFbFgl2KyqamPuL
ezx/ChjjKDv2WkXqV7+ILUQFb0wCiN7ay8jorIcunKx4wrj2NwPLnaCUbPuhhM17S3C2FJXI6d66
pEoglwfnwgvHNVIdvY8+XiTsU+tEZ3rCXgyQbUNYaj1oTQjV5xL39YjI86MAcx4AMGpZ5xpQgJxr
TXx9qJsInvmN71bFMiRxKK1aB34UgWg6sXB72jSIoh7TdTuFpMrCUk0tr6uRuYm1Cc2QHsP+5xJ3
eunA2jSIpRimq1Trm3Fkvgqk5egPcpLy4uf6PFAnwcDXWrFPFF/NPtvnlh6OgoIRMhC4UOXmY37D
zVqF54DYxVs9XcJ6VNF5hysVSxdrT9w7/kIEcveT7ucwH9kr1HiP6VHEUYShKNN/BN5FYu6E+CbT
sSaw3LzHR8ZGWaLVGjFC/lrGuY1LA2vyBVw9VQ3F4Kt5S12mUnuzEz0nYFEDUKJX99IUyKyoIWtO
M7fn3Y1d9+HhF7hwJMiJpo4OL0sfVaHm/KxDC9EvhrNIh3DCm3jZ89JY+EbB8lBUfnCyhLUC2eOr
WoSroaVFCzAePX+WVvBChZd/ZW2hFMqcI8oTh7puHuFh5zIuKIxZA/XG5cN0RKOZPrNLIzTp/9hV
8ljYsREQLR6hiLcgZRhPa6AB/1oRsVLbEENX4afYMCsLS/0C8WK/jl2YW+BC5l5KkkSRBF/YZWOb
W49O5CRuO7y6AEtprEb+Txa4I8QaON/qduMxFeTd2YBIjEsEeo9epkbSNhMgpQB+8147n/USALVf
APxHCO5Sm7pdv2MLeiWALG35EO7JFnc/O0wBfmZQ9+N5cls3B52cKnyAP+qulyCuTeUCEJYbMuDM
GAsGL5kP7x3yhA0iQAjCfitv/Q7wpxk1qDgXo4z8P/gy7tMbnkkhMovwCLepcdUGVXcBELxpC301
oL5OMLrLxQMbj/HIk/z5WjUC9k4gAgTKSA71daZ2r39w++QqIN2FNw2KZVRhn9hwVtUUvNljWnsP
53jHRj0Pcr/sVZMD/Q4OzUpcHjxoM87A1T3CXdg+FtEVznHs3orVtBgAQ2LfLUgxOeTedUfriNMb
JTgwFtK/6rl72BaknENE7iCwmdKaN/94znzIjebgEyUpNbmWIHciKPPyaXMyW2kfSF4AtEsa7zrH
3BvZ7lUoTzRLBRBuvdJ4ANnuorj262ureiTCDPqgTQem7vEd3gX+XFfNzp2XQ9+3/zNf8XIpQm1Z
D1gmcxIe2xJToqS17vKCGSFs3o4pAiLOmVbJpTZlndND3jssr+2izW9n2HJ5FseTcSFD869iGXf7
S4TvPEJ37s1OYBcHCN1p1IaiolDPR4wpVfkDdFkfU9ByFKJNT4RcHSW7u1DHFJCknhP1O7upLbYO
S33DlLCMAKoAjENTcOKcDdyEx0vFZZsPrPE8YCTbcaF7GDPILTyWMf1pKP8HSri80iDo5vRTLLjr
eyxbxBrHlOANWmj16mpcylQrts4g0OkoL7LKgcOym0JcsAnkQ8EEC0dyb4HcUp26GjhS+7T2OR+0
aq4wLZ9Ba13UUUF0v9YXIz5I90SAUjXsLU5sUXKUW8iiPGSNS+Tka4RcFaTj5aRy3NUtdESNg31d
RIZAHNmSAZwOGUZq+SXlWScCzMCR5VRBnYQ51jwXe3URcIzP3GAu6kdtenaNOnzktlkh0Ykpg9XZ
UiCjTq0Uhf8Liwat1v5C051rtj49c6Vlf67ZPXy2aMdTy8SqAuRMzDCVlXRbRO0UyHgndf8rcFKV
ospa7i49r7zezTFJ8eG30zKR5HtQa1PJHG2CwOR5sTwhqKbOvtiHnKsojhtpqKX8UXpuuhtzXhsq
kly+ThICU4uewOZTiGppkRSof98ze4/xG4NA7L2DyfpSesf9DeTmT2IRCiReYL0J9jVqq0waxTkj
bHdGzTazQBGgBZ0mDay26xXwVo3vbRo6Bj/FthKkArpmOFK2gT8zdwq4nrxyYnIfmdCdeqXqbhh4
zIwFn9B10bBwkaMGx6tIUAKSfxSq+mBcw7QB+GOWQBjJxZlyaO13tW8wHBRdhrqiE+zv/dMy0O6m
sb2rZTwh92QBtXQnSCB56fC3OihcqGHbtAXf/rWRB8vhdsbL45A1rA4nW9XRLEvOBKjqCf1ghCDr
D3SqVHKvqgf/tJ3uRE5v4YDz6OwObDLeGsIJhduJCmlaw/83S0JpV3sBYjwLr+MUetpUj7K77Jmt
ZdLXjNKLmoIr3hz5l+cRCiEZS2wRwTIo4BHDOCudGBKW9UFLowp9SdAAbBsDkkiQg8GAyzB1kklc
2L2udjM9cyXMp0QM9xFBXOHw09+5zstpEaL0DJ7mAZS1vIXcx2wBWP2yBdoerSPf7DdxIoBfHW/n
vhmC00j3yGqtMWOglY+3PmoAwPfav3F3eUegZZPYTWjdmZc+htOR2/Yeie3Z2bZV5vrYHFGkBT3X
dE2lj/aHzizB9gAV4/N7WbcmTjLIiVfe//hvW5qRzCwBObyJrHHrU9eP/1yo3d3dEV+7jnl7gCcM
hpcS0Znjicp1tjB4p+bbW6tkxBHB/H9wGqv2JF81bRSiINM+qq+RP71hrnKFyVzwnMlFbObY/en3
mx5wC3nQ52JiR42/Pstda9ULmzDSRXTJH0rchtDpgkDj+0y2wH83HduvDMLTH3iCnzeRW36ti6pA
bhdjP3g834KhBe624VY8p8/CI8TygjHUHCKvgJIi3iY+2/SByBunsUpdQHMsUQ59V+HaFBHkwtqw
bZ95s3lwDWeVAuUm6O6rlkqIbp0bM8fSSCwvFcV2dBdW2KoLAcZY7mt/v3EpQBSQfPuAu3673uOT
e4qqMfJ8BzkpUPSQ5wISzpZAgXxllf0VGFhJ1X2w8qGWrGCqeXlHVvGM9BS9XvfxDHGBbiv9a7WC
+11g5R3tuyNo7CBHCU4bB/Lq0lCRjpAd6XPt7AeCcToeB60PzKm14Z39+DMw3DWeNrpV7GisquBl
tjjMv2kkMkyOVYfWrEHrclHtBh+LAAHZOX9stnyZ+1YXQXA0rSF4TizDXd0TDgAKuaFXy+vIij8j
0FsuFhZSV7BjYYjNpE7Tt9KzzsS4+2mVdQ/QasJ75QE6nJUwcybNs9tegolB8H6PiiMDDezaT/17
/dl5zkdccBnvyDaZehmEC0eoDlVlVOhJC2CDfrMTmBQEbiLIblzQBbFL+Q3mJJMD7F45GGWJU64j
qMHXnKgDSO8dX/0Vkia0CpnAkJvFPCc9qZBhMGY8wcJibFNusVQJSXKyVfYhZMJzVlt1IvF8DEgr
BMH9mYle0PlF+LX7t6dxfcXlS5kB25TB3+0L5q3PlxM8XfMug1CBMTCw8NzN79pxtBRQlmd0jqzU
2ge39QRC3AMqfnbBldW3o487/Efa/aZBG1hqmRBEIMMp6RIn2GCOKklNYiebyfW+fckoQfeSj3Tk
1U87eKetaVnmLmCzWu5Fs42YN5QGAT+YmDQSmz3w/LS8eybKvfi8vZ0CXVRTwAQqhsts0Kw7g2Yc
UvAwr2CCL5L4EtO6q35GhQsbqVEveCuRwpJy0+gLTfpfjd2vxyKeH0uXjoyhLmvtp5nkDjbxd/TA
RU9ro4IihsOHc7YMb38MQdbvEBTlrbcK80DqDG+fjxzxUv3RKg0hf2JXcfxQlc9v/kvmyxIVXf/v
Pn9gDPENv6mtWVkHtw5uiNLicmCM0c3MdZDARYqWmMkEwLVpGSWwdXWQkYBFtye2af7ysDp9pyPZ
gz7WGxGt91GNkJQwY/+VWlNXihhrCoviga1EZ9K/f+Ac8noVDD043kJFCOw0Sm412JTLjwWjMZ+r
ddZDaPtr6MbGdZi0hzSuO+N6PxRnHAF02YIF1qikoDvS6rT7p8RDOqAuFMnMb/PCBSS6oqfFdQcP
3SVQpFFOpbpvA1pUql8/YCqJrH+fy92P1uCvbaIHj/CEGmoyafmcL0BYY1yF5N+k1KgN4l0abBqf
ADTAAThrG6MC1Q8esVfO/lJFR2dj6jYS4TMD6aPrp6+M/ZwswpSWgtIgiF7VXJC8+cFYwz0soc7e
DEX+8hP0LSFAly2xrwv2Gfe/6QD+CqlQA50WMuSI6NAPzB2SckFwZa7XmjIt+WfzUYTrgbzVPl6a
DF4LcgaQWREqSuSKDBV3/mYMhCAgpjA80GaVNjuP4t3GMMqK5afBBm9S5JMYb00v0yOH42ADJHYI
ERtgzvyi0/cPsk1KRlvlRIKhBsRhQAXSnHv/UT6nthR9D3mXUC35Z0Qm4a0e5eNuYcFEHXPbMt25
daUO5S4ENgSQXlv9f6jOVQoMcjWnLYC2Tb0ZYSZdsJqnIoQw7uCpOMz4c6rtB1f/G1Q1neTdxnL9
ngAbCTMxvwgZ6i4jubaBRdQBmIxg1TP+6gVgA2p+uPnacz1gFqgGYDlg1Hm8XJTdrGL01STD1BAh
HfY8vJv1/FqXwqRqqmeBgqeljHPzq4B2RRkmDNVKxBvgLgOMcq+Irp+sk/dOfVZRdggJfbBPlpuy
KGL6tYUEN+9okub/4oQlOu9zURFFRAWCSjtAsC1mGSqw/L5F/WbHP8eEU9fbZAYuWot1rfhk9N2g
DciAg9KVaF4RBrVObCxuKYol/hmA45oL78CAWp31OlAougNGyqePOOBy8ZnXOHQVgjekNj1sZuLb
Vi+CvB3ddHrTsD51hre3ykkKVXeZselnbyvDqb5v1AdKfssvty8hW76zsjoHTCZt4fw38xrrSK9u
FarNuyxJXxhRFcJyLT2gjM7vfAEQtJXaLgL+4qvABEy084YMfCeD0oe5L1IRsr3M5nFzhYK733Kb
IkYHuUPBokxE+lbYR7k/MW/dzCH7nSHzwJMRvslv9+SOajO4/181ID4HfT0P+gSbj6SJ/el0g6RK
xCKfQidxzHw0FRJIMaFTM8g3TTK0oEj5AdYe52CkNGaSINJuHpbHmHGA8sp8u9iAbcynxPlPCxJg
QDc6icy8yoe1baycRIyyEE/qiIH7IzQmOF4JpyoEeG/mcH6i6JE2PQUSPY2Xfngx2ivTalpV/0Ti
J69j4bJwreqMqHyduxZPfYgKhr3ezq+VqrMOuCMW7cwwsnmsNzIqFcUoARjMj36KzwkPvEqngBK1
3d43Hyl4/NYwqspEItYFccl76N2nHarSe+kbNvF5qw9dG+/2g7CpNPj2JRza4FItlHnIF1KM1u+K
CL9om/VTSExwCBqBHJ9RlGN4m0PRMEUi/ta0nfhH0FygrU34bos86uiL7eBYyAPttQ2I5AHjKbcQ
8OWMjs19lVIwsMcvbTpYrc+xpWBwukhadKlhFz0tS7MV0g8YOfYo4HxWX5w3luViThvcdq5tz6PF
/474bQeB8waXgt2aqPUr9g8cCY7KvGGUm/8dI9GE2poyTmwNJBWlMK9hFGqde30tQ8k+doy56Ea0
qKwF3ULptCntE9d82yefe1u3nKRSDivhRZUHdGDlVD5rmE7s0oCRPNkq6Zsuq1HG8PMwHAqq6C5D
p+/kz/0X6wpxVprXN42cbRSnxIliPn+DsmsZQhL0V6H8vIa+SVdqJqQPOqQooCzye0brNMXbewKm
144579oYaB+YEPbSXOYYu9BpDAYzkzoJly61GNi+N/j3scCFc3joWOMehhDUQYsWKnbxdXF2PeWZ
vRBTPcyShGAvYXbPmD59pfyCHUGs3X6peqXxqG2MX5MsHbPo49syUkoVqDg/F2dRV+ZjFoBX9s5I
r3svkrS6xz0Db6MYGiRhNt3vsypJ4lX1Coj/4VsmrNgip+F87QOveVcqHFOLx72IkURdRVQ9R95t
zEzmIqmhovJdB/LV+sP1C6XUupXc5Dc0sl6g3GMNlTb1tlwhcbhq8IwkiQgz0eCJTYWWa712aolS
UZ1W770j2osYJ1vQMk5MlSZAJnCFNpiEmkxjnqZZfjWPfXIc+7RsLC0XHkuQZ18flCMubgCMiOZ6
OJPh+1xgO7sQKfQQ6szfoPjjjXPFg3QzC6RUFkLGRkfYVzN2wM4T4qVrvwSE8Uq4W69DRCha0GIH
GpXcaLJ2TvjOx+dLN2FN8MxM3xgnYG/eCa6Wz1itzl2X6DCvYpl+2jBeQwSM6yuIzpvs94z6GVvD
pHZHvnfRxc1nhaDCiCa/kayaPt7hsBjAsFyBHMpmAJieQL5wmTDeXwcF76eS+f+8kjvC0hqbyHOG
BZVUiqps5Nbs3IZKHSfPLJHryNt6QmcXnVC/Vdcw6RwIauzNUfKIXFLW6Itkot8GEOIDHouG6c00
Lcj8vYw1876p5ar7+7vc/rWkecLeRLIJeQKIL+0qzSX93P6BWywCmxo8Zi+7+LI7rvpDucjBmZFS
Qtve7vDNxrAFr0KXdL84t+qYHJnAPhxW3TJ2LMggsCTOq1HspP3JR/Xu4lS5md2EZdgv7zV2YntW
CDLE57BMxqsdNyxlw8S/09QOoypK1W0ZuCauu/TnMnQNQWDiSb0gM/yVrpEzH1867Z5c2Co1ll2r
KG5TNlgGl1vsmWlX4rHOcKNdOxmhjkwEY5nctp52v+xrU36U1iFZlyt/emviJa2ZfeY6dd6IJFEl
212htRDm3EDAz6D1hXP739AFSWhT7j6uaPOKn282Z3ahsgjPd7bs82Gvgxnj2gdH6xAQ3F0CMKd/
ldGqlX+7tof1TAPilQzePLr2vMFsiOa9VnWgNNun4JMsUVuIg3aWlh7Kfd5u7+3n3F1IIGSxhGP7
yvRk5y3trtkeOPxuer/NeKZYf8DMRNhn3mnzjG0INCBXSKSbTPSB4bB6Aykscwb+Lt4mjB5XQvXJ
7QOtxUDz9ZGEW5T4YoM23jR9t6xOtaUXRXoVSEScGXNLLZQ9cfr6f5optk0h8xnjG5U4MeiTWRQV
dfs79oUHKwS+fwYOs2Vp5AUOM2jswDWKUXv4tsW7is2pXc+0LU9+W5ll2BAFW+Y4LYxiplZP/PJL
029NdcHw7ARY1WkBZdlrlwpXei/5F+UCl6LNecsEjntr37Kjc4cnJ2TrCkVqCo8k9kMmRQMQuYZP
FWAP5ihuitosDUKBZkcnM46lkpo6zcmM4oj7+IySwSQrbi0Fy6Yh3Ypp2BAQz5JdzIfzalKwIBlN
BEoPtSNwoXM4oqF7xfbtiFtVyQE4TnY0mJ1zpBhiwk/powMZFr8Z6pGi8H6w619HChQ6oIrBTJWd
+cuxPgBXpyZJwggD2l9atUzPB4ni81md//sIstFu+arFruVJPMH4XzPlAo2Sq1VLBWRNS0dfphtO
KdwysVCFgxbpYIedoHXMz7jTJL6HHgC/awgwK/S2PqMCW5PiKspEPwjw30WE3yQB3763c2+1uI9l
jmMPC3ZeXnOkXL+n10DHbVcpLFqDZuHTQiqY567fWUW/MGodzbGSs+qD6CU8cZCxtYPUHgXN/XIN
CY5CO92/i3mw3u+iYbJ3GOZnoCR2tFYsgJ/ScLnOjtYqHIpqlNUECJoX2QPOBBh0VutKiKhi2SXC
QdxxikDrkrhuSMzub3gb5ak+1v8+bhWBqxiTMDIXbKF6AGtISUJ5fjts/SnwGpgD0oMziRUeMzoJ
bC2Q5GrtdxawbzJLgdtYsnnCPYLtWcnZIKoCp3ZNuguBERTZGKWSRZJTxkBnsCchQzNXTow6LR1K
xmkl7SVkKqRJIETME1zEcqUvLXmi40gr6FSMYlFSw9Trf/P1qpbZTVM/XKzgkq19P2LxmV9f0z8c
rkeqXJWr8Txa7Z3qIgpokHniHmQWYEKRQFCbQsNCWb7k18VmxpSdBDxKSerInHxYzvVQqPkT+Ni4
lHJZaiDLCmp4QUiqPyYUZi52VCwoihag+Ome1jgDm9iM5GlPaLJ60kqCAtvfxD5hg2fLq/JC014X
J9nFca1roLubYuAU+hNsOpgQHYgma9QBlJ4NYY9NDAcYm+Hj/7F+SZTtVPD27QMQlG0NgPktZI+J
B8e8kHegtVNCOcoG9RKaiwLKncrpzvyzPBK+nq069Ye2EVKnI9SsMV7yX0MzcV5KNs5kiEe6x8FL
E817ufzUG/W9WbxDek/7rEC8AUKxtd77anEFNrwvhTaPDLq52sn4o12OHbfp5Lp1z0AyzjbfAC4Q
JKfkIAj3CSCrRP+7rmZ4UVA48jlWRJTzOGez2wXstXLWIWrRqqLRw3ocCtVg+6v/+XovjiGUcRX7
3ESXH1LezPN3iRtEMpdggYadceQUMDQnUZuxqMak5XYEu/8gVTy05OvDaI1daBonjob+GjBs/xGZ
E+KEKpU9WhUFdBzJKAvMnYJnQYvrhj/nEIMdOKv8sd0YO/7onkMsyI8CWC5i5wzT5w9HCZ5hBE+j
MD7gBwZ6Ax6tVFKqYeNA7S2kDcD7Ex3FZ5MaO0mTO/IoyjdQaf4vprCJcAfBJt4LX59C4NCeh1RB
j5e0gqHHHKSguoEDZotXfrVBIXLUoIkwyqgvCoFAuylXqky2P7WCK6XgkM5D2IVDLLC2GtqmJZuH
AMKoWRMP0YwB9gYe4uRtYvMf9uHMyazD0kEPtPTFTdTaiiGiPSTPHJr48+PPtnu6ou3wzgAmPMt4
9xI2G8ZxTcv9p0Psoiw+mAyC1vPNJdXcYKEHsVYmMNHwP+9fKHJrxMLKdyL9jDs/pU6FZbGLvlad
b8WbE2oxirydVMGssFx+Jm4Y6j+914neHMrtmHWErbuLSOB0eHjmvNDDB2AbVElF2yjbd5o7D+Lc
u7jXb5/U/aE28U2I7Oub/mCUZSmAx9navozJn+/YB7byFEllMecnpTHh+FN7XQWG7JvUJInVC319
Tys1ijCzl5d9yVCW32ufulBHbnsVX9NWFgS6jMYycvQRzKQDeKt8MgEaSWmK5npdyn4V64l80uYr
GuwEBp3EsgcFTO3hVBWhPvXxab+rOEgMtj/UC366l5kO8WlZtR6kIHQ8Vba0hFujRzsMDZ4FK0Tu
QUUievi0UrstSiIZpgT50oH5hUY77qoGECwq1fgnRkj625MPqZU3UQGcNsW84NU9+qOVflP+Bqe9
EtRZ8IblUlwF9t9yFtGRN5/Fqn+AkxhPLju0BkzIrRe25OV8N0STLsu5sKRM86I3qfihVUlho2tV
Y3TCaqKkqcSkbpmYkIBNp5R9Ci/4ZouZnBkVImBm3Rm0pqmbCoW1SFErsXfB+deON8jaPlDPpR2d
5KveSnCddPLIJEx9z/Jrd6t3O87SvcC6A5FYAtSlVSZTDhNWEhyrMMiKZEoYSNqYLl1MZmI6lFiT
IIGm76+lsZVP/0tpE8KmQMTRlvp/Qf8/fqVXc7dbDA5NQPMFhfH1K9Fr8GvYc1EX+ID8SOdJj6PG
E/Nh/8BKGbCwmhwigV+kEgBHUdFYxlUYbk9s37HCADwm19H7abX6ELVzlxy/x8WsNT3K5Ti2EX33
vB73w/acm+pQyw7j/IyIPmi/pqvOUA3C/q3plKsUMWiRIx/cpfnxSCT1pCSyiF5qU9F1u3w3fDEG
m8ckoa1toUIxVI2jUX68WquyGNNFNlVSAKn7ESTuXaRlmfETc5cWwWTMVCj+/h51BsnrTs/HnIdM
iNgBEbN+37Kqvwym/yaMstQO0KppwPBUkIbaukUqxlNIUDY42I8cP2N2LvBk+32DQd8niH2I8+lR
/fXlzETZv5fpwaHBHEaCNog4NBWoM7esn2I6qRwG0PRFDm/mEQsWPL6yonbvVYL0amnxIZ000RVb
a7gj4QgcDlvCkTfr4Jyg4E+mZZXzKdgEGidHYfBoJ4z0BAarqFO6xm2/8cyDqBODn1FpUGT7dDvg
1fN97we0qvF/DDzRMie+rLBIjtHvtgQm+VoIb0glmG3l/rOm3/JeRNRo9ehQfvnXfEH3neMlp3Ak
YFP+rzIreNBy1WsrDvU07UKviJKUNev4qzjAek+90BthvZHqVG+swNvXudOqOBi46IeiOBVcUCki
xkn5niIZxXjpOD7q5yIRR0AkuZhmBGCcq1Gkvxa0UCqTaBWbZGD93ADtDGLfJRV7gAdummeuY8IV
LaRDtBD+DmS4mPhch1JYgLLVOzqRupkRxVk23jZzPATqhv0d2v5fG5FZtSvou6xdpBumQptXQ/z9
Ar42VxYseLhkY+IO7XHHMJoEjt98V51OGuW4fU2Rd/Ry4NO3wb45fZFvprK5UOq7Y2EicnvbYZQv
lZ6FeYXK9lOHUud8qKSUps8igLG6qbXPTU+xtS3USR3QlM4QsTnwhewF0zJqesvqVhN9rrjhsrpf
bKyKFWzhUSnLkVnAdFEL1Ps9Us3BZhOie3DFqaXsqpjNiylDAkLyI3/bcMADqJHXa6gy7unhF85y
tJvvN2dcBv4pL2GZzLPEjDuS6sdd8FL8a0/vpojHgzti8vgtq+ERNnt1BBrJqWipnlWLDzzkMP3D
d+UDuC+0815HcCdIPCTQ/SuC3A4ly64x4pY88WCIZGzgdfR0eFZKGADMTmSUioPWBQpJ4CekSicZ
lNd80ETpzR9/MBD42bua5Gxvm0HoUbxJ8fS4PK5mmnZqFcNB44u/UfzFD+saCape1Y0hqgzFRjQP
77ENAl4BazokRrXBIj8eLQ2U+xxXLo9gDsmjNDmGhX1054+8DR6YD3E6lwmUxHNMZV796gdYZjbo
PE4jbdD0KGVgm5L6Ma+eqkExVA49m5lBL2Z0Na5k69/Y1gyiEUB5NNmhRA3BTGrFJ6dv5llYsFf3
7A5NhfFgIxPCJ/PT5rhVSdaFc0d/Y7M7Sj42r2JYShJbQJYL79LD7MagWeK4TDf1B5xqVv9yo0po
OFFFCjCRNeqOpL1t+lIYQV0hKvcHLbURGLpe271imhbQPHvAOHALOu692ymyJECRwwb4+P8aoyqA
LT7v+ADig6iLibEPuOT2EfKzFVZTRrnSXkZctuOx8PoYavFimCJXVn2O0GT20zZ+kNnu7cuG3USf
QJVAYh1h7UP0Bhk/pbgkdmbvGJHcnftp0DOQpZl/tAKYaQbLYRF4HV9t86vXrV1fmaREGZNb+1dr
nLIX9EY1P5yW/1ocLFuRfo4I7jz3mDPI1vIlUc2PoJltE5Y3Pm+poBkZPX2bu54TeLacz033vePB
2Mw5GlNIiq0MX9LIJDY16wszFVRSuPYxX1+43Z13yWuvnOqcVNfSucnrV+xfZTS+gFDo7yimKfCN
3TDzVNam21x1Er/vo0wxvHoG2dTzgkpt+qq3lG9CCe0+ALaqo47nk/4ERF1EOajWFVzzrjbHWtHK
QPSsSWgM9q1/AEc5+JB4SnR0gXlaCDSmXmVDDVtq2FQ2FkcEX2LGin5DYuffkQ7VxBPrSjHMI7fb
3JLC/qlS5Zt679JSeijr9PT+FmqKX+BGMzReXMKiAZp8FXCPL10Mzov/LLg+2Mi0z8L4+qWp2TcF
vvVmY2drL590G7xDKls+u4AQS4+v97JozSCFasm5WxtVD3wNeSwrrTuykw3rvPAbJVVIWkq+idNW
15YTg0fR3EPJ4hiyfI7IgeO7gUQ6+v8TISoXvxJsNqUKyfYsEhFuyEznxNw3ZnrGaDRdXyPkudnb
bPmjWULomfoUgs7aWYXlx0KIwq8f8rHgetOf2y1OASlymtBjpTuWPaVVDT8aIlMSFvaj5HICTLKV
VGF5EHdk2BcDSJ7NEaVIU1nZFMqN8P0jabQewgB2eX7xrYeXmBUBQDizjHAzBazEEoj/IVaEISJd
eE76q3mezYJqj0zitVBtqCUwjTRirr8ZNGsgv+r/iS+AuPzxZEhxDToH8H/u5OSS/4KvFpk9yY9v
OUPtpFgKbRmOlVosFCyqlpCp1Pq8jRnads0Kpj1FIpV+lACHtPWS2W4TRc01nfLYXmv4wx9vMwkW
q7VybZk1/4oWJHa/Embu9HDowYGQzq4aHP2Qp6aCFWoDeLhbHrIky4TEsSXpvj4Gvv0lqkoqR+91
uJ2FERM5Vt/OM+Z/l2En2nTdc4M4kW3T4MpmB13OCQPqpxo6ysWwi07BPzvBfDkxB9tLW0sj2anM
q46zIIALZGNrAhmS/m35gK+mkv8H4q/fmUsj/uEpjY2iUC7ew4cIsQsUkO0Z3RxAYWdW3gHNzNSK
sToePHIUTBWY7ZZ3ovT4qeHzJgcsFMRTjZcNJLnlSR7LrUFErLXhjyVRc9uxXbzZWAq/3d/8RbR5
fRVzwa6OcBuSRALSB0q7QjGvRUIaRNpIjZ+Rc7Lj6WDXMWvPr2RkPuWOlyXwC4ujVc/g+wUdyC/G
zhFzhuCNXRZFz9VGqptvKXSxmUz/NUMfnr9YrR+85uX+L8BwfPaRcCKNUCbfErMv50w42GVIxRx/
JxVSR8lUZKHbTqxq+8nRVmiZik0WROxA+fgdVhMdXvGcl0SLVppL8xu9wKyKM1RgQspuT9eFlMMP
NvMPYfKie3SvmE8vNOvdmx7MdusN2ViqateNdVggDRHfJykh5xeFTS8r64sRX6gLJoLVrETOE+SZ
oXioi5uiwAwZmPLmCk8K4zlcoEFZ2+VQ61WWn5PBfGqjV7at5UW6IrgpbToN32D9yRnKe0miNyD1
Ry2GYOkkMhfVKpKv0I1aVGSOA9ZU8Fmfcl9FOfZBxTuDzY96w44TrqvdU7rlahDzuby/gtSzBcuA
63TM2cxoM1alAdc5sqmU6E61vk1DutoJYm3oonxv4EjLW/y98OFY3L6qsV8TeJSMwUIcht8jVv8P
iEUMZryiHYyp2zVOItmmuWMGuJwozFG3tj5EFKxY6lo7N4Si/erj+5q1cUFNssqZogtIZXW8hiRN
OMd9H86muyWINxPxDP+3aG94yhsr9DPRwqo9vg8FfwsoGQUid7aEJFM3wWG7pSB3phPHf9P6oWfK
Yg3nT1Sj6ErQ4/BDkTXD0fmQQ+y1DdvNs8g9pQqBzBL4bN/7nuOkWV8ScMyn13GEgolyVdlmJUZZ
S2+RcdCx2DHzxNjyt5IjgnGJwBzA89k0wRgRdiiCFA5hQJ0ssQlKF4IcQsp6LNrkR5Klm8YYAjwS
TUCKtsBO+AciXW/i/fRVO2urazMMkWD8OAK66XXL+i/M/PgenXi0PJ3Xod3IuHQDpZ0JuW0ApeO4
4CqN0cqZjlH71OOcwJoVU2e0HhUDGG+jLNGFj+DGR/9KaodtetTZk4aTlqKFgFQjTUorQaa8xYI/
8giF1CIW8UG7ye9nM4XuRQGjsrd8PRE9JnDBw9ub160EYKLilC5e7UWnWKZskwIswrTVFjYQOuQK
yNHIq6+dDbIprJWojV8NSETYtaNSrc8n4OOorgdb5W9SOpK2gvUwD0OzoU8YFeB//ii3nLCYWF4Q
rQP1Zh2UReCvcsl5X79b/xKzcOmlQw2E4/TOY7oPvKzn2F0U+MKmCbtbs0z8UtLVtgqDL3RKvb9q
cKZD//1+urxGBS07rNMlde1F353hJ8DtyO3m+1bbvECgO7VnpasyEZBwmCG4rFpehAcWLMo6BEFs
NdptsZPDLEdtT4SrEDmCxry1cXwEAfSyC/f8GDHSNTYjX2DDUgwOItN6D01Zw3hj7u54zIgvX4ph
gHZvUUviUnB4aA1xK4DTL/vRl/e2cUbdl0hwH7R3A+6Tgxr6p52Ed3NMpHUFV9AoeHta9T5eGkLC
oqXEPlvbJl3XGdIg8cJFpwZD4VANFryQm9IigwcmOKVC46DCiLzkYKzadBOhX/lvMofkLnx3s1Bc
Bi6w0BJEtVZGi65woIdQXKMVc9jMK/JW7Bp3qsvBsxdGYP1UP5SwkeHNp/jZMjXQ1mY2I3r3oVcm
lMh9Z399tgIMREe/vFIZTP10nJEEe8cqMroGhoyullTg8cJ6Hyic0X7DtkzVTLzHS06P36yv9j5X
mAUS40A4RgfzKLHadhH4Z452BQPc6jyInJFdpxou8ddo5iV+1GjIFKwua5LCe8rKBZL8hZsSL7Nm
bMoS1IfMW01p29ovaBC1neU0pN5satiTBzaFU7Zf68rG5T9zJ4wIJ8keXshmVVNqGwTtaNiAHueJ
s1zMX3bMouQP5frrtM8jp7klbynJbhdS5yClWiH0DFmisCxKJayqUwfG/94opF1iK6j/nDpx9GFP
Ljvg8y4ta2JxUll7eLIUOwR6ICllGPLy7L/em2FKjm/qWPTxprB9q+UhX8wthqk/OmgFB+cSF8Q+
Aq1AK4vgrM9Nl9ZjyIO98Kfx6gCKxi9eHSd5Qx83kEg3pyc/mhcMgnKwM3t/ViPyL1iQcavgnSLm
eQ9siPfJHnJ/3tdiFbAhiqdEnnta1YowJxru/B0jJBJ75LefyF2thw0CztsmjqDKGtfPV957+dwh
VR51eoeG0HlGa7Q6/uvjEweQd2kfIZDPbVUvcBDzeS5lKx4komFKU40ZHqCAADEmluQbAsYjawcg
rVZ6tr/1qMptoTY+VwpouzEvVKXOPxP0wqzfR9nr3lsCDV2AgITM34ige8SaUt5MAB+N0VAz034A
NdJG3dFt/ASyYfaAR1bOjpaAc5lljf68Hj0l4Jqc9yEAyr9exxKr07BvnlKsjS5ZmKm+TdtAG6So
imv9EcmBWvaTRncbdml2sxDFCuJKF1McpFcQCHjE/Y/p5q33Ub/7HuIGGi53dd+dF5dsmk2mvLpo
HO/QfgGIfgD7ctymZ4nsMfnmHiHu0ZrFR23IA39cdGnYAHoLhSUFgenw1g4bZJ6Kq+9DA98xbYVM
UaekCOv3X7r10gj1UkA/Zvo5lfHcgp/gNSVQWNF+iIwpPIWYVd0JOhXdV6A4qGohOogXg5DJOtOG
tSHs3ucX2Jqukm7j8gRyjBrcrOFza14qmysUPM5hFfss6D9/QscCeGIdYJoPnHmSlX2fbPBKoKT8
6iBUei6f0lNlSfdxUrcIcLYNFB2zNSBOxPjk/tEaHpy2XbteAXRPp33cDeyf8WHebacM0vB4+G7b
hCuh4Mt+rRWxPV0l3l4/uz0FLjOzdRHdmMnP6tmppueaS9J0jseBkR3wI0hTTYd7KkxZd+t8rSVv
jE2KbFnpPM7mF+ArOr0Yqy/LUefNT4eMmGnlxtCmkB6N+fiyiIcS6xGTgMXtelg3pxpALnnNHH1B
vWbseMQWATbqjFrRm3nCPGurtfjOKt/Rfa8H6jQTW86dRsW/GYACdg8Al5W4o/zHXjnDPFyvEla/
vInOjWXRlK8WtZkh8KcMGGjfKCczAJdmEQTnGRuTrQThCtfntl5eqiTax8QrqBw9HUcVg7lfZEhw
sSLPie+Rx4yPOWpodJsRWAUJ9G3m684ii2iSZvga1MYw0LcXPHWRPzmv7vBSXnPlncs9hn1aSfTQ
anqtY5J148k/tCctJRrL7u1pFIvXjpQlcsf4czO0tMGQvn4k8vl0qHbzUjLhN4e03/MuoOG/afRW
4eXroAkrH7gZwv1eN3cmX+kaOpstI8YYihhP+WGW+GGp76aUs9tzPN959c7fylptGShch04+/luz
5GnrOxYdauUaVsB9xIw7kimJy4o3K68LAJUljtAHwljpu53VgGLCQ414ciJhUj1YgtQghKs9JI8k
SYbqROkfyDmsIEcFPi7RaxffmP04MDpk5UPFFL/kcW3wBLOV7OaTWfJju75Hbl3Ihp3tZHFyl/wi
28OwSif6LPRHb5nfFADedFSElDpSz/poIzTiHs6LGBTj0VwQNKtcbWlTfBb7C7i0HV/emDdi8YBb
VnBt1W+rASUxIPhC763rokc8YXyMsxsA1Ix4d9Rfe9YL2RdqbvtnkpC3jIIX4QmFKdTTtDU2OyrU
GFoNhhcPFXqD8Y4hh6yIGU1tFTJtcrGruw6G/b8WhkvyeVS5BY6D/eDZsKuWqY1UslXwAPRz8MTZ
iSR0nYt1HdtgexW1SHTze7Ly8U6+F2xe8QfA2zJzOz2h0ALftYZIOzDo9gKa5e1Ai/mOhjQ5swpz
brL5w6yTYP5Y2dZY6vVnttj0uDzK2qIbNDHIWcFJrvMvcDErI2iKPiuBl8ISMs9uuo3AWSvsNJxX
hNQAqU54tNDpxQ5cmynjoG4dpDZOSKKD+rBGVLHdc6LjHizHLw69LLBPLA52Kbo4u4X1fO23Nn4P
Hvq8R9A0A2PFChvnPcfwFJbtApgB4oiH5sjx/R0E01/i1UEIRQsGEfvX4gZhv3NiJ+VI3kMQfq5g
QR2InFuQ732SY3ujx9xYPbIfp41GAIO5TbmvtIDeDqhMyAM/8Qur7CHrjCxEPi9N5ODEjBCXD21E
A32vy+2AWoc5nYgWjvHqGZi5WIvtiXaxzAc9OSF80Z71YjQ0LADVjRDQl4alR0rUXhi/1YZPHXy+
JXZHdjw6GONThkaVEQ2Ed1MG3yl7n+/nY+7kkkn96TnGQ0hqittcMPq4BGgzUNb6pDbHgw99VP/6
DLYzG7lkG81EgFXcuC1Clhkl6uG5rC287XRQmwdsB1673JMYV/yDdjA8V3bTrxSTh8QqmXHiL3Pw
AfOrLIpDKimP81PYATdOwDNw7/4vvcJDQOENCDcwmJaQUffXgAlEg+XnCgOqvQ3BsFKiIUyB7+Sn
n7ZJX5tpsDVqoKelHPVZxdPS4xyvgO0i/SB08oNeKePUkGOGiHmfMcSFy2s8ZlDYFhSafnXCt1f1
JgpWurhO7qtSaHw1w0APkFZjKOzQ2/VsGW7h2kc4bhBUbk1rMh2ZUK7oaG5Ccm+19yuhYXCDGmZX
m2e3VVWZ16D2McEf9EbqLYL0TqtepMhQyrYiUP/bBIuVaM6npn9Yb9agORNcnFx0b06YwiCVxgNB
dZ8i/adXKDQOzmOcxqYGjsg4Wgnq4psFxTyIcpzfkBRdw/P/kECa9iPCfLKxNAgFQBCDMeUg/JMC
LdN103ml2Islsgu42FPneeEO2Hpo+e80qTLtEVuk2zbWlyPISnqU70A9AkaO9Mq9B6nYLKm2Qb4z
e1O7l3bU21Mzy7Ty4JD1Lpw1skDgK4p/4z+SYk95IjZoMSA14QcEqBe6ek1V4EO0HeL9SeFuCGTf
+t9JZQV/gbdSP+SC2GMSMJoDxhl6xnZdAXi8q8atCsJLFud4FueJaTFO2M9iBwzF5GxMQldW4T+j
SC9twagFoGgRkx5uJDkdqmpI/JnPH0ZYaTXlc0eKHg/twLYp9nbsOSUDj50mtdhlYDCo/iBtE7+b
TuPl2v+8s36uFAyRPbZZJ/4qmrw+9sIogqQ1Y2Biq5slguSzzh7z7yoq/7uVA72e89p3MPlMOslU
iPyRgPAiXVrJDvpaRs7I5oxkcnh2D5UuU2ve7NogUlJFdKkvIjgNpoCZf2EK2VdQ1qjWQnJffDj8
mIowGvD9FgZPgSQtDCjnh3NL09l/vWLPf6NM+gNZJ5syIsfnSGV7NtkRh4hjVLGnIrdKPCr1bVDe
DDmqv4/mjlvrynIfHgLQUGoVrN36FRVXVtgXASR2Gyayf3Rtk7eM/CUhx9ignZ2roXo4i1xmVFf+
U2P+NgZSNvCmdz0d/9tg8w9GMaAftvEiw80oHmgPX3vLeILPsmVU2KCUNdrBn+7XtWkU64FnEy80
0YWSy2sCzRcL0TJ2wn6921dLuEifqa1IhSjGCwkRXU0e81UyAIipuJYsvjjHZrOyhPz/v297whWT
na4yGTDn85QXE14heCY8y9LKd2EwjzfcmLX0bN7vSCd201AB48MXQB/X0ip5JTGBI18YXCo9J+pu
0DdYnpCE0jL4i/nVSj1gWgus9axgEd9Kpb7fhG2z6hFYGCuQLDCd2DHNdfBhgIL4VtJriFGgOXzn
cfFEXIeMg0h38y2E+Wl2LwN6yRwitcMHN375D/aUuKXQPZOOlYDC3RIK7pb1/XjgRaZN0dCxufIq
nYmMtDctHeglrNwRcoZqt3qxFN70noqmi0PYO8CKvBmoO9dChrnPJdhiv7/peIOHiwUaXjvW4If6
huounMwDybEO9i/tWxdaGHgzgQmWm61YnFbeUO2orqC9zjfyLPeG5kBfTJAJU2SEZ1YaVmWkJNJh
mrBrzWTA8aW7dbHc/AkJTYEFJhVgFJvIqQiSOnBUXJ6w+TEb8ov/hU4uiV5U3R/0duDSDF9Sr03V
eN3E7WmRce+VWAJ/g6M6MB7d20/1QN2o9gRTtjfRe0uyHsAOb0iBsdBnI98o7Fut06wgQeqZ1Vfv
sgF6dABoopbafGwmw0RVbV93dE3HHMr8cIqcKjWsnJoNk5nWW8CLn7yNc1IhUEvgfJ5v7rMdpNjI
2UsswENdDGU77mpOwTypCclKvrPJifRIYgk8Vmv6+ZrSWLdwGqB0y/KxoOgVLFMRsPq7mGazgjVi
udRYhtV7VP65OqiXjIU9CGofjWf1xx3IcRj+ml1F8VBGGQUOYxHX6NYPpoRSlpXt7D/c5Bkod5q8
gUs7jqbnGTYI3oN8dguSnkK/ALfDWjjmjO+52caLm1fa7+uoFKY+EfguitGiKQBQD1O8R9dDbUMF
yPPACBxnfkFCjQZJa43k3H4zB/Ul2uO8h44VjBouA2G3eU09yxygLWItDnVtsiB5Ntw3j16wNNIN
lYIkTvmNvk9ed8D1HkpJpLCfFoBRelSgSd78fyUPY4io58UflySg3fFERZzihU3R8VFHW3CAkk1l
omppkExPeHWbHqo8zx+tO8ss9bYfxqsi1dZFZnOKnIKsj2yr36fI94XyGVWiL1riItxnvlUM+V1R
Ie+ODkJ+oO4iYXXfyqwu+41pCsQbDCiOrfx3/0OnQsCITAfkvZMOL2wIQPUuh0QPeSgqxo9fSLz5
DRjc/yy273tj92x0NuAXmDZ+hd7pbCKo0QOswiKEb5NITUIVYl5xP0n9+7sU766E1s8zSFkBOgml
KwMvYKmfmvgz/G9gdP9YGrZRA4viRzyny0WurTBEBy5sq8wy7oKew16eSLO8MHt22vjgKPvFqoSC
j31hA8zP1zhx6kKZmQVVkfZr/UVCkVlmpgogFXMmzMX5dYYtUJ2/qKC22CXF+SI30YO5KxA2LlMQ
RjAeeIop5kOt9Ccv41C8VairUK2oKzHGWh9W+qKuEDr3qmYztc0M4m8tyKM/Ygw4bi2qKglrz+sV
+YjHUj7/inF6hG2DtIyzKooVDeERhD0MAZyW/+Fblj8gjO5QdX226QKPFElnjuSh4MypkJjtsvE1
YtNvbptrCMjsUAoZbhVFDsUcXQdw3PTLboRX5idiC9DJDd+Pbz9JVjAIQbOzAOhFyBaZwKBq31ap
LRaJlvuQi2yVVLy2h0ufZl/MkXf1ZwcameNMyZY01oP9kBPkqqHUwseFz6pZGpf+kPiGICGvQpXM
cwyfoJ6Hi9OB+f4qD9Q/zF3Wy9Va2zpEFKEK/tBGK/YIMD0rMbI5OTX5n40UABkGOFR9t2B7LJTF
nxgJ028RAd3wjxo7/FU4yPJOXGxkSlddmZP3bQTWg59yK5ZFbWMMaJ09kk5V0kGHaN20R/eqhGHa
Med4qXe2iLiIuUJKZRiQvez95AxnvA4YyZr4m57GwU5qA0aWLEHO1N3HQOiKSPIBPeFBGkS2FbJ6
8xiaSzAf4jMb6GpLPiGfbOFIf6Rro+RtUoFs3aIxxeHcZE/yIP/4ooUPS69kE2D77MroCEyox890
QZ2J1w0Zvba3G4aNM84j8/oz+mtLy5d6Z0jUEpUafIdxQgImUaS/fG5WUWj3Ha82mAhydFS+gtez
EeuvJjFr7F0sJSHz4QE1chr1LitPGx2+7G2/oyuYWd0JL6OCNPnFk8jYFC9CTLgCW1z6M9cDziR7
MEFHzhVzkxqr4Uk0fOerItjcGT7qQrN8/QvgwJGBK2J9nYOzK3WWg8AqsvsokVfJ5akj0hysSsWc
ZKO+ppxOMiiOJzMIYUUaAW068xxCx2LhtlJl/FwxG7zxJOA49YVcXiNtzgwrQn+XIqsTIZM6YELf
SRPECyXdeyOkYIJwy/9Sdy6zReTwFPoy5V6yU1VYBK9FKsvvNP1L1RYqH1xGpVkxiypPojxjY6W9
LiTAClRkBMkRVcuaidnaaBoCHpbSv+m2Og/WQe/pl91a1mgFXGpKc+0/7U1jyJ5yYxsG5x0KcXU2
OyeiXfCQ4Huhj7zFgQ+Qwk7c0jARFWR0om6R6EoL+I44rJeGqS8x2NiK+96lB+QDwtvKb/HZsXeB
aBLr7IraAyG2PdFFM1uPTJQsvf3SBubK+nAO9PgQRVdIZuHiNeoyJXBd95b6cy/hqf+lLMU4/e0M
HT2vQToRL+u+qNlyjIuL0fVRa4j0eIGrcjO1vHuwyWC6rWUI5dJ8jzkahmXa2iNT+ZU+Ri7vsMeO
/ppaHc3OyRs2v6YdxZ5wPasKTpH4XFkVv6UD3AuVw/wiZ6xPd3Hh1RhHOuaCels/hfEmyGIo2noa
0Rl+FbjBesolDww/RcfkIWWdNbllg5eEgPVKSy/SszN6IUORxBBk8D/XzfQLEgOFqcTr8rke+UpN
jSalXia1VGuF/o6FgY8N5zr98K6IoY1/fAK5uXln2YTQz2PIHGphG6OB2iNFv5LLE0nfh3iyYNQo
CouswScgPmRxzQVZ+EykreBaPXa8SmsqgXkmK2ZBlma0OPbEAno//Vrk59ihCRixG85OkPGQclF9
bZu9sSXEasz4KeopqxQpkr4NWFk//jyalTXJy3YJfOC52Fh05yQ96ImEX/BVdSDWqpTEIOZFQhOK
kzW3F4MblnXj/r9mcKBPmtqR/9xft3ExWCYojJWvk+26BUtLqlI4gaH5fcC3NU3Sex2L6sdqauU6
mOT+KCe9usYmNEyGnc5UW3Py6cJuL6LWphPd9qW3xx/2rNklyRiocktK8fnrL1ZkRIjBs2Lz/7Cq
5SFrSszfAr7LZh2TmdEXsSJ/NSlqMo1FwhInMcZy1svNglvYG9x6oDPKm0lAlU4DzDxIKzK2GHa8
CYtMSQbMbs5aKreCEuW2WC2LtHlb1YRIls0dQ0h8dBPkKMAb2yz5HKXCQknsc56uwrUgb6Dik1WW
rWR17icx5p9Gtf4EGgb7SwYxgkOOydtveSUOxS0pXQbPhY2IUKrrviAgcmv7vL1xI8w0+x8Aj2Lu
WMxD2n2STBXUGYrBuzN58EiBbYpr9AGOglG837EVoe+kJ0YAaM/K9Ydpq34IZE90p1IhEgZd7F6z
PVbTJwqrtfFlyz59syncy+gknd5KwhKeCYkBXEp2rOTgQXHJXWVfT5v7M6a6T/QI0izbfbm9FsCe
wiuJyHchFRcCDnRIFxoJItbRJXJ0gJhNbQKFjjjmVsFwJJkiJWKtFTiTY0c8v4dUdfxehKDrCyPE
nBIXUau3V9vL4LjQ32SsuDs+rr3rGLahYWcm4pRd3w8C3IBSGR261GUe525TPYW+ZyWAdtGWVom6
bHxsB284W/kl1jart9ChHQyRRzb4oJpseXWkO6Bg/PZ3pA/eMr1zm/v6ZocV2VDDolw/5lPcWDTJ
mTIS5zg8Eg4GPzrL1kPz1UYvPEfV6fiP9hnAOYI17fH9r+0gWbUWrRLu53xycXm7g6wj7vlaLxKA
lm8TDT0uTe8QQvuaJs9GN4n6BhiUDiHC/jqG+iO2wiKm0M4uoQeSyZ5tpuzJb0wYl2shoAUmYm1G
0tQl3E+vjNVaZqqA7iZaz6waKPDTfUVrnCQpHsbjEVdV/bHGtXM+lPPircetZKthPdyimtHM5ZIJ
jFdKqAglZxHpBUI8hOgjqeiWDDW3bCcZiVY4tf3OiMQeCFSbe2s0SYasXmfrepS+HpUEo13SdJgW
PcVIIAlIbngPjUdJwWIg0IKeI1sUihW6M0gyZdxXfXN8j+UR6cvlgSggcvg6PsHdhwboMUBZa78m
NUjLbLT/0ZkWMfKa4OxLFkB+uYQSZwzmu/nQqofGOGIQ65MxGk7kH9DRSTPl3b0KFNXurboy9zdW
Gv3mmYCuJXTo7mLqCCyFmJhQnyezSjJ8guEj3qIT2TBdSGdIWf7uMab3y9tHvFPgJbzqp+xX5724
rcz9V/XreizSvlnx0rhZwIdawKvnOfU047Snprh0cH2ZxPhsNWy1IJijUmTful8BD3+2xAatBOL8
WGM3iHr3CH8BYCGqKQJM96hs3KFQEJeTlkbd2HYE47mMjixUcFS+jSfNuZlXbx99CxcLdhPZEhOq
QNJEVLfEnzfw5Ga3+NoWBByQ8mhVqf7Q3alamrRgii64ZKayERZhaZER5cSZ8GUD3ctPXHvFPWG5
v+q3W/U49M9+w1eMJirdJm6wwFWEuY2/5w6D7V57VVtSKZKtyuGrPVuh6ayFrvmB0RVGSYZ9lpss
gRrT9vU824jWaTmmLf4qySj3FcqXuho5uQtmXAZHvggrDJbdUiNcYCPQQLPJbY0uuxiqjVYQYfhk
0Eq5JVlZ4CATscCHUgXJBN9+7jyJp74/FDO8FBdYUpHMG4DqO5R4IWTzXdF6J41+VfaniGgBq6Xk
dKDaP7aMk3t2RgtNvwm5X3ylbi1sGBVm7ZqciKAJU5y+tDx087C6nELcy8RMRL+CXFdoOS+R5gag
x7MzPhkzZRW0U8x7z1tt5N1iK3aW5XUQv76FYskmEjd6x5bkk6e5jCDLbPt2pLJLKVa5Ri776eWJ
9b8Ul3ttrLEfoldE4gebkJEwFt8/1whsohEsSRVA5986CZ8xNXLU0tfpKWRJSXa8tNDtmN6/JHpg
+Kfggcv7NoHPoFiZqdzsCzXixwGyE8pLnv6+zPR5rNz9bADOnecZeCycS/avFa/3GaTGgtxd670F
f4CppEzIy5CXRZZe6eqlzPXsuGJ7641KiqCypRjlP0Eg+9Fbweiz4e2PUaGDSqarKwe8UloI8Wmg
paww4xqxNF8burXq0ENxZ1SewaGHOV4a+iSkXiSnAlsmim6coa2f2JXau71Nsa4FlI41I74S/KSp
IShJwHUEv2vaxfvfGajslWxoMbbtngRHq66ePhEV7dXIECvzF0oj0hQC0eXHHxpsSsTOd5AZ082J
2DpGb3aO/Zb84br8PMbZqa2MV5WXYdgWDzMq1QkV6nAJND9afkH9RKzhuyBWy2zdRbiawe2v84jR
hFzYoNEqB3bGey9vcsFVogRcVPTeHrMkJs+xSzkDLMKxKsoFrLp1kz76Ynjy+v7bdBflUDGToMoL
/LfDd13c5GzpCAl2c7KLr3O5YwhB9TweYIh6pAqN/63TIVVjeCOx1IT/dzzqBgGL6dj8w0JH0VE3
nRNE4Ulbz7hoAnlQYPybdzkJqrFd32xVuM+FDiQX6tEengxNLI/Lf5gJ9/R/rF0JHClDFUUB8rgJ
hSlSxwhFg6URbkFb+T+E78o/SzQQn70MVmto53I8ABS6s/QfSd9LY9cghq6xBGnjJkDQS1NJevWH
d33zczNOaYsuWHbLQQZxXaC8agej4VkJMTXQN3sWSYpmsJpRsFzSFEpJRr9yH+x7fGGriJbSKRHz
fxMHVlN7iQwkJrQqKtjwznvG5BaM+ERJcXWz62eTBEFwseWWcdAmGW/WSM1CFvrejg/I1LXqZztZ
96Z6Ybr3AMx0vEropoQ/73kJeUNhfzuwXVYj3Cj2ytPcN/vikM3bQybXfWdkEvtbMgz5MqTMUgFQ
OB3MEzD/hBX35pAKuIGXgpNNLMpbtw/A7Y2qzQ8K5RKSaSckeUIpSo/6YGSfmtQcDqs+x9JKETX4
lj7g7gfxe+u4I6pVq83WOXaOphNWMQMFGBLQNlO4aR96ha8Z4q8mrJ+yin2A6wgTXRrGxv0c0oFt
zmMk6Hln2iIameECP2Bk6fwme+3JSmGqrtESs5UxYPWw7W282BhGF4l6f72he/2PituoYF3JRXjY
1LKmmCet+i1lUEPKRV45uifI47pRGpvUuUVqTlgPkDtC08UjgVEyQVh/NLRSAVchGxhz6p0HEnP3
CV6Yg+DGr3/DkXUqT8qu1lcNe2GOBaoMNd2uIc1tFdG/caknmYCK3enqziM3szo9h/iu1x5UquPI
kVCEDy6bqykpBlwFAkcHyUpqb6vblo2RgDZ0Pqm3GSGVPWuKUdxdOKODcKvVnx0TiyBpD+mC1V0O
8DsRkq4ywCN1cUB/VH8O8F+YSh2BPj5PX0T/BNlkiDMETMAKixDB0pnJmrlr7McGmUP8rW564khx
SbihP3/B1X8OJn+/wMEHgvNniyelNwoqUxPO3WR6O5w2qaAEeZSDf32SQ6ZRyG+G79VulNMUe9Ih
Vc6b8zMjT4HIkeSG2G7uSNMI8tm+pzH36u4pkndZhGcefwxdm7nmPV8lvddx1qExSGxvEZSOVom+
Rv6A6YNKvz4v5J49Ozb0+xM7fm1+YNvbRl6NpaRQZEwN8zMPeJR2c8TcuLXOMdt+FoaiDhOwILYl
m79k0FKLEaDstag08Fq7IvWAl+gPdLjazPqeKlCJW2m7ifgCp6C7UPm+u1xSGARNK1toPfoxu9z+
IfJaTfCLx737X1Foh6xFYrLAmhy4RosQG0OEQyehKyMSKz2kK4Y0thPCBADqAWHMUldbmVWLApSn
bL2tQHtXP/ZrUxB6vk8exZg6JXeb3hlW6q7rIuIhi59vApdx7XFLFH7taHNFRoY/2jw5ahMDPRLx
RGRa/ddaKFlRoI06SXJr/75wKcct6Sw0v9KhkNns2+PIbwcrmEO5v/FoQdovOFUHfTxO04T9a8fn
8SD+pdPwd8REoEdAu2sTx55cHs14FrKNpO4N/fhm24U194c1XaSkcXlK7vGcVURq40rUpnADYoWd
tf6iJgmHeXMQxYFO3SPS+IB43NjZihRiaTrko7P6rsgRNxX+zxOQJ7SLLrQqas/oF3RB5uZ6Fddu
L4rFSxtEcmNPN7kY+pR17Qgsd1xdsOH2mbEQeeXnmLNKZEOt3d6iCw261tkVe3UcuX8naN670289
uvG0uk1vQKVOu7f4NDcK4Xm0+2hrpeUl22F5ejZsDTkLXBpyMQ1aBzezo49yuR5OM22ApDZd/iKd
DJ9FtC4FIRq2HlGuq5l8A/Yh7NE6wz+9mXGyD94d7MFAm1uPNcN+CAHQ8h8GmfSXwtt4jSbK+bcD
nRj7c44G6qwqK/sorENjwF6aScEI9RRgzPdPN+RzPLqKsZdRJrNdyWXYZ+vvodyWLnK7yo9j/fIc
l/8lC+C/2rTC/pYvBOvdhCnl8d0PZCQoZSVoZqMwqZHxDkllOGA7CgyZ+6XPQEcR/cpGgHAkXEZD
hMuMLImP0Rws/NpFrb6JcDpm7Y/C4r05qQ73FgtYJUQwhCLzFZ95tADuSaP7mdGjWWycB2h0m5we
uH8Phkyypuxray6/FgrZ3CtAAb4QARJ5qV8P+GYuHCQ42mmlkJcL3uiDGKu1JPvpP8FoZNE6dK8A
s0VIGB3tpj0k2rj2c0notU6+nwKI4kd0ayScDGzssFkbx9FEFlBZQsH22XR6pm5qOfQBPN2oe+qG
jya0VzMNQ0VCweWpYqFF4HI4xPETWwXIxln5pMsCn5+SskQcEH3F0v2LC50y50Fw+jhJLedTgu9Z
gTLctDJbbf5BhHCPmFMCNdYKcJZhjzbacUVwE4qazA+keMTfPaLosROh0dMvXXwK8aQYcsVatLGY
ynSfv3m6KLWpQukzwdwUC+Li4GOerefTSlqOyXo7kFROfqNgbTXzq3n5oKyo1dOqw39HNsoDP8gy
V/kJmGVuQwc5jCOuGt9aXlZBqp1O+G9t9EDML0RfrI0nq4Qqt+pBYsfnXjjCMCR9ajsEyq8nia+c
nT57AvdRcCh6/8ZoBzPc+YbCk4TZnnvb8NIcR2SwkUjKUMAYrmjEpyG5MKpwSfTzoYjXcZnunyJj
TcyP6X1g0blbDNGh6+Un2YNe2Jhw/ed+kIOr7tvLM1byJiy4T1nmtMQ8kYrtQE/61M7E9SPC+jKl
UY+72CtGqatMogop9S3vJuESJ0y2hobbcPAG4V+CR04pImDDEu6Jsn5zvYQj0HOHcRvFYV/M4z5h
li9N8JtHUe2abvRE8WgEpbd3Ny6RIs4XklSXP54scQNf/lrJS4L2SNF3Pu0kHT3aUsqJLlVI+NYl
T4YrtjvpZXYQeeYKK4h2nH1EGQ11TliEzl3l16OrCxvbZgqOF6ChEABsulmdZ9IU8KqMHLArOSOC
tFSufFBJDpIfQT4gcGIcDEyn4iK5Aav0BRiVKIzNC1lkYt1QY73boWq5KP84AdwUqA2+l7AfNyr+
kWqHa914wHRhQ4oTK0IqB5yh4nK2astheVG99577JqSpfl7CnuFLt9bcpbCU01ISp9yyfUyJ1O/A
hR2Me5G2dR8lwngW/btVa/G/EeVFLzwmIfxzlXXhhClgqAurHN9Y+PYbr+EP6VxbyFMOrgjZPuRU
LrYAu6cqzpNlb2kCnFA5C00MT13h97Y6SxqYskoyyFvUftbrAIEpKGDlY6u8pB4YZ/0wUPbVXxNt
dmG86RK0LP1bKizvTvK8ykQ8rD6vSJL9ZVQhJcWBZIDWh9i8sH6UQ7L9KIPrzQHdAw3KXcAksGQU
vvdNTYCP1h8/ayQ6kkidlsNibYSMwTUWxY9ahOVqsaR2dsuMnOAAV9IhALP9sO0CdzaBxnlsEsK8
OFzToIRkyd/XmXy6i5UdY9zsrb/ZOPWtpbnqPqNbAHQaa1UJxjkqkf4t0W6zV5mMyRLwqseY6/B+
pPK2M3coEz9O/qBGRRDVmGcwJpRqxj3qtKC5GXvQ0dyiMcrFstZUR4DyGQtvHiBpbyYC8SHN7hr5
Vpf9DbiJqVJuhE+sO+llH4I4TSCn7VfISu9mdU3MwIiwU28ydx5mCEd5Bfba2vSUaxhRoIETYjZ8
wtaASoGW/MdSkXNxE37ZI5Lb1qJLrQXGLcyTX49CcMepeM1Mm9UUZeoQoitpY3d3f4/YL/BY2Fdq
fC99ykk07lqqNNH006MprY+pLbITArq+EZa48MhrcW/rzuT7dEWunmVZOYLjMZbRwWwoqnCc4IRr
hF8hSjHzqfzjVEc2UQN4KW0ErHVu7i4R+KbuaBvwLjZMnMgos3PxI6KB73lAc6/T821PXv22kCl6
8II4pus/5nZulu0EgsdXI/KC9693OY9TpVBg+PAWDHxe6dF6vaHqjixnSmQHBxbT0dSDJd7jXSNN
dsjmMvV6/xg7UldhAPQIEnIlCUSZwJvWqYS7g/bOe8X0UZfXtZpoJuEskzIgf/G3Ldg8SOuw80Kk
WgQ/3szU4c2AJTP94T696nVsW3dMbrRLnqP3h4tssyzPe8lC0+JxC35CTW/uKjfqDOilSPuUx03F
edv8lXeVkcga88swOZxrsYVLLwlgyVy9LDtCad1VYkZN6Z/HoxFTDwKjkILsBBpQovKwoKSITIxf
f2Hr3uJIlpUUPGo5W6vH4DFH5Fh9R7INFi/Qgk4WU1ZwQbo/5x2GBCRx8GgPHTS2nj0pHUBjW6jv
L4sBMP/q1avOejbo67tABr8vA9k3oCtHpUwWN9FvtjGci+hzPAOXMw9MrKejluKn79b/t2MEbeYv
xD/Ki6U3k9Pu17T3QzDgx5TEkUph/2GsGXcZ9+STvH5cT3/oBENEzbhVd9X+y8mTh7EeUFFsZPC6
gbHQ1x6a8omrMDeI4HHXVNxOaKyXV5VXtD1OkHQnrKLTF4Nv+f+XnBH6kK5QO9RnZzxF81uYHz7J
aQloFY02kgnd4T6o8nYWKOXE37cRH8ruZkm6EFeaIjVjZmPssJS5zKnPZxfguSSxqPa/OGwt4j+T
mrJunlCZD1hUaEuHf8g5zGp0uKlifTiuPvCQaRRHhWh2JtPMwaP9LnsfhNeO+O+dLeYgfVrnndka
YM22mnh7Ej4WyvErOaK2H4oxZvwlLMPGuizzIErb2bdbcc3VXCFGXDpdXNr1RPd/8912qgzqbmep
whHepg799BoIMqgqYqt1Y9FN7EAChU8JOna6FenLGPdjvZFBsmXJw1CFv3v3WaLuBi97do3waHXc
5iGuFXz7OP/etY82ssSzWUXEjYrSifWWk/9shawdwh/IlcAuXK8UhB/7TgQDwM8T3JrvMIaW5kl7
i4btwZBpb1x/nWNWMih8vYgFVEw54iUKHI6jvt9NdhPpiWL8CwpF1tOIst0aVp5k6GbxDWYlXjTP
gVkDCaFqfXaJqleCmT2ccUighnhDkTVF6S489NGJoBVhkh7kFqOVnkZ1/reieUDvrpV3VrLWnyIx
WWZeqpWLNwwSxTJWEfT21NKDwFfkUaFqbUTFGF9L1/86/FRHXGjhdaBPE4pDhaJ+ioN1Q0rehzS/
mY7EYM8XO5ofwhJtQA2y9l8nZq00DkJOM7Ux7mF38ndtAuG1J0pFca4e19LuAeYbo2GB/T/8TwCr
YQJu8xqspXc1es7HrzKPI40IvmP8DptbHoLXAk6NGFxdlpL4MIaWskiW56/XEC09NUJK9u0wyQIW
eGz5Qc/ZL0LTwefxWdrF5x3z2GvDmx7DipBrhj03N41uxzuNy3b5wlieI+kEJxSzpHzEdMXrgFcL
om3SAxh/t+B1VTFVO2MYHu83t2y6z+bQMW3cHzoteDrNJ4i5IsgR1BLJ88vGAI6KJVbgqvegbKdL
4UNt9jcOcs+9JQmLb2SF0Q4E5zmFGUpNmeuerbmwZxl/Ag2YARuJ3ZmGQejrQD49UbeGIFrZyHHo
2oJ30k5mv8Wqcr0ssiMswINr6Lu+r84pj7kH/IvmZcZxVGC93ZaRND03cH81NejcwqXM3hzTzOiL
pmYz3Xrjzy7PWFpEk3foK18yE7srFunfESDAQ4WHvZD5XFADBiz+KZpKMva92VbpdgkzHBwd/Mp/
co3Y7HSz/PqeGucqEQ13oKQrL9uLVzGJvvqdYUt85GlYcnq8wiJyldHJjkD73b+0jEyCPYGOVnAj
7OtGNf56Mw3Dee0xSmPVovIuxEbwV/YL0L5ZhRGOlhM5kdk/J0BOyC3rJIC5G7ffT90wECj+Ult5
Gq3OxJap+yyN0y4n0X70sUGwpeqRJmVE1cspDeBeEnmoO4AiG//MWkeMYSelhpRENHy2r0ONSn1u
Z5+ohQDZETRDXCnXiP8N6x5+WDS+Ft/XEzPwwDVZi8zTpDwqLh4ADdxlefuJdmXlj3sCE4ESg/jY
G/VYbgPd9bTI84GZ4cRDOvM3MXbzeVSbt1IRHIDljzdXwSz1AxpSdMHBV3s21De7fNkpxAEWuUxw
Si+QQe4DvX58Sof3taWDPQAUTd+fJ1iSwsMcG3mo9+bMZe1B8JjAasQMFagQ5WvYnhJuE3vTyb2F
NmvQ5lZZvL+7w5vRJfKUaOq/JxtfXAA5gZWlAfz0NxafYYBYtS+HVcwWzbH5VEMh6Ls/cPeOdVJU
srVMClDiH5zlc4d4dJ+LgEhIlG5KTplQ8G61kq+GNTLbeMzpB26kCYZKYpdw/RSohXez8R3A3UNQ
3jtMDCicnhrtf5prT48iHRtfbRQogsehCP8V1nDN73hYwky3SDsqgrcRs9j5f6mKTdayF7NJOf52
juwp8wtaA1HUgJTbFaRF3lm2f/RsFHpZ3fmbq3nqudsea2FxxFAnBBw5jVI5RPycKZfxVnFe9SoT
xNKktdM6J6YT0sOr4rYURycvZ0oMpNP0lCvuyqS+kHMcCpkBLqhSMOzCnUBiK7+wkWAmyC/2n8Be
IlQuuB/ZveYhGCv3E3gqJMuOgQM76bUhXyUpMvgjuSy86aI30miflLcullBVqpNGhoT87JvTpds2
GedWASlnNwTout0RaohIkcAs/RmDR2hIUJN/jpVgwE2gIpD7Wtts4vTS9eRuUwAxZZ2rybXgdXaI
4Y/Kmwu9Fxw3J+UnftLvFIPo//9xdWvBcS95O982r1qtdHv/Uk8Hpm6dcCj7aNcPXbejSih2brQQ
Gwbo38Jk1Qh1PzWON79/X/5TnvaZdJws8LSPXG0Or2Ab0c8BDrmHkfZ86BNJSSiJyZnS2qpoIn80
RBCItyoefwDM/wiKv89DoOTmlHm9HErbh5O5f3yyLr1dfsOyZR+se61RyMnKxsMmyuSf5pEB4XWE
bZqNsJdwgHf1hqYT31f4DlMFRlMK58/PqGttfXTj7VCixsUnU+oibyICyXSVADI59RDnkF278DnD
KPDX+H0Kr6BvBdw+ErxRARvMIPKfraUYMaBj45KCpVm8twqt5xvbcJxlZIJ/eamgCuQuAJaIxX2y
yVPMnfBbL5xzTR5Y0xZp2bz+GVS9JOlH0A75W8eTv6LUvxjggilakHP/NESbkux7VvAGi8iAk3ql
VkyLa3fbWB7lKNWHYVnT7s0mhTI885xak3KsMeOmjQdRU+6MV6IfNjBlu2cQuIGXFmraIjBI0QZ/
MYcKGcZPp/ruhlNMcdlnyONNjeqEwR55QKegkTXoumfwMa+vSceQfxSimG/ov0M4QQBrilPPtqUB
4PTzx/ZtkktyPZqlsEZs2+EOBd2ydtyIneHkFOWjyecScuOhhDuvx996CS5DBynbTtmQ+vbyNlxE
JSioSrn4Dbp5NTT5+iTTwnAIdQGu3uO3H+dmMMbYlNY9OTF+x+8PIOMjRRRl06pdu/L821uYJmUD
6tfNUCprglBwfAiINw4dFUF8vZCjbw8k9G7AsdqGLxKQdmcur16SpKP8TzCsxICTTyz0MT3Ekv/C
Trx83YIDin86Ip9LotAu0R7meYdtGcFaYP9EPS73ZsRfQ3uBTP9+NpDi5UopwgZPtY2MbY2yI79n
vqZDc43+W5laHTUDiR+JrTBvnCLFEmukpwlTFf7jDRtdWOa5kkmilrEjXZT/qU9xtjcDMv51bAL5
bivFQuk1/kQ6xAstKLa+wA27cpYzQN3pms/WrlGLw8gkZagXD9rLNi3j40XgQA3AJdC4brdF5B70
e8DxJlu6MuCsogEWXEupFbzc16xUvGzSOJyxXdGmzbVVLz1KWKMxBzPYVf3px53jS0y2mreXDahN
E56Aj9EIYg8znlUnbjtonaeE2kb1K12ewHxX3y5HH2LIfYukMwhoL38BGQsdg+r+KeMF8atE6zOY
ruPRGtHgNH02ZgkEF+CxYLJtxUUd4REImdVExXTmGoDrnDBWmj6aOCbY36QAGU6U0Vnpklhi6POa
m6p3FwVPIoPYw4Cogab5sJAsbQUhrHr+Vyk/6mCdUSnj0LuotLA8sbhZp6b7qoYlX8ZYp0ByZqUk
Z+oUvZMJjNP93wUZFGzhWnNAZvBbhwMyNHdywKt+DNTCFPh8D9fIxRLX9qxFSHshT6DVcag6V5hz
I0K1T8lENJCYb3qbWI7LK2eQTLQJVdzdufq8xXEqlujdaivw98YpuSvZh7o+oFQ9ZVoMNiCZSfTw
nfLnlM1+N1VdS49+1uUPfkN+D7crfvtrlv4iQPMdWzhCNa4bvCgbvy2z4MV3Wm1DFYufkDxS1Mkq
wznpv0GeU+l3d81m+8DrDQqwg1cQUb4rQHx0ZG+usjjKlPo2A5SVf0XqdR1ZjXU0I0UmKe8k3XwX
Mm9U7ar2wpiM8jx8Fsemwo6/MH93x074SY1jizLJGCjGZ1WoP5Kilv482GU9p8PCum5UutUrD3R3
V2wTWxhP3Td1PYzWpu4CPZ8nHxOHQKtJU8Iqof7lm7S8VsWOGQJi5n09K4NjqdI8ntGc8AJ+VmDN
/DGZhgewrzeMKoeLk821V/ljd9KthQhemrWbuzO9Frn0wO+ECZbp9cV6C5FdPojAS1jxacRaruGt
0uB1XYC/FhJVFWrP8sdxNMEv6TCXK6+CWGicyEUUbEgWmwxcwws/e7AQ7Nior8XgKHgVe/AFFHt5
DEMr+Hdqdj3wotzFN9d5NLxVHhPgWeDSWREScPMWJz5H0wpHXsR3mKMCJbssNdIw3ejVlzvA5sNr
l8swBqgsisFxhHJx2V58kfCyCmt1XZsGHkVJYJtkv97P7d2qYuQgnW3/w6jyxdiM87n6/SwK48/M
BpzzD/mJ87LUtd/rpFn8ew/IHm/txQq3Oh3wevkpk45cp9VLpQ8g6XGZtQ47/4wcPBPKLHeZoXO/
BuWEMvXKKDSYVNSeTLbkwcjDMaTtBvtRTr8/Fe7h2TNDkEnvoNyGkRJhz5QUFDzURqNR+U32vqF3
XO5iBK4XgP49t+Oi4C4wgDKvEOe6byloq/8hsUtYeLGyd2dl1g4iE2zCqc7dQuLr4IzHeY3cL8bj
Fc2yAf3Ccrq46LkkYw1/RSd06kz8SbtZedR8cArsGd/MD+3WZK34Xxe0F1dTf+/+twgnq/JPPXSe
t6OR2EvA8yNYcSdSp7yW+KwoaB1rcLZv2qVT1nrREWj5seU6CSgyvIFAwPwWdoEkSgXvH88Z8nYm
jdpmy3NxM4jVyhH2DbRhvg2Ol6BBIt5zM73dblts/b1oRVABdVuXKAdJiWN4Vf9/hWew327b2Cvi
M0kL/nvAozdIFddZ79lARzVZbAtart5Qw3dBixBhDsO3LhgzW/Xq3YISUsAWQBkAa+33evnEJcaS
8lec2n3EUJczMZeT3+bmqL+ZWAbpio+BspDB1E9FuAHxwdNZPrsY4zHqCQ/wmLWOT3Th1stWDpxE
RYarolaGzbjcr/l35KCVyuhOJtc6T8YRR8HDbzhbOIHfIQBXduCDZ98vVNDBG8rc7x9jV7BSa8AQ
lc6mWW5eO4eEZmjGU+L0rwfqrVJVC9bONJYZJ88gJFq6pIMcsY8IiQeK+WeQbc1OiD+K35McSRbb
5rC6U/7G6L1K8NeKNc70UsnRo3W6hV3tYF8nG5gU6Ja9HkWb9BP6Jj/tUuZXnDmO7tGBp+DobyxQ
gW3rMNe/vKXEaRa7DFL0BFze/lgPZb8ehvi3yW7GVS+7ScdEB+C2/1zTivY4Q5aPkRZNEUPb/GVH
jvIZHLtbOTFetx15mNg5tqxqUhIFD2aifE9lMrlJ4ywups1/hEToBKI3JBUf/F5Pv6SF+Mxh74w2
G0KQcjOGOAqLjRALT4vNEg7cUAB2gGEnyMq5Rsk9m4I9jrJORbXxjrCdpQd/ZodAcEibdfkbLmIN
zD6HRXA/kD6qWUy/WcqLHbs8yFjusqp8dR6lHeSoZLNeReKS6LwYLw+mMFHNw4l5vG5v4PvWclRt
tE0vokXW68UiKGqKd6hdOuEkfuQZlgGN3Bdi/uNM+sKq3/Uxa+sf+GQmMFfTGGefGFrg1ufggC8x
46D3bPpZ45kJuXbAoxXJ2SLQjAXw1h4k/5Y4omqeqzQWfh8Smakv8NJXMS+9YDhSnSgAqSH0b/Jp
9p7pEjYUilEmt97eBvPKJDpBfJ1CF1jH/4fsGos5dwcQNSecSYpdu0fs5UYq+LneptLzeFUBYLt5
aYNdnHYTycoAf9NPbYy+C9EODRxfK4m81Nka++AP7N3ne7XsVjJjjEyOLC9vE17HM1Jo0AtOaxGj
SH2KqvWAFefRBsyyxQDcvkEsYMHM/UwMBk/0GMvTajHIPthMq4oow+4L635J8XluExfPBWsc5ROL
KUNHkVOuC9kgDpfgNRWQ0tVKtKyqybG5/kWNokOoW4PgrtHwrRzUS1HXilZzGEOS5U1P5xXPbJat
I687tjcRJWY1/VP14c/p66WhQwM4LNRaIZVLleeO1Z57yfjc3k3TbAZJ6krGonXe0TcS0LTtghnQ
r41y+x0wFFVpq8HsuWex9M3vtPMiCu75WtBJRutwzQfrV4NhUQl5Hh+RUksfnzN0C/0g68PBS9FY
59pXMLcyHS4KgB+4j3DsQaw9VN2X6dbePhU7pY0/01TGLoJpxzw2rt4tDNk/WQZpY/U7Kvn47u4l
HI2CyNDAFL6aAo/3dQiJkVgTMvcc+HfqvsuUo3bvvwL+0BCA6XAUAl32XibdVRiO/ISnnkZTZY/T
VwlhKkpDd5wNWEcdDJvkEjMjhxu3Gi0Z6vAQmL2b5fIxyTUJg/6gxoVeAk4ud7xbGS8Zv/Wi+DBD
QRW4NqMSGfJwOLnTN84YMV2cLuoAzmAbHZa6KXRqTR+PLSM1X/v+DF8ueW52pSCx+N7PE/DkuSS0
4XTmNGMJwokfP6iwf4Ko+/LRD15W1cA7kYkl2lEb6Cxv06XmnI3QbaZ5G1z0TrCJBX9pkG/5Z0V1
OXddNvRKvX4Rwuo+F0xv9RdWWiL5NFMsuIGepNj/E1WR9tC9jj9auXcXaHU3IntA87xtLHS5MKoz
1zFYDgYkhluES5jGnleFSoBLenf99Mk0FOAwGS3SayYQ0F5MeTErdgpZ+RoMkEikoB5l5QKrj6D8
vhzxVt+k4W4piD0dTsScPoU3nrEAZ9l9ahxCHQv8x6ML2eK6JMkpUHfNYLtpVmqdlrubmJ01HsuE
wNfgkFobdTiWAUCk6cAwU7+jBrOe3sS+xOUG6wCJGBnaM14Rc3nzb2xJrnZRjLBGE0KvF72RhyBv
IhSi9iBeVly78ZM97cvEpbafqP9VF4X5xyk7aep07fKGMiNjgkPJO8an99KhrZWgxQp05yTBBEih
+OYnnKsUWh8vJca+VpneDrUlVdsPZGkO69sKolKqH2P66dGwZJtN0vlxmzDw9RDrvqtWbTq0oX6e
Szq7pg7Kyip/dCUeM3CCNhKTqXh1yca/tZjw8zvv25A6b/bkwEW1shtRX6V23LtXEXcwQOJG0/TX
jjQPXVIPosDQWLsy4FCmr3XnlON3iLwGx3Z9fE4UFF4BE3NeWsrh1ssLAYmmW4m7V+j7yMT2ARA5
gxh8OuWoB0kjWvLOmeTB68ZT2Z2o2iKukQySChQxBbFA8l6wYkKBfYYFt75pcOeojisZHznuKbXK
R4KF32m6yI5PRCrSgDacotef4rf37dH8nCFnymf2MdWxk5M1biLJuIMRExAUrLkOLPoTSSfpruSV
aQU2cxGYNN2DGNuMYBh2HF5aakWy8K7k9N1HSOF3fmZjAO3BqPmGocNglIONJDyqt7zH5PTUn0ZW
Wk3X8ioTiM63fEk1uuqMTKDGH4ntyO7eZLkTXLWlBvJBjFzzZU5RyDXWgYGsWqOLDZoNRmbzNm5M
7lOvgCtQAJgPfdFcGiKo2Li2uzFJq7CEJ2b++CBgMxbVawuUjTbcVDqFxoFYUDzu8l84IKpoB000
2c0so2USIlWxqTW9dnMeHbvnjdpNIZc7P8OrOahJBjAUHaDYjAxoiN3V/lQKWxCQSetmzvAZ5ziU
3/19th9qnb371/2J0HIXrX2ww6sOxc39/dgjmfmAjud1VnAOqtATXWNUU61KP4RFXC5JJpuOd5o9
zR2LM4d0s07e5SB4LsOdzTYeQ+cQVVQW+FTNot6TRAyYgZzx3bRbzz3nSFLg2y1gBN7YLYMO4bJb
KsDozgROIASEV3kZsnGaGiFp08gqOYGchANCowfWI7+GDH3w7HHG11IyrASvXzU1lLJG1U97NiGH
4XcFs+UV5GYAlNvC2+Divl2VUgml+7XujbjNy7CJfMy6thnV8sX1IW7r2jixUK29fnMnh24aszKt
63MMjsYU1G7pz4mdIrorDiHAscA3G+m0rqbzBGgMaC66epxl3fOSNL7t+GhTiu1APH4Fc3S0QssX
5bmQa8miqJwQS39E/lYlDNIGJXIMLAAEVHA3PSQJ/m40pR4dU9UAIzWxUT4VQlfKsScEooZN6GcJ
1RlgpvYURFDqYEemcIOloiIjdzZpIMagKVPGk+sODjr5cDxbEga3i2EoHXTHwqvh0Vwy9CVis3uJ
+FdjLYZ03KIOV76f3IEGFpnX6iPO7i6EkyejwEJMx35/I/vgh866SvGzwGa+kkcOigRljeE8Z43/
B8CBk2Fc3PG1qmnLPhntlYbqyFNp6hcNte6NauGOysz30qErqncRpOB4XNOjcS/AbwcR1c8ARvtM
2FH5oPlbJAXO2oJeW7Qmw2CTfThyxr21DhyTFS8We/Eka+U5IbbuZ+w10518r30pRkZ7ZcaWs9dw
ShhVs2hqTWuKPkB47cq9kfb5PPmhZ1KAj2JNtlwYya32xmvwvEzeFOKk9j+/AnVgWoAfl21lfwQG
vUF8fQYQLIscpRAIGwdaWFNZ9Wx2Sl9MtXTT2bKmYSv3pg0DqMgRUy082v/jErTPCU9x5n70olDp
BZ6VdVeQ6OtQwt/+SR7HLmKFaXr9VVTm5hn/pFZ84DxSOeUWrRrHri9YbiEhvkFxJ9C3btX7v8pm
wn2rKTIgLfeO7If1IgWtIZuGQ2IrtS1hy6aFtDHSpdh9XwYnwm6XLT3qO3+VZ18ZQW+4Sagy6Kxj
llA5H9VpFxmx32DHKexGxtx8960ZNb/frRSvq4Z1yzCHAPyxdlmbEHsOnCirg0eIGs7TcWzUcGwB
GxwfyAjUgzhpTHplED8dvqEjB6K/LSsLSrRljIWkeoh9afz/AYm7639qUbqNp1bJGa1EAGxrBWlM
Qdj8WVPfkN8okuzaGKVpi+ecy8ILk54haXo8kaqFieKBTzUKTeTINsiOmYbSHzg57X8x9MP7nWSr
c9mmSBiBeYLaPDJH/Hg+5LJ6b2Ew61svWVlV6mI9Yu8t7r3Xc7ojIAegx1V4JMCYYT98fL1NFLKD
8v9Aj1TZEW5jSIU3C9uBcOwEt8FcckuKHLslCv9aRKklFF/RgmVgGtdoUH8tWll2X2bYFQG1rTc6
Fo5rCik/NE/m/WF8m0oOEzUDdN3LxCuD5BeRAF6+WsJD1aceTUUtQJLvn5ZED3nAZlxR74yo6LJJ
NyA9g7Xcjy3XFaCjW87J8YBPiEyo4u6byQA9q0S4Kd+7eiLaETW+ooMh9QU5ZsommWOFV80q9oEC
umCt22/GW+OumzlMnQDH9g8UwQKa6hwej3VQV5dqm29AvbrhYu/v//1a8Ld4SthetVmY+u8k330C
ADD1A6ZwDGfTUqlwTeR13GmNeQ8eCRabTAIJD2dZwibWQ8X2U9l7l9F03/1OnfUGc4Ui1tnkSDi7
pDExl0eq9CuPkh8hcVy9T2UjEs0WNqm52Y0KaB0ThjF2eFNUh2xIOznQE98hzxa6md6wh3vFTihc
GKZmU1cyIEeUzvXGvB+QFYW/I3HY74T/OdrSofPIAtEWXLiiJ0bYWK8UHJuCxo2/EqCRES378bDT
X88KwQ/rH86UipSPtBmQkvgg8bO4UN2BcP/S4dEheN4v7IF/6y/h4oB98uSFHXE5bxyFy0osY/U3
6CWjRVUstJtu2+oFT6TK2SFUq+FKZ8G3Xf9TLSkdAD6nkRUzmGRYDJn/DnQolJPX8SCSmMKIbvDS
vDfSSa8lfV2+829dJSWmLNdJIoLvQgBA2cQy9882iSKvgF26cFS6pPP+QLPyjgpqrrogfnSh3guK
n9h6xLke1rlXtJdbGdP6VHjt4n6K3bzUusNfxvb9WY4xNyZE8nRjCjzN94JwlXqkZvc73x8ZDpSx
KK3UpY7LVKvNSrDMmlqycgWonq5xoZFavRYUEBDPyj9M0Yu+aajIZV6ugbR6ZtBza/MJ/uwrS8l+
/VadmNlsCWX8epXFyB4Zef5W0iyEFl1hGKIHRaNa90+2vOMIaSvu99YVT277Qrtr/8y5b3jLxMPQ
6jIzTIZl73Odb16M934vT7ZQHndXYYKMgBb5DJihNls3O0ZMkAPoS3qnH4aU52jwllz6jvllHM8R
LpcuACWXyAOM53nXvtIIB1fhTiUG6mPWytfTiagFGo6Ch4vUWEr9qt8lMkYLz+mWKGO2z9oumA9g
XGXa6kvxk17zgBdq875eg3Ixfj8NEBmR5KlYqYTJGiO2qAVv8ddH2EHmKRdWMMjQICG+kPzgi8CO
+hd3LoRfBmnICatqU9BTOu8llOAEkxZEtCzIsy8aQdi/5qDQAIX7pqG5c8/KZ/QGRKkCX8tJmeWE
ufQdRPMTaPFNoE60NRcl/PdUy9P0mTwNachVPL8V3lZHv2SWnJKS+8jgho2C6zNk/47zhnE13GaS
J3ZgLrj9In+8kkUNJjzDc4cTfHpM2pSJCoW/ORQH+nUVHdXg6e8rUfEpEqR+wyBySBiMgOVQ/fGA
w5psGDiveptwv88Beod8yNgWv/yu8MJw/UXbqG2/dHoy/wTNnsN/TX7TBIjCL5YgV1Uz2zQNGfRy
EL9P1esjnRcdtAy6PMJe58ei4lysM/5mXSyS5S/jXtrsickeGezWdTxVbhO1AuNLPgn4dAKlmjTq
BmeOnoLq5SXsbCS3WvzKl6kjJl9w+svFp/iV7kAChTf0WINJNRBIF8+wAThiIJu3Wfdxv0w8hvQA
GbYSZJjAiSptWX+eoEpwm2ulFXWyvukCRn0ELiy3jyoia2ryfJtTZbWSYFIKvYvp6M6J0djoZP1y
VPrjkPdihjDq8uJNhDGhqnxwvor1qScU2L+WXCqImgAVUEfYnfDWdRdVXYuWGXyl4bV+SMTQyMug
tqR3/ipJ1Irerwdt2f8yHuD7FGC2oZ2zX6oPhOZt+9WHpdc39tKB4pIqDi96JLklX6CVjdWll81m
CEr7cZ35WGmp99jIzjnO42KGdGOXyPCVQO5FgLOdgyBDVKu/XUUEp+muM8Gbh+3fmcLcgYr1vpFB
I+1A9PktcEwLhg2Um8dxNNIFJCQvbBa6pHGQVqoQ2ofLtC7R+6LJRJOnFuqAK/NxitxbD817+aII
myt13/3mulKaFSUjaxhOrPvgPPV0dD3X701P6a7aAB/4TKiDH7C7/b0/Sdg3/NEHQ9Mc/kG79BBn
KKK3ANcR6TxODu7jH1EEDr+r103E+Ve66zCuepNLCRK/rizBt55DyEx2cAmyGU+z/I3HWH7LELAu
io4pCep4btl4YkEnDZEb8HGGgvnVr5JmNVWXKcAEfNBUtlW3sixhiUSVe2VhoittdRZLu91W1elC
PA6BvJ++AI8AxvAGwsOlYzsv6AWbXLY6AVeaEsPvbf+KQImZfVu7h+x8XQYgHexaJVS+IgCvMKAu
lDOYSL9FQVzXIEZdD7xl/A9yN+Hmfj6wj3N66Y65IMFiglsAlojrw3JQgA3vJsbpNR3Cv8bMzFLU
+AIfTLaCZM69XG2hsVLgPHAvtHPMee1UCEBDRFImFfwWJI0Fy+FGgL2TpptE8ln5NjJxnkpGnMO/
OpbEcVQqE8Ag/ZMIGqAU0SEMVdxRiTY6RuwPETkYN56K21/ETkvQLiWzUbdp0Oxq5fFAz7BXdRYf
w6AYIxRB4VYQIKATciiTh4hpzZmHivCEDTRsx0ty9GL1THprs/i5bySs6ktmCwGdCeA7VCZ+izw8
wcmXS/5qFUdlIdcS2aAdi04eigi8iLrS6c+oqndhd66FeFDGzT+p5XjC4DUpo/0bfiOXUQSWuJZA
GCwd3ED30xR+Qt/9rdXjZ8aDa1MfbzGsl3XTpZsSW4nIx8uEm9f5YNlL5+NcZnKkZz4f9WFPHYNJ
vDZP2LnG4PlBIUM+4uOLblQ5/5LXLndWOwq0YRQt7/kChNI98IX43KRuEkE98ZlWen+jfmvmgFWT
RqszmUAGtL04XfXUBYclUoACwWoy5L8CaWBaY0loV22aVRUM27n5Bs0x4zCx9oy/pMyi5a2k5BRv
8UZG/h20aKVHqpkfhz/trFN5eUPIS7a+y61RiPRPiuia6B6stsi2XYQ4Z1yQBUqRb10XGF9/2QFq
uj/jFNIC4e9msnogzK8+omzeLCMIJfAoq1Azqdrs1P/1R8rYJ7Pw8DcdCq94EQeLsJRQnhPaa9oO
8EpgU2slUbLsjKpFFF7VQzdC/LCPz3Z9sC6Wn31zpwsjlHMZiEcCBxZSpMneZhskUu8v91qM8ucd
+NLw88loKCtM/qxoJR4NrusNo724smEkMRef6GqfOLuQE3RqU3AtVhW3j7Qj+H72rz/VHimDTHoZ
5oZxPb+sJYaOLUS8lioSsLdJEHEypeXMuTKUrT7EQZNxaM0RA8BxCZZMNQ9glIZNT6mFEiPw7iR6
FSUlzkbLx3oZ6EVrCa15F5RclhGu/SKtyrTisPse7d7X75F5fTCRwpuvty1vzSbmPL2LQMbMMwHY
hUEqggMa9ba58sE1Gf4yzGBMLMvnb+6+rgelq7sDiOPoIOE5yQuJ9oh3JSWVkpYd/sKJ+ccthL/o
4sYtG7aBwZcil8K428VWoTLVh93rNttFi2ukeDmgUz+ckXKkOqtyyky2rqHTekKJaRVj50Y1+OGV
NCZvp7yUWvvaGSRey0c8zaNA6gl7clU+Gk3lipKU9xmhtBmdl7leykXBFUEw/5kAEWN+R7JIlO8t
xBPYsBA7xTa16manWDJMo0SMaHABaFzXOCtrRGyTBh1D6biniJZb9T9+SgbAeqAbBWxYiRajC72y
jShOj3TATwaW4NrdzI4UYy+q3ZMJudwmJfndGhVPY+LWkRMYh+c7LoFXBRk9oQ89yMkvGJlUL8lI
8mwG7yYj+yE2l5YybrkfDr28EotehYweEyGg5MhlSBBpNjJZie+gHvvryb88m+6aVwS8Q7cO/XSH
75eof3KkoxAYtV68CX0p6hI+0d+JkNLH+bf4haPlf+QEYqW2NnsW5UpdbIU9RCKnbxybl9fiew7T
etgbT2vu6XgSVmDSOiX7decbAxOCcufTND6Rm+AkQg+PsS3DoPG8BxOpJZSkTNkVHbhZ0nR40oGg
kObZop9Wg0AV4ErOJlZm7E/kGvb0gCppI1hhxFupNelGqkbd9xmJqTBiXb3cR0Q3gjn89eFgso9u
nejrZHXMCSMPUFjRwAAjzjO22ksdO6/Q1pp8zJzKdPN2IVnFK6MIaLXGp1gzpHSq55rvnyQ+T1Hb
mGOMCEC8ZnHjcQG+4qsJoTnazzRHwTK4mxEKy8/+wYhKfZJO7YKfFQOxOUXmZXIyLCwyBeF+F4a8
cp/QBLG8UfDMAXl1ZUX4lILc06HvJUpaEOCIZ4imZ/299MgM/4GETgIZiPDuFDfLnkr3LlI99apS
GU2rkRm0F4/5jFMAcWIwrcaMRocDvTjvYaZDuZ1pXjrYxNlyIfY1BarMcRv5WX+6oGb/fZfdlzeq
f9Mrip8H1+o7uFNZSDni6MES01TyHdLa+Sfat0sNBqH4sTmr40TyKvpZvBK4GRXudQm1Lj0xUXTr
PalaCnXBqfwf20P+nWb+wZmz4BNi4qg92YlcG84aK+c6V0PW3MP4vH35fK6nD5ONawNrr8DQP0cu
mjtS20mHPHrfTVMr+YfwIfp4hZGk1iJSTRPEmpk5ptTT4tolPJV7wCLZwq+H9J1K4e5mUwQ5We1/
YEuIggmEyZUkVSG1as7ftnBIdPR034xkmwHvRpVGV+8zpjs9SDk+1psxYuOFl5U10YRUuIQTO770
lNjDG5TRQXWFM6Khi6hqpWlW7BZYRCYIC47Pf/Jq9w3mP+aw+f9lFlz1d7Lqeiv0iejD9E7+GWyf
A7I60A3kuq+PESlIvRwwt9hqIunISXzraOAuPuH5zrddHs4K3doYdaPydnr7BcNj20hovEfT+Ywo
MaW6pfw+Jd9f01xL8GGLjQ2OdxgUGWY7f2o6CDmSO+81B6aVxqrokd/bLPPZbTaMcEcnZ4lq7xQd
Q0IZCA46TyZADKD8ZDTlIriddIXAYE+CGLykw7HpM06+Uul/TwW4AIyo3Bp6xSjhVv3Rjh6mH9w4
M/TheudqS07suVBkQ+X1OGWbFaJYQsNHgBKTIG2QQOu+KMPOGFNnSXqA39TIyMRa7eWtDxAbdvLR
i/3fx9pSkqOlbBn1ujT9we0w78hD1/hZX5X6VIkXFLhdwhWQvKJO/3qHhvVHETsOffqv8fjNOh0j
H+ljauy7kD6HelZQamk90hX1NfIPGXuCyVMm3IVE90TUZZQydBcB20jXMaFQd3HvOTxW7UsMQuis
7Z9r7xbVhBmLkYOD3TRvYkPfyKGJFvqf+9QoTFoni35zYjLc9ylubvqyemX91C1hUcC53RFSx15q
J6YuZZVSwmDUQykHWlxYeILj30ErDi5R+lnKZbNyuItarE/+EUXRqSiwtlSnlFwbVLaCFffsdOI7
+07ggvaQ6EvoFu4/ywTuWcQmvONGjAqsmt1AztjpiihF3MvqX7dpz/dm3eHTN8YXD3msRNcQFVnB
Bmcl47ihJcIJxkZAYNN8KsuXQi0t+3k3pcFiWouvqrr7UAsMzWXlJotnb6kTLudarlk3ZX2ggcky
sbQT6QPQNqzj2lgxK7uYoMgJYGOQA+T5Tv0T0vTyCTRDVcuYL2Md8VbtoxUFevTDsfaUClJJfFuG
XWDtPJDvWv2I9SCCd7E0DKhXeEo9z2WnqpReBuT/wyQClCLaH1oh3LOQ8Bd9dgTBmfZ6rUHrKkeI
/YvK4e6Rip9Sy4V1T0tJ01I2vFNHUN/U5ABtwtc0/H7NeDFkE/5wu2I2vFC0ZY+Vz5LXJIdr0Si5
tZo9cWYmUD4RWA1BYHpuBP8izypQetq/jZ3hkFwfRPdQksTzMWSI4bWBzIVPLEBTNaf+J8Nwqci9
MWisFj6aq4do8tdxI5zxQakfCZIVX1p9d2xgHnHO6tgvMPN/ffIUX2Lgds+7nvVvOrdyxt1dRxSR
/ZzeFtnYumJq8B3U5M6N84D2Z6OjYc4IE+Psqpy+3zZLT2FFnAZ4ut34dmSwwc5db4XPyILFMnB7
T2HisL6Vt7ywuEyNQE24vejKGH/7/kQ2EK4ZKC2u2j1MmM1D41vUZuyW8eWPdEq+RlBjJbFzVDRs
RBhCF+VwjL0ByGl/pn2rMAglYDMk0BNime4f2Zq363Qm6zsgw8/9bZHF63e8FxOKX4EQ383GBYkE
R2SZfGyKBv1mDXt61GTunG8sksUlURLVBb15kkXDYMEca1vElguOMaXloafwLPL8TOfMWY0Lkt0u
CXv/re+qjJ5M6NWCq9nihjwPlnwZYvr9gQexY0O3lZ/RvE+8WmVByVEMbWGlz/4W6EAz4QaqChqI
yoFjwb0XPAXDjNfDmwef9l+kvNUdbVRc3rBUsb2UM3la3zU2+xkQtxDmgrFOJq6vD9dGT1aq1a41
tk6uNuu6tm7sjDGU3vgouupVvIrxk+VmKPdjcfb1Y6lsWgZ3nhTnpTeEsyrU365kueL7jETlm/L6
BCj1kv2okPROzAG/bKlebnL7zm2wCrwrLQdGXI+ztjCDdNF2v35XQENZO28j+yvsrzwpwr9yq6oi
ygZ4luwd5DgsEXz1avtCkLZd3lRuHduqOof7nAqARhfnAuhAEgVNReQfhpUBrrtqLXjxw6L4Y3mZ
rkluxYDETZfoWk5UOy5c85eNi6FCjNN3Kh4aYpaLG+rjtPGr4vH2duUjQ+EKrn77Ry1VUQ2rHyvA
gs7cGup1u0k3766MgPSxkdB4q/8MlBby+4ARSC1/54snp4Rq0B39vOctEsO72PkRWbQt+iKrIeJQ
07QQM/vY0eGS2tpOscuOTaMzX7Lba3diRgbE+o+m3oryU+sEdPQxhCsHet2g7kpaW7rthpV085Bj
82RAmK+DwZGUpstlul0lK7PDzNzt5Uqhb/vImYhTMXrvTYBcjubXX0OpFrI/yCkLSaXWkBwLJJU/
V+BFoyOZHFELlsrDi/0bZ906WrvcJCZytM7rUGve8n19JiP4Hgfae6mQJNX213QQzg2AjcjQceFc
aoVEj6NHHoRnz/pusQaV2rikHLCjUsUenBNvR7+MAX/pNHzPm7chs1fl+z7CBA3oeFhdFw0DAd7N
z/d8v9u7ibuEx65jKcSCYDg1le8FUItKZwSkoera28qZFk3fDkhtymKitCMsQ7ZG5H3fRFLo8YUn
Axdzul4gBOHIXX9oDck5qOCGUZFBXMjMOQUk9YhQ5yQDcEB0aSp/PgxikKBkIDdDsDGcDdAxuUf9
Otw4b33bgrWsRaeO7MQoHJphJjq4dgDb5CWcMbLhwbh4s9v1pdh98RiAbMKUdVWBN7ZqfOK4Cor0
KgJ+7VFGX3NOKlqIcO9GMAIVOocS3MwQNHbtq1LCKAxTcALgHQekereMsgGFESEXs8ZzSfbMWhRA
VHOCH5yWHBjODuCpXcIUTDx99BBa9Wg/rAuD6nMs3d3ICo6l+KojmudUAUIj7up9OplbFoyV4l6O
AwOHnAvBb7QzEuO4sdp3/NKiHeVKohf6zHdBQBW2/4ich2X+DGdMoNvkhj6wGlF9HKQoZDeqAb2E
3KbIoVwe7/8cB1WeJfNoOdxhSWfJdikdC5KfasOU0cKiEpxtudtLIIWwp63fMnhMN8nAltj8cfka
r0ithcc8ca6xLURQconlTNQyt77wuiXkrG979zP+xiaLb6bqtLQCyXmvcwmd63k3kMqUuFYPVkt9
XVbpLwT+XmpYcp5fptsgbksi/MeGJ4mWe6zWAclGpIJvi00CvHx9oP20izOhazubun1UwfTTO/JK
4RcuNXwPYaTi5uN7m+Hgu9s64nnu2bcwwl2bh1WARHW7BvCXtKE7wo+mKa8zYpgZuW2M1T35EeKq
vfvSQUz8EgElsu1+T0BQB0qvA96BpTokqa5lfMRXBhYMY1zs6I6nimyhc6jleWCSNC+PH3bxjI26
9lGO6nQ+vXIXxMZ6DpbhsWrzRuWwPMxiWZWYlVn5n1bLgCrpEKnHY2B5W6pJ1gLEgZQzS0aqKrMo
m2JST4hEozhRf8FL65d0X9wqBS/iNHxPdqqCaVABN0PQKld/OkkIqrlHVPo1xRkcVqScyFp/a5ZJ
HjJRHKSSMrVfQs8oD4kAx0aymkkHIhGDkXezRsos4uVu2/FfOqsOycjQ+2BRtMhcEZiYbHomPjIj
mi/6q/i12Nz3awr2bsuc8vQHNnpFvKvK9nfjFpWrP7dyS5rWA5cCt7Y1m9oGcc0iQP1K5C/qNlae
j8jnujuEdqhabvqUsrCJCPCB6DWpceP5dps96oLHlI9aOTunkPpNNfAvccR5KZ24daEPV83Kboge
XvZjN7+N0tH86odrJj8j1E9QNtsvwvCPFyzy1MDlKgWkOxwY3YmlkH6veT8/OaliAygSHqX57k5i
v2cyMXZfbkKp/9jAwAf6lkisJuNUJS4CdaJY9l1gOSAhe7+E1Nrx6LQ3Hn6lJ5O848PE2td+wmqs
Wf3HstJ4OmudX4LzipV4JpWZizBObG5UvrJ1DUgYS/xMUFThAqIIOR5/g6UJaswEwkStL6TA/HJl
9UAaBZuMHG3qnLsjGnxrntcarjClK5ZzEku8ILt4+H5J5J/8Ey33ruVhejgncIIVQ5jD1h8MwWNS
TacLbQjgA8a8m7cB7WvnwVKALgy/6ENmduO/wB6CBKCIIBubmCW6ePjMwDAnLvg38tG1MSxX622f
65DoBao8A6rcmNKtsgScTFfeMiBfxnb1lY9nXa2c0lEw5/vTcrjh85dLZfVrKTdhvlryl+yUiKjP
U7vQh6kqifwvW0YPq5ccPtG93Mn2LyKF6OOBXwUnTCF1oOphhzTvhdpgsYOUEtk05vfyB3BhEu1F
VleYvcCLYPAT4CloXErn2HN1hjVkCY36jAWovytoApLkjKh/ARbx5K3tZkSHiFz2/RWlxNNSegCU
g/dp8kYDBKs5cbLBPRfiYDrHrirLpeym8tFvH40r38JVg+ujgXS+nU1k/yiH4HX4tXCWoBGuP062
gl7qImPvq77EMHpK34T7nlHXm2VbwGXGXyhUO/+Pvtn/YxXZ/kiiUiLIkyISKqUAZBuL90Z5KLtA
KTFPhMCBQYx33smVKNSAI2vl28OCZdirdgulPkX+wgDojUmNjO6zuOXHcOqnftSNcgaAalXFTDza
Y4t54bV91t13iDSGnbb3MoOYshuG1t4iyC/+JuKgDjAoxKE/ec8U2+KWURcrYQ/KP8cPEpXA4OvO
BFd431UAsmR6bntwKbD9uW+bJG6En/3bw4NaylapsU4WHX9l9aRK0aCU2uSz5VIXY+QnDtXqnVg3
/zWaxdwJ0Y1xXW+QR1QIOBM82iNupbN9g5L7tDHUSLO6VXiTxBf4ikbOYcn7V7qiIJxNeDRKJSyu
9662D3W7lOHApbUnYQSRQdRN3NlKGjs/baE4+sqhxM6flGNwEEhC55BzK3a0ljX2TcyPspi5eGuk
xr9WBFSoq0D+zemw3bUkTjIBLicXU5toj35QJLtsCShexQcozD5wySt39b1xWCIde+BUUNO535sP
4BhPLn/tz5cUx0g7bnZofgoCSGdH8Nl68vy//nFP5ZDS3TGgSLW1izbcLL1Ac7uokD3aLpvvkmuZ
1wKqHYo3sNs0EfNu0jDQOOxiWtUnAiZfffDIthkrAgbPEb/T5EgeSApk+Y21el2cHgRNYsx9MRL6
u29DlzL6b46wa/fLvVbjmH7zE0vg+niIb9IL8jTo9vtM820/YeOjTY7/g0u0VLz9cjV7vraPz5Nq
UdVaeWqJ/ikiwknrfwejDwX9fiRunIlnMiCKTgkQS0IedUW/+5Hg4GtTKnB5D2o4kCrV+TeuIXve
RuokKYnwOpy6uj+FIe6GR+LYeFdQZD90yvPyVxJbd1qrnjpC51iAl32zaFqFJaPkhheD+4EQSxyV
qzPxzNWBXcwx6MFms0zcHBppAV2hTwYuZRZ5aERtEkXanMj0WiwLcGlTbJ6Wfr7J1OQfA9hBZWGc
LjYcfuqdp10sDx/DM6zvdVlkAyuMAWSGt1vdbtRXNkUBht298HiCz9bpFo/WATfA24OJ3Q88H84b
9sXUBBfGfL+nNXN72MC0pS88+yCNsD8Zr419bBwlZ1CBNql9MNvizSb7W8rc4HQzF7xrDFr1AY1r
cESZAWfbw4kGyJwaovFYna+RA+jUVjnrxATkXU0FYzpdfekEN+P4KiDqHFvaOagKKNbxCVt37h+b
C1KuAPQvDUfaI0MIcCe52RGYsv9Ht9EIoOP1E9Utk4VEIrqBEFGYyfsSCmOIdMDcgWDLiA5/4WW5
v6yuZBYqLf3qHyYRamWOusO223i2WcJbUZdtsHm6EYhbGG7mX/iHTktx9ehWkVhz6woq5/TZfUKI
TttuF9MQdUjKJPXBTi/A9dUSpYGiyx0MQBnuH0o8BqgY1r6zK4QmaU5ti50fdW41JYJ6CuMmPoMU
7koiS2E7yKNylmjuF4YLWfZHibXIMdoEZzbiH0byj4PM66WByBwSp7E62rb6yaNQkR+QwlvBi+8a
MuH3MNcHOkh495JQixJQ028WJ4j0ubWHel6iPivRwMElqet+6khRkh7rOK10s/FKv729VgWhQGvn
n6VpExjurVbGjYrkvaLPDjrbhpCt+wAHhxR0Y3MBXv5norUcK+PWXciuGZ3+nc/k7PAYKYPMzcrN
SLtkPPtKaXFNeQMmWp5VAu9wnKhsM5U/H1hrxzOY8/VfyiLeJQKMGH0FV1pG0HYl7Hy70s0Rp9Uf
Dtj1c7/lCk4e9KwlPJj/jYQDjbpHrn0zDZddCYwPculU/TfJnvIZMv/Vefyk4grL9fhXOr1Mk/0e
aqs5zvTj4GQpFIxJocy2zMc6I3KYgc9SIFle9lvemGOw2SWqDGHkoUcCmjjCOxu/ga2M7nH4yYWe
4vpBvSB8E1MX6mQFmVP5RSc/QnXqBUu90czi0Of36XDFNgpH0SBt9lg4v9OMITMQmoQA+bdlXkC8
OybOm0fPXd9HOlhfz/LPqzh0li4xioYimrxEDGlHSRrzLe/9LXVDr0feA0PebvYPNCzC1Lj1UQWR
PtLL9Ku5ozwOOwpPcnttKfcJtRTu33y08vvemSKyWlNgKga3adeBHo8d8Rrne0LNaUZ9eha93NG5
WjTirAFJ2CR2iwvCpYaYX5uho9nqUY0ub+A0HZtxYW7G9OMrXVdvM/j0Lt1Wr68a5ogvz4tGT4hp
LA88TQvgL56eBvDaA8RAEcesx7/Pv8APZfkLsFvfuMlzE7gKQHYiUVHRlbN9AqVjJoGox3VlKfjZ
giqAgqRT7h4Uza9un75il1mig7BwAjORz1CmLqn/2GPEfX/OyP3WdY563m6/4QeQWurTq1UoQmfX
tYYS76Hqq7AqY0RY+oX38n7EsAdpxr0uWpmdlcYSfMh2gtrUf39lSWD26jPDItxueeC40lZfoXs7
jEFugjmW+7pc7C/ahGSgugONhvQkzv80fbnEE4YhKzjS7gsvoi4jA2tovvBmspOwW+14eirivQEQ
m7MLpMCZllgNW7obuI+y2rd1mARLpHU4wcU1srKDC+BCcEjQAI0FC2jm04OalU0a3JqqNm96xg+a
srJ1eRYau5je1YLwNRz7EoqICjWklavN3Oe+N95J3G+CScEWL0qhgvCcW3NoR8vroFfbPxQ9xLfo
ZyR5PdGC6b+iX12Zmt3kBSa6wd9z0ntHk/nw/8r9ZnfkX6fwNKP4hdSQ8g07iJd+iogQZO0XUn0+
wpvCUTm8p9FQ6auu8lIJDSwAjGzF9zMusJVmheWEV3zr+7CWR1JzCMmSI4BNmmF/+rLMvbHfCBlN
3e0KrCYPezotrKI+a/SZogx1Yd/Hyr1o9K9prdVEpJXutAQCQURDzSeCD/Vap9/T62po25rB5Sqv
v7bdKqADk/qU1BYOzC7uFvdw7bLo3LwNU24xuWQu03ZXErQMExWhkbYdMovJq9BRHnkEmgpV7P4o
Uep2wuMBf5zkHrR/SsFqi3oDjVRqUI4zOesCbFeYWGEV7R7rWSjF8eGGkNs2osf9Z3NrurmV+LjM
0seX7QJTTb0CiRldrUxq8aKS0ykrXGPq/bvDpgXh/VJrx0dqw/4vBiVkfzsNY59PO3BpiVdgNhw/
4cMb1loXFHFp5L3Wgc4YlRNVWcG4K9hMCzb2Mz+/UhTilTFK4PsXDyxKXbM0ntLmoakmQ6xSMeKY
TWw5p6spkW3FkbAs33Crwza++rMBKSeXQQ+hQ5ndquXCAEHPNh7DTIakdmREEyKJWq/irw1QvSi2
E3u2F+8TqPYAZ7Cw+PHbwZPtyyIGlqnrQW4VGlY3AwDhZ9bA4acaDqRb1RFeu1147UGryZ62iGb5
qK7sqHPHOZrexpWHP3EMAs/+jlrg73px7RMhhawGzYiZe9YvV4iiRHiTth0+D8QgDEgnrNZPulQU
7lZIVqmGhcDU/HpplShvXFXs7an+7sxDmd31ehVES1BNnulUcdu14pezmdQ+dfDG9uQfdxyQ883I
TM+SV9Y70ab51BAEOzv878CBP2lKitsJGq+ZraOKm6ttVDA2G7yRx1vDLxj4URWcaWu9Rxl8mYXV
Sl7uuVfCKDS+AZ9WdV4X17RzpZJufKBU2z4pFkawzbRIu5fwl1cPLeme06poEdhC91rbaJEje8Px
T70gjc6clCXXNz/e8Dk1w9WP4q/W0USiVe39aWzFBD/Dw/z+NnHiv/Eqo5GOkw+j3GQbkGWI008I
cvlF0xnb60EmfFxv+Jy4AwdFaklZJhiLyCorOvIBOd4XeSs3JDTMy+Iy0Ok/lIH/XQq+tEmOQyYw
g4pdbg7K3WZ2ErC3TxQ9EC9C2STaAELBv/SpYkYKwtHMniSZqHgqxxgcq/EhIHudig8TmdxUD47k
Iou4Ei23Z7bAuoHRfjwARt//nLJIedvb717XyW6CiOnEm98qv5QDRDvLRzqhNEErO7D/PhctHxbb
vLC5oGUK2L6X13uLzXByDs4e/I/fYku+NLvLbwZh9utpmEYOuBzb2XaC3/mp7tyj6sePa2U2+VOT
HdWDiyFK3RvQLWfCmHAqSiqCX/KnfStggCcJyFr0pA6vzP5m8qtESRoa047WFR0FelQARzpD8DM9
RPbVnnzoEgcelV1ZySshsgEkFdEEL+l5bG5W0opY8DD8I9XnmMDBGvRFvnW0bvNYApmZZXR/zOE3
25D8ZM9xX66zg/oPUqBDLmMd/T2SGaeFpT9PoevUScNzJ/zVt+z8CRfVrMI+GAKD8hfXIUJMiNgA
qzksXsnYunAKsw2F9T2qT179a1Z+8cKfYrmeTV6h5TvAZwMrLDbFQfnK8mzQ1ZWylzlJcnkCI2EE
VONvVQZOG7pW7xmAyYIBsQo7LUytw2QqFs6N5fl3EcD8eUBwhaWSnTzEZr9XhqLwY74rzk8b1Ojp
8IYgRrJttDHoGGV5AA4/e8zbgNkWQbSB7gxeCL7wlzagwKZQCLxHll87cV8LwncqZP16T+AQRBrD
A10r6SJz5RYT7tfdmj9r6RYOeoIbRp74ymcmNVcckWKCSwnMQ7tPc3NlJ/7nEhvFL+Ixzuqcwauy
pKyVfSH9lpivopEXFIwmKPwwe7o2vioVOT2FTqmDSGunbSBmn7aVijm2WXSl0Bt58oWUWAHHBwy4
A+6R0pJwIbXiq5GPWdxMPv5JPcGS3gGOldHVG6qYtodrm34g4AvqcnTkgh38k0p4GWls4yDesz+l
N7u+md2+mxvr3jSoDY/W70Zbh1EPbMqzi4Ri900rzWl93X1CvRyW7jOi+ILltRz78dyrYNxFOXo0
OzxSD8KUeEnzzCU20wQuUyD2wH0sczb7c1X6MKOwwQqv8G6AXe3HW0nA2ocJkBCKH9JnNShBjgKE
CFswYnRLhr8Y/h187bS6AXDVhEkQhmQJXDQvyDPHYO3qdgB9q9YPJdMe/iQGF2ZnSmNnWvjqrw+V
RdapGnJzTRmotudBrxmPDm9GV2+CcMZRDE2Qv1epqjdy1QkRZ6w8R1hxHzxRd3LTQD1uaUpxZREP
/FSF773OLF1Nm4BgYk0d72EJs37Hx2B9hEXV6Qy7csIYNwCP/MGCkedRdBS2hP10XT3sSNLsQy+j
cpjRaGHiR/Kiydd2WfIObp1cRFC1+T1hoz8icTBky4YsthOS52ykqENb2Gz9/GqjMpkkANfYaY5/
LSXtQKlyR9CSYHUE896ILvjfxy2Za3oWxaQVDjtcAPu8IqKXppo30SCRTfmxARQ2nJfR/stmyS2B
7kTYAbAJBRA/CcHEvZtTra+3LYnQI9//g0odWY5buQfvTqDLgvZS3BueDQ/z0G/+yfwWjxCAFfus
Ua6JsWVgD3LAgUw5cOaHBOZuWlxTU1BUOV6Np9CSggjsqnCVTR9T3j85KiPHKy8A8pfN/R0Aw4SH
M7lccxy9w5fD2xj2pgzSEBqePLxw/lV+cOPoGLLCyrGDO7vBaM8LwSmXUchsoTjaIIJQIOZacHDP
1q4ZyY8TeQi17s9+bPcHdCz6nNNfKou1EPOSOBhkVputRInjVZdVkdFncasGY1HjNQORhBP8v1eU
os5bCuDkO0pcen4tOY7zgiALSlOgDPTbYRpDj3KWMzCxocIMkn/S2YMollqDvDoy6m5G22nvaLEA
wy+RXfvw4N4vm77Guzo8u5Spm0zrPoLRQBmQmrtOTU9/Co4o/ppw5ZoJmxKuVtnCIBnlmyzHESlL
jOrOXRoS5znBCzcZe+vuk7lH05oNOT76021IKJN7r1C0LfS4vzc+xYZKOxf5z72xxZrcBj5goLI0
sqztg7HMON23AhXAO4dBPQDDLzMbtabLMb32IsSaZdY6b//6SdPVfxp4wNugznV0NkQExdg6rSsG
ZPFSA+Xg0ba/yDKzGcnav0GXxxK+nfOM081ekrSxhhMIZXdDiqN9OYYdSDczfvmeuXNIb09M61LS
1wTzGuvz44AFpQW3gLgePhEON3nNLeReH7+Kf/82nDgexPHA2PP85VgIIZthLHfc1wEC+IGSCIH3
yfAnZzwz+4aap6raH83HqkdPgHomRn0MayK3SqT/F6x+da9ZUGL/wGmDVJHnBHJHTPRn1+EeyCQW
L+lHEIcqEcVn29DuifasZYt54HNL78JMMEIDOKbsXSaN2HRZcFX3gsnP15FCXqFdguLVqYSR9rEL
7FVkEg06O1ndYG130Hfpqpf3+Si9WjK1R54jq8AZgK/QERPMp+LXwpnb9p/Znitn/qekPBDVDvOQ
YgDkcGqLT0ttGWRcIXHmNt211Uc9q2qeTfC+VKvD7B1EfuEXlPEjSEByJ6ysk6CZOO1QErm3znAM
RCyzP/fWz7I5U3e+Jc0hmusENPu51lnWhmN7cwS5duBig36DTdeb/guHfQHQhaG/xkJS69SvptwZ
ozPUOKfdE8N0GP4nAp0X1lyxmKoSL0Ou4p3QPGlIpBpX12sOQuEbbLCjdxojMkviDn6tO/jkMJ+E
+F+PiTce9998yR/hi/vpUzeV0j+yLoUTR23h0ZijOAr51BEhJBe/Z5U37c1Kqz05+XciU5jWpRJl
XZa6NmXBAnsCe8yZS/LF91tjaP3qoQyZ0R6qj1O+MUyyPnRzzjZ6SJXo1WxG1aafyrEUm+1Srnd0
sXUoB+bbGqUV2lrnyaESEA1Zn47vPeNZNW7pwKrNcrStDKcSHUCfqeHjLlascgBJ5i3G9bbgS8bp
yyKC3KYP8i2TOlIXq/pdgtMpgbpQMAHSAfHgjoyoN+p9Jxf3Dp13cAXa86NPpDf20UCt7M6gaivZ
gs/Xtkp88WeARmD9/LBvAWfAdpapvjDfjJp/rAWg2Se3RYOwck7AyCfItEsYZPowCKg0FUk6Krlc
MhRCSR6JWZ+UVJUbomoGzY3kqvGY38hORpbVk/jb6ILrVMlKoIEjRxY9dfbHAI8wqlzoiV9Y3T9n
jQAfyjjsTm7GaDmYIbLq3RHXdM6ecPAi1szyuhYLkjUjiRFOS3BCa0Y1xTK1y5VJsVPrH/ve/oFS
kNIvukG7/9ILq2o6oKsIAkntc554WtlDyREtAVR6xLuAzVSJMz49uWNNNg3yG4Emo7Hy7Ds4rbRG
t1SvcL9EOsWvOp2a/GOBJNzcT8+l6J3uifWMTUiYMEupDObL/Na6qgtNulpOQkRIveZ2C6qmxNHp
Rup1+PH3paWvO/2lcLBUGKh/egtBxd8+yweHP7cNlsY5UULTpCAHLtPBcBv7R2HdMcAPfFgxQBlh
IRs0YqjFPKhXFvmlwyAI7FNyLFMG0caGzXRv/IWo+ITcyUICFE1pKzDbSA9Z8/fvhpjSBjuYtfnL
/T9oe+X+YrNi2uolKI33Q7Oiah0Mwjcx1i+/tmUWvo/JRaxu1auX4o06USn1BZrNJNjIRYqmWyYi
Zdzf/v9GXpLiVaNgQpuG/j1DJb+mM592kTKixd+3CGTbuwqhDd6e276U/XK/spQyydsLoDyL00+N
LGvsQJ6voIj80QHv0wdvm6h4lc88OYQAd41h5uqHoqa9/MHCeCQRz9hlcGwjrgHQcfsExVOD50qp
Zf0e4Mo8NvJbNwF5kazQ/tfXgu1nIVKkALxZ2re73EOTYbrTaJOUfRNn2RkYk6sA18TaCA3D6b8f
xcQhwbvJpduLpH9Xc/ohY6LaKDrs66uUYqduI9ue07tDj3yk5l1KxvEGVoBx+g5HkxK+nfANTf76
vGF5HuYAl/vuAP+Hk/XC68PFcDFkNH8K4WPsvwS6Sy590D3Hi5Et0eTi3wp/RISjFRzotsurHv8m
eiOFn2gpxce0lT1nQQTEPrYWtKigAO7lyypnekSG/xlbJxHtnIqFVJLjMNuJZ+ZkehLoLw41OAP2
wKSMg5OnJoJt2UofUGoMojURO8v25yvSvqyr+VdT8ygAd31lOAsdGyiB12cWij/BkRvP6vZNv4KU
p+fuLIjF4vC2wh5/GKhievBE+s/uhkYC9pad4S9briFa5WzNruUbvQ5VNDQOoXCvTzocZxNx8lNV
0cBAQ3qtXyBxNjrGUtuMmslTtj4XsHjReepwaUMLSinhSCTCdTdnB/nJi5T85BfI2eNxP4w7DkO1
+JJRlF4ApgUgTiPH218fcp9q+0iNsQvYJ+OsLfqgXgY8fBmoEGXB39ZMuDLgHRIpTOZmzJaNIM8M
9M9wT3/vHqgaEm59dWL7BVfy924QsMI1zTE+oEym2XYhhhSBz+lKT+MHBclrLjFBqVTtriLgmDK6
rf2e+nEqQNDeY++s9LUgSynqr7N1bPQVbjaw0f66zlSCQvyIB1ZSMR8bxiauh/aWhr1q4fk1Op+2
Jaom5H6S0KL4pQmkV8Jtbr6lanRSq/wVpHRkNM4chbxCUtKn6FV1/1FydMCGlhgQTH/l31+TshQS
/vM+btPcJ26ZB195ijvBrJhQW6cHhEp9ezj3XWajTvcWDYYEarDxxJljInXwPJc/juOcTtV69r1M
wcarPlEwDRwzDwW2HdfJn1mnqleR+VyuAM/MEvYZgzcTV4Av+v7kv4d8K7xQ1bRscaU14KzmdntV
S9tgTKnJ9dWRbWvUIt8Vy5pQxg4xgdsKjuZhIrWgzEG3sBLrE2+dPft/7iLi2Uv5zNEgOy82dpXM
vsNfWy2hMWyZ45dOzxnhdS6DYlsEjAeJTACBIH9YkDn3U25eso/Pgt2iMsZD9mP1ECTkRwBljBbD
VzdQARdzJkKPTnBzkhJPAABLb8kThulSCWfYl3SNH2bC0B+yTxXURQMY0Tv0DOvHTV9HaXwwHY0f
MkjhfBfLl/mPLoX9+/PNv79opbMOyFdrLJU3jQqmqhMeBHmSzFEIPQ0hrI8KDC367mBiUCjOmNJi
BkW2lj9152aZOF5IhatTesevVPdSsSwGLKnuZhL+FvcjDoTbMVrj/QCFwDw/U2pYb8NrRs5JWvRi
Is5I+zPmG3THuC8kSC3Bu74xXdDEQk2MhAfhefoCQq2SslZ7JrRq7MHK/1Lv2mg3HJU3PPm5CJw/
7Il4rTb9F1UkJ5r05Nu2W+r7FTI1qiMSgGw+2iIi30TGTjF+eXZ0rt+RBu4YrX9U5mkxD6wdWcBm
UikriX9XB+JxT+MeyNFSDudlXyxTe8olWOQX8crWBMxE2MtO6TC3nhBRkG48hAIwi6JRaMQK3Ulp
QE1FJAbU3+vdRke2kOgiTn5hBgUdpRBSMJxkqNjlgnTlSICnVBqBFnT9NNjfenT1rJ4mpJy3/wEW
HpNfT1NuRaypJvP1w6RWp4ZM3BxmOKdNdqABzj+lB3c3O4Gbon6K5DrVIRm6p78utJKWPwGHCDnk
rAG/j6Vrm+0Xq4ZSlqozjj5bRbKtfeF8aQRmF1t6SSTkEzWmQr81Ue4UnhVh/oBl0QqU7cBjQNpg
i+e0oOj7N1f7TOhQU+G779u3Ss7mcO7Cm5VNPUqP6OOWdPhcSF2myLRqdVr6I2uEPfWkwDNTGZZ2
3y2++3C2XxgA8VtzPhWIfvuzBzHPoMjmNZ3/mEK9oa27/yRP30HZrSmw4A2EprMctOeVjmvRk8vF
9pvi8W1NUJKW8icOQj5vAViEebRMNlKs/nC8Rdr4NG4ROZuJSaMpBgC/vGVh2lZzae7IQweJvr8j
4YRz9NB0JghD8QUiNON3uzwoqm+UFsImh+lMiONQSwP8KQwlcqnS1Ku0hHlHigIeLGVueasuKiNb
JnOfqfN/3hsI7MWt+n1tHkQvv33Cag61UR5d9vYfaw5apc81q0tW+8+ZYPKh9PV+/Lbnjbt4glRL
wZcjoNzBtDRmkUWUuIlu0J6HTx26uJpESedW68h3CZgjNtCH79J0mrKr49Rxkuo5r7iPjGWyGMv/
zeKEbh7d3OGTkEBEj4kykP7BdT56KhQZgH+F32jRWHXRwYzvrX/F0v71hdknZ6K9Ld3Cj4OQETbB
jkFNvT5R81cFnl/ILDFn+IPByLq6DEj3p696ARn5JaGuC7IcMU2NUzdV1Btuq40gX8TBiLlnPqq5
RkQMZwz6IoZLOauHXv1RsjREGTmDiGzKKzmSNsQ+GDJYgX/eZDI8wHDZJ3gI1LCZI0IttYoNTBTe
7l4My+5jzKCpcdUNzM5BPBW1SZXIt5qENuh2O0cMg0rR+AHeOAFWDBtwB73jUChZUlRmgqekVUhC
9vUtBrNvG9C6kY9lhuqb+MbpDDaoIHYJeiq1u9gtNmo7eTUjypV4VvpGMrYBJ9JgUSAANrWXfIIV
NeTsK7am33/sjhvU4rsJICdyXM3RVAj1gsWSzcaG27ivmeb/y0PYTF7mI9Kc3vvJQ3ATJRp9rhZh
MjOo6TrJuckqvwjNAI9EHZimbZoBrL2glcK2q5dSu2aZjEW+3WgZRpUgiSDAqsvsMHRaR+TEwIIM
rsfl8RUgADzUBlyUzuxscDMLYRNWX6z30OiMplEYl/IWbg3iVJFn5KKsbnZdCyOWLJ3UFh0wnCkL
6BavinsAbl2NbDM/+/Dlc2vgYMo1vXW6YOIvoxLruLKr71R/XNtoVZpHALyDHo9/vtTBnlDW5Pr3
Bcm0QvBGXaIVu71pnQHrXtb9Y/bybUMJE/ri51J4nP1CLNQqPpmyZxiPTpNFbaEpvPrSPW/+ZpeM
mefmrhaoOREGpSMT8P56PyyKsIjJ4Ik14CYXOvkKN1XAi12YvPAFU0bYIqEJLZteFXiHHx9lS3is
hPIea/Y760JX9dPoHV7BOAsaETGzrZ67omvo237RGMIEBspg5g3LgjnvL0CZnbcEzxZM4+sFJuQY
1uxNHrT91K4N0i4BgMzanAD23ajsEjiP6mEMfrfbX8abjEm/afEp5v5K6u/7aseR+UBsGg9b5A/v
ns7TtuoZTw/eB+RDsiMseg0JZSCea07oW0wxR+I9GCIjvd/ykwvcuG6YBmykGWKG/9oEPRi09dBQ
v6ppfNamMuHwAnSpTj8L31+9eqtvuoSe2AHNxm/N49ztIFX3FtuJg2pn5VFKr16/cpQJ8AEukzdC
4VGQVXjaLMIlcc9JFHY1KlJ8Bpc/CA0CePqNXBm1G1C1zGKPt7jkhjmZn1gUfb666SPphVKVHjvG
TZlgopI4H6w2Beu5BmhQyLsF5lkQ7fJCX44cXHG6Tyn5q79u7moSzqybxU3zskjK8sVnfiDmePE/
qSgPLzzpmjg3GDfuw6rEN+3FT3kNk6F7AR3j/PdoYnHf1es2kvZLAQwPsIT6wHRP3TNt7k3MnLs0
k9oCP04Z6pDq2IgGdVnRGEwmTunSIRUwyk6O/WO+DM9lLB7WkAeaJLr5TVHzHrFyS5SdT+qaMq2h
3Pjqwa3jbg0jRGFMNCyk1KYSceAeTl4+CCrVFlwmslW+HJ5nntThqX3cW7tHFHhHT58LxeUw51Za
7g3h4LV7NhkJ4h+5CkbxqSB8rdJYfrfd4mZ6UKh+T9zwVyYUUVBej0SlvXWDCQxWXC6vZm98OXV6
9n+v83rYkQbDhQF/3KE/dRjeU3HOqWj0QKgwK93EwRBlD5iFnaaspvxJ77dAMiD2VLlYGhQx2Jv3
z/J7xG7C1FJWwNcKRHQYLZkE/wyVoh0KbAwzzI3+DdDP3q0pu9795qI7zmWijqm+EfQ6jZ6Uj+hg
wb+cSZ49W1bCa0qFSHdVzLYSv8ww+svfaN2wBfSHkKxp099eTXCEOMDHDFGyB9KUToUpfXN12sW7
Ipdkpm9mMI9Nvd7W7Mx0LQXLSKgBtfFs1iXjlrQeLX8MMFt8tsguoHk1N/YCfhSl8kQEiWSNeQUc
W8owzhV3mI3w/tbLi6k7041uSvCbvLL44sYub79iIRKFWfwDM48pMV/WDe90p1Euhz8MGTPXRK9R
QMDUJkDgRQef7zTdhdNsSRMvoIj+ovKthbZ1Jh0/I8RcwWUejrY3U1iGClxdSEimvm+SYXGF394H
IC/RIbBLLVVbZnl+WVUycSRyra8RNV9Zy6mRUlTMY3F+WraDQ0AxwuLVMLnu6Kk5kACYSkHUicR0
9TZtPPQazmF79T0orvV8XxbZZqUI1+M27R+7vsi++GfAR27eomIbTEfcXqkAwUTF2ng++7MYl5Zo
4s4J2i7GMS3lN+LD6R5B7nwjWFN8ckwMnHPE6IQLkRhfa3bU3uo3F1VrW3MC3uvmxAZULYlT/ILp
GiyhtoMj2/euXTh2JUQQvSi7cur1p6DG3Dg141h3yhFOu3cjnqXLf2XN+b3U5y398j0xjVW8tZ79
3AmskiTmL7ScSVvXGHidLiTKbJwJGmwvsLRmxCHjqwAby1+VexzF4nJgeB8mWK9AJSJFKghQIfoh
mGbMBlhP8B26xjTMuB76fr9XMdi26a9LG7ofSebg90/9io7bNQxpCxp+ThI5srFnyNKvwoOp6asO
agDpNF71ACPnDr6oQ4ZbnxgSSXyMrBD/9z4doOjhntlE3fjVP/xz07EOFLseSwX+WebiVt2zrocF
Vp7lZnvLFQwCsNYeZfWoCtP0A0ddlzbI6xFjgDfF8C1FkiPmgfwbKYFz6SdX5OMo+8LQPFQ8m5ti
9M8xCjLnN7Z5AFqDh9oNtmWgCVjCKsakNZTzMNkmFUuOrPWRgO1yWI5pgeyGCTEqdwojZ1kFzRJ+
16dYGwSQRQBjeMMp/RY5CTrK9/UWL2DMEu6hW/cimqBAnSezqZIjEOsRb+15iN+Q/KU16buucZdN
Tx4fnWwMHAE7Rl5VtmbUbQ5ZSUwdsLHxkPknahZEO4tYiaenZsG2VSC24U4iY9h3k9m+QSpMKoT5
pPso40cwyneGN4/DJoMODhQv9bWqE+1kkJ8pUHGcLNdh3SnKfkqm+Dd9xtNf/bCdA7MKldr4xraS
CQuEHZJR8nFxwza57spBF6pkDB9z79w3gqBuvGdjrOC2VZzYSjfMqtaG6H/HaFvT00F9pVJRC7pM
DQEtEvzL5P5gsBp0fSmdYpl9XvncKwokSyWOIzsw8MXkLiHBBuQHICKYOmwijGjOC82VR21UM0oi
z0cJCFLgoxT8BT4XMvVe7hIWbH7/VVuBxFTOIPnquxl43a5s7amoKo9dYGqLz41NbJH2HVHbi7uj
AaEdHfYuT/7Su3lmfkzOqrROeP5NUoxQ6z9JKeNsk6pmstJJNrhiq7bJyT9i1GA7xKTMiH8L1tyO
iojVi/4VxMepj1+iosRCq+k+7HjL+SUqALwEGpZ5cFm5n6eWjXhP3wNotxbCVxyZ0CCT7m73Ifyy
9ngKClSX6+wO7cE76nWcOa0gMyN7tEpv9lGN2IH/Fyir+W38DH7qXXiq28OjCFiSzGLCggyWhou+
O108C7LKW/vvWNbyIYvCBhQBlhPKIOHs1YzrBg4rZUArQpdBWMUokJmVl3tZB+vXOYHzwqUyq0WE
WmHovP6cHO8jSd0jTdYZhq4DNIUCc+HFEPDMJNpzoXG8ofep85MAU+mJdBrdgNv7tgORvIFeeD4N
zwlh/Xtm5i3RpJ7lfY9zUKfmiq6YGZC21+TmQbl1ex59buuNwiZitT4nXVXh/pfdrUL9Aq35POAk
Hys82MIiVQPrILEmYpcLqpWBS/0/Ia74HjQnxIZJEQmzaV5y4uMAdwNpN1dZCmcs1o7VHVnfo0yB
FZuG37UOVTpGu4zMufpO/mskPmbZb8ERMMbFT0wZF/T/uDxfGHU+uxb+kaA8Pcu2H6sQSh2kPISd
/Zx/cczRSWq29sXLZ/9OV/yS3eUm+7exCGhELbWMhSQb9YowTXe133JphEo/sGNRPUBOh30obte0
N1gXRZmWW+BWMS4pxTOHhBY0wwz+9RG9/Z8P5yYc+bQWVKf6I0EZ0LGAHKli4pUMTEYU595jMJ1l
5TM1RVHqMSMlP6JDNdAUyjqZSBhxC8kgKQ2VrvdNo7Wy1tGEd+lQYcUjnTtmDvTgV9eKTwkS7vPs
ow1TA+1dQN8j2vs8K5Qj9dHnDMoVQk1oxhIrCXdswCIuOPG3FcMnJm2Ep1c+AOcsrtb8455cnJdb
QLjilA14IqW7RtQ64Oxn4l4eLfdzOX1xMljnC/r8QuM8e6SZlYoWmNpMi88CY4ClnJ2djbYkYJLk
6e9O2SnFMG5gDYxvMprF953ptMKWtLqOKvEoyJTgbXVqtyYmscLFzrnfkNnYCmi+BhUPg3zCMdaL
fmQqVh6A9cq8jNNmfN7GtifbvbxGeCwuKg0Z9E1i/POMO06PXW85wIzS059ZPd4BDesmH2O4N8Up
6K0vwHXj4KWVhZpEmnbGFmAKjegQA52OpAIw3KS/1EhZpey6QnMwCCcHcfHzMj8FAe9L5CnBNs5g
KsBYs5N0ns6z548FSa6hcj1NdHno7kKeTnynpMcdWX16YDxG9EiinAvM5vTfN1RBWOKxkK6WxSq/
8av3KxFsmCqTx6UvMim5LoIiBz6V+5bGMH4XLUQDyYt0fn6C6hNfVFO9ssio9IgZx0uOjhEly5fl
z4aoOqCfM9XI+5ciIy7j6npicl9CSNlMHeAhO0QC1ZpYNd1oyenQu9cbIhGqmaCyUrWH4OebUNzX
79cSsS5zDLd4PCvEHK7QDBDEKXfSklvcEhCn18mSA7QNW++z1XmNWd6rSXnvBmxXIx8vA9N2DLfC
CdeA6dxlD3/2zGJ/DOe3DK3OdEAleN0V8t8BxE8hVTFFJlZmegoLPQaQKlj63c5JSxTa8FGgMQr/
x+PtvyqTdbA2hTl3pqjanKsxEqp5tmCbn26NgW+jFxSOTf2fbvYmGALNFeJkeGk4+RXUPWJAepuR
VLAqiYZk8kV1gvwZUifuDluBboI9QmlNw2HF58V4C7B2b7LVkrREZCQsL7IFvjhvIMjvYr8X+qnL
33rZ27FqZWBLBwgygTWAhP9kgrm0Fewx4E9Sr+BqN5MNX4uMtxWoNa0B7v8LAqoe66sQPSiMF8t6
59AyUYxlbdhsR8mLNKk0jcEYoEqy8mKmD/iJhk5yDds4X9doSh5yRKv9m5otvrByRxli6fzrqaoy
07hmf0zOF6ZQsWcGQn1GGjih+SjQSkxFt/h9VoRfmZ2WiX+F0lqlH0r3zU13I8+ce+eOjWfz6otR
8/a1hxM4OJS+w+YbHJ+2aatw0LcN2LxAkqPzXcDsvfHS0plvsd2mN6vWzcSUK6f3nglQzqA/FlLM
mX37e5mEAYajHOkUtTFLBNFMJ/hae5hT4JIbkYNgiO+RZZidxzEM83CDBhOnsRkC212+k5jDDdVm
U9LebDZSXmoBxbFuC1M4ZrLogftCIxb2jOLN0llc2YbTxroql3q4TuZNYyAa9+HdZkkRCWK+hweN
ciCLFC5/Ds14FPGdtpbqzsZmiv7atQl+q9fQme4xo1YA83Qq9qadrRr0jn+V/IRAoSgbS/x3kUQb
PD2LEgrojmVilo2bdkgwyaH7NIIvX8vwWjPHTdKciMy9//SqyGG6qgyCB7Aoezw5yu7CJ1+9yLb8
B1PDUsPfWNhuLAflxshxTocwmHdKdpWLOPL9aDP4O0A8UgKqwXCmrLZUi/pl7p0Fgq6aRrw80Nhh
ZFnqce0lb3ubSpNuoAHcafXIz2VA9Zin85QzQqqTTUznppdIb3MwxZNCY9BGZWOzYN1l3DvXXTzE
OaTcqPo3RwSdOfm+u98EpPUXzhu2hfSDlmk6+wYwPJDIzRXM2oLWVQ0cc00G0dxR+w1306lYTxtf
4YHfM7AeGeHgbBumZdjvHssRK0tkz7IqVvmmEMZHr09QlGzzWC8bTeKqXjIDw5gmENmbPCYWmgx2
4Fq3z+43BAeFCec/qXVoD6s1B21d9IG/UTNGqc/Y072v7s1I7xqFL9aEoTGpjbC1tRaJPcBWXgSb
DX/TJycqO1x3vMkAXLUVFWZQdHB2UwhroHT+lsNKIwKFcOB1CyxggmZxT0LdoMqiOJpQDCYQefWn
qVHPEnN876X+D02Mj7H9VJAoBeuPohfXKM2nci+bpoyg8RxhCB3dVoyctTA2WPaWVj1ZEbfgfFih
eY0sN8fpIkAED8ZmqBMS1iRAE0CmVWZqS2nLZF7FDD/XGykff4Cb2k+6ual1ESWvTU7iCEXc8udd
PzqodZBshIG3pUN/mQZS+3ZWQGx2oGEEmyWCY5rHqwW8P9dKCs7vWfUmD1EDI9Wx8Jn2MYGRlEwk
D2RMxI+CxiZhacsj+id7d7Y8uA+jOuXxdqGvXSdhvE16nKOT/xEW2Bcl/Sj2olNgv2k67PAD3ndu
MYO0bVxK/XiTdA42vsjLyV3FLIffzICpr8pDruqXBYS+SabnQDa1FVH4iCyTX7OaTWiq0U5h/OSU
iCWedRgirvQXWS1YkHfXPPNV+wCelnQb2ruitIJ8rd3IRGrEbju5yz8RPMZmOyrIfetOA7bWq5s9
7ew6+lbakrPH4MEM8tisNOZHQiMa6rj4dPQ8wnGfjKuDvh966kADS8UVvcZCeV5DX7L6boPtchRu
PECuPG8k3GmmiqTIj51chYqu8MjRyWQIT63+K0Bh5ehV16FBW5BxjPiW4/WxK4x5zWdJi62lU4II
YSQ8aufNY6X6eYZkPKSfbs9Wr01/fRpR58nCnFj2RdITGLAOrMpiGqgu5x2/x22DskG9YULKoQJp
llR6MuW3RxQ2Hiu30QWG4SElYjRGINKRjGyCHsaugSy+bsRUoKE7Fkl175TQ8G3U1qPcAb6oNKMC
xW4+XXPsELGqXM2KtDqxwBKNjsNwGIdj6ChJPmU3hEMKXRmCBwzDDrlvljBVFuUWhe4RQNu4RZvF
ztcjYP7TTpRj9a5wux0nRkFPOT30QWf2Pc72lmdaSM04mQP738aF70IUAYVDRYi4K7vZbiRNQBnA
euJgvs+TqCOHltb3FRg+UDb6b1yyC5yT2gAChqNnlH61LV1231rNZDmcuySwLBWsiVPLicq4jZ1b
qUOvCFxmfptsNT4Fdot5DJz6xwDbAYeTkIJFg5242YSlriU28htsnpIiTaoXH23SUE68ObZwXAie
RHwkRj/dyxwYdHNVsKRwuTPdsQ3RCI3H8+X+GIiy5FOQyPLc4Ml1o252RVc7HeEfPh1QwDfxvS50
O77C1bIjFuaeMLY6V05uCk4WgI4l9sBDZzqOElmS519VIULiFWurbFQkIorbSbh68Xd93SETSOyA
gAkOqWCQrS7fcnJtNZ0z4fCTHjgj1cjKw1ZdnQEhUD3rSs3Ooa/cZMClk1QpJ+bEOUJBpAcKr4Pk
up012szN+ao0qcq739bPzeOGRJ1ltKMCYueOs7CSerwA7GrlU3GLV1IkEG27ynupLvXK1QzN2NkL
drulK5++Yr7nIN+W72EHDj4vc214jr87+dxF/maar5pxE6JNRfTgvMSG58me/0exPHnHMEZuI/XF
0xjBTk1Q8JQYxuFpAGKKUTtcZLgPrqfrQNw7EtJCj0z73TLyM+N1rd2pGIoSm0cjBKY+HLGYS7+c
SAklJ82V0Y/o+ICSJoGDO9TrUpjyKD3jhCPudCymi7KpOt9R0YW9quv/YRD4dj/I0OaTsbcsftBE
cNBcI4s9dzkwDpCtajY88KckKSvfJjc1rI32ySy8IHDRLuYozmjAPlHdz9cjzzDzQLz8fkJut4wL
wbHfiEmwxBDHmQoQ7iMgpiaamY36o9Ixkda2FBnMg7zvazLFHHr6vDKp34ZK1t7lvAfRwq44Somi
nWXn/njusEjCJAuiF5VQOy+x0YMdCVTNFqKmZh5djqxOv1IIIDrlNuguqGHkqq8iZAU7pAHBPbsr
NqhFzVpEMl0b4r6Ukz6zIgMLZB5pIyrranT94MBUrCjvI9N5rt1JQtbvzCrhVZ1sYG43XzbDLYfS
EsvyD5O5QJoBqsS8EGIQDyx9uj2Kz1A7QgySfsSWwvEpq3WYKu/86uCBaNQqd5e91M5S/AwYAQlu
BCwXHls5Bfi0A0PZ0Xa68wmiD4b+BEy3A34eXfvjUAg3SdwUyqFgE+XyltI9LLAvZlMzIK/yv3mg
tazzU5oE/k1WLx3IkK1c+KcwEHP7IYMoDjPhl/Ro5qcZ32/L2aom7xwgggr0JFTyvA29+Y8Gf0PD
XRXo9UCEOxc/OHedmyrrg5+MX419eejDWbdtZ4nWEokjpxnB66ejUmconq3yKmi1zXWjG54xAgY6
Fcxp52qaBC76Jk9vcRfCWptgX7cMolqH5SBGfu/qiGpDlPHRoSVfPUTJq1YEJbZQQr57Iz3Y0qz7
LmjAh1jz5EXOwEaHCM62c7phBvft/YX+O6MCcW0zjCRy2A2qL+UTZ5uB1ctEKPRd/h4cU9XAY//L
NEBV8+n45S1mPos0lLhkx9Ip12PkeSSnQT/WAmk6qrUUT+tHn9mlcVVN5tpEibq538R7rwqYZGiS
sRurtponpiRJrWxwKbVAgs3Cg9GBiyCTQWWcu6vlXBYHs+wEGoANXGInpJETUDY5Zjg40djUIUts
nWLAe5euUHFeykh7dSXuxzQZA5WCST20e73NYnX1V6pt6wons85t9lS/Iwow/EWNHeFQGeddV8uX
SFZJM8GnKo59rx7NIvw/6O145IT2FkuQf9hqoe/PDMOJYTVYjf7k1daXc2eZxtcgiNsWlcmIV4++
Ic6cvjaT/F3+Ejov+5lehh/tNRGm7jj1jwJDxDhLOaoBXl1/cDtioE3ey/ku7+Ib8JbEj+DHbrkr
xlnQfr8it7zdrpJy9PwSnaHARvC0Dqabvj5xxRszjLTu220rGE9eleMYTn4V/lGMSFDjUPSdlg5O
tD6ObQ7d4MqwANAhE/UPkXDgcHVXdBq1ZsgY+ImRZLmLFB2MMukrnZJuGLgLDfksKOUVV2jyAArb
DDeFbXCTzkqFIMQQwu14NaLWykC/QToQm9iBhu0MNNXrhSr2549TAwQuLZFZPiKltV8YLuZke5xR
FC8y5hdNAjZDzRTYu4dKc1Wp/UTyih7j3guJ4BBrKhI03S22GsNDw+g4tW6YmfmImWrgp2f9tZgI
q30mTPxQyqAH9cmN5pC5pBYyLMQm2Yemq2ngonJFrRiSiK+XGo7uXyptpJZB09UifyXBN2BpfBJh
mPs9Po8/37eGm56k5KyEanp4TOYoMEJWyOG1MBOOywtxhMCe+GYt1HrFKZrTFT2PfvGa7hjDIyYD
OeAlG7fR8mKkctfw9F6WHBc8t8byRx6drG/xmyUAxPlq2/8o/pb5Ntllcd3IwOJetgR5ygx/qlU3
aoB+xTdOmZlu2HOZnBbCVOtJy+13WdGvh5jU08UbyzUf2f+hNbjOJVaLUT4kpNYk2rU3pnlYSilr
7YDSYOwJt8+zRWyNRsALFGUx3JLz9ihYDKpcYlp7Tl9HJkOUYFJvkPx9TPFBqaI6pDyIsCC21jxS
A/14QI+l+2q2ig9nKL3QHDpOTDtZuv0rCBSwcvhzUIBN4mePqROJF5oVcOkXGfrF4YQBPlTrMmoO
0gCjum77GZP55HJdKQScLWh3mnbNu1vmCpukjAR4iwCP6KQEaln5KqLhCfF4/7ffXGqHhV3CNOPg
vC3VZTnJmGYfqnz3FK4MHY2CSIKWANm3e2nvEpfoCEx754vggnSImei/DaBXhXE0nRTJFxZ4qWib
GnAJkxD3pJg9gqpRpN9VpaZ/en2rZd/B3l+vjZGZLzqlTZY2CCkaDOSxNBSR14BHHW5n3H52g5xO
ASQ7WRF5x5rXbllRFx3wDFGoLKAHZ5AcFZGklEVVmog0JURr5lp9LNBUvU42OliHjwloBarg8+u6
JyrEHwNrJZFGPrPBbKGJRuza0rTeTjBLuvPTl46jOoXCFiRfMKVRR+Z+yu9iVsbyxb6CpWGk8O19
1sXeQlNt9awE7azjmaU0ojaUCLM3BivFbCuSg489FJtzSTa1BhgnOR9gpEngibdXcmneZkke5HDL
HtcH//RF3yBdI5Vhsr28DKlXv3vXIJnKorMU/mMuk3akm6gspdQCbwXMlb7nMYUa/4pgJELhamU1
T0WV/Il7+bVDRVv+LEU/hKFjfI99BohnvzAdpkV5UnxHWw8d/Xcvx2GYFt7xiwqtbuIanU3mYmNG
KkiHmq9RjzqQMERVVnY7YO5BUezHTtjrOTvmRVDQLYp9PMMFNpVjeMcDp5ZpbcccBZet2ZZLG5PE
thqvrPhDgQIrl0RRG46h1OT18FnxjKLX2/aPKreBaAeVdr7IXJfA/Wy8NVIg+A4JQgjshUXkS/Lp
tlyQpq2ECpCnsdlmvGvqrqlmskJz1yP1Xo0QEpn7bKIs6jX4h9QfHXWIBdxMDVGBFM0xM7qQ8yom
0w7/PCd95XcZ0Mb3odVuvhhcaR4LbjFY6vlzF2XVHf1nxG52mtHEpylI/Kb8zwvfZY7NENx+0WIb
Sc7NOjkb4elewZhc5BKI8iJf514W7WXWbjE8NI5uPFy62tfLhENGRYMOE78xyciIf9YbiUe9elln
icJwv9djdZyIr+uO/dXjxyMHFCGhIrz+zWr7eFB/ogsjIpEejXXOVzYE6JxUa1qrnjVM7unJA7Jv
PgqshDW2OFv/Nr0Tff7ja3XOfauJR0DuQCbGtpt7OayR/eENCX35MnF2f3KLXUZtX7BbKvb/N+fg
PqslO3hphq22ODvmWRu7aEfM+MNE+IeyQHrqtgACJ5/hF7TgpGgu/KoRDCmLuDBzlzJyf6i5lX/B
nPly62ZH23WoOGksKvceVLPFK17gqDYGhekO9HRgcLI0imdBBxPfJGYtmPflK0+gjZmY6OqwVt9F
641akY2oybUdQ86ssVSwJCFGFn5YtSd0mvCh5X/66hBIDLbU6RXFFrru0/eerwUDYbWbosRxLsRa
ZhMQIykmCrSibRjN0+hkhMjfRfNcyyBjF3+ng+go6oK+q7j5FtmGXjM5EBPFqpH9gCTtyXTBh2D1
90blEcWtBe5wD7Dfti8++jpM8EjPskx5RPpRmTQa87ppmHbB22m3y2PTPuVQGOW2SuC4XGCIl7u4
PIY8pgUMXwlXfZSWMkruyAYXh8x2LI2vRyUAEPn0F1GEL3m8EYM6vowPu5PhMXs+hvf7VtkimFU6
oaxIZJ7jBjckDy9O+jwlInp8ttr9tKXOmcnL32dR5bNA+JwLIeQD63rJ6JfH2LM3YHKoEFcSCU2S
IVM3k9c1hLLoQNKGg/MQNJWphG1N5SgQqRYhuraVXwZB1Ab2EekImdi4RnnlDascftvsbdroiciK
3rWhrI5ABDZNITDNMNoFTyM3DsxMERvvPSqYAS3VaYKptw+71y6weeQkZdGTr1X1hATedtx78hle
zizSeTIAq8HZYONOjOGeTePkIml8twUpA6PE8uCwtrMLnRj2YFoqvFBUgtFx0eQ2F7+5tEGmiDgp
g7TO2d+x6QlwSTLQbr+A7OsIQic2eHsimC5tOh6dpPzyxmEAN6rgBdwv6FS5HKZrXnmpt82m5Nzi
extQjqaoNilgCHdfRQBDdDNytNsUPKIiL49hzwGY3fQoH8lGfQIwv/n9hjxKAqa5QEE0LZdMR1cT
D8gbmRpOpvAXvkp1bqOOq6BERjA1m1Or6rvnjeK/FKBx/utQ5rO2czUraMxub8r9TVd1cA07byxT
RcO4C4h76fS8OStK8SCqCTRWHSrXM2YJ2+jaSfjcUhXcLrPx7xqiDVfZivIZY+KOZrtvZGQ0+/ci
qcQOQiiqW/8k6rc6iVXCa9vaCEaP4cmt1JGZfKWp0/gwotZnbC6fm8FzeqseZf0wezDKdKhIEone
MpOZ/wf8cFtGCI6gRee3fKGh6sjD1JX7zJs/AfS6SyDzibJNDRj4tYiMgWP9nssHo8iiKZkkt7ws
Upkl5KbA/R5BkH7oNY6Il2hn3OAauwS7KTeCSO9mlH8yyhO9+cPR9QwuXif8ObqiIuI3t8ylVf3y
VfiYjOzNdF/cA2ZVNGFG4BlJJtLYFd+9WbXBS5x/yPyHp3WedeFBGwhcuBkq56UGoH1nhFZMQAZG
l/rG67HIiI4Ui36KvR7FTUaF7qzYNuNJPDX+aWtgkEE466JgXsB9k1PIzrH2kk/56dFWrVhLn1uN
evBkk36/uh+x3yKtaIUWg2DPqr5aXuXUiJJXJjFyJB/uJdHaesnAoV316xZ5qS7I7ndCuMn9tYvK
XRptMbnGMyBmmavy+vKtUdjnGvllqk/wFA6iYR8xGdctesgq+x2BqLBcWBPOnDhOKrK50UajQRMD
55H3tykmcb16mduoFvL6W277CYpV0D00DYlWHE2lnaO3TF2gDvWY5lFySVB4KmEPg3doW2hRDH3f
PfsVfnbrYrGmjNfChhS60/HkJanywkHaiqccbrUg2lnZ+myYAMAsn4LnIk+Srd7nB/WxMc6qzr4e
PqzxAWO1eyCdRyzUHBrWjwztXBdLGfeqYaLIK8uIvHSmDimPIi9oK417+VG/OkJB8VdUMXvDRg1b
1aZfck/hjt1CXcJT5N95KUlKb7NJQdeJp2F3l1rNsGIADBWk6QLSr3FYvtsS3I7+RIJci0haNrqO
mSsglLW60pEuLVNoc7n48b71dhTfI3A5FzTmqyOiBpyOxo6Vv3cKJG7+W+z9SWoe3EDG8Jppbj4V
SmgkgpHHZNhsJtkm3zXLH184tzf7ADwFls/XcgBaQp+w8HdOdOsYRupHA5svGwTJ+oA1u1IkTnYr
y246BCb5wLvF3rKLDyCLPgKXhocframED7N58BzROm488wQoTrSyAj22O9Sflk1EBj2tevc+wkIX
UphNUCPhNNJoKejKr/keKndQnDrwQNFhA+UDqM+AXKPwGgaiUXnK9GL7hMyNi6sipCkDvUV2KlA3
2B2V613hoYIhrLjQ7GS8Ce/Jbuk0CvVxpQYuHxiXRaIVYc+ZqJ+IDG21eDC/TBylDmmr566oQxb3
oRY2yb/5rv+Bw2PlZOufuHPBz5fuZ0YFBqRhnAOdOBXIzds/2SEfgEJ0AjZ3v/Cem2ojziuZj3SE
mUY3uJpUAF0Dc2YA8LQMiflEQJKMNK8PGP9/H9gcXjEv58/dtLEBf0etGBZlmSj0pwAua6L04pmn
o6kgd04AvPIOtOLN5dqhrCj+GhNjPIervSPfc4t7UBcetbRfWjy9dallfeQYMd9a3Q9s90+nrLux
TklXbRVRaG4bGZJ7YhQ4OOKDr756KKdLCbsXP+kMW2n2DjeJ3hcQmb15ADPjWRmbrYdLH3b5Yfh+
Am6kCANV8rN0AdSEaG9Z1hMU//NpbI8t8/OQgiaz32BjU3t3kdvnLzUGHPCBX7RhkvlXBcKTNDPY
2sXrZ0zAas+W7aeu+0tJvWGmWIMBbmlf5GAYm/iv04e0y9aEunWuprDfhscAR2Y3LZcL8Ys+b2T9
KTJ5mni39BOGCECx+Juyj+fBjUkNxi7vWQW6yiA4T1Xhw4uuYVy3J3IFbz0vt9/1funh/6cfJFNL
jiFpjm/cwO8CLNV0XFmKaWJhoYoaHzQ8BKvu5PSiqyBadBN0X0LN5kv1Zn+sInE7khc7+INWVFQp
OTr74QW6Mv6zdjbInG050azaasihJXQHCdhBcY2xmfhEapWKA66+sOmdpdCQOZ+qVVtHbVoVuh3A
fbylBtkP/bQAQaQhOVocyf2HEtI7cQYu4WmVRpoaG8M32DPf0QexD1cAzz+Tl23B0/dmQemUqmze
SxumnoQfH6EJnCzbRfQkqSXsbyzJNQP3HdC58L6K35K14lCvNHJ6TtSiFbTcvbBTIfLL7mxaPSgi
qEE4BZ6Nl1tA0SnPGi/mMd/2p4+1BICRIExf3l4+sKgefQyYi0deIdtY7LtcxWBWwkOGp12BkC+T
/mvf2jQ0Qi59rT6Dhll8FGs1FXghAbCfiQK2WzZTtjs4+gZ/7IfZHVBAXyrGwBzso8KDoDdfbJ0b
4Ik7yGDGbNSYj5/AHzbZxe3JzLJTAZUUvyrqe0sARA/k0o+die2JFKLQfJdBLBCOTp302Rwp4ZEL
T6x7YREdAt+yF+5oI4N3vIIkUGVBXnEqVMR5dgY7eiJUeDlBR+j+A5j2YJhBwtsJwp92Du5Gh9pG
OD3kZ7Yb8YjeOrZEKNA7rPUEMDnY5BeJ3UX5eZNrJI3Gf2POE7IC+hbNskkZ8/mY6REzepXkF+7W
k3foXNcD2jTM2KczIlmtIIPzPiTI5Vtk4XwEc1I2CcHHowhTKp7Oe95DQg7supPtgLXpM/iPHfqV
0tTHHzCZWCYcWoBZ16a37cYx/D8AVcLIpjeKL4Pr8oOhsubOI7vVjGcv/Tja0pZTgUXZMvRe65k0
+UcwxGqeyYDD73DdS72mixWj1RnhhTdIAo6FCVo7YpmJyQvM4R3kM3ZB+MdVAnN8gkY5URf6/IyL
GxJEcL+2YXCb5JKVwSojUui+mzOC/tvp8H+I4ku3Uky9AUg/w+66l/La9lixGn8pqMea7Au8UBG8
ef8T6jPXeaOpDJ5ApD+ys1kcCp7zCnW8n2KcvMyFJTHLykqJ6FgRlAR+Y/1QFkVeFoSEEsP3RrU2
tZzw6QzNsi52hk87n4T9uo8TQnKhfLd7YcFniZwBg/w4TCpUcGrCBjCaj3fY/QNzLXpghPUvtp3I
u6aKZQvRdbrh5R3dee+LyRAWpyb/UlsAv1JAGcxoFhccRRapIri9k10fHso1tcn13eyAZVPDM8sZ
MlCGwjuLSdZKM1aqHi/YZJvN1dz1oVp3lKfgr66V93exiA88QhUlIsNNcb1yttKqDcOiQoLbAKrU
HGk+40GX2aHpykGRwt+5VIJuROYQ5YYATUbagrtA/X2SeuiwscA3wW7fTQCx7AUBAws326D+iw/3
g9EkdmA3AH9SF1V24sxNbcYClV6jYuPtUBFW3QqTFP6+lpRMJsmvHyUmMcsavm0mgH8H4WyndkxV
aXCMyAnPSTd3ckGLNp48tq6Ry2Yu8S45jAqHQTfjlHAm59pxh0SigYnkhSwrM1fEF766jznEH0Zm
TY+Q0w9oUTdYRJ235N4eUzRbdaE0e+zdsBiDLb4tRjcPgmVs2vKFd8Yyhiojx/ETU+6pAuh8e/EZ
QzehcJ7vPbS3oQXU3jzVqV3RqZIZBhEXZR2cIRpZU2oOeeAWmU9kBEnAvKzCkXo3rG2b+fRBuDFE
Yg4ZOrv6rHzbVqeX64IVEjvzbxSuzYQXDzdnEdLcBrhiC7GetdmxyK4bLNI86/3oBXxSCvaW5QgV
54Xfza3hklJT1tFp70xESBrVte7DimH2mpdB6rvrP5SRI/L2PCcK0YB/tgtE7qvElyKLF1XzLyYm
0rN/7Q/eDaDj2TOrnB0WKduCEnNAYQmXNsf2NGaElXrjwCLPs6+dlkKc0RBDeIHaJlpU+XahCYDf
bSJ2FgMBpndM5vE9TS2pixIv4wrWqwfEkOKXKznUZr/iKeoerltYS0Bo2FcnbayKJK8RJkT0/T04
NAY7GAerZmjS6WP+an8bFoZzDiJg1aNq56Sl2s1LG5J9xKCtOjWi/8K/Y4iEsx8wjGmZiMwVTYgg
tftyFUQgdEDYUBJSaKz2iNcSiyLofmyfUcHT+pU/qgFg/uOsuE+ROdnDOPMb9litfjMz+xkmE4QP
zq4AU6O2DVu0CNy+NxkmqM44u0tIw3im1H/ljGSBpvFVh7xSv/UXHGR3EDnap11yvVOTRDMkYwKl
j14zcnVItYfzN4MnECkG2AOwc6oImRfzVjz/EdNFIQdlxKhmc/4qETwlRJJLkTMVhk2Kk5hFEIXO
Lhe89uxK262Y2TSmgP+vOoJTFwHBUZrOc4qKcNQHckq2NECh4QmvkL1HTHV5qUeCJj3e1Yyky8KH
WMlWFfjKYMiqUpkb8pLL8GGxw5EE9NoLWdlLjjn9xpdVhD5w7pE78bY/ARLCPuJdKgGNvUfuAOeE
s7uVFObilve+hdY4iDkir9YUGcswk2O4EjtrpA+v/sRh7d4fE6MuKfJq+2WcyDdpg3oBEszrHPZo
yp9dm9bV3N0qK/Ns+twgYYqGWfPZ1ZrCTEUUcgrQ1AqrqqR40Y0mneKi5I2Nw4rk6s7WfLQvJDDT
eYNfKtbGT3YRWtqdvaCZlDGZYonu83BghcvTIaVhepWipFSAl+8geETlPkFnk/XhRQsboU2eIXmT
15lKxUI3OrqFxAysofqvhOZf3Fmji4+01BsDnhcuRmZE3/iuMJFNhzlDEuhhH/SXYnqN8I1WjAn9
d1G4BWyUZrPIUJ3jJBJzekbwBIq1AuDN860SiLhXaKTtQuFFu/acDquC8cJqaz9+roUDJNWFql3R
T74vnGJlDp2i65o5Tw2DqEPXJ6O9QAEk055bLL1mGy6oAR2HgY9mJy8kthScPsDPgVopbA16kmUj
bva1x/i5J2IajYVRl/lb6Ngfa9CjwoSVTowQg9iLBDWCorO2xIzUt0pFcRKEsd4QkgVerp/3tuk6
RMlHkCNB/XrJmVmEFumH/yVafBMMVIM8Ig5uk9Kdcs2CVyWrvdLfCr/mxWwpkDaBUlZmQ17eZ9x9
vbPXNrh+PlA//yLu2lvvuBJzxyGBTqqQ8c6F6knns3Y7oLfRg5Ie4FsQubhlOdL46+EaCWM5N6wV
nLQ+czVr46eVS09MXgtTFGW7+uJ4bCbXurlxZKFC3uKJl1cbvamTA+rn2FqLHtBipK+oV0TPmWBv
Wqtw2OALD36Sd3dJ3RUPfymehJKuRXHzX32jVeRoAe5wHFeOfdJgp0fzUqk/pXH+AvX2BD7yquUx
vveEajwzNV6Hx2iQmUj1aiVt1+c281EM97t+rGctYDtypB+ZVmPgQRJcwE1VuUL5+gQ2Prgyqxpx
6q8JQ7azU2cfJMS9oU74pbNt7A555WNzDmHS67BK1SxJyOWlLJm7NOQlpXiX7Q9/wsBXrreIQBXH
nIW4n9kZgjULTqpAxxs2b31cqtBEG1URCanMDwuLHHPv14/1tQ8BNpq7rHHfOfKkDocFctymGG8Y
8fH6r3JJs+BzArROoSTLqry7jPjMH/BuS5Reh7YhR1Kneya7y3+UgiuKPels8g9KI8OefXtqPc0w
DzTqvnxhemVnvfiHRMf/Wv4LHCVHXfId/UZKZE64tWcNwCnJ7G7k3KaXE/3vltLpLqXUcnOR2muV
vIbU5jkxSx+WBgH04Bm3BnsqRTQSuipVubDQjwuP7NREhrRd0ZNx/moReg3/XgFR+1ITNPtitby9
h1FYaR3gYr5wzBqBoQYMBkF/9sCfnr79EAaATFceVVxWP+/GFfANYHLL997D5VklBZMUe9ewNAwf
/47Tpgs+6+iUuHzVkFO+6pAJpAuisi/Oq3r4+CdPtxeP16+FNDUep3Wh0TtNrJjCCLkMWP74CAXN
kcaaGFqnvkD3CVOQmJsIDnEWpmreaxjL88oS7Ys/OVqk3TRVni/gXzjJbfpDZU1zvzge1TwzGVPF
ifLhbfb7cihH4plsS/D2CkPCHNCfAbWcSWUDgmPVDVebEbDR5USMHB3bBs0QlEkRTKrr9OhP/Wn7
UrvJl9g8oSHKgbMtM6Fpu7Ikil79MYIfHIJkqx3xWz0jcJdpMkUTjyaYIOdmnyj5J8XVPs9fmhCa
9cwssqeCFdvWZw072FGUPrwVHzzrn9HOuCcjdN78ugQJK/KdX+CwBs+s10NM0cqDjwb5BF8FPoEs
x7Z7VIy1HRCLaU0ejbpN8yw4J7GH3EHXQwPFo5IR4Ov7WnMz6ZTFNkQZAIUZL/e3h5+Kk/qvxUGQ
bb7k+xw3jhAc5oLGZ9pKbqvtsXeWp5G19oOgbqKkZCbQXTNIZE+XKq2AM3wrDzcrSXS0UDJGn0OB
cg+mdaeCshV3d06cLWx0jGY6wZ5+hsGpUCf4Zj9pg9mj+Q+WlAto4iJPitSI+g/DLmTQv+rO/XKO
2ODvxbKd6emUB6KWULYcvvXezbD7kFySyfINzLAOJVLg/E8hc+LeI4rG4pI7a/V+YRRdA3JVY6WC
eOAdQUsr6aGyF4pf1qDOFjN5VRs4zIUXTzxse8aRfPmOnlwP465OvVBbEoW0HTZZfYOGS//XpfMq
NdISFgDyhNHM5i1mOGQpiHweke6Ej2QeswszfpUPFU7AUk2QcFqjpsR630h0etVxwbYv7Nj/It/C
wzdHsodLvtMZacB6ITYTAe0HHghnMGFlvSHbMPa0/m/VvOAxk7C4k8dcpE2n/zXbJU7krwjiYA40
1/f3qlOM0oTGKBO8Berb5pBcLe3L5k2w8IUNXZ3fFB757DaZHQywcsn55IHgKFUlOvAbu1WP9lah
4IamVi66SyyFp/SewOcpxP+ZWiFNNlbDu9+RwYf+NifUZwdeWwSKR0lnmZPcTC2VAotJrs5TifBi
igJc/5dXEmAeCVunySjghsooOSUhBCZuAXHjaq2ef6dRfOtwxJ5Xw9XIZkbEoUmzuLcB5faZOJaE
DBVvCqj3TOjNchCNXnX9TD7pzdKO0W69p7IqR2g2gjbUvGdefkBVIS6eZE+zyd9MWjArvnYMTOam
RirrNRdPmw0uS+x5V5ZfxJuwrvupbxNZCCM20e8YiK0Z1w3z6LNVRkJxoqc054srqjpSQDJHW0kP
qWGX6wjfkYMeYjkm0mG2q5gOyzXQe2DNGnmpip71VQacbf5En8kHStc9QDLv+bhBMKyuKYMonXn/
Lulssfm7f+Lqm9Zg5xyyzJPdZXim1zQp+EZRcLan/SF2Ag8n6x/GszQiQouYcKFlHJDt+5Lw7exn
syVlERKFRqtXQ/vVdgft28fQxyEXs1OJYD5YgEQQ4c1yIXR+JaNS62Y1WxbNBkmlYTvPgbXYBmFK
7DTPfatw+KlydCAmZL6L54HRcMOVJQcZcr+n3zj0g8rcsecTcBnXm5vcihiLX0qwto3NAaX74WVn
37BO+78dzDPNtTLc/Y5C6pPx2zVRfuqUlKCSh1ApiGWV3oUvh+4mjj7QSD2jJsnEyXf6RgUpbx6d
Y/qvvUaVOQIzquuCBgMp0f1/XsYZdlUTLPBd8EVdjV1W3R9hLK44D8cFBLOWD2cgcSbfko7+gYKy
vHsUWJo3zfxDpv++6k26yk9ologvZmJFdz22pudMFyPmuTqWebzn4WmfU6/W7FLHJIlC22GGPDed
p/wfpjH5/FQtca2eTunUxE8j+357YhDeclae8AThWonfkvA80m6h5TpR4YMU2trtaBo7IceQnGle
E/gnLFj01QAgrJusUMxV0oGwan7OkRT8FmVqURzzT5+JnJVqd3SRGW7ypm25sW5CVvopfLLB1ShK
tCHKrxXKS/5sAb3S2GSVWtBWUmSgKI7eTgKBT6LuQ8u1tXW4RpgXKNtlGWWxQf6wM8eiZt3qrmIY
rn0CsLslnBzaso+KPRLenUR9GGlsEk9JQ3o0XtDCJ0cMJOtGythHNTb0aPy1MPKCYm3mKHUZHQte
kNChSNMJFaKdohhCW5af9AfAFukRaWf10mvds53xC6mG+pU0TiMfLm1tEJ0dKQs+fFpmawlCBbso
qtbtdy0jx/ZMbOGvIRmyqoH1EfyouaNftcMP+WFq3WyyR4adwKNZ1TpV7YTtx3OZNv2AFfNC2eAA
90+zQtXNX7I8XBpAzCsWEHfcoYrKmn72vy9vkLzjbPVEjHW1SmojBUP2YMP/7swQOYlnWEvO3+jD
GoLu7ByXi0p5iQ9V1pDpv4yBdI7JuGz/BYTUPFPtKqNfJeGbUrOpPLP8X7Fy/cgpf7u0kZ/6jshl
UnmbRXTZRAau0Gso5wCwBz0AAcjuUNvYZe4wIXhXe/tPLqN6gG5m9rotPZKOR2+tVGoWt5TSzpzp
fUe8+Rb+AqOtl2tL5WC0i+pQIGfe5lBLYjhWdKYWAUHHD3axTt+RMqJWz+JGNaqMD7weUzFjxRjZ
INoENTmndqK4tFAfS4AQdTEUnGv95ZMQQ0fUpR6f40rKAhlbaxMHtoYrwhq78UYLb5YPpZ2O+wm/
IKTpV+GOPeMIJefic+7PlNkh0XsN128WJqQrVggJLDegO/yt0JVFy0Rb57Ln8xReonwx6iRu9HdZ
V81o4VK7Lz96JG7eqMDRCekFapSJii2wiU9nWg6U4UfIhhwawK5dHX1SUYsS0b1irmzSkWOWxZZQ
f/bJdu5VhkKVjSqC8d5jAV2ZqGxUmas7e1336VFx3MzBVP2K3qlmqQl7kBtGFZsZ9i6eEA7ZO3Dy
A9UQqMXxYLMOGMWI6jhS8yeVypk+Bcm2q4MbQ3PAYfKwFb7t/HtbOA/tMQ1cPxZSsRxhXzD+jIaa
YG9BQJWl5NwknzH1MWN8TaXfs9R96nq1R4fVbPNu4j6y82UUHOguvG9YGFuzHdeYcd1dxqYGvx0h
ynya1nGnVc9PDTQVEdMZWMTulgNziUzSXNxcg6+fvh0QEGqOqYrxiZUbrC9nVYkjsTXlfRoHYe2R
aN7M0TFVaZay2bKwjK/LZkRVUQwXYVwc47b8Wup5P5Km9bDowucGEx8ogQvDwHWKhlqXNf3P0o6J
cEa5SeWxOls/O7W0DVHFlogOAzel0rFN0xrZ0ehI+UdT4ExmQ6snE0XgeRoYbHpnnXVGaERKI0vS
Zaps87MzB1q/eQvM8bMSfv+qwNnrFPHH0onbpaLycvxVHPsjZU9RsHL8AhZS2C1HdDp+XkqWp2Vn
1GVDu7bn/7cFQIBrlp+X5pqLqL0yohDn3lp5EFqBVtiVGs8Ptg1kRgYMHqzVNReLTCu4c8qIpjYJ
JQpRZ/+jmIW/e6j1bwMseV+tmERQLenGz8Hk5YbvHE8Cg+7cwZwA+GYl52O5pY7FzaPz6rk5pKxd
fnA2fql4QSAQF8Hm2jS75wDevoGWQMBgdwXyErQKScfSchCn+g7WqIyzIczUtUFnvs8v0hbHflps
Xf+qjoi20WZbtcCETIwneUWjDic6kLlsoGmn6CpuNTf9o8zGe5ybJPUxZnrk4P6bV3kLwPSYoX+c
PmMhX4Y3PYdzI6HXYKjA/mmYX7TldSBoForv2PQByyRyAmlqyx9sPgmj5uH0PjsSY0rWJYIvk0jb
nIkcdSX4bPeWpTM47kEUFR6zEDa7kWfZadJeGEo54yvo2LcA2y43TeLq5w9RmWudT3v7Pr/GjmVv
K/lXuMV+979aenfKdCLl657/3GqTyEx5Vcfszd4KIJT7yThvaOnF42sRZsKhxg3+XfpzA+YGN1mf
286EMbeMXtl3DbvOzCpRK0cXgVyzoVXpUWL6zCZAnXb226TSICMUJWXm/D5iqlWUcthz8tQxr/wJ
eYdt5zA5N2IwRKD3wxKaBDY6wlnNmwNhcm2etLet6w02yDaDCC6ySr5GjCLhH52UGcPOAUcFVVid
WOhKlftff/sd3JZQKmveA3FE2FaWP4k5vuH079ZMxiQsB+x04tjmfM9skDwI9gw3HETM4Cv280Tb
K9OVCB+saKmevQ88o9gXZvqB8hYTJSkJS+hO4S8ptLlarJI2CpDbbLVSTPaE881yqqdhXrMx4dIx
cmk/KdBI6vgHik3bMiERUGC7lP3CW7qyfTT/FkPlegrJLgxKp3Zrk9z0zKvukK+0AyKQI27qpBxp
kodF8SU0skM7ZEe8If9nBapbiZJOQwdLNuqVlLbALIE/HuGjHX6v+LgL/lW1nDLbc1LykbdGioB1
7k5k1rDTiuca0ASFavfBOO+vHmVLTSdW2rywdp2NOnw6eppesMUQBcKiQGzfzRHDHSlKzXAsRpdQ
P+c6RYumv0zOlx4f0MqWGFEh6eNnkV8+19TA2MNogP86j1VcgAPRbRLIxw5YVjR+IApN3h/h4lWz
tXhoU19DZycuEngcxtnJpXQGRb3ijsD+9GHktSM/0LaOUZpFTlo3uYp9acw9dUfXSMyfHmZ5m9Fh
euUTM5olqh7kZ5/j1wRtfM8Vi1RXIyFcGLCv7/sLh/VCT0L0CnbMQ+8qJITihAAwlwpv/AtY5uzQ
rAyrFyUuQj8fwsn8hfU3izfGonl1m4xmyKyWXYiE+sFINiXD6MM72V7yVJBdHagfS+cbHWqfvMrp
0sYbwWOxqxMMYxFmvUe/E47l0GdoS/rqohot168tstO9YgWHT889FiwjUDNnTwZyB5/8Qf1DEMos
fmc0H1aBHnuXW1nLcLezg39Bln6jJS4X/x95xmaVXqxoshLL8BG/MQLvqiEe4Pf/rjz4yBaozgZ3
NRx4uVRmmzHN/xZ0FHitLdhKcriLRQXnEgMSu9/UaaYuci/IBdGfe7U9NjoL++7/SLfiChnt71w4
btKFedadyBNZfk35jXc9Y/Vsww1dY9GZZBbYoXfGbGeErmBL94i9K2AR+eOToKSE7tpECiRMRXyB
Mco1YJzG2iF54T2hAUbaJHpIIQzyYt0K/bitN9sf8c+4QM2UYh3WKtg60Kk+R54F55WMN8Sazd5S
51OzrBhVdEhEmG7XJtsCMQSaHOJ6vc7MhyUG4qiGIRnxkqJ/Eqhm57Hi7NHOX6ch1knr9W5oyi2T
jj8vC5YMXVqRe0WkUX184xmTkf4vpB0ctd5l3TRA7CEch0gSxA1DCNoru7vIrIjHw+Oup9pdDCvN
5cEqjRCEB2HAaBwX9cDcKRSnO1UMOrC79e8uUvHD5dlvdMxj1VMiXf4n79sqSu2kVNBQMcMyI4iB
vVsrdhnjqU86LCsscIZjiiMe87Ry9uFHd/1Wrz1lnW0A+BYoirwKMLTOcOf9lEfBSKzgyVT2W954
ZfNsgz456zYLepg1r4BS3WNT+ehfVF2cWF61zq5r5ZzGwusEtF7RU1NCToizHD3DA6jjXH7oeI6Y
bXB6wXiLBZwzXXruAa57Y36wweKB54WLxDDkql2HwDQJhm4WwBuh3npJRkXoIOa8ds63yMWXtWRI
ZFqLX5xMRs3oUShIzB9lfJb9c/mEG3zBptC9veMyrQEqVfkx2JsmzhFA8by4QwerXA0SJgGwRXJn
W62eryBNmC8mLPgIoY9g9PGE2QdB4bLHFZt5MdCg+xBVoy9gj73pAk08iy1MDbRhBmP4+dVUQJ3Q
umfBPZ7b4xRxVY0zHSeM8IAXroHxA8cWPKPUlZ0hDTyyHzhwBXmgB0S3HFcoX25aD+P3ybLR88OM
b7SBHZIvnjpenjSt6dbevecE3iMMLTFj/METy2QCENox4omAFqFa4JEZCSe/r37BmWKNf3Ee/xxP
60HpXTQAppFiRefhKxXI1IWVihQh3bjfsiBD8GzTcG1jGQPyjKxPAb5FdlYGmuHu17KiyWiurvQ0
Zw+eE+DNXVD+QxE+PJ67pSGKoK+Jf41c6hGomjBJmnAbl7V9VZQEInuDPwRCGkceQlF3ge9e4RJ7
IV9OQK2NA179aRO7lXSdcGL4/lM/oEz68Ja9vgAzHFJ0KHBxJZucO9WTkvNCTrFsZXl55vRCUe9O
g8kLwHm9R2YyIV7XNFaz1UFrvtcqUoSJ3+5cygXICHhCeNSTuJMD0U7+ewMlRTkvZ9svn40GevVI
A7ceBytuYyyf9+6VPdBn0ARUyxqlnENQtiGJ+8U5pHvZEz9VcjU1/Vrg5BjnszEw65PL7r6rGqVi
BqYo0gD9FIRQZe+SpoSC353r0wG7zErzYdhutzbMuzFN5mXGZeem1CVVF6gvC3bbgR+V0wSeG8nl
JLrwtlomc5F+XU/lHnLxpCexp1xp/u4rJNoNx4zDAF6O5FZwE3tbbKuP0AVuZQ+ZtxRhWOoYWOza
Gt1UsQXBynen6TaGiiXjznRcKv8kJmVW8MoIJhk102EBH8TMdtDYMuGH4ZPqPc/jfTmvkL1gVRIp
NdVGAhx6gPAwzhuu+hN8fA2CpvwiAy1HgCMjuSVp2j/aA2sBGRMSV9vD4FxWxTa68jjeiT7gcA+e
FzmaJiA1rQZUy7TljSgwZTn+Aj3HH4p2w+CQDfK09m0ysMmhwkt/4M/MeeDSFglaoaHuf724PXX0
BI3+qzb+wOY0u0G2oZRxz7VE0eJgyQfpCi1vSi+LqjFJIX1N2YScVZYTgAn60gNUDg/zEhw3dylb
zwwbDTsQn/UmfLbup/KoVUOq6CPQJkjFxpXZz1E5T/D+FV14Tn05lTW3aBkntrataGP6CSeLxvuC
sNzNuOtDYY9cz1tuYfTFG6agSmz/5koa+3Hwtm0VYzxogGdELVEj2qsm4n+Nq2fq+1uwRwiDkUjS
2g1sfIOz6cBwdAoKvRGubhC9lWdwIyx650PmGGISVhbJ4/KMOb4eHBs5BIaUQ1XQ/oyKzW/yIei8
PVME5qMO+KoYptRXq3Xr6qJ1c3Cm9E0YATyD7oioykLsToBS75Kz6EsAiugcx2SOahw6PdMoqEzy
cVPJwTLtKXN7Dg0AXJFdWhymWTgIM/JIRb5Z0WQzQ8o1BapHqi5PTc20Yoomgba0DSnsefErfkz7
Ae4Lcdhs5F3oJYAvMMrhtWpPWGbQyu9EdZVcd+0mcr4wmQ9dgpazxL5AXC2D4yHgD+f3aRUF29S/
MZ4/EXyeqYW3PEumBo4lBOBdYEHuU6opa1PElIWbFLn9+GgxSydOQxZ5xF8vt+HfW31aFp1xK6Mm
08pp8JNK0lnoUr6wbAlS8gccHtjO23jgmI/rULhqYSIisl6enQoLAb73gG7nwVyIzy4suROk/qv4
v5hfoMsOPAiz5t7u7LPmqnJE6aYTEYWMK4vEhCVlxduMHNzheYtaBPY1RG9D+936x0EQp1GmafVM
MXGwxYPUYO8OyWTy5xUkw/iUiWc6aJ1ryRW4S3umbrdhO4AGwgPPvgV5lArhZK4S+1AQIMNQXrh5
zUhflL/r2cBuCVFr/NC54n3fuJvDLId2emtq0K8vwMea3D7VW1S2dt3jufPNIzbC5ItOGsXZAW8K
amTGO50OPueURoC75xeKrI78UMx3UfvmPC30CDkb51oA2l8u2iz7xG0a3F8vSBztEhZpUfb8A9RE
cE/ehwq94/QxTR8h/dBk2lTAFaC2/o77AuTSuUcOYauGlxSvmh6xp6LuE5KQPMzvs5JbqMKtWFWB
g1s7VIhLI+cgxyktqWtjvkSB0XHD6lhtJw4bkoVQhv2xQzh5ql8sBzK55+yRnCCOyO4d0GvKQTgY
HqdZzJX1V3i35771Y73QwRe98BG+igIPE2o9qkkfP6uUijEp9jBnQ8Aozc7g5/fqlidgz0QLyRki
ZIoT5PayEMXdkAyqsYf8mBcoBXQR/yQVDYGuc3jXL7RBrbIWy9vQanTZr+rig4QcUNoChDdL0VIf
11O50aSJvOWYf9L9ltNOdDkGyTd6NtV11wi1Z60hrG32pWg/Zi40KzoyeATNlKi4rOMkxXzNty4w
pYvB6Dw68a+fM8jIPHjcf2XVTS1ajOGGRLFr5B0TyaMlOICZnMgRlvPurmF2C9xNXb5oZ7j/6OnP
Mk56ql3nLxjQ0ThRwwmdONFjfQXil3HGThYg/h4tTJJOMjfmxfMWBGG2VV4QvZDycsBrmp6ggx7y
c6wtBHpwMCm9F1db9uN4SaHTtuoOHXSb+zP19lvMAmfDG/w1wbobHO54pArigKrsrrR6SD33Pl+a
dlQ3xnMrP+VlNdeDqMO6jQcxdZewABcT+DNnmd9tYnoyPGq87yNYnIxSCrJBseGS97F6hn/gIZsw
BI1MmiJeOwig0s8Sojz7Kt3Xz+vIAdKd99EGLomQtv7Our80GyrgCofQ14cbI/Ed7jhwpUGqfNIP
i9BCbOFkj8zqfxJZ8kSpAiKZLxvPIMbCnzlqKpn1i72tzEI0a8ayiF0zchhZ/XnhknfliOKVZdh0
EeGwAq/ACqkfhSPXsH4Mpr4u3p1xAmSOlQCjRqCTBUCPHmJiJ6TNxl2vhMOjHK0JWlxJmE6dOlcS
S0KtjOW34BIMIb9uuEAhlLa0M2Oc2MpiVj6o//Yhi4mvZpeOEly5X95JsJNk1pG1H0IxLI5reCDn
FcysZYdXEt+RU7GgOI67mRBmhN7cGZll5SAOcnbAgnCLGr1oTk3mye0Ttkvki4Zty4NTBv/nM1NR
GXunCNcJ0iqJ/E05B6EpqFF+CKKkk3QYXs32wtlbZPwZ63bOIhfANWnNd7bN1oN6b46dsxX/qUEY
gzozmoXcAQWoQpnVFqLrgGV5Yu0jjma+mi3ACpOc4qU7usQkrAqb60IswhjV45JJtyQcH9LIxMdL
xuldF1QfNSdpdfHY4e+aLkT5Pyaru6I/2UU61lhWWTskH9WlD3fFUtnLJul34XdNO9klhaOxlXQ+
vAPJyyyzQQpq4T1SgTMKiG0G96RXjiBaEbZWKGy1h0n/HVprCd5CBVOz8fNOefVm5fe+4zyMQvoy
cRZhhmKHvvdt7FtL8jmbEJ6l9Z40wbvAZwaEOQLavU4Jrfp6d8sH45ZtTfPIjuoH7N0ynLYABriy
jXS2kLTcU3LnWI9DqUa9n6vOVaEAF1ARy/ISyQxVHdpmnRfI25CHS/e8cHCOUcBIvR9DKahzA+N7
tq1a/TACEUREJ0EzvpUHb1dIG3Z4udIxBLrqlNxLJKWlQewXL0ELmlVhWIyZej11sqEUSetqrkEt
tfms1k+c9mKFnARUZ4CnpUo0KmpObr3rZDuKPTrEeehZcgG43eUUlqdqe4thVCB3PVa9OMExZprH
ev7bPrzHtT1LbSZNOKjwV0vcIGlx4r96ld/1i2BmC2GkDTZiQdlsMIIGiDO7xJSkESV+yr1hVR07
9xbCI0ZrK1y5Wos1s+1CyY4+2aJU8s7N+EJEnJ0W3roTvqsPzsK6Fx/XeqpbF75TSup4POcFGimV
ClmcutrA3Q1i+F7+GsjYJ71psdFPMI/qDPSA1D5J5v88DZvjnBeHyTk83BkCiLI4PnCi7kbAQDDg
q+1GCn7Wf/NuNQ7VjPpuQ163dHGuFwmde/gpXg7JPs8UxOKuxmPE9GyPAifWNKsDB+tC5DFAw0vQ
hMudCi51fR1iwBZTOo4l/Z/GUIzI6aGinFHGVoy1DOQx0urAYRGyYdsn7qDids8M7BQwtx2lUIUv
GyK15/z7ZAfK+88R6j0jx5oyMt/kBXG0JNfc95H086SWmM1XTEX7QJoS278OkJGF/lRdPzCIxbcR
AfCn3A4kG3Yz0Buv68Wn0PLnS7GZzru2jLSQ7uc423cV3gxcmOXGR4vIw0JKefcHqC4fZTTt49bq
dFVpUj0uzmWb8nYBY8cmjEq1txv7/kB+48aMOMGxNfLKEXY5w+mPFzq8p1m0uVLi0Rh+bV5Q0OaN
o0bL1wt1j5iwt89xx77DC/EucJJgwm39oDPPCdfEJCdEaEIzHpaRkF9KdICf+VNp5zPm4ofiINY3
eBgqlcXLMsdKJNQOaQEXewZ0ZsgpPiD3/pd8sIPxZTSAL6j95nZWIvaqaxH7mE6qjZgCgbglA1n2
wdk6LewedXBvZd6vzGJtCql59hHnIeD1rYtohec/c/GLjC8HUyv9lkUKI1s/yDy/7M0276P9R/HY
RagO99XcmNOmrNU2tjabNsbh231vKmYK6m9eTUxTUOqFNAHcU6bn0/tiUOs2No/I30MJ2n9MlGTd
ConDUdmC3adTEynspie9gj0ws/nGn4EbojSV/9zL4z3offTrlml52u0GuIMtHMSCcnnPr9gOB7YO
EPvKvkBoWRoysKA/G8KyHIx9W/iu+8E4cn/BxXRPAuTky4huolnXC7P9gFkKv8HX6HIkXcDVCwss
72x6cTfiatEPHCvxDpbkxL7gGbALh9s4ImrBISC3x42Y13LBRfYRSbXYKXkcuY13UBtOwJ8yrYQg
SiSDZp/NVK5dH7meXCdioMy3WuxbkXLQqRUX2LiMs8d5hAgZVWUJoOm3uJnygTvhRmy7X8EPrWW9
7CzyaMR3kZAm8WilSrvM/nfXASvCFxF4AIIIurc3N5orMskTfRTUOSYDZ+vXf7Lax5H9JD3o9nYe
JnHNXJZGPVKjkwmPEThp/KTKotBFBSGVjghWzrnM4qPqUPalF36iFutQurvZhc4T8zvbs5J0QNI/
5ALyj5Ai5AW1RrjSUL86ixUNMkt153ibPkbN0DB1GAnEPcZbERnPagnTJ0hUKNljA8sJW3ThiHrt
/6NsEO5bt5IBmFwzVYy6lB+urLzeD8umTuaNCgEHrBmaAHAKsT5nCAZhe9Vf/s2n308RXybAT9+8
MdD9SID8ZAT+W2GlfTblOLyVsgRal+Kw+mnV/ibsgIIi+1WsHZLAu3OaJUTPajoTDo0NlnnmvNgJ
r8Mr9qAav390w43AMgMUULnv8kdW301nn8VJRMu7wwouHKP/pdAsX5XpqMYYk5Z3fEtuOyu7OvKt
Eah7ZRdYor0jpL6dEefHCvhMxCrtEd4jUnRXGxHdlcAVr/9K68rk5G+27CLkqKR3tDWygDI6hqth
x7Ka73d8Q8dHhbTcceRo45dJvvZjGmwPrS0yTFXxe6/Qet+nw8XHV7eD5A2Uu7rEMGaO5qPZ2LoY
Wxgxudsjb/PbGJkss9Hf0He0eyC0PPh0eWtl2/y9f64P4qur9DSte/zY61JXp7Eb7P5NQd1RyTpP
Z0Y/4mn1SPxBwF/pQWcDIUJKqrXT1xL37nB5L0ZI19X9hAy9OBxrheUbu9cZ52Owb8IUl1TyVm/I
jTgGt+7BEG6cQ74+yJNUZLznaikqYus6DmHukUP+xLUQyHlWquLfFuc2yDX+1jgj6dQywvKqVg1r
B9z1QT5UoEbbljYJCFBNwX8Q6eDUmXJjjnC8FfbKLXcN7uyAmQVpDXEm2GeSsFoizOBXbCyZvfXy
/3ceoHF6/9Eym4/nXw3Ot1BdU9MQR02Z5T/Uq28RHEbhDBB7l7C9lqwqTyS0SiNzucwmaO7vTKPI
jB6vEaZRJfyLvl73WJ3qFoHjiOzBeM7CPmIgvxSgXB1l2ANuWsjkpPF9Y7//xDrXjJiFleLyZ3Ik
4SRNU6zxn9yyMJqk+8zF5/XCl+0Zskt/QQFroputzq/+S1B72fIpd5yPSYMW6jNwzOEcXF5oUiDR
1bLZ+5Fplbucqgcne0nyEhgf6Dre9ZszSnhWJ+uqiOy5/CyoPkaGqj5d/j9/lTBpWI/A6FbgT3OS
AM3MlG3VoudBQU8FlhBoXPl228bIH//GVFRbMM5jMnGGbOXV2p2NXwVISYvGHTK48o8TtGkucXoR
hiIdaeluoN4XXuWKxsBGRVl/LGKGwokXwmJdT5uLluQ4SF5CloCG++OFCNadmms5aT8bytJovsxE
J66VT76hrvq+HZVPaVr33QK0RRZcYnQym9VgrPY814E2W7JM40njzrQKSLtVdAhv70gEvyaDxmdO
s93Mm6n9mHomk24z6dbSa1dDRIdxjU11VrIKX4ZHkT0oltCCd5ec9YmDJc8bacJz9UFzdZvLKPm9
iIQr8t5MgmtE+tsyy5bHf66+3vDogl02/564JX40yhHAL8EzmaU8Jptjt6lhq1letYlUzXeUQVLn
z3W8bZhMyNgBsWVB3VDunpkwGq2PzV11BXo0eGPXev5e2EbVnIvEGLIpVoIfBt6tPfNr3dSgMvX6
qtVCMHYeI+vOwoXT1FscdEykIyUErqDXIpQPgdxzqi8qT5ALPPgBl7LEjDpoJKiAyHNyo/f32AVB
J0kE/eaD6BjeNoBd3S8QBAYQ5eRXiUsaxafpQYnXtN0D7AScQ+DhhucALvnAQLighaENPNz4mIqh
QrwAMEi1PS6uJBthLm4+MvP1PjuCRyEs8bHxkgDhS0F4tdAKfsHk0ooRrSg6OuS1V9OlsoqatddI
N3+w7sRuj1mogTLHcMZSwkZst3gq+JRpLPhHQwe3JBPOHM5CSC2hwJDX3mrnp9CJPs70UQbHQYAT
vzidmogd/800VKKfUfkB5XhLL2h7aDBIYCKTHx60elZMKeJkCB+uYu+Jj7lgBsYBQEgN16GD6lw3
TRExi12nUe6RuugJzKL9l6/r34hpguhEfE1S4LE+ce0oxvPzpW/enM7nox1VdI6he2YylwCKJhjy
5kk/AM6grx/Mgn9auI9e2ylhd2pkzyNvUAG+dLQlR0cQNSUf/mRXLmPJLxn1ztyFqgN1O8OCq66r
0KY7pKZ7VmV0xwvNQn5Aq7zZBbVfOiD6C6I8nCA+XOfOqb0/XELKYCSOOT668NyI+j+kyhu7s4tt
ZrX7UKUmJ5Qc1HS6oyjfESpLq7jbzBm/lHIzI9JHUnpTXEIqWc81bvGtiod2jHhOeQgbnVaK4bon
nY/Mu8D98kSM3zFOwHMmoLD2soh2KBE0uA8oAxlSDYd/wLj6OdlGclR2FySoDJlwUfB4btG/iTd1
EEhpewnxgFqg/ZbespuOqfunbIzenVNCZ8qBRVYcNjH9A1ewg1Ida67oi51jqy9bJTij0O77UHF8
BEwi3P/cm5ljRswYq3Sq4coY4DBM0oaDcCZEq9bcx8Sht85IFME8oxcIo85sdVJDBG+1PGxLUX4q
3MnYOSD3DD1UMEI6hxTPdkkCX8tL/3dxBtC5xBfUQ/Q2HyJxrASRDBUOBNl/sjdmUGfjBgUoI1uz
ovMNMRS3GuyO0P/LZoWTFj8kNYDF+SWOL8xFLsc398nC1JM48GcWVtuZvqXhlEMwbXDAw9y2Abbt
FnZ1V/J++KeOSYbkMhWkEn48s0YLE/NhHZDdQjBEz553nD2zvZYHcnYaI9FCZSbmy9R5kZhEniFr
rtG6Q8J+/s9lAx5LT/vjtRtj2IgU2UU/AibdUn6+IKc2zuOqY9e2GGGYxEX2Lh8KxhzDq6kpGPaS
Fs4JUTBqBdwB1XThIG/7eQ1/mimNSy/H9DbbOfffJ4b9HBnNLnZFy1jUYgl7DJXJTtUk1fq+U87/
u079KsEsv6IErqBgqZymG/5ySMrc4SOquN3hYAYSFvw5M13B38sq7YrebT/vMQcVn/0AoWPZpcpj
tgJywtdO9QUOJuySAi8FnhA6x8H04/ayQTSPcl6s2u3q+11FDIRULkpXJPXTIWtftbaAyojP2ckf
KPzOv+4+KoDB00E6luGf615KwnofMd2ipxMLxBEaWPPBHvmoAFcOGwa9AXHiEfls+cqHx90PdfTx
bED5Q2aqAc17QJuN0OZCsQgFBljvqXR+/ts64jpxNL27kQsnxorimHVnUO+r5Htcd8Cas1b5wn5G
fYzK2wkbkHDPvRNlj6gnLkZb1UrRKWBqXHRUUX1wRKQS8f7i/9aO4DP0r/+oW259gxTpr4caNBam
lWeQQjWaH/kRHtnIpK7W1PdE/JaEgdrcK3IpHUSNa5BsacsJwYyeUjZd0Vwt++O+g+hr+dmAoWOd
WQ+9OcVPq95OUQ6GXxkp1XOsTW6NvEC5vBmq4VXgEUD7XUk/9kitXZ1pszqv6eds+pyK1hpnSgPy
zIsSoHlCXPJ2/asiJekppucEdrpgJbStQ/T9ImpJ0ulmMdpRow1Z+KCVXprbvIC46ym+G1/cJK+/
zhqGvt5laCJe9aJQbMFZxj4nYPFGOnwgLH8tkhC01ArevquZAgy+O072U7esWmBoAy55173T4Nsm
9VkvGRKsjEYHdpHbIyhBB//g0IOjqk+E9x8TA5Uvp8HHcrfCoRp4gNQaUcoPErsL6Wf39Axj0Ex/
RDvjxWeFtq3CyW3LThXeUTezfKcFHQV/HbpcEPWMwz/aj4J9bf2Pl3SfZcE62aqZo0c10TMGEbbG
W4pgRU1xexbrN7KjvMTim0RX3OUAqKJeaddOMJ1ZEaVQhh/lHcv0r5eecMwc0kFrQvNsjEurkWNh
BLoPLpxQs2iSbqoHYA4ERxRhITptUj6LV9hOVWkfOm5xMHJyOrI2Vatf5zj7r4Kb/8eUqV4mGO8H
WuLqoC7gPSvR4PKc7BoLxpjBsyjn8fmvF+oL8sHVEURHfHvq9WpRHOWkOaYLzU07uiRXrfqwNGQ/
a0cU8UaJlVIjNp1Kf02LZYE5R8SYmXLitJnzpoguDn9+wjM/0OLVKfEIW6TJYCnIiRLgplkja1ph
IXRes3XrNlLr10RHASzBGOa8msxQApK+wVBQ9QAmCnZcPbyev9C+4IHp8VLZIfnk/wg/Z4uNzFGi
wiKpVsem9qgaJvkmnBPqPGzjcKV0eJN4ayHb0PRJHB00QMJkzGhopzTS+EUgXvTKL6WdtqMYQIMH
7TppdBXvRNPio6FZCgt+jYBoQ237mQsUJnbJpz3r3ua3bPl4ekcMJFnDjYWjTFB2IUjr7z0icIkN
n07Oyg32h1hDaB2+iYGNuCPuzdlcwysUt2AYFSU0BQU56GPQu+sl9WQv0s6CDwa0t+O1Vril7sci
AfAATHlZRIOihnXsV7/49IxiWnRceqmLiFUYuCEpzwXr0hgUqFIjxBw/apb5yyJifJXJucXBSl0A
+lIG+bNTJ6hYw126MqlRkxPWdCL9y3XwiraPdXA2BUgp0WxqbKMcTXyjuGgoIit28tK1NIWizQOh
pYCLudi4vEZAz9wud3mlvEPJZAau5sNWhUz4FCtNWaoKG+AUmpk526rH38TxeAltAQUpG7EAYdnS
rzg4XHEu5eymYuvG6aKtmVlqx5LPUYw/0Eq01Srpy39bHHH8iRj27M/Izn9te/r6WfVOvobVaNCS
by7+SXoeTXkBdbaZflsCVHzFjmXpNi65iD4zu49hbLqKyiyjcNMU+zsUdl+zZZ5Uo7xvKQI5BfRY
5lBfnzqrp9tC4AJbu8Yo9vhgPyuXRa2nFyd+DWcVc8gSNTCCxB+uqh6F+XmXTW6DlLMl1/hIL632
hMPrU76bCLvZqvHK1fP30H1rpazVZ8vSrB2S3CsO4KOgMMD+zrHkBGHtBInQuTqX4Ieedl1onuuM
eKXUfb0WW+KR/pI0ipPDJQ3YMnNH2y4OapIC8lPV1oB8QCmei5jAY5zmVNoGfeXeNylUPLZ392v1
CDrDsbty2ExEO/el/aOgUM9iAestpPeOSQqKq8UHSpBr9mr7W1uJS4AHsqDzRZhnewGagAFB1GB+
SzddovX7o1bAFFABg1agkirmK6kENLJZWc3/FkQOmoO3eN4ckJhcNpAZvmv/4ElB3IvRisO23Nc6
2hRGw8KX6NSb39OEq4fnJCezt2A1KJHvz4ETWEcB7zhXqgnnoAY6buTxBLz9M+hnegn6lcAHw8xh
4MMRR4644cyxje7shI7l9+MUu1mBnOnQeDNzk/g/GeCGX4tVNjaSaboQXESkP6ADFH2T8mWvtgGU
/dXJUXejzq8fQzuFXVZB6rSkkU1VNz0zRJAE7DDiyns7YESWiuWfZitw+rcs2/Qa93FnBbEGd1br
12nczDLLxTOiz02EfgG1GtpelCT+SJ9E7hYjO8l1QDTaxB3i0/A9952lpIAo+S8g3ZBvIycnhx/k
MHXI80TjvGCnsuOEplzhaguJpWUWxuE8mek0JKxbgEu7ZFQZmV1ExAPw1C63fxoj36045hJLKHqV
BRxsQryU4fQNAMe8bUbxl3YnzY1d5DKdSoH4+wWzqFUgDSEeQ2l7ekndak81oGIXVeVp49l0RaGw
AiAcIDb2DSlXISkIwI92vwvQU4DR1zA5TC2v95ODf5xlnXE4m0V6iJ6q4T+KrwTT+53rt3z62vB2
KcnQuXUwWQgSGJBtbPdFcM4pPyH/YMmy8bNrvqKo8tCo4mdXmodIhjsj1lSQHNbF+GqjVkOl6BJL
7+tjVwEYr1qDpN4rXdSdxVA58PLIIegbap9TuwJBG+Vhy6hUAcX32KnXbhmv82ehEAn2EAbJ0ljx
14YbXZ1v4dARQPF0Kbb9pxVNeeRYnUH5nkgdPiJBQ7YKEGfHy+ZkfHlwzfS3CEhKTR+LYND28BIO
nluzx6F7nxiO7e3cmdhqJwxwMTmIgrEnnSUfHRPPrBYxde1s3fVNldqUCT8J5C6nHN5PdRG6aTiB
UUTom/Uf6zYYTpsv/yJBAUrGds08AT1EvSBmiobszBdLG4oT4PVWlldwhAe0k98AYT9aQ/m7Z2EQ
EFjEWNkT+sZr3CXZGmFAJrNXqTnk5iHG2PcKW9NxYbd0l70TLRx632cAq6YipExHnd6sPIS2CM6a
fy9YY+2OYjE+VqADRDHKyyRm//zkB/JJqwIMToC2ixvQaByQ5GEJY2LdNNMvC0CXi1p9roeAXQDk
ISb3+9K4pDkojTASDghUb/atOcTqdTAtWF9JOpUgz+g4LGYmIaoME4qqGT6Y8PUPeWW0ksejY2qz
KFNpB+SkheCfS3NHjAUyUp3mDNYaDt2Mv2uuqoeMoShbbedkO8/0/QtDEAcA5iGInpkoDvfG4wZ7
Fd3zYtCN846216Wu4mvWv4zUSDzGlWjdAKbH45sQWoNb4qeVpew+pCR9H4UC04Jf3OqdlPWUuinz
Rp/OLf/MQPLzT3MWIo5s4qdbUDJgbf46qxiu7ZlXTTGLA4cTw9DR2hIxDPn17SVj7SnDIASJx20a
o4OCp5xYIX1glTScp61JPIZsnJjn7PErk9Iv3kxIpivsPLOFBtOhQ4VJFYaGYG6bPLNrky4NRZd9
lSxjMbLIoIPz3BRNES8ZDMlcv0CKvrDNYgef5uDvH8Oua8eH6MD2AvF5pNY+IMoUWWi6kBS6AW6C
KEEbhOf4+v4gMjmBaOCyvNaxkScxDeSIfBNqci0Di2qOokZxwk/NmoNhbRtAyypnw7NFh96SaEj4
gm2U37iEWCfsczCsQ/jlqJZNdma8nXaD3i5ADRTLluYbXFfdKMy8/Tmn2cZ1ammGDeBd69xKuiOc
gFi6xEvPUhYYhI6V1U86zIO0xMmdxyxfDPT4ro19EpCNH+rre9hHYIlzndrmrQLvceKve6eKFmi/
5bk1xjqnp7u7tUPb2WUK6Mcev29x0InQSLAfe5F0GMRAW7JMco9WaM8AFGgKCaLTh6zzp64gpPiY
7JpH7nKmU0beENqbnZLr1uhSKTaD68HdoifkZyd52NyiKC8VME4QONhQ8pj1G2bfFSQn4HgmSvgQ
Qdk8wuecgzcZXriRARuB3VroSboQzY+ss0gl1amknyhes7cUYGizeqhkV7UgGRhFqBfpCy2Y1kk+
URtLxu9HD9VVWT/QFHNxCKz9aGWbTT1uMxqWj4muK8UGCQnL7BOeXRZqrMztcI57lffXPbvbzUyQ
5kF+2Qc5yaERjx5HUHpmF9pohglU5i6WWgYDkYzUf+d5M6DD+59AU1vDruaYUq3q19QvH0DWMsQg
RbICq/AeY2cBFZRL1ouX6/EQ+F90KMM2X65tFV8zwMRHmcEkxxtS4sSy7kRhdo+MJwv9SdelaZqe
doY+LK6sC7q19JtiIJPk3Ke7h3UuMAH5qZtxDEzvszOCr1k2qOxS5pnwxEePVMta7UvX2oTFtvaa
E+RW0+eokw0EbbbOvGie6T0KKdR/rW0d1xTyf5UbqD8s97V9NdxurqNLh7W4dxQirWlV2L4S0fUo
Lo7o/ho86yCKpJw3aw57zccizqfs5xnsIt4DU2qPDmvRJT1uoz6a92IGuWqVwyLxkK3ODVf2JKQt
m9GFSBKXRI0zaL+iUYkmodM89mneY48LRKnLxlSzIEYn0imq0F648vGj3pNObrLqMyKBAIucnoc1
+FMQLFET7KSFhFTG+LYXH3xU0yO0xfzcNaw44iyMyGOzopT13VW1nHm/1Y55IFapzpkFfIJAjYql
bvcJsLGE+5BFV/PJK35VZJFQoh82AvjQRfuHleE2S3S2AbQ3jYppBIYStmyCQrnP6m+lDdzL9any
js1arCp/sBCVq3tW/+DCwH2X/1LpO9fA8pBYYrAM94CP7dkRQ2OaQdtKMViJdw5KuH1KuArA+vv+
qsGAJdwPvgA+mf2so7kugy+1VxUzQTlZD/k2UXuI7WTM3/kA0NQ6l62j24IR/6xVzlH4frziPVS2
IVUhunTgLs2hYMNH8O3OFHtXXiV1hgjhuQq/tyicbxMJtAEy5tM+njTw1TCd0TZwHCi14Dd/tB+U
aV+n+1d7TXo4K1lTip5XgHybYUxDIBgJ9gtoPAAP4uuPoCknek1/i65negLjlK7wQ6fqLVRTkSKQ
0HVOS/zZgCZia2Ufo3hfqwVzqm4t662cmCmHE1s9MmPwESgskeyc46CgkYbI/CYuMH9wRfnDLsLn
hnWH+o2y+B2trWYr65mU9YqN64yLQ7FBeAWZVk4mGyKGni3ce+TLmY6IW5qylxG3EcU21qvZvtZu
qcB7XrxOa8epq40j5BdnImGEcVRAxxKBEE+0OSyZcVvD8q6zpQ/F7tlIbR9nKa/12KJec+FHVqi+
WQrIFQTZEaYsj4r9ck/IuBMVAC80Gv421WPmaiknxdg9HndTXYvMC0hd+/B0p6PEHAFqyM43aym7
pp45CKS6w4ZGG0QaJ9rflsWaaB9mGjjjY7MDXeFAj0OlA/I9w0G0M1vTkY8FtfWMsRDGgXkSWWey
AGVh00vitOj5DJdZXE5yIYKw/MFmYQf0WxctE9CRtbVY6OYQVCWo1PlNmbMLLVAfnQV2XIdzZPn0
W9y5dnSH/64FlYMKLt6t155YgbTcY9NgnHMKjMHzfpAZkQDOBD+AHy+AaKD8WrxHhErOrTJNrtfp
dq4nnHAbnOtwSDOENuZeQK2UEs+vFDII9gjM92ZT6+Xu3ov87HH4tsi/SYu8KCZa8IaW0OP+2tmH
R5+JNc1tBpmD1w7DVfT4f//3MToe+U0KJHNNXmIF/2nkzXkAd4DV1oZNeKGcEmn9XjEtvlyGNNIc
T15ebaBFLMJfC5eVtFkr3vc8b2KRpA0n+qjT8991vj8zhwvgu796gCXxu48cQIi1gA5Fl4RSc+5g
gUnZqo6HNpvK6tE05JXoBIIaeIZHnp5P+i1VwK7va5KGfyLoYgUncWyqG2gtIT9XSvCCC3EUpWxx
DAjUPnOukY1NImoM9bjE2/sz0DHVfR50Wp7MYyQT5svyW6j/mnvQnq8mK5QB77C9KabBIkZtYFP8
BnGY0MAp2ULZB7NjyrIJR3STuwuNbKnUcKtbHV0XdiDz3gslBw8x8ApE0MqnmwweNzdwe/WWg+bc
2Ud9rccpf9Azn08SmAV1TolhMb7XO8HW3DncA1QNh7Tgo1mbSBQy1RbY83ghRrXGI+F/V/iFSSGc
CJpvnsCqswjydyFni4r0ho+I9gX2CzPDyN7YqJLJQCGQMxAzXw8hbalIs6u3Skr1e3fvlbdAgaHv
HUdlwb8Zfl4hf+usgG7FEXfHACKxUG/vTzQoxKjREWMZJwJJf71lfCoDOCax/mf14bldEoGHTwdN
2QxT/jjzoMQ7ue9+l5fUcGlZj5hMdJCNllsE+ffTWilF30SbFbBcbMaHYpo8+zAh19s99h0tUbO5
QfBnTAHy6fAws4T7GHTyXY4CKoctpuuVuFwLFHbgW73Rbr1GC5toeH/Gz3UmQYMpreIpGniAS+cQ
bhmWH2CUZiSLANpSrsD7gBud1rpcWEXmk9UcW65FpsUDZp14b3UCRUhmUH/ZfjwBEza1xU+zCp0B
7ntWvbgxzinP+ghlKwo8lneHz2V5Y0GmNdE6d8h2GVZ1ImBGJvpxsg5RbyFVITdzqe4CFbub4+mZ
n0nG4rKO2VRkzR9CTcL4gKZkuYSSlrZH5yJ4WfB4kOZGibragmkmmtwNk0efqAG+tbzxachfw2th
gF3Tigpn5v1ltv7O56jKcFfLucBFsNV/ef5Av/KGzLQeBysMn7eKaLXgJq7Pb+VnfAWW0FNpRVJr
NVh+pcEcL1O1lBLY5hGgUJDTiy5XAB6lIswUuG87gK8AwTMLlF4vgk2tEydeBAs61ra8K4DIllX1
A2nnHsLEHZi2P0C73J1amA6DW6YrRWqqAYndH0EB7vT6UAum1ArYi+FgIMuLO1a61c9Rqw7xGB68
BjTidZ7GUhW6zPBAYdzI3vhVDSVnCli94nH9SHmGaWToQ73dgPHj7KIzf0pHkPlszDr9klBUlJTh
tn51Vc8QSLtDPEYZwEZ0cBrLyGI0O4867He5V9gFgsteioHpWe0sDZm6AtGXxrSNmAJDKVyGmBKJ
DMjF3FTvNML4egfbxpNUGrcaIQg7rUMK/oDCVsm92nNPPVBw8E0M8Sc6ZTV04YX3IL7h2OYjb26s
aijAb4eyMue9XxcO2uz6gWlJG00+h0HQWNYGh+C5or+p2loy7RWOdQXWB6yC5UML+GMll11GBj19
hgbPmZjVm7RlnKrHHNN0ukmfXWjLKimewiWLo+MqZoPMQkpbQDIdhReRpwzrOArSkVk2zK1WaRhx
EQQfQ0OodamzMOUu27x5wHc9tcmmr2O3DX6RhB+CsaJHLlVtAzyr0OR6M/6NAVYNKQZrbtljpz/+
rIzmnrDL68SfvG9Zji8OMrjMjUJMQtlgzZy0lZhzlpSuZ1WN4keuLF8oXktnft1cmwwQ8u8nAEcM
rlhckNxaNIOUWMlp2ngo2QF70meR3bF68ezeajoscf5J6LxAyoucubs0TEvFw84N6dPh0+NIV1lU
eI4dpSy3QY+MAfNGfNEvfQnx31itsOuY7wkgYELCcazsE8AiBQfDU1irNRRRMY7aUDCicedaFsnB
EAROGrOEpq9DvNS/svk3iDZi/dWzCVBXkZS4mxrP5CRKyppDzwAnA2/GDlx0zApdU5DP6hCNVdKK
eRmxUhJMc1xqnBQlhZm/emru4CuUYb6BgdVJR8CsCQWt/XsqZoNl1FM6NyotxuSUmPcQo9ZSiajO
+KKoOHfP1i7JKSh/NsV9Idbu5ODr398r2XKlDmJyB0lSs9LdVbkkQMxILeJlqcHs+Mrp3O6WdwQ3
wQSehpwkGpELDhNb1q2iw+ttr/oxh3I6QZ4wM6riwpe2Y9LmUJmv1ZG8kM2KToXcd0fz9uBHG9ZS
ygcLGRrunwywYyTV5Qcdt/yCnGhciRVzfkuBKi365L9Zo14tvde5Zpyt1pFu4K+DKeekpJbwOs3I
x0eUsknqkCYKBJUjs+tNYuHN0Qmat87ORFhCYPWeClLWm26izU+L71aO1NvsMQibimzfDb9E+Kqx
124SZLfIxCVYsHadQrREFkL48bcFuDAcsfKqblV9P04etCq/0rUfcd1bLIevXrbKaLPbd+EjRWdR
NC1e+EkNAV44XL46mLg9QDxKT6twrQne28WjQJxSfi1qja2EqHd97EQ7rfKXZJaH4u1Mb92piid+
KIrht1BF/Ns/+k+8ayY22u1a/6lsD/9q9OZD9mSnhFD0W5VlHpO04WarLEIEoKmRscnAfYTE0jDv
gXYiimf3OhGxfnETICm/pTkk90XeQBpn1nNxso4LyBw0OdE4bUINI6g9brboN7IYxK98xgAdEHag
tvXClDsb1loj+jiyJI4fF+g1YsRtZm3lukcGWc4H+CFDHxq8OaxBCQ+2E35FCvh2Wc2BM/Cd27ql
5L6tXISSX35z+PA3H0vs73hXuwiHAWhVgWai6YtobG7uLs1bZYfno3xgZ6gzngR/mKPGfoSav0I5
L5H/dLWR7oa5n+Im4M6U+fTc7EmqYPvZl93KzIuDcf5jdLH7JTW2tX7qpCaSuNjknexQemE4yWze
AH/vlnshGKZ8IdoWnttbp7sUe7JRtnaYSslYrMIqEapiYnIyCzki46TTO0daz4VFhqwbhnnE/hJ0
EnGTuNVbn1oCitnAxnmnkwi7HwwQqkS/+DVposooBkrRV/9ihhREQRcPRZ7HJvuGbs/erE7rt4Qg
tXZ1nwe6qkTB8VMXboGzld7KgnZILYZD2rmbJmNOAptEsjXBfZu010dwB6POWweNwNBbMLNEv/Ln
JfFWvuIjZTS4oyJ7fpFxZloIjlCNbHN9mK2O2M/UlpSjuujzSw9X0KMUExWfoSCmmuzXQPkaOHVm
eq3LT+wYx/ookbsncyYylwWzXsz7D4IGfKB4Mq7Hy7xvZ//v+0BtTE3c69xqSOO1FngEDrhp+drl
dVpPRE9P7dfePtitRTo2TD4mYhY9tsIQ5MKJ3eJP0ipw43CLUM3LQFudvyiB3h2kIxGcXBolovJ1
rjruH/2b80cSt3BpeXJ3zeRfMRoAEZo1N3BNH3ikcvsQzyQY1k+OyDF79MuUYJS7ASj54UlFrECh
mEVkZMik7243X08i3vF03vSLOFlvFYS0eeIQjI955MzZgPyRTIKFkK0R/1G4fC21hyyP5V6gva8+
BObHAWM/3WrlL5Hw6uETXpLOLwCy7j6tzZzXBhNjoiJbhb+8Wl1CvQjQpFi6inJfVzVxpVq5n3lP
0A9PYUMzyIqXsJHOxbxmh+D/4+xNR/hSLTiqzezPFZQ/ROub47KVvv4Jhob20+uJUCfQstb5DimX
I4LoXlKQkFSVK+dyWTX3Jg93bwNUKBhetfYh7wrSlIc0RO2QDAiwYQxkHyDMRgvAYLJ+vaU0wNLb
dQKXjHYg8du0jVpeOgeeN5dzmzlKK/JiYvigFlHTpbAWqjcWgblyqsQ/lwZxLmlS3R/SBiyR+kxn
CzAkUJL4vAvZGaf/CR4N5ev929+xCzVrmgciEDjBe5shx7/40r08MfCVzLlQwn8/lmqzHBe+/SDa
CPjQAZK26iCVIFZ9qy0xWa09kIAgpY0HRUeODaddJ89nht76E1jlkN3XshX5FfyjXc/hQK1fevxP
5fUCXxRcnfgJSMiXgHcvqDTE66Qr2p43hxJurpCcfD72VrxAFwbWDI+4LofvD0LbGjzPwbb/nl/o
p2GRblLA2jeAQsWz5AI1N/YhqMLzKi6M4b5zBqQJO6F5Cd+s7ipi9CED1B4PiXNbgH8qAsLDMhCF
/+Bz+/QpQ9XC/ldCyNyfjlue6ay7MGBdpLWerHCn26GzxJJ2xuz4R95/cBlst4GyX8vkqNulaKrM
ZFCK8npig66tguwqbKbnBSkt03MrNk1rY/ONMYVhK4K4JxVIt4zkBOuv+qlYUdTwbo8redhvghNO
n0J/Qs+cjW1jyEM1Cp7T4mr6pM8JaHxy31/2VTfYgzvDgajEgO3a4ia3PTVvN9vQh+JpCjsDKgSP
KURYtQFoiSC+iR5jMwGJtnoKKgRDzyGvw641bnTbYl/ZS8wjDeygMJUFOG+OoebgpjMBOE+4Z6VZ
Vg6a/OQF7DqOPht2miMyIjJPcxP7TT0rvU5K4lf+fa3DKd+usJyNqwFa5D+L78YC6TvM8QOtYcZi
yR1YmH8+RA4WJ/rPegXZakxcR266yd9YA/xdjCDZNQKpuPPwvDC/vqNg4B3CgVNbn72f3zdf2zQV
tZ4eBQq/+FpmWJym95MZad3NCoiMS+75S6dMU1LU0IuYb2TRlqj2nH4z83XMOsgx9xGHff21zX2L
ceYolN4/up52IZJMmaomaijcyfDPn7CJsI/K8oceRKOc0Zzwi/L0A429Fz/0I6CYXZvgnnzAaEIc
yDVCtx44b9iTK9YF9B1Iv41HWbGQT5VZQRmPCy/YcK0cm+HmZN2eg3Kb3zCtErA7hrkWqzkK4f60
VsQDnpkB5ONsj8sXntZ3qmc97VIKyW4oLdFdEeKKnH6hR/3LVqjaUqP0wrvE7zXKFxrsb1HHzqmv
vilw+x8MBsIMlP/FvZq3xkOL/ItFp+oyu86a3X/m2ktcmb4fjwoV+JxAsrSbEv92oXH1SN7HTDEM
bXXlL266gGHaLIYwW/Aci8wa2QU0/Icf0qeTfDybzPLYI16XBbwFUPfuTOQajChD+ow01QbOj/Ve
brhgHsOZppouNYwkkVVdtrmpT7m+icYeGhwg311Ts6YJWOifMH+MVyMZlleS/dN4EBQ/N2HAwZPv
lTTdBm5AQ+Na+I30uXgzWmTUbOdwGFs3O3oRHESVtlq0RuViCAxqKP4UUNZ2gAAjsdvXDbp1aiJL
cHJn+e8bZqYAOTsoPKPlpN3DyP7xz7Qew9bRg9Pxwy/KX7fl3+1KvQldQPFqyHZNDg9SSK5Bop/9
tChk+0HMoQp3r0GDmcobVFExnWc4I2G7weJjyqeuS5ZNcokOXwF/gZvfdSkxDos30Vm59TdfHHQD
CTYYrYQOfLmkN6gVmlxF/dttEmecrPvB1nU+f481j8u5KtHN5u+m7qxzBbD7z2zfu/0khdzdxU7k
O/pNqdPZZakEz+HzOSWIgpsL1GJoAJApuvC7cMkrpEtk1+mZgPh3jhzmQozIRXaIF8Ed6etNA93D
1nl399myokLlRVbaynPnwBmlnGgYRf02XG0BJr1+b6Lxe2WgfyxHLhLB2QYDSzPccX/eBEgC5za9
Cg2VsiLDRR3KRJU9fjVEB98doYUA3viCgynJ1hGqeUEtKIgYwOdRa0k5d5hZr54g89JNoP79oxdW
eVM0wD+MqlDdok2EZCnzVZd2mhJ8oLYuyEAgSs0/MxSgdySa5N3Nv9XPFSUSiHmxjDmKIZlUfAry
UBWp0lnnJs2tZ9DQUYhfx29dm39KiS4FXgW6hj5pmujZhjcwD/Ccv63bMm1gphVYBhFQXfv3EgSc
jW5QPN/cPYj+uFAUO2AEb47rtYqcsb9s/9zZC1M04TBdPyhUki3nwHGQrWywk4/y8xA0KeExChGe
bzMlbh8QsDPVByHSkosEGLUoGdzqVxPUOm6uz/Inx77onMSDdWYSST55opcAgpHdaJi1VMi5RF4U
dfSBp2YCAfyvqNxv+QcMlcO4AwBmdkWOKzbu/RPxxV9nMpE6DUw41J9PglagStXEhMylukf62686
fBfmVZgDweMGqaSKPmQmJFoLP28L7wvJorYxXZArRti/lVsUNFFd14CX2jFqNw9Wkw4dnzfOeBnj
O7TiB+EB1njhInNXplAH6NK+x9tJc1CygCmcmhEQvCItV/y6F0DuC0vwMxUhwUCXHKer3EKXqPd9
G2yztn/gHwFKK4Jk7uPhKJ0UYI9qwDi1eFsrL2VekkgGtr73l3XqknNqju3zgtJVFDcW46S6SuEV
pcR0d0Lw84KVYhPjuuQ7BhSq4cElgqG5HcI3ywS5TkWHqwtlNFia7LNyCdcBk2uG9Rsw0kdFUnf6
O8nLfur4tFqMdv4RFW1NoF1w0JSWvHhpx5EqeXX1/QAa8HgFxqY4ZY1eG3gedrAusi0xn/JXS8tA
1HiiNMmn7ZnpohzAN+l++F9mdX0bwbUyf3R6zoIcg5t/iMs2eiMO5wMA7Z4ETJMXDsA3d20MV5wk
bxiSMwypQ01qx+GAmoG1pts5jX0fxjibGkJ0o48S3WLFxTq9pGeFFJveX+LjZuYtyY1xX2XHp5pS
Msmoxce1HCpcO5/21XAX6xnCrDwbuTBsB2reMy7B9PqSLPKHLB9SPWXDLl1UhhrYItKGbRmiyT38
Zbulf+Q9pRY0p/+6Xhhnudyq3r0pR44X6mkWlGaIFywC4/x55sftoxvmmZjgXuGGnKF1JBVH3TYY
8xZT5/4rOuFVKvqy/dn9IH484ytq30FCH6Wh7sx/KzEGJzWOTG785TDt81PsjZBLmyHMybS/K3ls
f/BD5WULfXj7CWGtauQ5167ipyPVCJeU9Y7TqO9PeLS6zEsbS0fUEPhp7t14fhXVhL1MixtvsTIl
zCqzxSPdTS3Al1ND58cIG2n2JuzWTL3u9WE6cy+4mQALJU/nect7IQ/G3GIiDyr1FMuU70dJv5Lp
q71kbhCeD0gkNVRjHFsCBPI31mrTsu2ML2iI0V11ogz6zm8jVVbi9dfGapM6myWe/KtPQTaWmrKP
ChZEp0rlyATXPl5xkOqhp7oQ1nzEit6hdvPkG0p87tWJgm9l6Znbar3Okthpd7jwrSiY6Iwr3O0x
C5OOWvSUtTSuTwIvciAQZckO3zub7Y70Jn8nJUqMd62I2GCavFvzNCgj5LM2c/EPbQYeAQRaPIbD
K1SlvcfKAMHQHbXS6mSR8Phkzw2XzjVl9U7rqSH1Z8AM7WSVkmaEKYA/OknlDuDatXHo/AbpofIj
WvEqbJqqwI+E1aCkUEMCaQyuKLhYINID7tHRKTfazzudiefRQ61jrMvz66IuaiqlbtlFWUQJ6Xii
aHka+oqsnosBHboSabRdkpVtG/CmGXnCXhb07eLvdxDKtzpkPg6Kj9neIClCn4tQZTUsVVGKdHom
R44IOg8e7d4Aq6OD3qM/vFVP0EmchC2CdmrItd7lLasJKI2G9IBeCflmX6yqNnbTefvO4iSHEzBK
g+Z6uqjM6VfuPfxdURzVp0M5+BidIak5K41f42GjV2x3YywbIcvg544sWT6ERsqiZXV3X85S+spA
Eos6c0Lda7eZmpzr85jDnOvAuJnpGfRUWkjJn94ThoNwXCrflyhBFGMjeJslvE15J7GgeWO9RkM/
IbAp22A15Y8tMQn0cueXuouJE+ns+rlejQrMqSQ6dmWNGNLJKF1tlOA5Xk5TiIQ/lshXiwArSsEu
h8Y6KkZnyHyLaFcI8NnHaGYT2oiUKCE9FtQQHNAIWmS+rWARgEJzGfLblN7iPtm78x0xl69hXjbK
1ethDd8kOU1icGhVy9782gs+vv8RdK6XsG7eatEnHYm2w5v1gZKqVKOX2I7hZYUQ3ngXyCNxgXad
FV+0d4vQKp/PMIDay5v+t1uj3HxmV5s3pW6NfhMKMp5rbJXZU/fZHVAvCXHgBELxvjopwUXfHVGj
C2OUi9Jal/t17QqUFVsk82OokNAISs7sKUB9IMvFQ7xwKoTqdXNfKB/u8T3amox1IlwunpPn0uEa
WtwxGQX3VtgrV3ipHdqHUc6rGmnvxmbdA9zggiCiptNV6jkc5beHKj2xrCDqJ99wqw8U5Hls14f3
vf17RPSlW5mZa9it+iv1RM5G5NHzrSUCnjUcsRDGRBhLRaLSok/OZjHKQ9W1CeJC+SVlOKrwB5u6
vxjh8s0Fx5LhqP0WPZ/QkQUH9Gfd+GO9CIG4QN6Cf+2w4JvFyKdROs4NyO1rR7JqSqGEmrnFo6Aa
NsP4D0CGazct8DW2RT4Fp3VOhvTU25XRLqwxLj4rW7ySZxoF2uTV/jgwkMX7eMPhwzdYeOXG3zxG
j4ssLaS9wBavdt8xocTCMUVBXb1ybDv/TI5Y4fVeKm4rrXaHontxC/PCcbLZFjCR96PBskYxBa6M
jf0hfQTmwmUatx1StdRyBApwsiYdraGYXbP2ovGj92tHUIckHM3xG32X8Qj1xY9jngyGjNxvFqKA
fCtvUqRc434kfzZAezc5JuZK5GudetjHkUc0Xoy1dh2fuwVCgSFylYxYeoDmAGS1o3zHyI/IjfMz
4UbPfKM44BNIhN6DDOPiolydRaRuxlUhBE6CNju4vE6wOwXWT0llQp4g7u+i28SaCDnR1isVUGed
0Apw2Z8V9Bf6a08aHMPsynRUFoWa0EiLYxhl5cMK6jQQFubxWvUSkNQRQ43PwbB1XAhqTvf0P3if
9p6os/arFtDVY9NJhIugceH9EyCasSSxmBaQqEmGMnbcvYi+NUFBktoAZ0YVJ62u/RvVr/cC9RU7
l/nDQ9+uYn+ag8ZB5Arw6EN5dnGtz7rjVPmmmREHkX/3IZAa5TI1tUJIUF8MuqKKnS3Ccl56MhKS
rJ+NImN04DmOhrJy9uCj8IEmzsrKqsE4kfSakssueNxCbUnfYaxGbouW7b/dCWXCKfbyTPm6KUtk
ZxMTBh3Sx5NReu91OU0coD9+AcvVUqswvob8ylPp7MLRxMB0i/mboxYadN7LpyydvayYfGaBmqHL
iMVODhOzgj+RPOEyBF4ir9MF3326ztGeyXwbX8S/4fQryqVLHRBOysgeIlNLaLbOeA6K/PhFy4bY
dl2GIGJmehHIb9ilRrE0k0FPQ6yMqmYqePnZFcUrtlVIy2k2syTV5JjfsRXWJNGHJ/HCERmlvNw+
XC9RuNiECVxT/8Lu80KcjhXcim5jBMB8uwPlhLbBnxPplhfooH6Ssgefkz3eCjYZPS2dm8Er6CTR
swQDcvNFo0JbdPmuB6WZQAa+qwWpPJmnA+4IH1+HqrHVudazyDueWhX7w7OWgZgpDQ3CJN8FBVIX
cN6Yuou4ewm7zQ8ZHqhwtnixGm+6zLiOhfvVWOnKL4VBzM9hcfNuRlW0a5cQ/W1lIE8mGXzLoMob
RIDvMJ0feD2d5RYFUX5SYy9mbuNgpUXoE/L+VR0TWUG28IkkAqTdtjQL9E42YsoFczMltGGqyKnh
VAg3kAwcaY0ivnTt1Ry1G0eMlw1LweVEp3GKMSrGy8UzGTcR3tN8c3X9eyUEyK41olTgmTI5Z8Ck
+2h1JAYMCPxmhJDxZ4dUhWM7/RhKRfeR6ZJRAZEf+sAzG9fNWDsoedpkqdozL7i8n9wreFhd/WxV
NSaS9mo0gp6EmgnB0Xee7SuS0/g84ybhBXjIsOTF7pcZckZJrlx5Jx7Sv0zdRUDR3Mu+ZxzB8bQT
sfStAV1iHFrIUnlvyCY9TBKbyv40/HaFqRInBLQxA0e5nU1HJtYgapP8LIh19vSEufwrEByrBJNX
EQlpikxSmq8vW+CORIVVR9RKZ6tLY9P0GTj7lxJZsMG2LU9q0KOrbQuDIbZnCuinXzQ8zxRTHdfw
QZJPVwiORHtOBtrCW9ZE9qctJXyC3ftJoaHEe6tl1oRg0220AxhPdoDDtHj0nnyrtBT4YfqvQ2KG
aEVER20bOHzrzlBzoe62sWW6DcuYaDRbzS5fikYdv3708da/66AZEBAOfnTbfbtZNP8jJ4j2C+SE
feUXLvAbsYqvHyDYpzlOfacErzR6GNq4xd+4Oaxq3m1+uxJCCaQAFNstX6xGsXysBAF/DOY3ArXO
fULFGLPpMJD4uIVMhr/SfVB7aeWq1ID+2Zae9R0reb7I5dUI1P6DSilaiCrIVC7CCyz8sO6NQQoS
IZDU2jh/M7RJD36HjNuRuOjb3EjBApgKpBbtrlShgSngBZ+UiuN8zlRrTR2h/uAq9tx8wQAdP0am
3YiknrD0VwuNUxJ00jawmsV8jysurdWnIinEz7gPBsy9oWoFNZEvLxK2OZuTpDso1c2oTKawF9JD
7E40VN0W5YYrILe7y7IICTukXnfdEAxRgqYq8DGnB8tVGiroWA1Ob/Wi81/ZZ8u+3wIm7KMto/fv
Ts1IbrCcntf4BnCXKzgeZkvjDpU2ksVkaK89r/nWGw060p8GIXvVrnRidOHDJ9YbJ5yYbdnjepBE
CQ03GGw2fK9WCPdjea3cZ6KpF2T+e3BIIBgpnMkw6TC83rI4TSHuxnOEULmneL7V5c+wvlTJyqS1
ddmJ43sDzQGVVsoKO2PQSLsu6tF2JR4KCAblbccPN4HG0EwiGJpAVuACMza6HbLILrZmBX1o4jBF
sVOkgQEl2Jqz/knqKbISW3zIuemXcRI2jpo7C8J11FEGtlXzk+bPfmnQEfqiv7FOpDOcnJr01c5f
QUTsXueFjJytVHAlzGt5mBveT86zcEGiq4/UVBFjRcCxEukZp8hKUUvFUNfDEcBIJtwfipHKaSGc
0Wqf6/7HOpjxYOsPuhXH/OPkg9v9DToZESEUPmXqjb3VHm6v5MR458mw4H/1iDOWchnWYiq0pWlt
XI1QR+7k4x7fvw3mV5rpqeb1ORCTEvDupyx89kXwJvugPQXISdbJyOP77Mbzvwbql2JiR4VQ4iI+
J/XXZTSTRCphtvUSxehtYgqLNUl7dNNDOxzKGlDZS5hSjDeAwjsf/wh+sYUiJ9WSEtz94wVwNOPE
oe0yx94vduG+Z6qKMA8DOauV7pp7bcoX1NrQlIUe/DtBcOk20fj5m75pFgS40aWjsiUGhkhPhvF5
JURxxOPfL/0P89md93xFgAZ4QGAQm/7sjlpK9VnVQ91KIh+tDWprc4Xq4KS8IUeqZMQjHtZUVq+C
CCmCfNzFM6RzEGAEldER0Ok2ej/Ak8yZwlD7TjUeeymBqVYvLOZ0nxL/u9Ee6z8Sh/vqWkAYEchm
PBpXmXXvegXfMQVTaF9FwH2uHHpMdLHQ3E11Q+Jb8p06izcDr3HnZOd/D76S4j32MPuCJ7OZv1gW
IEzDj/dnW1OYdOdcMcw4afiNqYQu9RCp0pH01INO69WAoLj6jyLreVv9iTgskg5GvMRVpDctAe01
mTvOaFxAu4P7Pm7D3iNURCzXgT4fA8DE7x6f3Qrxqu8ywoIiHLVhwQtJ9z75168TaCExP2Bd1TiN
uA0S5crS6IESH8xkB5q2KbkHQi5cWS711Sh11Ok36JEtC9yw9L0ufv3TiaI84vmX/uWg3274GbaG
+XMC17KEVqVOURGeHfpBi4cSSey34X/nkkkBaAZm21zYMFrLo8TiQc2mKN4KJPvj2XVU0lywMXht
JGM8Va9BqlPf77phMdM+W+KrYfOvLDTFKtqbAAQr1ayDYSdKZRU0uaLiWblqU/sblXUyF5KI5VHd
Cy82BXJuR6y+fHycxX7yv6FzjwLK+Nn7E1cyMPGk7UtzakRUkBSnRPvltLGE8LJnau2nssIHYkMj
rlDJI8wKo5xOoEewAK1HcFSSIBXGMyWzJUOSdH8fhuQsE4GjMiXRj4Mc4OiY9RUHlFa8pcKeBmHD
P5FuvHZq8qFJD2Ne0C7bH3UVlU+8W/ptEl6C+r9VoRDz+i5aE7PF9lUMRqRs+W5V8hZIZzz9b8jd
gKeWI0iNHYLuBKOvaWrAKAN5wjNTd0ZwuFzryEPAzuprqwjkNtoJ0h/0F+kqa8iNaS0u9zWgI11v
+XrVRX2W9AcpSp7eVurwYSyrmvJHO3Fd3O3YXJ1/IFGoQR60g5IZXVqWK8P3IOpmEuS/yMEOQ3uS
FAawX5rmdSiG7X7eBIwJi4H+1aar9aout4gOSlJ0d8SgXHqJzFUnLv72NrieFV5xBMD1RovwvV9w
IHGPE/uwTEouLj+9lpxBJYdbewxMtVHtGY0BbnjJH0+D/vmgrCJllrpzZWP2yjd+C4pyuidCzAwx
SS82qmhva2BIwcq4NfIBiyQQqjYLCnffDU0z6ivxcmJW1MR+sBYigStqgKEEpX+yHGbv8FtooF/N
kDoaj18S9ztKI9/fDs5PAd3XghbhB1r8zjxWca5bCjsZOFlwj4ZeR2b5B8PzRj5yj4qCUlZv/8OA
1CWtzXu0KwMX1QpgIn0s5jObwv46CcrndK4gt8Xszu3cUUG6cl5RP1VFA/EYLB4NX3GyxFJj6BVo
RUGGW7/RA+aZmp1JcoiHwN2a1ii66y/JQWr97nMlVInw/KGodHVVh1aOk2Ngc0ZuF92IqD//xOTo
2PtEqU1nWHfasSE8CSMqcgNr/ICSoKOK+iN02WSIvZQgYzkdeCPo2q8lxhc1iSjQ0qTx3B4S34ZT
DNoIvV+l/RmIXrWFRGELjmScZ5Kb14hpFQ0E7rywOohEKAJmmGJbYwLpqiNYKHzMB2voJWonZVeD
fO/2KbrAtaHln9fOHT9mvURGJrKk8xaD1afNc3eFIfbqUS6EfRicevtaY567gOJmllI8hgfoU0tc
HdSfbf8mE6DkFCCeV4a2QZGIRM7BbgNv2X7W10jF/zI7xdMxV7ApmEaTeKfLILVCvHnZ8zwxf/jS
rpS5G38uJnYV+9cS41Un/5giZDwcSUqj3CsBBELgJZkBm+SzYew9pvZBJ8GkCNqKtsy9uwxHVNPJ
dBkKexVqnmwuwRJbjHg80KmwxJLwkUHAN0Y+Xpz342AH0MIzntLHdvAeW/CCZW5K39R2gY5oBqKm
XTHPtQbkoeYHT85aUFTQStwQCuMdfAxRU+Ht0ebgv3YUDeQdsJ1tDjSorr6rTNyubx8d9maaGq1l
eedVQNgxjf49h4E6WpUdJDgGeF4bOpV+c5WM7Plg02KbRJfHIUb/YdxB/tZMFUTyWlO9cJi+f3m0
RTHFAhPwZoAC5RlpXRCNmBOSECHAEIodBPadN0UH1GRvJytPsqJHJUM/+ky8zPbqjfrFhEoAQ2af
Bj9bBn7ozHyBBMMlRFvZgbxmdU2jXv979XxAdiJeTJRc/gwyuD8JDhE9uJBQzLuIWbrawA/Hl0SB
BUMjn+8Eblia704CnUEhhCcFfWxJyNtmHhEefey84gPZCJixJYFcBdqNlGi9ZJtkDtfLyOvFIctc
t3OFBIVuwJRgN52IV2/4K7HfWJOrNi5XI0E7lFjEsUCCd/LqbK3W+TPHYfuOYLoBSrKl7p6V34Pr
PCwUscYOpZALZ/JbbCqW53cJwGdfTq6DfQE4XVQVMrFQlVXttaFbbCq+QZneKrIEjIXxhmdLbG71
XiXTkMI0/jFVzLNOiMMVdxK/AtyR0ZwIUYql+6LDPTLzemcRLgqLtXzMxYETzkMACy4YDWRez5ar
2mlkDs3wThKS3GPGeisSHPN4Og4rnQCcT0Q3M20gCRQryGZGRvOiuF6d19iq1egJjhB8u6HJn6VU
T4UAOzmfK/JkFARpTBNGEgyAe8US/Q9i+e4Wt4MlhdWzJIo3Taflz6YidaRAb9gidk9PKHQmdaGm
wTr9lEeUzMaEmBllPpq5WzHZtgt3vG+q1Q08+fpcLjwtY7JW9xXQzvj1pbh7AvrfZe6+SkJk9jmg
pxlRtGE3Ib5upxei//XziDwTdSYEMC02QQABVa02CpWLg4TkepDxqrulXmC5NOjnwSfE1xbFdwy0
XX1vWT8PAM3mYRagOFw4HFWEf+CNMe603JitwaHhTjY9N0cYzj37+nAHRIuEAcrlCscZyJI28JIw
CJi8yTdIyaE0UngGu4EmBcoEBPJCb88zzDIbKivjkaBBFH7/BGG98WAYDVfnXZIj/AfeEsDm7EIU
PWnLe0urAFe+K7zcIGS3sSIMWe09nPyXBvd27M+nDxnLVxDGPAr4RYUJY/6DM0yi887rbFUBZ9Dr
0kIsg98mflFOpLrAGIv5/tYuB8LW0yMvHe2IuU7JcSmPEr/Ej3EVYlR/fmXPayOJLl7aR/dV6Uam
vDGAlsFNMIhYsEYXMNdA2GrUD0Vu+4ICL1xtQZpMQBi2FsxXrAA/QuwY2z2V6DllzRgPUSCd89Zb
B53vwksIWCpsI1xPTeEf4Q2vGseMooo0lll+w8EQhay9Wdb4oRfKrPBelHq+KEGwik5IXAATswXB
ECDCzEivxpmbLrd4UUuTxBWUQP1I5laCo+FAen+Gm7kWnOTPzReB91M/iMzRaR1eIKc70amNHyd5
AOyIITzxkWGNdEV/onbtdvfwAUA4sXKovVQlmdoydmE8vGk0uIrBmUrZTsv1MMmcwnqND5477YB5
1PHfq4tM/L3RV1ThmAGnGMsEle16UG22/QvnsOnsODbPBieYt0ljG9diDjjupMoQv6KsCCiwof/F
ODYu0CZDojwq76/Ipmq94zlsjQKPTuctywx+rtZW/lsfMt8ex46wS8eRZM0OV99E5Wq80eQCWAlE
ODhiMDOnuUza923NKxXIG5DZSK1OeZ74dPt0deCbdVPAUbi3qVLZ3GhV4eStlA01Z2k1KvVS1s13
XI/BAYxJDN2tArUSLmXuJSFSkp13iUuaaV+z/SrFEKAMecR7wXbfDU/O70dmFOkIz8Hufk88h5r3
n58mMqEFBBKcaOeU9fV9Papisd2NB5tYFV6qYKOCvIijrAwjm9mK8LhW+hBxLaDJJdzAsI5klP/1
jlA/2u06FLjyRyq+AVAUZggqNVFwOFnYIKwoBUpEdjs6e3ehRmpe5p0DMTeVJdzhM3OaASxU2pB3
Q9gwbc2G1eTU1ndcLNlva2CwZZo2azVxXeCrGymZdi8LxbhiLnUn2yLpYzyzqS7WlrQQSh5iACZ9
81z+hS8ieAQY69TAWciH1aMYXbM0HcBsJY7GYY8omHuutzyNyMYEOWfEEPJJcM9+uwDpwzgNgMqP
sJZ4GMdvMRROmVyAHyZWcC0Dap8sYhaxATcbtaBk6LiKpz1fo7+itP+owV2/4QNQOCFTiNOiNvUv
AlDdCJBGH39j/T7QP2kmvB/yJvuB0et+NvBlu45DHjawXPHmlhswPNzGwci8f52TKMv6pPlFoBnl
CJuveXhZ3fOBEkUG/uXJ2dBB8ctUeX+n+kCgWNM6qgat4xPDZ2k8jLukJW2yi9HJs8WJff6oWcuL
xQP7rJmiVaLh6469yBk3dSc47VU0JMArlQchdeaG5OqznSUplZO4iA4+YQtJAb4N0yyzYqwxdujg
vjCu6tqzXJ7LInOuxvWpe5K8Pz+FO26sWjPL0hn1gDfEJdCZHiZFwceyAxYNFvA8+SLS2O//gjvX
mJhAjRa2ymuMRNxn+R53Z767e+XT57vstTiOw6blfvuC8tN5OZpuT8KBbOt5SnNhBmMxyH1cwfE1
BvDVB/VMg4fGARQZ/6JuyGzWPySoMuCjnTQu+lpPycTdC0yJgaD10dU8kECyrQbr26G94UFjGlVC
26j+BUdfCNHp/byfN+nZrEpAOWhztWe6dvqZG1vQANeYoB1pNogiTtVw1vRr+ty0+48+1C9a1KaI
xv2zoN0oVpO9vB+91egbuQQrzPmOutwjf2xTNN/omthmLBD4rXtvf3H30HbyXx+5R1ZefQZ74J7y
avgNZj9EyM/ATaWS67FFJURb/xwJJyH9lmQy43ZaA/mUtiaVuLKnzsPMgYAixEAfbFbid1YRMW25
d74vp6HglBH2DuMHCCc7QOpo6Lsorv3ecwNwkZ74FgnDyQyV9lPKutl9SYtGGGyOAV71IgcjQleM
oU1Tzcdhz9uC1nod+FQlGCpFUBKROZxqy8ZV4xJ/Dac6kdywIS4c1FJ8LKuyGy5iDZJ7wIMJB7M1
jZW6gOb8nhCeBStgfKRoTPRy5GbatcRQTrOLwKHrt9GutJdInD+be2Ajt9llO1ha6Ak5DMXLS9Ej
2LFPcMbWBNikj2KAKQpjzBATUF7BIQppTiSyHa6r2RszjLJOluAawToI5JAXLLVdG1PBDk8o/+5f
4UQhIbBL8ZSeVHew1c+TCPZGFdFHdYrBSTkN+9WYRJDFbQq74Zw1wAtB3tZlZWfX9UK2NvYB4cid
6jFmZJqL4rgLTsT2ug564IhjMySZwz+oM8+xfjG0ojsY0O2rWOWgYKY1IgsfEb2IUyg8N2HdybKh
6ZFXOG7iwDvkN3etYRfcytREPSdePnLwOkrqQKX2DZrBDTitLkAMoeyUYqGZC2WRK6mUMFIRPzvo
UONOkjOhi0LLa9iNbVxtotAu8kYw3BVrmx71OH0QiD6uK5FZIy49qObp+iU/o2AvpjwgPs0ieYGK
p6IZapDJZB/TaM6e3IFNhJEcfPSZis9vLe9/vQiCNgVoP8Y80OlLKH3v4/bhYJUaNJbzwSCdcvFn
HG6cqteO15yD6RaMSMKqwN2h2qvUL/A6moj4DmMeVnUEJR9slU9iQDUux+TxKuuEiizJ8zMpG1CW
JTHCDYSux/rLlFMaVi/R8cAf5TITYpsp7eivz450RYN+D5M44IixNW3UapyC+JzJW+ZczpgAC0Ay
DkCeYyyvtj7siC6sts5ZmMZqOZeAgZol+lgJxJ7kvnH+BxzNeJP4SRwDxVihnNp8nHixlNczTq+F
o+kLPt6gouZTuuvl+SVKSgD3mWesZ1kjmc0Gyv4nIuYFkzi7q5w0nldIgE1P6ydcQj8yvttj0vGX
KU5VeMbuUNEwonxgpTy63dSXcmEs14cX4IF/IbFLhT3E+qfdhma2Y1ZkCsHaSVM9himRUI7qZlUK
kPTsqXQZhx2kSkX2oygrrjFD5G51MjkqfLdXLX4ZdhPUG6UakdrP1uD2ja+TtroNO0nUXBVO7YJi
eqmMPOilokAwaSIDXlWmTC7Y7qyC2sSloKvO3YOfj1iPYmZ+czb0fMJvwbHhRMlGn3Gj9CdhCxkj
opartaUlqoGiub8ZFIlPZtZkeCwxs+ajhyVjjb1PVHKKLOWIwN80N7aH7P2jxYIq5IIm/orAMetw
qVUAA0KZKR9qWuhhz+krMcPoRafrdD0sR4AGGzNb25NcqaSPhbHQl/yJrQGlp1iEADD8QtWU6Yzw
wpyLYW4wYvlMasklGjRkDIcCMM2aQjocZtlOYgDLVpufkIGBp0MV6Rm1GUJBwPOicjKp8lBGSgUC
fFPHvve6ZYt2eFaLjIvgwBi+ntDf6Im91TiJNdC6YuEesJVKb3D1R1F1/WHZ4O/vfKxXyiR9xyAk
nTaaZ/prqhVzcPYnFhIvHOuGVzELIOP2bBs2hIxmxqqDAS1qOOJ36Hg+ChHqilNfnFijqvUTN4g9
7DZrXvBvwv5Bqlho58NtFgXVXDfx637RHFr4OLEcIJpC7eMOyXq83BaKOx/YZ8Z/FvsbEaX5HBbU
9q8njy46rpbyk4mBsUi6FdjqpuMa8vV1HM2oFR6u1rxkcE7xFgmmKs0qXv7UHWeN1ZPxq/DkRK+y
6Df/4fhyIj0QDXXahGx8H7s67EDqKYj5pj3D375JcARZf4ZzrWd6QkTCu22WS50Huz9ZC4/g8S/z
klblY/wCW0mWwcJkaFZBIPd1JSwBvcj0EjbWD43gisp0rf5kMy7zdl+/OWsPtV5Wi9vZJYKf0HnB
jjObTZsW9dYdVYrFLHB74VTNrLYXP26eA16quIJEdiapW+VIICfiZExwlajtJGTJr6y/o0E04pxF
TT/DYFaBdzeR8RsNf7fJTQZ++XfgpKZaLOhoQa3WYrU6boMpTXWH9BQHzglg8VvSV+ZPdG+ClL8B
u+S03IA30FIbkFqTBvxqNnTyiG4r7gS9s9+EN14hzJBoBKfECh3Meh58gv9CcvKvH8L/tRzAv+Pz
ro5a6c9mc5KmQYwQaVis5a2hqXtCpWbQ7/84IagjnivE4yS4+BVA4wRBEbi+wRXT0BC0fPs3KxA9
fcFp/vCRKk1GZrULJ6BtNYnbE3xpS7fX3E3yJcdlKAK2AvS2kaN0+5Ze+UFMVkzIo+Zup4IvDUsp
9G40aSwau7nPxzKLJIq/GzHaZXT203upiQpY3ByB/kUPX8zWeHt1LvJQ0N3Zj6TJ0i7vqjXcxnxk
t6iDxCJ1JnWpbSgLuhKEO06UNj7C1u1kLU1ANSmkeoMV5GdwF1kCAWQCkG6DJrwyT+soVyzpqSdG
2sH3wDpoBnGWtEfXD8odQ+zpV+1zST87B/684Fc+tBe9JYy39Vw/86IoGsU5aIsEu1HPz8SAyIiM
uBMhGww2CQ9RD22mnNvC1Kz/RJpRToJBI73Pz13/TLzZZWFev2quCu6bqNT2gZ1SMCyQUAigz/Tm
RRWoihMwq9s1emk4SMfp+TRexT5PmwGHY1nXSQ+I24VYOU+NZZwi19toc9XGC8I9bHntMZVhqXvQ
MtBQGxENfuWFznaOFLJk/RiomkEPaU3nRzQxcfcKKqBB7dTf3lHshvPp4S5gJRV3BZlLhQT/kTgw
ks9CitJ8kGYvqtlW/oSktw5ZuCJJ99BYIdoeUbnJeng5wWFj8gGBw9qy88qaFWrTv+5QcRP/HxhF
86UZE+VWUlVsjUclWlrFFkMFPlltIsAIxkWDzLgZ0XBRQGqsJjS4jcseYH8tMk0GKk9+Bomm0eJr
2bJLBIgg/2kmLuJaE67JaEzso3ky6szw7yBg00r3TiXeu4uRu1sWZV+1YIYePY+33qNg0cMNi7KS
RV7CnZKFSJw6mSKc1GgomivflR07Rr4o6bcmSRoK1bIn0/I6fzncoN2+hG2RfaIYqCBvIw8HvheD
09zUPTlr4ot/nP2D0/xeVyeq0eCU8rEEMA7VcKMcBm1ZsmzfYWp6zwbep5fiBGPZE3AZpfqqtE0W
FMTIgQWui3E6Dr7hFPG4VDmiSOhO5REAH+DdjBQo8uQRo+o3rmTwBOhHxFXuzVG8QL58CLGLakeZ
D8fJjTOSdfUrF4+uVaXHHrid7yAM+af+D3HLLm3NI1KmzXEBr6tYzoVGONhjGz7v5fxnruWDw9+O
EnBNNMO3UISBzAQNuT741gRnrmiC4yfGq/G7K7+6kKgkkSvZGSwq658hasS242M1Q/ZuEe8AGBn9
z+4OraT1/eeHs7zN7oh4ThShjd2vmoDwR4hecAu4/zwOLWaW95Twa2CrKOljyv27PoOqaItYni+q
P3L1qinGoPFrumi2PbyU6hS9rjq7q8h9lno1lZb/epiLn4nqxuNU66TaK/asACP6HAVb8MSSUSc8
fyAVKyGryf2tuh3cTvxyxO+dzip1llJs5khtxS2h3ItmUdC1/BBAxSLlkgbg/0I5XRhQBQSCux1o
fgym9VxX4rDX0Mk4sYHxLYArMNN+mIUSSMqnSD0sSNBCCQ6ZsF9lOLygoA8LH5V7v/IuYC/YsBmb
1et05LZkFgyTxLGW+pq9BxZqhR8X6OB0pbC3ur2FQn+0v3E/ySYRSLZMmWEz2ZFW2oNYNgeoF0RD
bYu4Mi3sQL4A/VTz4EZrvTIefoYsU/wV87dpgTKvdCfsJin81CgKrlce5xbXXtxWx4h9xQ3HTRQR
kSdBDKlglLjc4uG6+x9RA+MlU2fXvfF5jFMsOaie3nme71QP85w8nAkRpPhZI4sSTSTIEdOVt6pt
I+ntOm46t3itN/4S/eThRhaySk0Ixq9BGrnxFn99F3XGZiTM1gFkwBxzsAj/e8CoFC6t2fPxQRSF
IsL8dkEpDn5IWub3NcXf0zGykUi6K1p7h6c3ivgkLDLSrxxBxy76Zz7q5x2IFhYm94FPtRADkAiO
B4bMp/CQxXYauccApvlV9ik9DTPbkjR++dgXnnuf/22M91qXsulPRLMut0u0fgCDgCRglIH+gRX7
RmhxNa95w7cf5GCtlLo/rwzQSV5S6GHsjc29edsefV7eflYsIuzgCzXAxudjAyIZUBFwAQE0sBlQ
mGfp+EXC9oY+vw46UdFYlLC8FdzeqJ6ju88HVAx3onrw7llSk2YGSNpkhAjt4pqpdnpK3tPBTRw/
WGk9Q6SjC0VEGw5aSr8LnK0aP0L+XB/9WG7tDUhsn6cbTotuJf0bXKpspXDTle88sFPWVDynY9Xa
hoj9K+jCib1bjwrzrlkCPIDZvK+SBxAN8euLgb0a27iK0CElLdlp8meckC7Bodbbq+2o996n6Afe
JrgBPLoRXgGna8O/N8J7ZG0H69EmxnEYZ3b+12QVkl3nmo6A96cmBK9gAGRyrucaA3P7eGaTDAAW
85BavUUnmdI9rnBMJG0IPfb7+oxwtAaYGMQhE97QE6VEkfXGIYAgshkh+S0OalFSnSKefiZykHgp
y6U8ZpUue+uILbK99iNuhO7oHy6eUoxi/i1unkPTZYgpQIdCOxoVmBNxUaNG0G3PlX2r3JcaUZDC
Y0us/JPMUyStB9FtHFTOnFQuzLm8BtFR9d31eUUb+e4N4fEAfN4EHJN+ESYxsK6TR63h3w7AETRR
hEV4GxulHfF7X0lwJdf3017+k1yxELdjksFQEw54+qBb9VWsLg4piwgYe8NKDaQqegmD1KSD7D1d
IrekQQpSCXHFSUGUnEzYnkKsaNF9B+0lY8HtEPnTHUop43z038/Vqc3RKgVqbLZPOgkqHn0q6oX5
q4/k0IsSOwSiLxj6oMUGAG63JHnJXmnJN4YdeQu16JHzyoSnD52Q8B5lHKMc7gpXJ3JascYGH7oC
p3GRswRnsY4dw5MHrDB7fWx73xSHtqlgG8NLyGgVyL8m9mD3cD678siQSExvbI10Lhzu+VeMrvm9
KTimjkyHFrr3yxVb1odcJ9CsG13mAha8IocWiHOtufbPzeNbXl4CtLso4BKb7ODKdWv8m2z7uuUn
4U/TYUAFFUuKQ3zqlaT3Q1cgluQBW/xsS3ushDHrs+SA6R4SsfougbBuNjheBDpsXljqpcc2Qiw2
0aqy+1XSqTL0xjrTPCd57arKCgopmLxE5yS3ojZfVcc3mv/P/DG6Wl10Q3p+7IuFOKwpIHipKKj+
Yk29eyYGPoCuE+6yjFhTID64/kCzgGgt2G4SVWe3WNZptXsYEXW+faH6fdrzBDN46A/1H7DmstN2
lDuD5aG5ZURflWzPrGsiRbOrMFMvVXJyW6r6EZafsTwS7vg9rrsqNi6BQrYrnTPpzOQ6+ermJ/nF
+gi9YK/k6C2RqNyOGk/BLJjQt7sFkWmsXGyl1lTPVwZle8mMITv6BVGSP0NR3Joj6M0cS3j+Njsn
f1Kktx0y3Aqw9G7bv88aXoIxDCwlaOK3rHsp9uh2PBM4sqjRvICCVOQOjF1sCx6K/lj/28lpdRsH
jL3kj3sgryjGAAwDQRgL/CXSp9eFl5QK8KW+fFSA3Xox/rtG+5xrf6v/62PYSuTnC5UQpcS/QUAn
I84t29yeY0iK1b17809qxM4BfGoqKqCcfG+jJ1j0DHRSwPNJcMAHkpze0eFlndN3Jzgz2mh1XBOS
EJ8JouuAuSq4uaWPNik0Jbl57qItg9xDwAdWEfOz3fFb8E3LX5GU4dwBBCWt6v0uXSYPUQycwCPi
vtyEv/gR4HVVYlfhdzglFLvehzVW4V92PmEfWhO0yb/1L/SY8+G6N0O9B8gRObbfDfHTmd6lWbFq
tWyQs0dBOrEHPA5ii8rfp/hPpw4jBuTFy1mFoQcUd5RnYTjU3I2DpgUhf/rvL1dvAu8s0WuzsloV
uylEhRd1ij5JvzzkAHD4gfLArjwUYIMmogwsAutCD8pXRSxOR5tQJDq1v0LZfl20Zlaxo8eyHCRs
aI9SfOuL2IYOPjytvVUrJ6MqcZQTeuedbSc29oq7OzD7wAFUTWiJkbFsgfsKmbtsSBONeqVBAQcc
9l+cx31GjXN+h43RSV8a+gujFAn+u+WKr6zGex44u7113bVCuHCKIPf08FMKBjljO+/OC1UtzBB6
w4dvYHsmktqix+RwI+5pyuHfDPa8A8nBDtpow57CGbEU9eq8jnkVdasw9mCRgLtcsmFfyJ8SpCxR
ykXPJNGho7vjYA1yy1sHK5mba5fFBBkNDqGluPMW2yO+Qjsiw54x8vpNp7iTJqu9I5tvLUoOMmOp
dx647OdoT/AdpAxWQUfSw9UL2G4PtMlK10kANZk6hepDT4T3TvpQLZ56B3L7lfM+Vxf3m/Xq85vm
CElk8DhEqwLm1W9sIpumBqoSxC0ZIlwRns7Q6cQ56UF9YL9MhSJe9OiQrkipXlCzcFoJpBkgWnAh
KWAaznRR9OOxuMEuc/E/1mcK66BtdtNbUb+Gr646iQ7e4KDp+qCD2yFhpyoPPU4y2KGEXz5N3c1o
Qe7OO60AiT9q4xh9J23RNn1SXC68Bu52/WP3Mt1zG6ArLLrBbiPvsU4JZAkbMshPAFNvo9LpJFJb
X17BJsVE9m8y7EWkGS7VqjFmfDWCsr2De1eOj3exIfmqjoOD7l8T7Hou/8vG1PB/iS6sUFD6dMMN
hvUfWaRCdNexsElW+kIdqlIlXKqOdEycjOl5gd4whMpgUGTNcr3QN6kU3Gb+DmWqbWevEjbaEOgD
7Y606niP0roy99OhPX8wtjNl0JrXoLpvC41QIZ1XAIohBtt71IQGARIFpJnE/wjZAxR2v0XzeCjf
7tdxwPcJVW/CAB0cXVCCOYzZ+QI9R+IfBMIRmy5nVYc+qBFx/sRUm7JDO6vNwoM2kTGWXgWLCDBp
oWWZwh7pT8OZRkUCDGuyDxx98Et4A3hxOb1G0ucekgxu4a4i5BOfi2Sen8mkvGJzBILEM7N4E7mT
F8Q+3AJ0abKLMZHbM09//eOdB3KFhoqBhWZ5a2nm9bZ2DibVXMy44cnN3ToQWZOdW4hNGale/lHi
5l19DaiRnFF0DxirdT0VTUCawSZ7Zk92hTGT4jBnhScHOwEMTg43lPKmPrsbZ5i6DAB+x6TRmktU
vA+7PdpZm/2l5UABbccz2cwlLYj1DMWSg/eJR62MigQfBWV0W8diEJmFBSusaNw3/t/io82jxyYk
OgHcMjSXv3s4rbhev6fYrPS1mhcjEZ7KZNoW5u+uicujnkuqgs4zP8z53C40/lKmClKECNMFVEZn
0eM1MyCq8VsQ0p438mQLxYRnqOmak31rbLgllM6RoCSthr4yi+LZFrQ2qolbYbhsKcYD8caQxCsz
ufDnxowUChvJLkwLxwtfyoglmqwfgm3mNirg7cW4WNndcp5y9b+jHcSn8+mOjaHIV5NGnycstigZ
65KGNghxXXzpTD9SzQvgSCQWG+hLmMsz972cRO3Hn5yn7JDmnb55XvslXOvA2EnhbTTcoebsrIbz
XMz4/KtM1+75HiQ5tHQP6tBs89CR3vw8bxzCPLza51Wfdl44NqeSNhfjAMc3J3jNTzlwdVZWeLkn
SoPVLMffoSBqLr6A4LLjS3YhjREiIcMmgPkdW4svePEDCTmqMCATFFekYU4WGXqENpMQNRU3Ij/9
ZwhtS38h2I/yribc2SU01KfzpmvsfxTH64w0rhSje9e/kyvsw2hLdli6zPuuHTyeo5VNGk9uQK+w
crG2IgITDXM62evl2+WfOiSFSZq+BBQKL0zAXi+NeAuI9sjpmSt/IXhZvECM2XY8dL6NE8Ft+1ha
vZaBf+pp2unnL7aaLoMx5PxzTMUhzWPpDXZ6mEuoU17gPKuvYfuOQphz3GQZkxwn7bGybBFXQOr5
tw3Ayr5c6i9eOC4yOp888IQ/X2psAH80m3pCiXKq84I89a6syG1FQ991e0pHsBX6BcdInI5KMyeU
jFOrEeQYKhqK11aS8+BmEZXBx9gk45udpqL5sNoJu09pBaPWTjr0CYFgolxF7dvGcHKTbb+x00gc
Wgoq/C78cBOH9gH1yfwi2VUXYyvU5aX6neFhkxBRZVSozuGCkiP7DQPr15vY2z8J3HSNEEq0oH/V
gcpry70SsUrp0N1XiRcGOnm1oEcdJbN8EaIWIF+ohboVSx4i7Y9i3dfAAC4jTbJHXQELB94LShiw
dwyjEDPfJMnim6NY7Jw/0zV5Nuw1VRjE0ThBOInZForX5bvyYWUI/51bGS+PQaMitJSQ+Ns0r4EH
2U65yo2FOV3yzrVq63AtGQ6UNXfe3+saD2wqm24crIBzD4fhNvnxKhLgqIcExdEiBHHN4b/Qqhct
DFyXGeT1vFgZZ0JSlwzEi+LqcKFwIokDGlwJYTDbVSqonGDR0PI4PIiO94jEUS+j5kEYn0lZ9/gp
IL/U0R0oDlEVkltHtoVvNP5wFIBlOOyJVwwZ6SM9+WgvoA39GE6Na3jhM2ICyEUKZR4yWCRT1Wv3
9PtbvPX+tBWTxZaS3RQObEoTc0tjB+I1jov2ZzvR/tCbNbMnqGKqsEbQQ1DF8SvJcJyKRv8NVYo7
GX5aKctSJ0Y1jF+0phTUfMv7OQG38PM5/ndfEFaqOvTk5wD2kCOFa8YGWCYZXmzvKeYuXAsHMgOZ
hT+ikIqMI9e9T/jUIbVcAM3R1CV9D1mt5l8pFmuuCYvBaP+wXKvYGiQEpg42mGsX9H2pUN/s76x/
+fxfGSt8qz+zNJxkQdGDSfNtNn/qAxNgMExkOpoOF7TNyYdpivKErtezCJgTNr/aHZ8ZNDklHU/x
ZBCXbBRaWVfIgN3OOaekhAAEhqgbEwxquiUwYtKciKwTN6df4OB0g6HUsKRnEP7KAHu8ItCxWquS
r48R+gxl2qL2gLwHntVMrsloey8dZwRCT3/jhi/ohDidrsMrAMPpMSHKAaKG1zbNbWtOBrNze+gl
mpJhaH7qNAtX6ZqKhxhQLhxwsSUquPZkVrZqVNbNhZIWgfOC3a6iNeyk10LaMZwQ9ROynfwA99lt
yd24GIH7KyBy7Q2AEB/8bE4RD6JJ8D92QqcYMsMMLX+2XsyJzksjYDUxLxyMwVD33npxIwA89aHs
bN+mzG3ZFSwzj2l4WmoywKJaSB51vppdWesRbM+v8VssDz8w22Ftixjys4M5osboEA3emvVjlGpe
dfSiCbJJDLzYshFbACDNPJcH4gvP7FclJHaBMBb/kCUA6xbaeFc3uO1kC3ujg1vPnNQ4H8nAlDoP
aui0dGCXsUCyed5Lwsgj4+36rjWRwP3tw2QjWwRsb8oKWtnempsyvTSe4zfsbDJLiWzmMuN6s2nH
Z5VfjH5SaDMhKj8O73mDr7d4qHZ10IXZ4l8URfFHuac61dkV2ftKbwT9vXLVxjEdpkYniDeCYgOD
GFHdY+VnTWY4elUKQe4AWJj+XQ7Ou9MIUuFxrlE4aPwnZdblt78/xGMVW5zdL14TTJaFUYf6BA9v
oQlVwexr6dhSq1w5FjYmdO43EIuCBSI0UEsvkz/vC/lhv0RxIcHZcpUyGqInL35jZ0Qell5VOTcK
JMIYKd5pwAs0Z72CsWacspvXzNiy878BgMLAv/Vi9uvxyNCBInIJ/hLmY4qyqKlN0tf8R8YDjVef
fyBCilb3scT4L2QAwKThYzyrIw25zT4yvFKNrbiMo9vEGBRDVzuTiYodq1QAPpPhgRIdarrmDajj
D0vQeF6dRMqzvCD7eq/sgN7sPrVCM8gngTsAiL4KjuwLfVDw/R54Gq0jkVE+nky2Y6s0U9VHIZVn
ZR/Ua2a6sc2a6gcjzplj2KLW4ADrOV/yD+gN2U1p5/EK8OLurkf/ZCuxtdy9U2yh+h/ASFueO42g
UV8E4VVbPhn1V3gHF5weas3IReOieVAvxAD7PKOC26qFh01jGspfeHhQXkmzpDnYpaZkvTNL9bPK
Q35zhs9URbq3BGtofGmoE6ayvGdG+89kjTmuPcZsu9AiNKsOM7Yc+iwbWNh4VqqccujYlrZFuTan
X54XxW3syr55LfKP5BbVEUW46jE/Dm8tcU29jOf1cBagYZmXVMZezW6ybFyWltOnnTFPZZrNpsia
X1nnTkC0pqdctykw7JFbRJiAh+Uo8bI0lMH+aRkTE+X+R+0jzQdXqwphdnsfQvUR6EDaqCNu49hy
aouVVN2SZDCPlX+BcX0GPCuhlIjMic12I+lyVyGbM5y+l8r9tDI82VBOesw/v+5/eZdpv7vK82d3
jSiCCECcinNqwv+GlMDsgPTIwwmNgN+AH6ZDV4aq19ryM+w/3LcE17LI4JvaSD8v5FMxfik2LfL4
uB2sTZDLRKbvJsQYf7KP3GPYcnbT1KEfMvgxtIXCz9RMGImcSocvzURksEJ986MyWK2B1k4lLHl/
F5hcAF/PXCo28dKI/2HTtqTu86wpZTnS/3esL8DYdGpWczyhlWXjdIMtyq4FwOG5T0GJAOc/Gc83
BUqBMNVZ1wxd9EjL64QujR1yd64kvPSyI2kIEMLtzhywCHL6QY+9zCwl+COGuhMp+vio1ZiVAOl5
zsp8azp9ed2gX+sg1Dq5AvSf88+NGC+VXKHOCw3RaSOEqaPTTrZe1bbHeP+ktChx/JZwmeayKczE
Fajels8phRQyTARcwKC+Msm3b2oGDSDm+u9xAjPIhhhTzBhm+M7hPI430G8CQEoyQJIFUbh7+7e2
IrIq/8vtqRcuqdm/mfhJDcJo8MNvYwBCsz/o7vzEPhr9Y7oZtRl7cAQSeROlomjDk8KCCg5yFtMi
N5+QludsfQChpz7mJPurGUhiZ+2sy86VJtMnDfc9Dgg5+hffL8aioVn0IaAHbvdTLBlwd6qe4cFJ
Tic7OsHlOWklI2nhvU6Im4Yhij0MyUJCiKfEibpYKTF7o1rw+jUfQpWDz4zWmc6XRmJGidrUlD6H
ojJqJnZHMNQUaeiHP5JIYna7Y87qI0KPWEzJrj1HHIH4ucsL0KfuoA8/T9AHQOkxxHX+/awoO42O
tju9vpqc2gnLRyzk+5l6euwz9szS0/n+IGeSnrhcP+7YTZp4DIEAb9Q1CUIimWyhF9ZAmOnUy7bV
tw0kPk354TBK+gwKDSvd0QBQW+DHP77+J87V8owOb7RmMaDyYaOKRk3tjEU4flVU+pK60A5xuXfm
h2FVfEho5b92GKsgiUrcBbr8Y06RAXAzFBYMb0Qq9vwOnrx88OATjht8RxvXEoSKhNStS2NhLQZB
SHCX1lp8V82eHv5MoG++t063Em90DQEOy1e3lzEzxI3y4EduxJogvdrQSx4xKmrfc0Rj987MDJxd
x7uLk8xeBgkBiwJbaBkkkBT6+A4ZYj4arDAhBvrw0fuN+YYPR3PO85F7DWmlYhOZR6sQmwUqYWVg
IF7khFtE0baBBUK9Do0RhlT4q0FnUcMPlmKTdsBEWci/Pk1gBXTO/Mdz+82Im97F2BJQSl1YJFTV
bztnp4Zl9m1JHxa4qcl/DTz2qpmePkhEJE7kANShkWQvTcl2LNDPmDseaShLhGItp37GgKK3YYBh
SjIVZdE5kZnclTyuiSvJPIVvNz2O95gCfZHv317C1mpogjH9oL46qcOp20LOHEws3d1zcp4Tj1yo
X4IqExsibucUryvZE4+MtjzEqxQ0kzv169yN50hm2QReondUD7SAdzU9hBOUY7F+M6YIf/2ifxSd
0IsXDUz7gIliqFVD5REVwLTb8Q5GiNglvj3BX1WVVfD74g6PtBxvD0gNYUvpYhqxQi342sxzUU/s
Frbm2uKvxyqhMe+JtY4RVxZwwLFY2puBmUqUZIfoXJxRF3e/21dYHK36rz3pr1kttjGpQ6lRSHzD
HWjo9bY6TIY8GRNl6yZW+kY77n/eKX384cskeNFoj26yxRFW17GThJ7lYoojhcwmW3UnuUzHxOZg
B/8P6gcGsbBnvKl1Ciz9vR8uWD4idINxPqV7p0LVbW7iXdOLAQSpqZ3C9gPXIseNdyecXLnUDvdB
5s4HC8mWboWQ2zFbQ+3KriqmUgmYEPLzJYivqMBYA8t9uJ6ssx6zH3xwR4gXwZ84DAcOMalhBy/R
/ux9b854ID4/ZWvfawQDTicWXhJS1n+pjZR6cnQFhrhmptacUzSYbi3g0JBR5BIB5m3VobV9jnyW
JtwD4cL9PProNbMbWV5ydVt37raj+Kk2ap/ZYH3K8zX66xYVJ4M/okQ66xLHkcpN/0+SXvJt3Vwa
He3xtHDJrCjQHk3BwzVPpAvJ0keSVK79mNn4+oREvRM4gVs7v5lIYH99QyDfgwbBBwV3phyRImH8
Uvs7vCFt2a9xRRqLKLFoPG24grF8hOuz3Up9dHJt5z+Luo9TUNQ4kxB1bKj10w7G99jwuO1Uqqo/
gTGyUoegTUgEKh0uqwwaOHzLUmGBunl9Ec+mKxk62M0Y81288emxzQ84ZO323Ul1j7a30CNgG6jd
d/sYplvywaVi/fbdBnvSqml11RrCOQCttkHfOJkZY1XpyFfLLzOuzOik9Il+t5OrPTPxIDLrYAO2
h7M33OlBIS/m6d7tSm+D+sVuRoAY+SCA8mppHC74I8oDG3LCX9sWxSgdt637RaEuAG0IFWbrnwXD
cikZgtazvk7islvixh13+2d7fjBhP2xFCaUrb9SaSC3PASuqRh5KWTpOG45O2ptgNVSOMbY8UaTX
pgQCLdF3WbKitC6n7UkMXlbpCB68uHU9EWQHFAa1tUPJ07Lk/C0AKnH3AQfkmqEwl6JdwUuHn31T
iiZWchmapzb/drewR4iJwWHSgTXjZhAtuoptpB7jSL/av8WqGEcp84e6Tt6FEEC1GJfTSsQa//2l
qbfA+au+WisJbaUWkbJUAGDI07pIoC39xU/fyXTIzxfmSW5W0Qudr//uWTKCdBg+CxKhwjCIJkG6
inP/jAi1aMc7ZymKdSog2WZzOQ5IbGkwods0XU9Yfyq/1rnP7VQBRJ5XDtQT03Y2sw84UyscpmlI
3PX5Y8yI8B5q01UPHJi2u76H3FpgqoA3mj6tNFioMUqtA3hxAH8efK4VFzi38ye8vwNuqh60IIiM
FiKz/ERuHpRJLYN98HHXGmRzliPfm+pcxpl0CdPR3Ml7xIwuYSXFXDUYOGnrn0SifWj83tac+Bi8
Xg9Ab36l83WmAgshaPLKKTDDfZMqyrNsocS/SNZ+bbsBEY5aWDKy00ee3IQGpzHURIWFby8Ne1wK
H7tcPpoWFttf5QNuspc5uxfd/X2GyDa+sXrz6r6ppgOMFKCALBAqm5hDtiKnL18Y44kRnSUrVqPK
uJtv5CwN+Me4qPJjguZVoA4pSH010ShpZpgbTTc8ke5mJLJPL4KHBaZcqVH63kY0rJuXSszhS3KW
HcJDJh2FwpeptqXKSCrf9g/ii5UzNpfDvaazDZ+u22Y3ElpqYdQvdekVqsr8ms8mRHbt6zo4b2YC
ni9xbO1Vqknai0njS+LVQUfm+8IdPoaudIa+CfQAMvsEjk6OxprMph/XUtUcxJXFUrs67L/RfR7b
kLSYlrn8wyP5JpeZ3q6EBuMvyQAbR8gtng+AOyzhZwOr7cu+Ow7tU3tMvbCl6Y8ssZBYTdtMoii0
0xTvVziXdIpBYbAnM4gngK0JmVN/WiECrHS/dSECvaPX8oQVL5wh8DR3/Rg38OhNsKZ+PkyNzJlg
5yt+P9gDzY/EwR3BCzIURIgh+b6NIaItxWGo9P/uRAnqIHQK27+RnaZ7+3XqjLC2fW0dpdCMJJQO
9gbiRUAJzVju+weguJsHAz2w2cIpB3cKGqThP5W9DWUaq4IEiqeJ3d97M3r/ErhVeNP5tmvAC/nJ
PRBUPBvMsMcpq2s+RMiGfEM/y3zi0ZRZVY7o06Jq3AAUBmk8+KNOgcMMp5zU7YWH/0vpYHTaTySU
SDJryhEsLvVGSz2ph01ngI6IYsnCcE2BmCuKPge2LmajiJ5tN4K+USjZ/hNv8iBvQXUDTogdVm42
Dg1s5iw6r18GD7euFL2A+jpMFGwPfgJYE6Vax3KK/JEUXkZxARYrQYoIoqXHrwn2ji/ULFF9dcct
wCuocM9/A0KzJ6eS6dcu4WSnM0FZbngpzMK+0r6RA8HqYiu1tXazqBbe2zd1PRn2Q4ep/oTQlD0D
k8oCl4Dzw4gMx7Rsw1/KOCrr12+M3z7bzkoA2O1zxyu5Cxd29C7TsWmdGWiNygzNgA8ROExATqZj
y7wkzwTfzXZPsbGW3iFJo04PWH+Bqw6sa2oSi1KkaryU/uB3o6VRWlYWc1zI0DL2LBC0rV34L1Ak
1sQQV5NH6dVaCwzT0qt7LT2jqLLbEQju5y7v23Mwacq8ftTi4HXUUojAeiCwh58a0OyazHdwtLPa
bIaR0GwgWIU7esFc8879sr+YoxmcpybKnQaZ90MptvGkw6MoehiaYvUMjyV00dpMXd0+tKqeyLuY
/BCtwvzjZBkkEojaF4VmbJUhX79YspXMJ0jJqr9MjXBV+Oce/bZqXM7SBCIGlZxudsmnxNFAIMAN
J8LAVayyPDnffVtDS6e/ZeLAQSdYo7KTpXQ13vg2MJewzkndjOVA2o4nUPlcwNZaMu/oW6NCzaAd
9l3r4CB2LqlgSxuqkqu4YXkAajxc5WAS2+RMgLvwm/BtuxHMLaBaD83KuGmvAtcSFkXUak4JWqAP
6jlTPCihhndPT0ZR+0SAYl1/8/R1goqGkD/NcJ1vm2V0SB6HlCyqDwWDBUK+6LyPyNyrxpnC91D0
a/1jFjN42pjobBsUVWGelvupw82Pcjc0qz14Ikzpa4KrzTC10tRrhRorYkyYAB++EYnBu9LVJMIt
obDYm7Zgph/bvUv+VftqcJRdCT3oyM0SsaXliaSbwFHzS+Yrhxd15DLSQOyKYeJbM0Ge79DssgSB
toHybdDkhSplTzEPPigUmdrNhI5lY1EGNrL6jJ82Yh15OJ45h9TlX6qbWEjCwSO6UhH90mg9be1z
NGefa3Fmext+W9utOXPiy2Jf2PL3AGVTw8ryE1s5BkMn9hiZ3+AvNNugXsaPqDw6IU2OkfDTooBX
vProCO9ILSMIFNV1e8zmFn5d6wp0OZpXUGEqLn9hTA49bYIJgBv7xGQ9OE1+Gk0V5ArKw16rmi4N
clspaMLPXb59p44VAhJQj3t98JIThqZiRhL+QEFzniNgE8jVrdPpQ9pbS2phmAAnw6RcexnXDnr/
R8SgUAAl4OSfcl2fzm7md6j+BPte7cjR61yzep4+jcwIxzgTtXU207RBg5ZxSYDcUlKHpEdmmxuB
QuTb9oO0QfjwJTo098FBhTy6IfIdynWtU1cP7+xw6eHb+SEfLnpCdbLYitnwDfTDsZNQwXARpYzF
a0aEevBR5y1npVbegMriDVPzU5S54s+TAUaC5bYFjoDrbaSbZSz/UWDUfJ5jly2Q1vJ8+YTGQUny
q8/XpigQZ7IObWKd/2PkO8rJW92TVuFG1E4CHRFsqaGmSO9WZrD1igmov2tqngKYjQKmNeGapD2s
ufPhQZrYsMFlqzsdtV9WwVxdbh5/imlpH6dbLSUMf6jJkIThIc41h71is50sUoMmKZf+yhmY4+1Y
9l6L8uHzOx6IFCZwqOUQqMAJIPsvRQ8r9QOqH6ewugCvm4+R0FSxe3UEwcB1On34ZxU14Ol63b08
pTpIidZwc9LFmjToM/AkXwP/ganxSDGiZ0HVFuR4wvnjQYrLgzMZw8a8Zg/ipSwVeql/T61TB/yQ
qIRH4GBH/Bk8FoB6WWtZtB6Y9ZhDK/HW8ULsul2kh5wkJJaB7MsIaSSoKQdxqD7zp0wnR7pZhPEW
553qi5UiH8vaFh4IX4e30ECRBL/Yj4M1oKsibPq0bDo+InxEkmYza8lEJP13MusEfmXqEQj3e3hM
09CIfHr9thfyEMEiodim24lpLYvvIxgt0Wdesrvb2Eh/TInVe+9eGlkfhP0avKqzyUti+mkGITsC
OkoW1JAFG/Y/u4ICREcn/lYbR/6A1nWFsu6cFfmjP/llS2GhI9c4rYQxbBL/aY86xSoYm+k6SIQc
ArQ/hmmT28LTBF+UUh9i5R8KROX0+xnLXF3u0xXS5Dce9S6O2KqXaRuHorHYU3k47PCD0eWt3RYF
SGhysB04eR7u+DifSrANbqVdrD6hXZL2vCHeVaFCch+tHbT+n43KIyKrIsHbs7h2LLcqR/dcEOvu
vEA/GmmFMpNcRONv1EVXkRKh4oF6j3EfZvJoqb6GGQu35i+S/tXO2nG5kiuHaqaashlqSdykOu4D
4KToWwRbjPOtgCdXBwfT2iLsXlZ7YcuPbXgS1Plj6DG9n+o7A4jonwobe30c6+n2bsFIs0tMjs+E
2ybJrtRZbsctGnVKyftyP6VjDO2J2/CTyU2o7qW5oI8g/IsclTRIkc2OFCrdeIJL4PW2R+Fks0v6
Mebi+POzrCdgAgys1819U2b3v/I4c8z18zHn3ZZ+/YonEPn2XdGW99dvohc6YoR9m1um3cZU5LWM
MdRErXekGEqUU3sl3Cc6S+LYu9t6VRkItY1Rn/NJrtcOhwiUa4oEfLMYOcmEWGsl5HNcAFTRG+sZ
0pee+AwhD+RhavrtegPeeOCFrLL4AS3mo3wqeXZh03r9SKX/2dK59GO6cUFu+yJcroIhKvTZojfi
jW5rqq0BN+uT4HhYfVGGoQkBVbWrTR/63PM3DcH6q0Cwpy9mH7mbC+Tn19fQ9rZuoFCRgJccFwBU
+7efqqKxnQY8wgiRDkWR3Z3lpPgUG8ontD+gus9lELcuEXrj5Uv+dDQRjip5JjApIhMOO29D/axK
w6fkAaEbjDL3RPOjCRjy1xf5V4iOQU+yOy96ArWbX4DPcK1huTg/9mLsE8ML4lt1rnol2uCDFzda
xdNT32RfEkqgHUSUEscZEVTWZbCWcdvDFG87Akmr4Tlsgv9stsw1U8z7NTenoJAkxIV+W8RAK1SQ
9yL7qIWtqy/thZ7hfukO0p5kKAZ64rWH+lH6bLMt7prW81N7kXNPAjG6CScdletfxGfGWlQQ9k1Y
z39pu+t9gRl4P1GYuGz+uziFFaytdMu0QQRGPcXCmIuFt9EyFsA/SFgKE3TIUWvmGRVI7QjIYVfr
5K3hxk7vMS+WyA1xzcJxhN9/yn9CoLwcvm6DPbuhU0gN0gLmhgCfFLBzxflXG0rFYm7FEZHDrE21
gYO2dwqP9dAKCPk//rOMtWibKy416w4Gqcqw+izyb9qt2BqElhn+du9SuCFbOg7PKscZvT9NEppR
Ced2P0+ZmRy6CggeLZpmArsNGyVaBQa0/gOuyPJwWpMWUQMQZUz5lPzMrEP7RFgF99RJOeD4CMBZ
cSRyh2bGCjC6uR+SRTXbuttsf13JpPnnGMDAlSwMujIXVXv9fT/wO3LAlHHF6aSjdzYvPtSluwFG
seMculwmHItiItDYq6KcktB8K45Adot9Rb2t4eeYiAHPRYxH6SfxritbHvL64pJ5d/nXyMDpzv+c
FECR4il+b3ax6uRjigBCZyOT55AQ3xtEv8LQWsqmE8+qLOwGOk9TO8NcUm/2C/sv4S1s3GrHayfa
1GJMXOhP1nL7Cf5dOuueAVFndEXljfTu+JkjxRGYtDDTCzKci3lqAf14oSvNjvxVQCoB3e3kEm92
Fa0qLgUWXt2VMTcwZtQtQXCWriDZ45rYuicFnew02qLWNBfpz/bT7zElzFNro9pcb4jIkXze7unZ
7D3U2GUmLtzReu1T9JkQJ56xGIg5nwSKv7mWW0iDLSVjcUgxhz0/8J3eVssE2Pzib131kEL0kgv5
/vx+EOy8BTpDgJ7PYunXhf9tETteFShp6ZZpAFNUdTP07a3FjuWAzamz9oiD/hpycRIvnsQEf1xj
R4PIzvRBgTSYjt4rRJ5Za0sP+bc6S6nI3H6eGLk2dAdGoe6bhKxHrhzDRT1PeAmohExrP23rkC7W
1/3aFuxpV4RE8fCP18xxFFmxBjaNNJ0C4/JX2X3MCi+dLxZhYOsWjt5IvwnriVosqhAQ0EoTT12I
FXWQRcdeHiTPkblIHFNkZhNfI8fgWEZSMPU6ffs3i5/KazKMYfVeiaCxI2+kkEXGidU7Y46Qf5tE
oEW4MannqcTKf2IGpPc2arHx4o0jgXIO4Nmp3OD9lYNmtpBs/G+2ovLvSU3b4EulomiPYlnDiuc7
nvkrNdA9NGMWMvb0eyy9VsvggRdkQBmcmVmrQMr9N6OVyZ8O+/5QUCcI6HXyr8nxmVMz/b/qOYB0
BxuHgjBSsJwavJZBqR2iq+6b5bXYGfGPfsFa6chRIYsXXA99Y7G8oa8kvrsExxIell63wFz0fH0I
yyotCLvM52AAVHZuTJaUX/pYxcAzNmuJeLLVC7ALViKDSsWky8t6IAjI8tapOlAMXxNiabuNVCRb
CaCtnsk5w69Bxo4AWvFmodCyVdxFVFoDv1/cMYQ+8N2dp+R77LmiEUYMh9+8oqgFKdxIJs/mbb3v
qAX4pDia/YUeUX9IFv8EVFzik5ba/4qsUzRmLvCv1vI3BjX7j7iffgIpcl8L9YrkGvOUVSqy9ZgH
wSvQCBZZeQlUyfoVhGc/fULX8bNJG6LjFv3PlNQ/56X0f+LFuGn/nhdYqbo8GxkckhfpgN/pw8Pj
q7D87pVCqe7+ruxkvxob2Kr9nWDxgPnyMp/jK5e9lTzKVQnFdWT8R5GNFLnyvnogUZJXLsSIC+BN
zQOXZjenaeeRCMNsf07iACs4DuWpIxZZZQ8Ir6O6mh11j4JOg4poCy8C5Ak5HDAQQmd35Y5xsOoZ
EGe3LuxS77CbTvWfEiCJQLnUfjuLMsjQJNQBkB/bCcFjpBB5BMVpOo+J1JLBvKtxosEthy1ANhYn
CzH52BzTuYLMe2IcyH1EUEqxxnqY0pMW37+ImiJAZVkt6c1bpPqLBrrUYNtZ1MnxtCKOGs/WvQ4/
wHTyC5HIJUPSvw9o1BG8DS1MEsidmNz3Jnk4WP28WeboIrTnJBPOVN/nKVw7AwvWFcLFBhqVFeBR
DuVWEUxgWkFeqyTEUFZaFHFXXUL1tHHIZKCeFemB0yOhJp/pF5iKNMjRw39fhbl3Gac9dUIcV2Hk
dujJpscs3LeZ6VgL0DBTQmgPOH/q1DBc2VLkEGhvkb2QohDsHjB6ezkW1vimwJ4EVgQOJXNhKtQ2
ND5zGhcf16Cav0TkcFCBN3AavpDQMiw3KMioZG5Wr4QCAlcf5MrDUARMH8Zcz80GXHjkAnCcB3Bz
MZW3rkYpb4+UYaTTPsDzek/diMe0XUeQOV9xuv5XOCYUSLI4+aniZhnV5f7wBBNLRSEzOZOmQy3u
BDWv5iGIOXHF0pCGhJgIFR2zEBpUXcqf21QTxIKQXREU2SgQSaROeXd1VrzdmHFYd3anaF/Kfjb2
s8DL4AM3oEjl4NmIrPTRh34IcxA6YY98W5gpEHTiuT1xSAxHZ6T2m2LbETgRcWWTjE3rYZpkZOJy
A3/7S4/ZsUMs4/pPQUIpKPBdMNELIUNpsQkgOlVNZZi3/WW78uQhr+UzJgv3IogFprS8mImKg4tN
3Gm16G/9+xGD1YKF3hnmdtJHmjGzdeiS1IOARsPMve0fWt8qCjArsKkGhG+yFmrLIotSPvLwMy01
SvXKXkUQwQvi5s/pozLfDxuc4hxycsPEe/RrPL6+D9h0Z2iQ45Z3NdLWszs6+pgcCFAn2oHXOSot
BKjxtFtEd/xDOVxEZxHbbspKdkRWe1J1vfwja6VUgDr9kSYL3XsaAS+JSwWpE6W7NFXcyPCoqQPK
o7OuzQ3VqDV7eWIUFej8zq6Y2bvwXd6YKa7UmASEnZJ58utRGUAlyPDaCcd0iyvY5MmrXCk3dkjl
/NyElD1d3uSgWgXZe3qffNFqunA/pYNE47Pb9RJd2yt8t4/LYdrk82gK5uRN54cVcFBSSBk8ij7K
zn/+L2Nq9JhyLfxZ0uaxMNgGbONUn9/NunK3teDC2i3FjLSeAJFkV2JYPm17dTe44Vym4phZvcup
M6jM3Dqf4Ah1gm+BWCMg5DKqtEfElqmSQn9YtFBhNkPjl93PzTvrSL1szFYQPfNvfwNzAxUGRHnf
9qyAW8RhTVKkQ+Y/mB1o6ydWGziKFDG2tDXnOqzHstf4Kwji0Spsixd5arSgk5o2ZkRogJXQE0uY
42pLN7fpNRJ8YD12nUf+IO4nJEUSHf1ZI9AvR0BrtY9q8f0rJ/VZK26t+mR4p2BUW7qEd5PrqF/A
PZfXZhD/Q9FIs4VMu9Pg7el92gnZWnGTqH0+6eSkNzGmDSo0WbNQETG4uq3fLimT+O9Lp31Z7t13
gZafyDosChHqp4AgVWdYd+4Uswq4H60DRQ0h/KwWbIk9j3IsQ9nPZQKwfOEyA5PYPAO1hCF0cFbV
I3V2cAmHUMJuBlbtPIYDdirLqnbBNyumT5cDTavB4QS4QdZWmTcaA7KLXsYDZQOL/KT4aZDYLxtR
7o601HMV6zBbGTq7W+Hdmf13153dPeTERbM7jg9SgHNoAxxQ1n+5XPgO4AENHSsZXHjV7V6ZgdAQ
3UNCMCnLV4whnGn+BjXhffjGKBoNW8LiUlvlkR62v5kwrpLG4P++ISGCDFSnSOQZg/LdWrRORGOS
iNqX3hWACQu0Srpv8gttJZZpwmUVUN/JW6F9HZD9CWOUxTzml/7A6cYE3DFoVcmIrIf4Uk7HpHFh
DTuxBA/9GLa9q/usLi+b1EosYKOY6PnFyb9TFTHVEaSEkxPdznohdpSwZkMWAsIphj9CXIfPthM5
GE7CBjpv5aDWpxKZpE86e8pbJR6WUJPWJ957WP0brhydgY78TS1DnumDpCXW0lMffdjj1ndWFWbG
HpQNkeqEyUxa6E/KryGWIVQxtWEF1PLxF7C+DpNt2ibtzXCQnvuJ1reglebDp5YtpPYVh83jrbHv
Y/KSc2pq3BL24bbLpj2sJU69GUI6d1zWxTD+xBsUgH7UqDldQKn+w6Cwd6rSWq7O7IcYonNVaZc2
QXYNewz66qp3nQsxGeh5taVgW3sMqA/SpNW1yHcS7Zz9xC0ZP5hwByK4Vfwiz8zonk4p4VCQlecI
8jPFBCjMZKrG4Oxh3xi/1ZtYJOJl44ZUAJbtO+gDjqtzR8pyVfyH6lVyXLiRDpPoxh55DJoHhJ5H
hUyyvub21AaPAYyAdaw7s53mfvutLyfe+sHyJHEtRDIN0ZNWRd+veJ7qS8U1ktW4xz1XWy7qX1i8
1uMxUBXtXrOIhsAwhehAGXEcDJmwz7J0WP1Ru8DFc0zp9Yxi9NXkjCg5ohX5QuDAFhuO04M97Wxr
uf8iXTDOPxT1dY4sIx53ka1IAneygWIoSx7gAobxZOn1z0lSkvJKvS2lBNrfzx75T0GJs1wBCjWC
2pCjjm1QU8RzNFZVYiKscV8aEscTpRXnirc02w27bx7o7fJkzwTY2EFGCwvBYQ3BoMBBCH2YWraa
F/j/HtPfI4UpWA7Zbnp/J7ov2SsGbjC9ujUj4FriJV7wvF6nMNYZeSvEooHjWrd+H8/WajxZVQAF
NQ0Uxwh/GaaazdSPkSe1ZVHp+K8F3Ae+H8Vmf8JoX3mSeqaGFlWKYLeFMNREwbu6KuA7DISgR1/N
ky85sLFMViB6Mu7c6vMz+VJV1fe9E8hvy3fU+NIdQA/646dh6hlGeNA2nT/AA9kW9WlbgZZTvJIc
lwS/hGVmaBKRTwp6MsD1HO1u6/qEfX0nRyhgUuc0tBJBfeQTJPovj4hMG9qvv63P0+aYTPvtP3Tm
MnZPGDyjFNIvuL//NhasfGEkqisHcKvm3g1Nl+L/we2GRs01iltj7vqjzc+KnsE3ug0i6R8Wfunk
4KqHJpwRdjUJRMZDrFvLPqwYQLYVfozSVgHmJIFZTBVbav03984I7oBwHCTp0UBQZmZk7P2ajCrD
UgiIYNDZkJz/VLILBsPIDED9/IJIpAVUduovhexjks/XMCr/fyy6kFcjeaYoVyk6wuxBWboYEFkO
iPHTpZYRPogz8/dlGIkUlXnAbA0Jv6SeZxdL/PmOGOFDOwWpkP2Ya9XcW4wpLGVXYRAW5eR+vFUL
+i9fKBP4OspvAUcOjzK3kyy6+no8tPiglzRnruNCppvJ2XAYkxUVUNgiIhxyoxUSNLAu5cKIE3U0
+YE0gZz3OIh+AZE1534a0sr3pv3zkKgXmJnPDI2NtSRTaY1aEg58BRpQU6PfF9YFUiexPqk2yKgw
+Eju7FFgW/QoKIILCiWdFQEr6iEUg75ZHkVLKG/a90WR53sH7FX3Fc3/V+deG4C9SfFsekRDzMkP
EGn+IY1hAjJFN5PKjBnkrrTf0V1iSWDsv9PRUvDmrQONy5xU0ki/Hdas+137g+sVymVEMxE9381J
TWXIrj3bjV18ImAW35pvcE+laxB8EBlm2IU7HT666yqPsfcU6bIAVTrBRyfqxkBGXlq7WOiYdS1z
X8KPOD52rVupqF6r6Ni4CQihE+4WvX+mG05EcvIO+1cXufEsdoeKKq9kDATh0m3zZVEuzxiEuJuX
xSdp1NvFKx7Jxd5QjB8zGgD8HzQb3MQkty66f7MYAlhu/Wd7sY81e0eGxj5pR6f9P4pyemI6Ixa0
RPq4CXyUOT3DiWF0tKyo2+ieFpqE/IAy52lRI4qclMJb1KopyQdbqkFgM8MJGjDwIfv/hBazRWZY
U/S6mOMVsAO/+rYMGsZbnKu5iZa1xPUYulVL09RQeCBonJjMsM988JSwOZeDDHTPWUgEE84K9IJh
FEKkCoqDzriUEIRrWYIND/a88AQUUy7gybbXtB3QEEC0JEtcpTw4acIfey0jTXmKF2j+j154aYg+
+cSzIijKiF00MZ1mCU4tJ0NwUIflxogNVmKH8dR19zunGaSETosPosf1HyeiCzWpc/a7ebcCl4KX
LHH08ix9QZRw3e6WH6VKJyIeVh5I/F0QFj2y4msZnF96Z8B/6uRhKU7xSu0c6mrnlThlcTFZWDcn
663qejptsLVmYR2pqKZ/wW/ScHO5g95BKJXdJTlBHpeOpsJ1hz7EwgphJC2/yh+gEBnXMPvxDWnc
cc4xYw9C39JtPTO0Tr9eIdKwh8Nu89sENsrya1cU5cEG85oBqtY7qSEi1i8YHLNk+j6sN32JMxYz
atvC3uRObmvz5xDRLi59AJ96VLU+ishdKfPf55q+TGryKdkK8feMEPQfra+Y3lRRqVN7ySvG5588
zDPqTt11rJEU1DVTUUMuPuTzbHUad1vTbxvIggyuiP6/F7N4fDmQaABMnvDSg2B5kJt224YJeHqV
t5V01v/moSWynyKugGkqHRpjGhGd2FcwYC7pyJJZ+EwDEsD1Cdtkc3ahLFkS/DezO4pX7HvreLpl
ys+sScFoxLThxGG4nOv8GJNpX/YnW0EObqg2XdetjGM1yDs+5cvclhH3KcOxBJan8FwV4QdWfcZn
MMNahr2lsw8uKND+FImeGUXlJEtQAcBzmqN2Cg13UdAzq4HSd/yIgU3Wo4VZAk7hzEoe5sm0VYbt
Cyt+6s/o7cu4gWUQCB3xXr2T8yK/j0zl4Rya8VXoixHShYLxU2fUxos6ZozcYdDnDOwSLhiOlkW7
DhbDMzavFe5L6tu6ykxTrbXleqpscpan7Gzoo0DA2VmRufUzw60RVlcyIL6e8Byb/3I5oBg5HeTL
e3siqv2+M5a9P8k+ZreIlmZ23LdBGoAeGHzM8q/tQjOe8Lt5KInb44a0UbcBsiM4+KocElrMfbXB
FpZYE9M+ncoeHLArh/GkesRBGA/M2imN6DLAK459MfyTFEPU9dR2zB6+cqHtAtoYxkmoGpWh3nqE
feWipCBv4Kz2vY3evkLl0p2+162bSsWNdAQx8SSAJ9lAQ0UDptb5v/rVC7C+RXmc1S9ESci3kB1U
1xzPWHgcEQe1CR5E3mCSKLAD821ywMbiQ4mw+VIog3y5G6d9Xnq8m1zdwxke3V6ivzs1b7G2WuyM
RNiEHozJ2TPhCmqOZoP7Lg9BfV/WHx+Fibz32vF32cNlh8EhikS9hxOS5bVVqg6Ge626JTdBo787
O+3TTwGbcKI8Izh5Yz7MxgcUljwVRNvCvG6V3uxrCPBGgPPpRKlcg7oKQj1LIaIRO8TkXJeYKYQA
9pAt82as8RFvLPMYbbttPk41rS+R+9+p+YmAdIcQektQGSVSFqg23lHMUNymnANd7jYVVswrcQRa
HnsV54hd+5hT+ugbJGr3Jsr2QMw/qMkiNOexuDJZ3cpE1veh7TP5TcKpncivnDHLyACTvkif5ibH
NJohzkiRoPNxtj4Z+jRAStUJNuEPHXUN6/agmaoxuw28mE6IUrARINPOxc76B6IZm3NaNLEVXK4L
1NZrNulbi3MbsaH+l4VDBYMTd/vIDFl94i/skY8xEouZyzK8PqQa+WBBdzbd22dVIodN6SEdowxV
nblbOLyhUtI48cTaEjtdFm5wybewBaFfrJL7JD6HCLSV6EpKS08H/LTKC7sAIAMXYknzUuec11c9
ZHeDK0JpYdoc21tSd0pBIb5sE5FNcMDVnLEOuD020oQ+Wo21Jn7l+BOFAVayRavYbBLaAzNw9cSy
j6LkQal6WPddFWC2ns/QnkoKoOy+sDgpUvgRs/b8YIbcjzb7oCa9XCtM8bfjYIs/T2OQ3yyhRwRP
5uCMr9pyfrLaVYG7lRlqicVzYyKzvI+PJRIgtKtIVHzLa3LFKbQg57Sxb346/mtUnDZtJHJ9yzgO
wkgnhu1UZubOMxWSkh1lrjIapIj6lkksZlmo9RZWU7aXvufBi6kh6uiw4wxiEB+Adyx07NjN5qkI
Cm46a2JHw+kQKP63WmJp7gDvE5RI8E0GTzPJo7B6bDFEQUenr95HBcnGPp7liE/sr/9WUtcUZ+9R
eBgqYz6U494bY8r8qYEvziwZ2WBB9Z1LNYEhE/QeEuatTwUJDo62mK0ALqEuZkQqCDKY017RNh4G
AEzDA3PH3g/r6tcXuHUW4gC8Q2P9OPCkskbenK8X4gn/Nu9Dz6h59NfrIEOJebL/OmM3fwR1uHA4
Gq0HCf8d+Zd5Xofclm1UdjBYKr69t/hrQ8hBvEUTH/A0qi+mfNU0EkA6AHJVTDS9I8AG5biY0rpk
rhnGQ9IWsNOf3T5AGNLFw3yBTN13jwTvs2UlZG+MExeu8tN2JBKeAlHbqrt66maVQlna1CJ6cFeP
biu6kQxE1wD2MEUhzz8L0+2QIc6eDmav1RFEpZib43+ln6feqjI2kKvRV7x22aYtomDEtSEIHE8o
D5DlqlqGxAa7x7MSDRDvgoQVnaWzMT5WUIxDF2jPmKmYCNMySuCiy2Ybjax7MGvVrnNtzDV6hsFI
ec8ebzlFQfb14W7K+SjERR7M3A9zJnJjH1UqnIAN7SYE0SbL2u1QFIMrLscW5w1PcaDxYFX5ihTh
0CgxEYELz1O4vaA9/B8IMavbP3HI8meimnbTOfbvE66Un9bOZb2a/pzxJuyZfgwpOeK/hoIUoJrg
6s1G4t1KfXkRaxH9suJcHshi8lmowr5sNmrZT9yZtJPutQvYdAzj0ge3DOSYkFa8iRdjeSDO67gU
UQbiCrFjd/lWfwV9wlEyYB6ZbSdFBFItpNLJOte/BlE9xk+U7YqOW8Ldsp0eeGZgaeIegcjVhQ1u
kbxwSQMSGBLJalBAlJGnk2pQHdxbpjKFV938FSAcciWWRMWR+s1kgBvX/uiHQGvDir/TEIVs68kG
opCNir9ZHT8qWXEokbniO4hTog9PKo7bPq65fGvhjSSKAoXeKbDQejhIfSEpIPzsaqDph4hyoGnA
mI5lS5bW3VXQ9jKpaqk6teqwoejehUIjRgRqYYMIuqDhqbZ6gWTaeH4iaE5TnPGCHd5ZVRh4eGaL
Wz3aVxHG95mUCFCAfvGKACrOMj4AaCmQUP7ONLZdxMSmZfAOUFgiaAfSDQSq5CFZRLJVcUSjz7LG
XwM1HrJ2xoKIReElB2YH//361PvCoXNZ228O5GOj3V5lr6ThYmmc3fYcQRd/XDuaxUkBZROHwOos
PemzWoEE3CxIP6RyoCpCSUE4q+nyBhKOGo2mhuepJTwZjWV+M/iKafhMSIfChTMXwTqiX4dbhsp2
3V/F+K03z0Z+5TQcE4E4avduWnvzVUga+WMNvAH6/fGJeh2TP2hurqrTrB9+eFnk0/9i1Gcr7/6r
TyUNd+YEZrEEfISTxZfkZFLUoV7hX3XAGreeqATVpm9EvFa9g4KLe18LqQ+GGnIl1Q1lNVHSwc1H
TpSVSk11LQVUGdvETBcRGnSuF0AfRiyM93Mr+Qdfdn6TxoSdXFxq+CClTeEIhT0pw12SMCY2VfNV
nsXpLt+FL9bvbX8i4pTEhsuycTmdZtcjBwTP+6PMLjjzdDCLhmsnjZL4HOUp4Esi+IYf3UXmvqyB
FafQDXqHCXCf+ntAlivkezsP9YWk7W7tbGoLRyiUMlzaUws6vL7/IIevZ+cBcvnqDuB/hs/8ma3e
l71IW6QKRoqpk2VnahVCIDkbJLqJ8Htvy8NnbSKGP12rauJNluI/LTUjWcaHo0ckQvzOVqyGJ2pN
oVi0TpF5aCdloaAEdBZHChRE55OhbR2tVtxhaJGWb5IhcY5JT2AECY0OMcR/o94EgYhPJsr0PcVW
wbuxZMjrzMzxmcdo0QieeJGM5aEthnNPjuBNhGKJ9q8S8bv8VbKXZqjEHFtYdVaxLtWKaHG4uVkL
Fs2ipULiyrBsD/X+pbddzSajgt7aFueu2vtf9gQTrHe2yQDjbVRIWeNq38W47JYoHqYkv8IlYg9A
XbyO9pMqMutF2Etnpv+HCpV451D2NHC4lkLRSBZWwbFeiO/LeRJ2MspkT8LvMBOefDj91Ha3EKnU
QBmzXNsF/Qpi4+26ND78wdGnBXec8n907OwWdhmTGGA/OFnaAbuDmMfv9JcwG2atvVJYZrJW8Aq0
wMx5mnts/kjUrmK7KyZHdWbm+AMwCzBnfgMQojqTQ33COlIm+JgLjxfcNipDmxkQwalyQi46VAT8
54Lh7y5/QmMJenwy4007L1VSUllzkK6Guvuv/dFpwQi9lTXoLlB5TBj53CKOf6InXBH7HEp3bf7j
cUP4LHuImgdr395IODlDUcU4lDg/lIPlr9ySW9Z60Br42iGwquVmbDMJhaFNGjjPxYKiD+GYh99o
JzFehd+I8QPY534mXDNrGvECylkOYnzWu2MB64x0A5/e5BLJNsj5m/qYZeC4iN1XmIFrV1R1D3Uj
avtx4zhMfZamQq8EF//w9nHPcSr3jPZwogWVaEi3QKFsjeJ2yLCcZaLehrGMI+4gky8GcZirbnVc
8GZzPYFYrgowmnn1jRowg1Cx7XNSNfq1liCuRd3tNE+I/yKZp9ObsnbC4oLaM0Umzdj5phZ2OPAm
FbqLapxNaY0kXVuFVGSJQFVDpy43dlb1HDmAbiZXzY9JCXYzgrJxGm499tmg9SjKnstPzNzwAxJc
5xBQoBsC9tQ+vytI37JG/TY67MW0B6HDzG54f8+QEeqdj4gHIClLdmYNeEs8J8bHKzfojdTQegsI
veIpxRSXjYMAoxb9kpUJz/FB4vRTmKiIMedox1hah3UYFhlemAsFDHYZ/hloOrR2KbRWwauolpxn
YCyA+wxxjAAUN2+wDAx2v+j7byafbxGazlTJQQFAY2/ZAtzYS2aoYf/G4efsT4kdDm3Md/R6kUIN
ujxJd27ps021jDfBp0/bIywNtklbl2vBYTB3g0AUoRPHcgh0pC76VxKQmARDHhWbvix2zK4jEuz6
+kyHKk1nUzejOx1KG/ODsk9xn2psUbZGTTA8TNO7pebpo88PiW5o1ghOkpEqFsqkoZ2bLC/5DPhn
IHUrRQEVgXCfUtVe75QEH5rdlHuzRSrBjGjT3Rv/Mgg02dBxP2vFlkhPqZUH+PRSeYhxB4rnGlVe
slpfLmkiC7/dl9g49W2aMGSfI8HUaTg/FZ2prnCWuCG/Nx9HwC/h8Pr+0roGQ5Wijh9Z9Ob7lmVr
FvFCA0qN0ty+3ziUlQ394+9MTuCsFZOj+znOkISLpc7JShHTrkmxW8ca9fGKANTZs5WojNu183qj
4a3m06ts3dct1Uaxgq12xi+m3Y1z+xPXIG7Gubb0eXetaRBe7g1dxRxLihj5CsCzkwAHIcEatsR7
cCN/4Q+DWplqY8n5y2TqEbmldueLe7XbLVOtKudimqq1hNgkLnrPKO8zh80VYjx332OKwJXn7D1o
HY/XXPS7vSJkJ6QqhXMZ3I8XiZJwiVurtmNG8i+o03Ci7ij28AkgycZlvho2SSYkLAvCh9dyHcLP
mD0MacaquKD7h4NpFahAGDc203TKQBDsbIRAaHOLV7yLAXKNbxnD6NGrnsQ1Om/0EIiIk4vzaV/L
aZo22nkEeYmRJkHFEKMntlEmjDd4SomlNlc47ok/LOXr1IOLtqUanMc3GWDSMVX4BxeV/km+xJw5
u1WUJJLPy6wADXqEjP17idABESFqxcnyMSpHYGrpKBVmMU0ptLkw/5cm5L8iwEcChRJ5IODIdY5g
/H+SlIOkflMtkvbYITokpgopBnjImZLgDdik0xkTSKqQOtObUpqVFxl5WxlTnISAgnAvKB5SphIs
DeufvaKCcSrUTclZLNjqrf6PctsI8oF+Hcm2mtI4gv9I7lOBfVLRvL0vXxHmQ64ctcvnkwLCmogj
1qyW0R/YmRU11Cb+6RXYaC7WaZ6VXRbhPD0uJ8w0eDqJWGcfbtHh9OhWoO4xeJJFxt5btdxkyq3j
yhR6520sgkP07/7AzAKV16QwzELFmTDHo/Kj3ZsEUc8LM/CZxCnwaY5bTat8Tq6dCuXHYX2QyJoS
O3h6DybVOeizM4JYtdLnvdwLw3eT0lO86rZ3MZJYeSeI+m5ZOJLLOXDknLpCv6txcxTcOnSi/jb/
133K3QEXdQmCirX8WQJMOpkugyKqAzQOdIC7Rpsc3bB++aqqddQeQMtacrqZshd3JKpp9BcxQdpr
lw3/KjAKfQpFFBbqqjThSEPTwb6hUwBc/lPQ3FviuSOrbnNs69Biux2Rq++lK6qg0ryLrzQ8gb2y
2c0ySbCa9cR2yKemJNIX7BbaygI6wycQl+NpvPKy+yBd0XkS0S9YHZPAlRAmDr/OwvFC2Tp9vOwP
2t5mxEd6MFqgyx2gWqx3/zEq7F2LOv80mxnj2Uq9k3IYzudtF4tz1DVb0yi7fJnIqCBN7dHS3Vhd
+YuheWubj7UNDoD5Ecb24lUUhMKElEVp1Y6id8oHKtgW0a71AvobcpmNxaDdiOFxjRbMIJ3W7lZp
GR7I3Rx5/ZHMgtrDIdefGF2InZNXIMqticMARc+mZ3p2DOnDvlb4OA7UTnj4Uouym0ujVOi1+zgh
untCokTMQkO8qn72b0FMGL728azwkfqrtxbfOEK/Z4mLRZter0Y1DIujzZWql/NezraI/brNJZW9
ydwWmtrWn/WbvKWgBhPrIUXlG11t+E32MUtxI4mU0m7EkBdtKA0RhAKIjiutfe6cb0gmAmwEZnvj
l4d5Z0vsc336io5Vyt/E/QGZjfYrTjZJZxjYg4E4TlGjcd6LClZTrICj0V1DEYgls5SBiJ7MHC/Y
uG0tuLCVjXWvMWSyB6Ud57gIbxaGqQlJNh7JRRXKDx4FoUUY0cz8xLtewRqps9e8yO8NWbQrOAzP
a7qmq2KV920mmWFjTG506oMnwfbm5T69KS/Wo7vMoL1Qcr78FVGUaZn0hYEsDJ2fVmSIWOTgisH8
pLpiL5pbarIEdrBsisc0wnRqXTkpCN3vU2tJ2iUm+6I+TT4zrp0n3wOU0TwbDjUl9GPYQfAE3eQD
bOe4/k7VLX2x/dRhKSCFCwjV7nyzJ77cWMZBJ6u3gFZvts/mMLU+VDqUs8Fw+kY8JB6G3nxxjzWc
fJPjCM7H3dlqoXTXMDMT+tFk7+Vcue6xvuhfzauLMbnqCvg3s9NzfXpS4hYHYe8JI2eu0zGCzslE
1Z1gVbS1E0cKKT509KX+tNWHcTagYDuztvKWOf7iCoOmazm5KIE0Vj7PZQMwZFk8YKuy1rzfuEfC
fr33jUk5jN3zOPta9TKLPCZWo8VlbOzY44YoeY/codH0eGBmz7INKOLRr2IHi/8AdoR5gj3UWrF7
gwlO72jfq+VEXgskQ5DnjBgmgLDlKAcF6tFHTXC/WiXiP5QIum90o0KXZSxURjpGANbLHhlCjTT9
rZKWEVaybLyy+oK8+97Lo3X/mJoKZCiul3ADfQXWTBgEsiImr1F3TJbUpsqsl85XE/7Bj5XLcPBs
f9iqKBHuXawF8e6jKf+WNeg8wCThAdcEkh20Rk2XZfcBX6rdtTUXxWoBSc69JfmDdCJKn83mDSHO
7MYwkw7ZeFcGyqOTXuOviO/0aFoucbRy3JlvQwRRP9EoHAPOyrgHE4xAs6z6HuvXW/WPnlT0svu5
Mh6z9QNk3vILGyzoFWjvVOuKV0E2FJh4R+RsYuHbpF3b5mR09jr+twBkOrGI8/fFvT3Ucris6Y25
lPbCA5Tuv7DUrCtqgal+M3upPTQQM6u/Hbb+ZqLaImHKGPb2QcAD6bI7yz33Ee8jtU3VXpxezjkt
qtIJNFBp/a9gg1C1BvOnyvZqTwes7vAv1jOSarksJYayNTqO+4Jw/X74xFqBI74GzNKOAbRHjKmT
ax78gPno5n1xEDK7YIKO1Vpt/LfheVDJNsw4t76J+JA2oXvx0CYg9rFISPGkZFb7NiXlCNQ1lA80
jxfEWHaZIIz/9w+SIbogeeFI6IaObuENILVttjpc7Lg0/CboAGc3V8jY0bNksFC83X6pbuGcR3nq
Yy2nWBQdHS8NxJtmt5lOWTO/QyIPGT1BpIvfXmNPMWza+cWMNFZ57yRo17+RNamjHLgcI8yk5wVn
szcIWZ1BIk6GO8sS86ov6Pwh8urxtYE/1yQpEWCOGuDxcbEP00NVEAN1DcJ0gi6dJGUAisCNhjrg
z3uVMi04W/3hR+EF8ez/qECUKcY0FW9mEdS1JQWe4ztKkDdq07wV8Lbb/EbfLx63mhYU+gPGZfGS
j+RsCBs3YNMwiADEcHzfhUVzLbXVj+cqkBeQrj6sNnh/dwPBeX+YZJprmnbgdmg0uCeMjXpR7cl/
Blf/yT8khWNW1pbZ1xaPwiJwFME/Qn3JOz6OmUWzKDrVlZ/lRqCvDuVIQkiGiwe8Xet0K3hNPHNK
N6wAWLvr73rEJ/3ZwbwGjKw9m/s388Lei4NNo6PQOet320PIOJtyO6OUitvUFapPWgttorYkTl7J
s5Ihq9DT5qYaItXR/nz8XqiEL80iKoNVU/dE2FdgFPXb08xMnDQR7VjihDWoOk5vbidp92LYdrv3
2qHyg4EqDvORlszytOGLj2UrE1eY3j94RMa1t2/G2IPlARSCe83M+2DD2R6ylLPlv/21u2NX/iI3
xsKihXo0Pi7hQ5KdLA207blD7XsVxW9sde4dOkvpxnxmq5AEoUDQsVsNfNzsmuYoXRNsU8UpFs7o
ToGSe9tbqavV04Sg+V3a4mkcmL8G+vGtOME9pAjphWnORJoKCSqqW/OBnCNxgZL2Lo03gI5vRQie
NU8JI+IO3NNTzHrQh3z5PCZL7iEAdWqyfj3fMkapdXMvzn8PA0MqiXFO3h353nlMqwcki/q0h3H4
sbUKS64w8dwAnF5yv+9IrO8ma5BAf9fTLXwN+DEbI+wqSIBw4FqzfBhDmuEa5/uk6i7iWWa/ImvV
IONFYMngpOTA/Nl6M0NYoOHoizHzwsUKtTAO4PaOmQUhW6l//DQVb9Ab79MmfBYUtnK0Wan0sZvb
aJUDc/muiby/a/Ni3V6wctfHyAtL31k2iAg6DVHa6Nt1+4p6k6tcUlwqShS6wjMThTAxoMKRKvKh
wxaUbpEsBicQeTYZegutlbij2x51iH3vTVZvsPGhGqh7uVLLYsB7xQcb+vK5+X1Yxl5j4m3IvU3d
FVQ0Uw3mjKKapsdJG9E0iY5R2HRyIPseU4hPpqUCtG8vZnnG9rP9q1Xnfq5rYVweHRDnKOUJSUYo
bGCV+lIO9awkw4/N9vDb3WntH4pUPVkAKDj1Kw/cOCeynp3NxkycRFQzB6d7/VVJpWwx96uW9rJp
TNYxKmWskAqn2OGvI7hBrH0Y5WqjljupXPVAm3cjxmaRmgPpOMdZYEIxLZ4b5EyTGfaF1aLRGYF4
9QpX5nXduDBo1MR8db5X3QldgWEC220m5VWFVxWtr2S/lFxv1QKl3nf0ZXseJ+qUQiKDyr1eea7P
HNXPH3hJIALFLWSMB9IM7+4BG66spyvucvGR1U1v7f79VAJPjyRQHAtzzQGGv9BGtUxtQuww7j1J
S7djq6NbeI01kbrjKjuHb0FomQgJri67377B25Gl6X7UWHf6zv+amHwLTlRzH7kTDAI0pqxFwrMt
wEdfxEUmbqofhSFxBZgsuul1qKt2aNDEUI4kJEEA9Nw9pLs6DpqcvRFbDHrDdWzDbLYVPf9fzoSr
UJ54vPqPXy1rjIR+fPtTmlOLs081JG86859RJ4qTS7Kxooq5INN6T3fuQbqwn2YJrPx8sDeJJFaJ
i/CZc0YPj9pzamxfwRP7hFC8e/Pd/Ip8KsG0Ck056QzhzkM8YQgd6F7c6VuNc+AGkTSxcKJuZsHD
dpZR7I5eSrRkVMAa/On1ijGEreF38mK7QANu70aCjATmZyDFGXEbfn+ZrDDp2D6HA/xmaBZTvLCe
qFAMKj7r4S4ZSiAdlV/PJYn4bJkwQBI3W5bBOoiHjMk1JZIgtuoGsEClgcGfI2bItAVorWL0pGjz
Qm2PKjsKzflPy5VfQmF0I5xm5eDXO7M+aI/G0NaJZxJsapuyoZtbyYoSYRfAm5O1h0E971X/oCa/
h5QTFv/zrix37X1hWL6ILtLVju2r79Lfwu4L+x2Ew0VwqXGekCnAP0UsjYSDMXQVfVmNWcCbUjfA
guHqf2gPh8zLt0n7WXVKpp3WkuYxDDEqBkQjSoxiJQnz0jP3tvq0HBRI9ZtmDtB3kI/2XWpq9Hl/
rsFVZjESYZYzrRRXXG2JHO+oRFE1JYq74CyOZf2lrF2qQyKBaQCHiDouZrHtJqh2pz5JczbByb7x
ClP1UeZaBgb2M52ntFesTFOAnnbEBDWT2Gbi/y9S3UgxJbjYac2q0ZnprJo0oIh3DBuEhJHaFm3P
vTX9rX3csmp3xkvTxUMnbWI8j04DoPxxq0Gn9BxKqU7z8sDE4O9bprFg65P5Pd7D145xZvEDlVDL
pAenfC+mk3Ost2VDP5FpQBk4HCqBgyHdMUCZk7sDfJ4+etS1/0ApolKMISaik5kdFPotuD5XEeEz
ciUFz9IWzbqQzl1fIc2vwERCVD4lthyOgX6clFv6yL/zDMJjMbIws7ymoeNpd6iZVYOIzlKdAqLj
Lv3u1JrJUa7lnEj0H96G1m9pu7MnHlLO4vvHQgYzQRrPJU/BmJuXjG8j2vNrs0IG7+Pr7injghSQ
9cLxmGQpBj0UhU4bgOIa93lP8W0AxJ3rmyKPnYCYHqo/0fEDnW8pLGX2w8QtVjyF208dhZlhiJXw
MoCeccj3JIInm2YH0ELs3TE3LHt+GPOt+eDjYleWmDclEzX823yyi4UCxGeryFn6n8iuBJ1xM8D7
51g3Jm4lGFvF705TzGKqrQXijFak5QFYLC72E9O4NT5bsyMjO2O22HM8/bCjSsdSl4gvSn+W4uF9
/e27TXjld6WRjtlQqcEgwxRXdSBqLBe9kzhzLBe/ww3/P5v/ma8CE7J3sfsGC44M56JH3agU2tNN
MRbre/3PDg3o+EnSZexdDkNlybUrZ73wBgN3NM6hd6IkKpjaI3et2IUI+Iq0+09NC4km1NyJ6UJK
57PyvoMaGIugu2bYYkIMS9o1SMig320rZeieqhDWVksheQ30Pq18450av4MxS80V+EYjdpkKxkTH
mBJXKNhZgyIPR3z5CBtU0Q01HLZ5bCllCbuv8CQy2utcJIyHHgZPnaafaHi7EFsenkuS82oJ6cLl
B3T7GJGs/Nj+PcUifobbhERz+O1QT3jKBEdM3nFtqMuFY3onIpODG/F+vCrT6wixSvkW+y1+kiN2
3MIzv/sj8Hp+lySIk17umQrOZ0uy5zM+hPB6oodd8lTsw/WnLlO3Kw7MkiGhANat5vXmMe/CU2fB
b3XmXCEumrCzKpaAVJYZWe36ItG2hY+9nKBzaElG2gNL6Cp9s+NoMFWVU3tiLGG4QiJrtt6iWwUy
OJ/ovZ1XxNYO3JTt9BVWIbiZJr6nCZdFFANYYUsW8QEs1/bj4FnChvo8o5X1ua8inytmPmoI2uVb
suwMxtAhKcTSCYpYvxwIxH5btiARlvr3wk2Ms44zidZBph5Z+NlGlUEfXimfruLECCj0bhjvAfqj
O0tBFLlAJrZ5JG0pgMHzLgZMV1IxDIDvaNXKs43hBKaYDhDYh4Dbn5tSFWJ3IKo0YyTU9elIls36
R0C2lWYmzgdZtwFYbLvBp1PMFBGkgsAQQp9GWryMj/dcNCS/i0ZGainpj52P8ENv2kOwPuG6lVTT
nkIZ40urcKSt6SDz8vuH7+aeIYU2XiNp3vBpZbn0Liw8gXLrHUO9v6UEQRRKEtgR5nspTUUbUDO3
eapU6oXWc4ktHnBFDgA/IdIyylpXHZyLWb6w2UHtBVlZuqvOUwS4JMKcoIi3zPgewM/X731KNIJH
cnRi6K0zNijP0inlK0OdL4mRwiDknGnwDzVyLGyyKHrek/qlnYfb/lcVXORU0uEKbffA8E+Tqjsa
egAcLGqDtKIyh+aJ1W0neQlrCCjwlfWC/fl7nNIbmYwBOUxx1FeNCoAWjDnIOyBllJgsTTLAMtSI
FVMkt2aVLTPIEiF1AvgUJFJeyn1RCfUYPzYgA6hV1rY57JDALD5mJoLyhSOacRws5k55ziD0eHK+
ptDN4JXen8zHZxH07XimQEJKqMfh+zlFcW0g9EgjGYumf7Ap3eS1LZ3ES4pw8fxXsmliCSqN7spi
BAXuA4zxCvA6JDaymBixg2zIbAxguQRpMN8KM09ISxkFrTYWmR79E6ukMl1VQmLTYp9zH9OXfttV
840bjP7XePPmTv/jV3xVlm7wQZwlGR4pO6aIJd9MqJMajE5WYXr1ywBg9hWcWS8tOo6/gsW6oqd3
O0q5VFDE70p3JOZgtmtSngpTOJtyW9ghcxusdM9Xgo8hq/UdPZWpNDgl+W2jJcijFqmmMMa9hNG1
rlWx4Zj3QmU7ajIm9dn0oqOBNC5GUc76TAoKn04/pivQ96Zfi2kVegg7Mr6T2NIMgf+C/TLz6EnX
k2Ti7stXnn2aul4qghSYvoBK8rWLLWYHhvPSCNP5ex6DwS1Jz+Pae6/MSOJdkMuyJjTXibZZgX4Z
YeM4qWOwO/AObluf5rRHQDAQJy2K1c19Ayc6rmNufjZBg64GWIe1DVL/+mn/5ItCLhfYXGHLobl8
1OnMPAJ9noeepIZquEpsGybiXkzfSKRArwp8Tk+YKaeh98O20Bfqo8Vg/FKZ0ep8Jyx5Lfr8+KoI
+5vniRru9d5XZGUUHaDPPXgJvBo2NOUyWbgwoRwdGCRWZDwCdnzJ8VcFw7QrFn3Kk/xePxNxM0NC
WZDZ3SWJIJtEjwef4PG4Ci0LjK4p7kGCMID+Vnc9Y8wh+Ua/rzWRHPEy98GkalX4jFzd83aNj6wa
kQoKoO1i40Q8nbt3s9ifzMKwC6g4xdxY60DBB2dKwGjHq00yYEpI0o/PIK6mzYKoID2iSCsJCWGu
g1S3SLAcMQF6KMAL2q8ENa2BLBS5wyQxt/h88D0LqICBeHD8MyyXm/CAJS2iknG84wb8ApuNMnKP
mFPecPswaJKJOD9gQ+XyXWb5XPao3YaG6d7K/riWLaxioS7lSkq0aknojE8afwoMp1aMvA/Ku4qN
gcg+QDlZZFuYX3fAtylm8ZciReAvQ92CWf5mVmLm3LUkR5MW3BIL17jFg/HhZwtOyVuHk4aCg1UW
ppgSneCZsMqrEaiKU+i6SqKUXzIgEcTDBettdk5SpS+mhCBdnHsx5YGFXS3+xwe058najyepD9LH
i7TBeoyMvNdikzRXHy9jWXcWjuLzPBfMvC10ZaPrCi+qyudRzTq5zeIpf6+e8pLIfib9MjQcCk4y
/YqS/bAPJzIWI9nD1JeaRmvjGMJ160tw47FBdoYKBbTHhGnaIFr74OkLJtoATXkjrcWDKyFI5iKs
UhimC07gsjmSqwu0LMuB1nTsxtlEtYRDbHjikkiKqNBDPHNlgO8FKbeSRtmzZ2Xsx/G9yeJ1SmNS
JEcGKymvZqcqy16aynfmxS2b0jpx0vmPHbf4H85ALYIgfyXUtv/BH6WnHqaT19cli4QMhibgtIhY
4kGetddApYe/0TSU5bZgPGD/E5U5mu8fFN7SESqRh9ngEOSav8oRVqDBELPLlWWX/fURvy6NobzY
a88YHQlhM0CzctT2aAr4Oaf5SIg080tZ7huBce2ktu1C6HxS0CGUGIF5t2AwJCNKw0GfAeZV2XRZ
24sxgcxQ/FC18uucVmU3UmrCBVvmX9IwhIH2sDpN9WpD7pOHMBBV7o1Q5b0lkgUAztNYyRD+pKTL
sly4fOrqn4FMgo1kDBiKnArHu/iMj9bXli8s1D+aXb47s8+jullVfE6eF0+7ssvHoV9KOepQRh/d
yuNxq0jDqZ/4yY0jFj/EswoqfmewJlp3fCw66C28kdMcmiFI7o9JgyzQ5nN90E69cJKahO53gvH2
1sRgF3aAuar5mI5FAA4pk5P2NTafQTV9mtpKi09rrc1G2mqYomkgiEAd0XwbtPOND2552LZeGggm
mqEv9x2IIJraSUluE0rIVjqZNnHh12G5XoFcDFT7qnCPoIlbnFpLAIwuWPDOkLjbRmstrRyPN1/m
PKFekAr9i018cMMLSrT5ajAs5c71CNc69VqqeaxRB2wyooguQaOrIY4rkiZ0lSXnm9adQFg41bPe
LaYrEtynCsybnWMSd/UZimpbKgKstGsHPm+107D/s+OzRqZT91T1FsUtWfeu/IfEmpbr45WXD+kO
bZH0lrHn5gsvGyXMFXyYlf/GHixp0PQ5GBkDU11rX4fo2ueKR4a7BC6yHDD6yvAFUQ61yi8VWs6e
98u7EPK8LMzex3ZdE96b2U7PdgKZlm6jPpiX/lduEE8OE3phDSY7E/h70ng6G1FWK5y9BgbyV247
9K7LsHW3o589k8RFuRFyIRe3mrSQ9hAxZ4GtHpMqgtuSdtLD3nzEMyG0sceLFjbGuDks0pZ4eZjm
zyjl1hCtnlheQ+9HAK913fo1/G8t1R6VTPdtMWKQYdP+z/t3aQiYgY2cEOUCdOVADBqA6MheL+SR
u5k3iimE1W9+9vwbNLtsZ0nFuntmdeN/+wvXb9ENblhSArRvRKo2GebU1joSg2JVXZSP4q98hhfg
Mybz/WVtSYZKg9zhFzupjH/x2Iq5roTvwruE5kdhuvgWeo8a5ywlP2/MyWGlfHcFSeiEhpwQO0hj
RPIkoDf5Ffa11RA0ir/frGjwdYRvRxpeSBZDa9kAyHyj4wV9fCckpo+tayhGuQPc4mhJ6eb8hmbg
hwrFHr3NRiUINaYWxRhRSNuYu/7zJNArmPNzAhumLORPnVpwGOYFNbhEwpkCXSSlkJAqxqdUZXCz
nlKpUHjDPhp/4XfLc2JFGXNMrnO8Q6JFYJf6wm1y1TQjeAgc2ddLbUfI+Zbe1Px4UmvedDUGJFTl
+JVauXPaxUeVq41Xf100vqTwjm8IQPjJHWvXWWuuSE95VDAjanJhrSai2xxCeJTd6PZxf+SLJDn2
JfK0IrnLFzXZYD/lHksAHSMhrul8FqiZyRCVgKO9iJD16B3Ot3msGmnsT7eXCjxwhGxxMPC2CVFa
VDsNSj9UldtfKSExMX+16QTrYvDw4CGDUZsir3PLprb9NjeiZXYVFwcqIld6JhFdiG7nV4gncL0j
WAU0io5lnyukHVDQRCXp6aKJWewSW5u7Zd7olkMeTroUCkt37SPyJPTryleIEHyw8L2DyRN430JG
lgMSGaz9QKFn+oFTqpzDQckxvAwCfVpW/1QYa5et8NMmkhDJUu8xjABSV3PIWnL1qcGPkWhNahxx
k7XSUz+ehTsOj6TTEG7YcbYRSVtOfTb2XH4PVbWsdcm+2suNK6fZTdhsJFxU9hGHRIlKlhpRo+Ul
7IGCyFtTJdjbRXyVMN9bYGQ3lBy1xx55vJ1kSlEXyQDW7KQqmXrmaiDt3ONqFmHaHcsqOi9RHQ9F
R6ZW87mnZ2A5jNN1s5WiJf/fM3I7dTawA0M4QMtEjZYBiUcQHw2OZxJ9UgAOzBDsu0JYTu3VwNhE
tjon3rbP+zdwS4niEQYYEM34y2hoTtTKLcRwVxlAeZzg2TyU9KuPAj0Qu5yqO/bMaM3mUXmvAibq
AQIy7JOxduv55cYlKlu28Qfr8EIJJUUFc/QjtnQVREcsp5FK93lVfndpDUWuprh2KZ/Kmz+wRGEA
VM6FtXOnqUQ4t6GrngGp5Vn4Wr4QLIu6Y3lYe5RXMArxpjoPmW2A+FMRfnD1hmkLeM7rVCARKOLM
VFCJ9f16dRlh7GsWUj89+OrBGe5MLRevfQBuS7fAUq4aF5TzoTibgQm9+3GlS7Loi2BmsgGNZLon
mbcvn6M1XZnDyKS7X7PSE4OIHfGZgB4yngEgtHq73GF1I9Z1NYq+EfCs8swhklaGK/2AdoRVjsUi
xvk4C891Vi+KC8vTUG6OEMIRaLZgFUi6V4sGdtvYkOzc+sZ1AiAKxob8mjFjeJCRhFZ5gx9O5v+u
6zcyPwC77J3aBk5yPpkGsw7AMhKbCoabp/oMDlS65/zlSHZiSaa1wmmly+aEoN3Pt4ekvatcVSNL
2CUDpiNHYzKMVMzNrVtz6t1Vwhlf5FX2jWAgsoGYa/7jMjv/YdagBTF2Oc0G6Tbd3g36b0URCoqW
7nEpQ5DFRfn3ikbIvv6QPvjU9vZlKWEhrYOGLlZVjN+lfHUo/dSF33PDgfecOd7d10/r+3U8aX2y
gys25Gc4PF6zAERZMgnl3H334QxprAY3zSc4d0BzEpqrydkQFILAMVLc7uBO56clDOz2nZsImPei
siA0PAFiO0YIVd7Vwe0aZmT3g1ZInIDIrucamn4hIZWF+8fzJGOhGbg37F9ak6lloqKoohb1I0eC
qLYJiHYoHeTW8SjNLEngIW2+LC8CzIsPZBTau5N1FUTgCmsuokjqpsxzaURYbbW7Ti6HSEK7UVJX
cMmNjceOfN8dQYxYSaKVlVmDW3N37F5sQh3fjb4hnWoFmehjpQ9H6jD6m0+pua+rHFPIuHG2BB2o
l7Boj9moHlLo8E6BhWEeh5U0rEprLcE/dDlKQswqYsLwGRbDYjByJHokdKMknlPICR/6jn+KrfY+
uY4ZatA3f5A+GUyrsN2TLSvrB6U4R+69Dl3VQrgmZ8+o7JPv0CE56Z2eHarmR0JvGMzA6LIDZgy4
ZST+bAksoQEc3PxgokFWG4artgK7cZy7TMgEab7039efcDnUpKJoFwDdwrmJCzvucoP/8leqlX7Y
P7bvNr2SdYd21OW0OJmpOuLtT5NKrw+2Xn1m7YLgWE/gK/R53q0sEPB/RU22l3i+Hkvn1gDuORFj
8kCHmCPZ8SWpIp+ewOee+XBrhFg5F9C3+hyVhxerCkmBCxqasnvTbGVyUUH7RzeNr8m9QkcQYsfe
kK2h2587qowo2yJy75AhbN11HODcZUDkxvJF/rYC1burd7OAW3kIWUZJGXVuUOTS3ZcGzD/C5P97
3dZSAW3XzYG8rQV8JCnFmlEj+ufPX624hKTKr+zo/0u6KBHe/AFd2SfRVKyZErEDA9etwCjRzwI7
dmq7JV0wqQ9IaZBNAo/OQq8yIpSC1NNVE6cXw5EwAzW8mf84KM+KQCqwrK5VbnJEOe0suHegNGHt
on8p6eKYHmtsIGqYkzEyvQ3hyHqcvvhSsg9ILVB4MSbX0BvNrFVoBcohblCBpbiGITjHtECc9Qcx
0LnlU/EBtqvgUK72YMc5JBAngCv6g6pFLd2n6BuZBY/F9BzbQXN5k/TI1D1COncd6l/j9dv8ILov
TVsnsJV9jS/b258wchB/kK8L4/U6kB9LdogYfMtZW0p+yijyytnEhpadAlLTUn5wT16XVr8CsPct
Eyim3M2GAV/t2KOfA2Aewm2WU0rIVRNOEBXSfNZm5vw1RZ5o2gx75H5qZqb2jjVbI7DhRdiZJ7Rz
1wtyrBuagae68IkfCCMDjbxfrbmbVkp+vSZNKfPhG14jJkYeTPp4hBIUScDBixZg6dBbVk4ZmLMH
qfnYVTXMbS9BBjE+Q5PMhCZ9jq0/fLHY7FoYh8sdOdIffLs93VaVnDkB/ssNRMIfst68KoV2lxaZ
5wVcT3ganFnGwKyWLdpopgoQfY0ghTyEhCHx0msDfngnuYuiP6RFuAPlDO5OmjXd9hXR6Ic9J0n4
XEKzfj80ZksIVjIVUbgZUlSDlSzddwccJJqhZ9KIarSdjrPXR06rZ4JXF8VdYPymexCLRomYzEhJ
6Y5umKYAFnpmfJuge/6FQZQn6VcXZ1QphoKzl2DhsxBNL+A4x9hTgYtcfGFiUoL3s7JMra3Hn2V4
Xh1poYFbQjVc8KWUzlyWzsl+tMrEFSXTyoH+hQUjklkjV84/UXD7EJGR/5o7k2douaUldjnvaszm
RPCMNG9IngXSAjozWocCDCayY8IwVg0H9MHhLOO4ZaaBvIU+qeW5Vf5Oxe91UkjNxFToZPxf0wpj
kBlg/7djAN0HzQjD3EPq/ONfMVG/8rmZcjez1fM6gjVdID3DWmHXvuyFhc1D1ZrqpenPhRURn/9S
MEyuJxXy3IM6xSl1KX+TCFzKBj/Lq7vGsmOzzVW94A7tbHswH+m7qTTbpz6+EMnU9q6I5WxRLqSv
LLu1pQmtAxyhtPcuo6+DJG07NrdPKrbwMqGm1niJcT5hKAqy8yfgk/nDmnVTkFEDyIdgRHgKotd1
yB37XRiZrYbVHA6MtPQ94bcpJI90SJKr01IO2mouQlrQZfVQv2/AHcvt1F6TwCDd2BVH5bVIcVPg
MpwkhKbc9q9oRDmIXANZjYQ800R988FihxO2EcsCTQ7KfGC/PFu1EqYxWC6k8TL1l/PRwI8U8cMK
Ku4U8ZBblI/Xw9Uoh/8mKoM8+2sA4yI0Qb6GLs/H2KnZ/gAzcxk8dvAhG+EHDFTGScQhaopqOg1E
UadjkuDdqQBoqdgybz29P/z/0MF0Sm/o18VsfCxnHJMWeOSY/K+8AsfXE61JyYcCQ8+GzM3qe3jp
IpMijaXtyxMhrBjgoj2qoBGf5jTS/y50SZ1Csu7h2uGfC6viT3ezr5MrymX1210HMkkKwJ2pM1WI
j0Q0mjWHDxMvDg5jbxVbK4UJ7dLjuayPK/ubLX26Eae3urPu8OXgENHBZejwwsTZO2Zzd+Jmilcq
bhisC6PAPTVT5KgUiwHKfR+AfbsnRgBjoN8yfOtuG3NKNl8CalIzlbXci+82Scx3jtCGPic4Gb5K
qWwKmn3gncGNq0gIA71/v2THONkUGktMJlsglvs2YPZSOjaQslGSQdCZLgQaE30WBQutYtyyZlkZ
6+diaxkmqMk5lVsMjl4RxaBlYd6y7/iQ0xtpYCAEq2laArB8LU+ehRhkYlXBqDaygLgIiqwE+c2T
1lW9oHUPzbG4LXIWo3WQV2clVzZH3ErBhNGH/00Dsk/FPVehK2A0d03HxEfpgFpqyFtiRh2siAYe
TNOH0yX2/8QDlMh1cuu/FpjOOgllfsr7mnzBuEZ4lZlU/aEjGPS5uX2GTH921uOUfaR677lYvRkz
nDN+Jfy4FkIvUAnPXjoPwVFfQmK8E4iXPyhArMV19B/RANYaKQEz7Zskz36J+deXdH8pueQ41Kif
aQo4TQHKuYksrmdZwY0zSM+U6gzzY3R++ZoeDLyR0/Or7csOraTNx4IF/UVPyr6IU4jCKMpVqFNL
HCgYFlsON1/gVzq0VUH1ICbsvmFWKhAJpoxGDGjfY2MVKBYx6WX+/V4nB32zwKeNLlLsYjXqqmbU
cwDfGC3tdEu4aQtf1kHEFinN5qpgTUlWOUWF6LYNVT0iH4az77CpYkyUbBaGaBvxbwOqAZetXPtO
fTEz9r2jUC1FbIaeFx+4GLREfHma4eMD1QifWjeTmCTkX9Ie78MGB3gATFcs2snzTVy2DbxB5E3z
5nTUT6RDLJdOivBbiGh8eRLNwz4lORGV1LT/Jtj3dDKz0LKKH4GiOFNQjBCsUpOxTkeU79dqo4CC
wpxthmCexWPZJ1Jrzsm1HszFHHaozsfetG9rvSbE0LY78sbi4bnfaXt/7eT9a/XmD5DVG1DBtNGI
xt5VlgbEtJV3357jBRMQTiNpcyP2dQRQMcFfroiVOCnTC2+BXaLOHOIJmyP6R2jgi0UqTlPLnZGc
yHodEiTfcVCFKAGKboIp/GlhnbyOV4EhqrQp6KoF5I7xVWSx9jrv7haV5rlsSQuaJrL6i6CvL9Y+
7SaKK4kbnENdvYqGYLM+PZhzg+ofU3C/9vBV9wEU8WUaTJo/r4B45vcoZrcR5WdkrX7Ipt9TI2Os
NV9hIabTvmrE+E0DFJ0yVh3asVRJCll14xcw9gwMP+6JcMg81yxxjGWakeJdFOnBjJNk5ul6zlZw
bcJOltFOlqb4VkyAVYCX0X7yeZy7KyRI4Wv3gOsuC705hC7H8n8Mc/IMgImc5+vtfJ3eAYTIqx0c
sUb2PPgG6Wp17+WnCkVukMNTCK0VUynur1fdCXFcOQNB+PDBa9lq+WRsDVjKKHQr4g9wL5Q68c6u
hSFf4Z5KkX5YN3BhPMFOaD8B7VVp2l/KM98z7OBbpezS9Tmd77VDwbOQqtd5LwCT9JIgBPAEkzHy
NToxRCEnPhxuBJ0SUk4XEQVZYJWh8Otzl5xL5yUqkS4R+kccl7Di93YSM8CaYZhIGhUBro0fm9ro
unxcV2jIpe5mNuEBnSyuWhAs1wn/8XQxKVNSqxuGRSx9OvOhJLfHfOLl2Bt9/EL5YRrkhO7kmKIF
XImaZNWcIvU8tdPAAmGh69JRSO2TMNaeQHbwqk3WqwWgm4ViFbJJidaGfWDRiMvlMQh9ILxqW3xF
0N1u4s7RqvJccqGZXz3m1C/XKF1ts7+iwIiUKFNxxYW+pfym+B3DMCTR63FNibvoEm5/1TqvWRkL
nIdRzxO/NURWKybeOY5z4Z4X5n6a70WSC0Vq9F+tnU8IngfhY+JMiPN/GEncMiIXQVihVkC+cntJ
12x/eouU5TrTHGGiXvT+q+j6LqUHhHEYXtc8Ehjk47W8PCBwq+ARC7L/crFE7K8uKIl7X0FTEQFL
fbs2fHCrAfe5H9v9f3jWNgeyRbfIRN5+VnI2rF5hEhmKbZgyxl/BbxbtdkGQzJR2SUz3huuvbL8i
mDJHW5JKrR2PsrGCSMaaGlI790czbGaE77lFAAKRWahaL9VY/2ARH7RKoDOoclQBVrQ9E2I5sQV9
6sVcGsHmv6nJlObSkuzLPeeti48zA1+S3ffqF/vGYnOqstrdIPH/1o3DSut6qiYu8vDwC8VHIe+2
ypBuxQZtesTmpqsRWwlZJlBLLe612WMKSvAemtxO2NR0Bc1FJJwHhfltMrvxzRQW9NFR4qJpeD8G
OtYoQwhaK3J/nMntIebydd9XgKexcU8b5UAHPYhKJhTtuZkt/P7/wqKrPJJJ/hv0RkBnFstXtF4k
jrwlq9gq5OUjbLOVvbRzbjYNFnQfgxV+W/+juDb86ZKtLS/naIVMNW4Rs1jgCI2EpENJXyjMPLGR
4B/e9HG3oFVT5wn1BMuHEre1QTUPWMh/6XNMMgX1bJtC3q+Zw0sO1k0x4P7OF3MVzkbu1FYXqBJg
lFWoAAnoymBAUAJooODWTjPI0CLfFIdCXaraLoqtuyS2x85SoIMSC1sn1tjgaeFh9npXBb6VmkSe
075iOK8n70MDi+om6buhkgMlc5OrT8+1xI7n4RPBXzIXwjyURwbOxbHnko4a6LV/nIRy1OUVzzJi
1uioTE0b1DHURa5oi9WcmTLozGzFvfnyH7UN5+TksokmMgr3ZagTremQP978f9/u+XS4f3eqigdZ
7R7gEkryg1kRo+oddtxHekdf5APpo8jepgyJdU5goAUGp80ahAXotDXPVsy19MdofH0PYYzucIN/
RsQaLTX6hFa6VJy+3kd+ekqXB04CCnxnKq2E/eP69TS+hb2bX4GC+QiaCyXGQVtPUyhbQb3iHKCE
Drgmx2r8zfspFj9Woo+Zf5u297myzWGnD1A8rVQEvJKEQIC2/TceH7jUhZ5LS7nN9AyTjBeS4gyQ
4YdRcqEs+3gKV1zbISGDkgf4gTNWmMQ5IHjvYq3773capnczGWndrZ8VYoPXWpHL7CXGlrQd6/j4
aTpf/5WJlHcSJXj8Gai92L2EOPKWCBS8RgU1RyuchFAdYMM5VdyKzZAu4z6xqsPU+FT01LUczil9
//iXPQ6ILSUQm+7+FADR9X6E6oo4pdjwI/s5KeDq7h4iOwwSad49BveQmBJm5tiOtnPhK7p5D9Hn
SaBVKgMGdGxtlWML6NOm5Iq+cnH8FtMwpH9v2PlYawvmbhuFbYx789r5hPoTezSQgSVz9j8NZYev
baerudyiXlqp4OXjbOwTenr4fai7f69AK4wJ6OgfrAHG6Qj/Bs6PZFcCrP0VMJb+eWypcDArXnrp
1k//l7RUJqYZCNYqn4vK/kAK3BIyGy/RmUKIFaiRrnv4g8nvKLu6ora5GbJ7o3zApTaUkwMNwkNs
wft9MGARCEGHZ6ho8oEZb8XFUbjsDLgKPZdPgtJQX2Rji63i+d8WcsR1oYVC5wxmLKhBDtFssiff
Tqdolo7i1MmH2Pkv/k6xTK9gjKm8nnknbLf6IOz+Sw6JxhB4zCjE8faLmdLullm03fxobjoYDZLV
mj//qkLMr2T7/TNzZA9ddA+GYCxVKfp4RR1RGAweKSP6V+tacCQb3goB3bLZwygRCf7gz0oAjYHP
+Io6rkuGP+DW2tcmqqOJSXPLpkR4WE5xZjwiovVGfx6zVbrVhABQ5jxbLaPsw0y5fSv2QEtyOknj
eBLR4pKo+eHZR70mMT3kzCPfzLvnIMGv/CdQ2CGIC5FpNetdq7MK20CfI7hChh0S7UBAJ4i5cFI9
P2imZpKOvaoKaDkj+16QdGRl94/UltUixC0tSs+fuU4sjyowcBoci5Vjshym0dlwg1I+M33/zXRf
ZnQWQQBPKUTHailXcg1T0UpbD9z7b/CJleqMtTO1A33iXMIPkR7Q/lOghx+7nt5gJrtAxU3WIM5q
dnpLQnUkbzC2ZaGrEkfHl5UIy3Kl+Q3AXG6M+HeujO/iRxmSXqEd6v5QcgJz/EGSpa5J5xzrNGjQ
Tkl6ptSjmsHpbZcaUie8N1fQq48F9Px0bxhBlJDnOELyE32mpqW04h5swATO84VErtMvXJdV4Un6
ygWKXM3BXZXNClGG0aJalC72HIRtMggjeiEy5Bfw3/OzMx7KPmb1EqdgJp46t8WOAX4vmVHqfaz6
ABJOXWjpnTn+8mf+sopY4Jgs04P7Bo+tfTqP6vaToeSLON4alJBpcgHAydI0+6/AfMoQCfS5TFAU
aIF95dmTWu4xW9Na3PkIx7Cb4Ey45TQSfakj6xb1Lu/fJME3jqHrUBFSyH/SIgG0DcLuO464vWXt
GSVI9XJ7AaY5UaN+LxcEw+DCeR3yL9n6dvJgRQ3xlKOobBglzczYb7TLcacsW+ARPdBSisMSAhX8
nrO9eGMwCqzTIBUe3rV2spmbnA63bo0q27OJYDFiu9JqzrUIt4Uop97HmLR6k0ZLz73gRATsQcHM
RhyQ+mIhrOSLcDgkpOuOJEs5vDrIjCfrwiwNFVzvmI62MmhehOvtEMvKc/QQZ68hZgMrm9QGF9O3
ZDXUFcPzcm4/5D835Swv1bnn0O+T/TPKZ/VV3yoDLPelPgyz/ntpVpGkXNgSo2F5QDDY0UcIFnJ4
DzgCrOWhLeAaFzB6cUw6JCs15AnWh56Sf7B9rN41kUEpwxZ/7+WWUbc+U7iLNxPqb2uRTwSyxIEp
Z/q6a/1MKk5ZznTrk9m1ubnjzECa+oBG+GLHJEttIAQnRoGnZ5YcnY7L6rQcRn7POntaIDhZY340
sdVvN3jmhAMg7GFgtO/aFos4TAKKdqEceTBZTsEr2e2J/3QgqRFQmISAdvlZrjGKlOHlPbycXU8c
Y/ZdVMCt0GECiZ4nuuFZ3x6pAhsfosZzzb2PzMZcOpuEW7rcgB2s3lRkVe50fw+e7naAjuphyuEB
77GbRiub9ts17eq0n0SfKM4bbbljWYPmiS14Ss24/julgnzna71PuoygX2ggZ9r0x9zSQQbMDS+G
zWjD+HlhElNSXKaYfltC5CqCpXT9PzBwoYc8JhVjAPyCfTiOe2EC31ivkhO9Go1nV0XM3GdUmooX
vfkDTXkA8AMsKp+6AE9P/j42clsZcBSx8eosd8I4ILDxaqqilNt/jT2tfenWpPvdtACpOFxjlZ6n
amu4Ep0K+VzAyfMYOjNGV/2UZ680s/r4vH++OTAxtWvhKiLksb0xhCj0zJ7R/CTQlG0+zJ26F3G9
9Tl0t+Ic1IcxWOlWFJQS3CWBDyweB/x2Nr/Jt+CzQUaI0Ow9cQyMU2QbbapNaAzaetT+5P0es1gL
/kmeXCRt8IFl5suTiMid3cbni7lkNGDjjQP9PcaReWFn7TUjfOcvZzWeRHGrKsPTDbOE/t8rJ4et
3x9s4Zda8Ah8Jf5u6DXpLlzrCxroE00b3zJfLxwk9duG+nId60wN3zwKYzBVV18UObdsK9cnlWM4
C3tES2LE4OToT2j3wBX8jMlOgSsdnlDkckzTJsEcni5k2GROI6U6YEVWVdcmxMorT7wzLs7vJelm
DgAhqZPP+hzChmWhZH0bLBOYbMsRcb/i+5rJEQI54Wba9SNxGrHq9k237sgk6wUo3Cv/lnYD/X7j
NPMASBjwDTOlW7Nk5aN0SvF/9LKNP8l1h/kiOT5VOsM9z9nLfd1LVG1he3bUibBI2tfUWTbNsgFJ
T3o8tCw9SwnAe/HsZ7sZJQE+7J0dt363qk69HQfMYK7Hnsla84wugSWIy6fMiwnCcmU4JDmSZRkW
mcpS0fxXwHJ28hKAjnDoNER3YnyyKJfCJ7x1K9np6uUvN51r/ETT72NpdbeXxPtB0gtejOPtGwAy
k8RsAM9enfZc8OElPRDAzlhH367Td5uIByTqEeHafG8JjICDJag81NsuzxFfy2wsQzXoXeB3y3ZG
uQEpsJWsDnK7GjZJyEcWzbs/BUMpz1UVUHyyZPXGv6sv3WuhKO3pPQIRuEtD2KNu4qknQpbeYB8V
Ahh01vWe/G5FqBUfd9SjwMUGQ+vjOOZK2JOQ3Shi0sFN5DlZHK86dFg0y95esU+vmvDGkT5aszsm
STys301XImwyMNtYUoF8IJz6Bd38R6xP3UN/TYbYdMFABusEgVFnJ/iVMBsV9mVGciTdNoxmlNBH
oR29OhLdfHB3hov4y5sMB2huUzAF8/7KRZVjZf3chYv+GjZ4pqKHtdXkT94Fm7torhhv+trejO6X
YYtAHrDPBv6O+Jzc14T1rZBkIL5nQxJ9aApsQvWBekbifq9UcwNf/LtGXeScPDW9nOrK9d65euEs
Jn3cIlbQdQq5D0GIbsroe8suytIn9ubvx2JC0yc2PY3u8vwkiwO1YA/umAr1j4CEuH35X74GEx0t
2E8nwz0YN3vFdTjBfR8HE/Ih+olfupxA1lTWBzMZYO8ock7tRrLOfE4vXhpNDCA0ADHko2FVQXqx
rBOtwij7bb6GFOOCtbl/VW9hTcvr25VAlKjtkpVrd3P8yeVwBaivnyquzenqVhgVeyyJaOXO7jP7
vjL5mHtvOBdUHBDn3VnXtt63XCbysb6QgCpA1b2TnsbckL9KCFCzeAWgKAt6YlnMEUdXmqTEpuig
3AFGgyps77W1XuB+M9ZKkbCSrPJGF6gqQBSlr0cUOYhyr8f4SwAaFAdV4ZX3MtRevrK/I2sSuvzY
ZZ0i1TB5BZHvD8WXarvnVgKRs0LFzf0GB3GaGY3SDmW4TLauqXx08HJsiRZIClxFWqF8d5LlpSSk
7mRrplUIqWT8Oc/PvP6LxRppqiQq73wMtJt3nwJ0y4nfQCr72AsAaNTDwJKY9WbQA2HZxfO5+Xj6
33FP2QLe5r3WBk5+YYR8bldvMW9Pk7aBi5WvzVUh5tje0Sje21PRGxkutWOTnI8F+p6CsZX5S1+R
8y3NwbXeg9+QM7ohRPVrintiz26JFMy6G96JJOSFdwT/smptlkcLRWKSu/zw2bF/SNaMdNENawRi
EEWIgMYMzfxL3y/OjGRRNPkqZOgbpC3xhT7mkT1IvwK7xRJN9Ud8CQReblseyjTmd6WHhrfj2dGh
l9DFJLHjmB+VA1PBz7418txPJJ8LjlWdMb9Ooru+P/uX0H0DiHCgty3BTdaSd5WKBaXwVQRU8GLL
RAsCw1aO4qVPETas7o6x0O/wlcWP5zGHMIvxyI6HN23v6vg55Ysx171sAoM6xcJ0O8/dNiLb42y0
VK5wEjzQIDlrzVJOmaR93o9gTpjXwqYhWFizbucZXnS4JYazFMjZ7M39SWLn5iDAZfMrwowxhvSs
lp47jbZar5AZZ3h9CxMsdHDvk0v4LQrOJiVgLXC7e9KOnZevqzOWUpvBAA4FUYkwLL7awzyjg42Y
an3clzYvmv1+1z7LbYwoqsSf8H4pi6lRBkl105rywoXopydTedARC2YG7wihPIrTuXTBsDnw6iX5
FtSDFEQrHREHIBwiL0tSFf7qKlDiOGVJIad4CPhK68Ae7NwJ2zBRmkM3Mtl2nsLRN2wYypYpW+fo
iHYrFvdav4Ls2I8MdBPzQ37zlW1+AbEUHCLg/UckT2pPFN1Cg9f2yVBG1+ECQ3cC/q1uoVv8oUhB
E4Of/slY5T5Mjy/pMlY+xnZodSl4ZcK0EHJq8q0ocpqau2GBY+81/1FlZ/FBOlkRBQcLOXutDS57
2qsTf5JmjUXZwgsk0OmiuUXf7LtZbtccAMO+ewrUlhUK11f3Nt40DcMiD/OFhNFcl7tuAyfdH8lv
wSsa3Yfwq5k87QbPOwHvVEf4nJ0m3uscDwn39pR4uKqCczo/f7j7cf4FLZJzfYrwpvNfwjBFE9kx
Wv3RMR91P4Na16C/nX/sxImdzGXfJiFvC8bf+EBoTrzC7oJFGgV86/4uSTEbvB/DA8PSAoUTBDAY
4j2vJw4yc39ONi4NeLaEygfIKnM4tLTYjxeKx0Q1HjzPTXAXvTVDbbJDQsKfwSkLhFSuRVLnZft1
M8VwbCaZWZCsmdtzQFZTUCtEu8zvyhK/BdZ6vd5IlgsuVFFtwM/q55fL7JImS1V6+tqFVrbE9jSf
iElSUNCbxMyf823UrDNW4LXLCbM/JGXIeEkOhV6sZ6cyJ5DfznT/HJDhRvhpDtcci6YV+J/CbXGk
2hVIln0T58g+GMgg9uFhqQcodq9xAcfpOGp8vfyjoMs8DqYR7uHYJSlG1EZ3fnYy83axx9DF4J8D
8CT3TL2TR1s1+meOEQ4x692H7Ru3n7HnesoNQyJlwCyh25A1+E6dasxeflnxhvGl6vICmhbq4fDT
EDtMfHcNsbqBnpvZZhJlhcTXAo6Id0FTb7CBPoAW0vTyqOQDyz0vQhvmfaLtL2gL94sgMTKTNvuw
fgrxEYXkr4paFr4/qNolFiWh7ZbBJptiPUqSMLCFBDZyDT6ikCXdw2mI8c8MkZ1tm1YLviCwSAPy
MPXuRfmOLO4cQuB74nr2hxLwm3u1FOC4ueVDb8LPCnheIg0cXSvWgBA+HIVdOm8bl0pjjMcq5WSx
9Aw549gCu9f2aaIPzumpHVKLJc+KbBjxIu8jbqJt9VvJL68WLXuT0tTsleFTaIsbIh/lSAAd5fn8
JhRO2OsrL/XQp7CWR2HjpWxp9p39f8Lg9TP9z6iJVueJ/vaSieKIE43b9CW5dbEI8sqV9/Xutz9c
SXBafCcwT2PpBqflxY9fGcOGWmbF0Fksgh4HWCdXpyaz1HC9Fx5ywOIFZ9NDrz9+oLxSxArhvHmX
m1VyV4wGgjn/vc6l96sBOBfyzxwNxp19KLwyzIneMmBFOPhwPwbbGuwtIWAMzWQyqA0X3g8IwtQI
v3T2M1EMzVQhVG8SEVNl3jAW2cKWJcCtXnRGtp9kPHXRnbgDGGT/Do30qeavGmHywBCZRIcHOMhT
EJWUzAWHkfCuDTVud5QNX+GYeF6qDqkJ01qyaDBJ/x4amMTvA1VMNuvt2sMoQJNizF91BABoLJcx
9s84DS+tKf51x5EMNJuBxgr9ANlwQZdeLz5mKuK4UMKllLaTaIWvRoWE8is4MyZC4DUT+OQbTb/T
Vlc3+1OxRTE6cxIQeeryd+DNxX3hPpOCSni+ffl0cjlF3SnMoIM9UvX/NhYYs2zcbnGV2nLkH2gv
A/UfyBzwWmmVkQ5urPCB+IeJlvOVy2M4cA9yP+DapTU+3QgmoWmRuimUGdU5W7Pqvl7qyG8MUp6+
gMem3xLSs2lkjM1P2hzvE5otcCpiGq1OgAqNAdbozYG+4bI8Yl5s0J9knRaTehwW5CQ/omf2YPyB
B78ksjoLOZ79kWKoPpANWdKH7/bE+tIm9hkB85Jk+D5S5Xv55IT9lqd4LM78MVawzdkg5thDbaBQ
UhRi1RIakZwJ3j0hHO1FGvba2A3yCZO2uXzafvscGixgxZp1Tf99GVxup+gQzKl8LuFTuqjTX064
g8+RUxOcUVadcCccSNOYpmI4cck2VgFMB4wDWK6QUsxb5pNmM+CP7b6YCOvR7yfLA+P3xva0+c7t
v0vH52xEoAH39YueklpSPJ9NOqq5+0mFDPimqAeYOpithf7WNi9cuylj3Z4Aj0pmSl1DDU1Z5nlJ
Gygyj9YS0vbiQu27cGDOFxvcGruwQVfBAew+cCkyeurBm/tTXiB2Jz3ciI80i37AfbZAYGniBDB0
Pr/G/DaxZciJ1izMCMZwfyNlrFIsiwOGdVXNs4zi+LTjO2F3vsuMRkvVtdopYyU7aPMJ/1jE0BeU
nQkr/CZnEZKwGtMrElgI/ddaoXXaJl4HeOmzorQgxsO60mIlWiiQGOI9NlQv4xUpYOWMOH+imv+g
SBEuR/lQjxoA2i6OCGF0M/oQMeOjdJxfCr2uEC2Hj5kPTO6NCFmhje6gFcw0euuq5TjCbPUn1FmZ
bU6Kdtv29lSfWGBNkKt00iCBiUiVU7gLLA/JwD51alD0cQcXZkJE6lLyP2VYkCTfRQD39tFATch4
2RkPX76idBz1p9BPKVnKxdI3jWJJm0bFZYe00iryMZOwymNL/XZ/pi1nA7/d4aHscVWnT5J4Y8to
3uc4wRBy37050wxllhVvm5QLCYeFPru24FaVlwCejAd/9BQ0iel2aMWtRWmHsCX2CuwzCJAAI7fP
1Zmx6jnuOjWhkx/HvPoKILeEiL9GM6MkB+Rv46zvEjNoup6N/WglXo2JGZLFfW+ILX6oLyB64lkL
zDa+Tw1SwBrMOSceYq6qbDNV20vrPU5UxWZrsWnC8SFc6UKyuz43YApyEN2s8NtqtvuRQYFKVX0s
pTUC9tlUG0+nkqsWRM0JAZfR1gJQP4qUK2USLxzBJCV1WDcY06Qf33Io8En0eOGvqG5fbzwDHApw
vnPFcO5dmeFKxp5/zMrl3DLXjMXUIz4YNdUFb5fSbJJcSjV/rfX/paUHbYjdIvIyLtJ+pb6g5I77
+TTP+zp3DE0cpDUCtIA2JTjzt0QyYKJVXBEmfgBXhafiPFYGK8uskpGEJ+6bbEofQUwg/y2m7PUg
ipa2DGqaMB2+eiw3FqAzTFrhuN2A0BZO/y7lCgMO7HOUmQPp7rgMpFP7d5jciwLp1c/Nt4F1ilKo
HOKnGtLUGjfmfUMYQkAleWCqco3EPpHyePb9sgB1FfLJdCZu0cWDDGolTgWhnmaVvvgFfDMAgN2e
d4NmlOjad5GA0xGij3X8Cvppo8ZCh5LcUT9p9L7S9jR9MazYbCNmrG84o5e3LQpXb2ErcKKcziNu
56Hl06QDBfC61PSsIfm+uu9RHHqNmAqiYm4QkV1k6DTikxeEPzlqsrR/1BgGzhmxHPOupyG55jxr
Ruelvii2Va67o6NEG3a4QG3fzhqVvAVzyh1mqund8LFi/jNGvEVh5vJqxXGICZXW+F805wiPsNA7
9YU1QLX+JBDTnMPX59spTNrqEqJkI8S58KZhQ5f+R1we2RU2hQ787LzYt5c2QUebXl5aiMWQ12LG
DVEQNlAtBK5XqcSzWP9pnX+iYDvNUhA8+ypWuL/P31o5OrGouq1qXCbf7G8VW97LYWZ6I/+8KiyU
JsBh1WShnDFp7kW4sD3mDD7PDD6xcBZDBLhxqIwWd+K1hYktVHkk2k25g1hAL6osFHNvSZFfcH5X
zPLVQ2nv8IyRDK39OY+OhTO9Tif9GjMaNcgBr2GuNhnDlSlGER8BwmHfNBuhB9NJcbvmwfqY6DOg
kN6870xq7kHWE5MuU9B1c+BeWQPUoxTGqP8JOoKiksyCPW4sXaBRpwSMDaOk06HxSWlazGXqkUtD
Ej9ElrqZs/qDkwxIF74fzO6flyFpn0tBwwa/5b7OdX8DKKkSv+L4RJAAgeE+SZ/Ca8qoKEOgEm3c
WfegyDW5rImtjOmc77fVYNiBywXxTZEGAQMt2WPlaFvqufBXQZFH8Cp/XiC9YkyqqfqHN17TBey9
eR443fAmkOBlaS6yt6pI3w1e+CfovLGktSqkZXCOhYZrTVL15a0GxWb34jRsgte7O0FeYcJDaY5S
z8OIdeEXKhLNzKl+WrFJGmu23ibiQUalYLE17rOFox44A5Lm3qLZkb0XuutwZ/u73rPCcWCsP8o/
o8pofH1DO7Tu63DBmg5XKJEXHVSVcV2ZsIL3BCq7ZvOFpI8GYsdAqLkAqu4uWge75c8qAw3YgS2S
ZyK3WY8StfrsNOsvjB8XRx9VDYxm5oKIcIf0HzFw6EwTTJuSv1Dyz80kGWusNHdRvKNBW/tVt20R
gRXVLSmEeEPpiRt/euqlUBFn5lfQmg+MAYxgCg8LHWA85SePx0mBFci1YaNLMKvAqB7uFQ82teQY
svVASaG5KHk2FE3orDlvVd5Bdw/RE5g7EsNWxqz8zeJsmHXdmlMqxeGAvxVUPYZS45G60NOtPcqs
rRolMOC10P3Fgu2DGJ63bj7zQgWq+YVSndtgDwQ97kbH5tzLOP3lSvQUd9W3OXgJyf2uo90YGH2/
j/xckXB/7k5BPltdngsfiN4qRJfUHE6Ci1GsZFYkJtExe5WzKVXSKr4Su5aG6DosSbYyYYoefcsu
HSFG9+YEew3CuJpohOTRJfQk6XaDHg+5FIEk8lMYZya8jyuiOjSBmHIYCxk6V5BnKa94KOYIkzok
8fk1GbLqckJ2CWf9NlIH9qO9OH6J7quopEnQMYzvExyotGCkb9kZnKbI9VICdfHU65nmV6Z6aax2
sNPcilxmLAqJY5LxVzMhDExOKGlvjFRxbkKPixKvJEf2AuMTO0wA8kiZNCexvEDmZ0lxhIcIhLWB
UrUpYLsN4A9bsuARntE8ndXrQnpGnmfYnV0A048j5LHRwTxmSHtDhWWrr2YWO16PLEy1qMidnzjE
5qNsLp5akKqqQ6Mhz/l5t3iqAgO7E9XhPucDLyzCbirh5i4S45K8iBkQTAfinZjxyqZ2aJHDVXrr
Ei5LP0WerIefhQVahSmBEeQ/mqHFTa2hscUbWN5GWfauLLNQBvc8+rT52ak/yO9fCbHZxAPXZfYR
TeF4OIoSTm+OOJDi/UW7uPswLp+P8ugnKLieLLxxthwXKIFGflUbjV2e3Ia5jE/x2qLKYGq2K9mF
AzEkyyVyNrb8PWjqPmFctLl7qqwHUjgVxxG8x8Tjn2fCrc6ykDXQJ9ZxCXjyS0tddYP6KWpgHVWa
3FimBRCBdM1W6ajFgIQjPpRHN7mGbnRfXcQOJTjWRNYMrer7ocvHA4xVHWbKMgB0k0yQ9FU7HfBZ
zK6IJVRb6/ndzrqNYyptwOc55IE8pf+wZxuj5Vfc3RvRMmQZ3MWJExvEl8BBD4mj95dmk6SiIfxd
Fls2nblMbRyI4izCc4uUJXITljY90hnUOluztj3GceAmdfT5P+RgNPBdbnNbSJTTiIo4AaK6BSjY
lrN4GgIKaavVq8Dhxgn8FWYVDwBrzEBKch3G8t/Eina3hJTQKY2sx9W/+qozv4Kspz27edZFr7Y9
xHSaTOGN32uKVkkCSBbsdNC/HD+W1s3Uy3g+8WKEwIRsMz5okvlf3dCAJF4kLTJAqX24oTZe/D5D
RZaq8tWeocFkCL0uMhfmSBV967RJx0Sqa/7/zuYowkOcyDQMLblvCExMvGPIRi0nUj4Z9hREnIDd
Q+ZODDTQ7vZsUSz6JgAsezDDI1pWzfRGkP5z5saFNOfLQ9UaBlFRlRH2zW4ASGHM0hUmhi4mYxWN
SQbQImG39jG5NGT//N6ciYlou4XFkj1T18rzDwQN6ifU1TLjDudDQ0sjqmpLh8VNciphZ86v/FO/
bdNxvsJHr5wQM2K5fOADXvvh3KjtsHSdGVn01pg6uQegzBhdKTIDo3PQJm+c6oqACXeQwKXzs4dR
dRCK+jhGx1H2HBbyLHetZ3ltSmYBz4dWQ39qUpMZVUf01KaIMWdY0d1aHOQBMO/KU9S5mEtD8qde
dwB2D6WeZOJW24imuyfTWGGjTT3v1RjWQFtwNWt3BAtuCJWf7z8VjqskZgBpnSQDdsGX5HpWBk0M
M+KA3dvydBcEKg0luNf+hF70AXEYgcm4DK0wXrtPZS24zDZXnTFzPYcx+sqNJFOKWqsEH62s2KIi
46y5/19CA18jpIKuv0sOq5ZrR+Em0bM3+fk2qp630M+eEOWFESqrj3maPM2tM7ytfm1Ir7e+6n+C
ObVaOw40+TRvEU8CyIMA3r3ukd9l96R4ZqKk+ubWoDqjh+e2kXH+t/eJTNNwQjSfU7zl0ge2rLr2
SueQRrczGqDj5PB31NfEFfMIl2yVPdJv+jtwivHdeo79oktIKXTbz8mnHqT2W5LlCQjayAjtQBJD
44OfWNr99ku/l+iRFxgl+IOwUXMReL1ncxT70BdErFuSfu7c/PMgWuSFLirL2ycRkOhnKyEIyaBA
DnC8RvhO/gIEvLgPfsrBlB6gakBADcg7FLTwvCCWcyJAj0tup6UQbOytRvwCnlmysjysHGaIQWLz
lMa3xcWUZ3PeFghemnCSmEixwxgt3pkWLmoibfyMUDJhuWe6m/WZ41AjkSVTMZQq1XVYhsg6easj
mxEC7hIrZ7odJkjqPq3CPLWPQNLXoUL0HHaBnjE0Ej9QgWuq3SVnSfgyHy4fg9t84MBQRf69ofn0
ZsvWcv+DchT/A8vzZ3MQoTZ+UlZXRpSonYpxtvdrd9N6vVFHygJyB5v+8s9I6PaAcV8oUTyWxsFe
nMbaCGQidjsARjL0TexkSX/OxM9TmAMDc5NpaFy4QAsw/CpfERkVVQNI3Z+7BhVsp5zPkr8fU05j
vfHkfdOSPeqdxLKnvLvviTDNKyQX+C5c2A0zcShrgHdu69K+L/HhnT2FCPpcIvEVQYiMDKOW/sMW
qdzUNcCnAEsW6NMpzT1IPmbT5rcINtvyN25OPf37fqielNp7KM+y/GAWYg6YJGnSYnO+0LThJyDJ
U8OlDjiT+AXfyHonvRu+77+qTTs51ENbQzPfLUNl8qUdYox6gMaBMu1mpmv+7JhsrS98jSCwkkTf
Z4n+cBC8dlf0+Qx8a3vrtrT0sx6tXKImGtOxMcpob18de92H+mRzP4Rf1hnbhJIm4fPPrVQT6Ceb
wxiC9AsSq4lQlMKFtR6yCJ3vSVp8GN2/qYb0hTPviTOC488058E/EoxZPmrpx/bYxCM1IAP+h8ZO
yxT2gzlO2ToQB+B1uTNrx+QeAUw5X/00iMrQyCb1ki8uSxj4qZGXXnRu8gd1DBJcm9Lp/raA7FxA
5B6SIdH0xUH/oCUwkqf3dU8aK3h4fS1A2uOpUT2cJAx/R6aEkGBeWPN+0pDdxYsi2ftQIToHTyMV
AWq1BrBZZcoV5oTO4hThicDigSazh2HDjB11uhiQnoiznQD8EZd9LBJt0+f2QtCeryKZza3sLefQ
pN0jc1Tg1vhswrMHLRibe5kgsJSqLUzIfL6Yf22iZLuwoehJMcQKTTUH6pdvwoK4xuA645uZYYw/
7ytwwgv58QGeI28+37mQlRb6ytluHrNgPiV2YhNzUnjEpmN8PLcJYb8v2CfD1RLRb41k54u8uDfO
lOsCbt9SMnEzKIpekvXMVQcWeIWhRzURx9STBJ2GpLR/p90Rw5+RG6CraCextvnLIawPVti9x0l0
udNmogHgGraQEhr/EPAdtCh4oo7NwpJNTzgaP0/PUBtmu2/nWaQqR1ytVFCJF4Gl9BiUsE5f6L7f
QYG7U+WlzBYBkLSvv9aB/2x3juxhjMzapth7Y19uOnWizCA/NgAN6J8c26rScSal+snNyj6gAMo9
n4EKlSYkkm/+gIMTX8dHwBJvAewosalSfo1c5dqmjSeQjd7RqcOJNPAnBypQtyQuX0+ZDOyOyrC2
K8WSpyodw6zTPip22Qwb+GgWuxDqprUoA32DiLMbyU2n3PlhaYRQo7Z7f7C6+rLBi8B+deX57G+j
d8TkH+EUYproZv1eKb3/670NidOonVoTNUIhs+HDWDvC8sQHFQlgpktMDyeGIVBhHZ4X2cskU8gA
LrzOGvh3D1n1PcANZlcXmI1xuqhcpHJpZqRRikRk1d1h76QWO6eFZCGoT6R6UIbxfqVgyhanLECu
m/DxPmVQt47bIDKy+YeNnbcWepCwdCpeOPgcwky+O/cEXbsz7Xv6S3691dX2IYPIEknA3rcqUe28
X2rROP9RGBausv+WHnO31XsdxL+XB5Q9tvGG9g7xqH77kRIXvFXi+ESqWzgs1HdLdCCp7aOvdFr8
Ax0LpA/DXaB/St1vKGskvyd/Rf3FDHEa7z/rQjMo7k93wEeWVNcaUmVDYnhOdWjPlexsl+8Ez78s
Tk6oxsR4KTN3PU+EgvtRzMD356nu8FPVQJJg94+k7zVBWqnlkf3hnn3d0yjP1JG2gR0FtJ9qpDJ2
g8kbJuDXvcOSIGThQyzC9h3S8sqb+05uPIYGy+Iko29WZeGO/ifXIadDUeCfRQaRXY6RgxkzXJv0
K3DDtiTdmloD6rYQy0jY8Yw7p3/3UX2+y3cpS25w9DdOVQPe1kfcVc4+CQxgY5z6+kqS8CuTLqKO
Kv7iB0BeGOpK8NO6MtredZbs8xrHMwG7IZc+DKX28JZnI0Y+1KIoh8IjQ/BtyebQgUe2AK/9aC0M
OLr++BZ6V5UqP9W7koAe9VuuMd4H5Cca9o2ghipBIgv4/ozssmMQDjdPvu8nxxXZbz6yc0IIvbsG
D06i8+PADagKyWdTtzImjdkjmHB0AaWBNcPCXovFQ9eIXTS73j4hhG2BA71RA3SV6SU+kZI+y5n7
b7ukx72b+5h3v/M6MpeIhpnJzfB3nUKG7Ko52N5VD4/8A73mAHPVmisYSHCIUA/83dm9oPxrNQ9E
ubyL/WGgr/HmUE617A1E9VguOUViaVPbEQFC0Dn3sYLb7OG3uT39TF4JxRHe6Dpy8PEEWs9Ctwbu
/Pxw41j+o0Yccp1un5STDXJHFaEBQniFVZpmiLH3QQ2NiSuN4sRqhWeYnSfsNKLV4ztzLR4fhWED
vokVDOhHn0nDER5QCpvFmoPF0ItMtiz43YnmyZ8DjMZ1jijv8lfZuOiCJ6T64gv/MdyDio1EPq8M
ISQICk9MYwRP3D7QqNFGQ2R9Qz2x4DGhRQ4Xydud+fi1E93qo716wOpIEfODMurgjJW0TKVWC4k+
El2dMVEaynU2H4Xn4Jkm/rEq8FULPU21n8hBGhIqVOvh7ONKo0mz7/dOCERSCFZrmdHjb56KoOO2
To5P5KsDZ+BwzWEJlbF4fXXO5w9izcmuUnXD4qsWEEm6aFik5iA8UClFT4ylEKtObs9/btVim1sZ
OB8QuCtgCpGvWm95ir4+9gys0CcBJfD/GU8fsnlnaSmABQVvS661Mha8c/O2r2c0OdupGM12F1bC
D8zeF/FwAuJM9E9ILFR39goY3bOuIDcNKrccR4rSrmBGMhfU7fu3YDGX++KJw5pxzaNYrebm+l96
h9wpn4cbTSzs4dy9+ololLCFEeH40cmoBttXd3B2Hs6o8WrYQB5CBR+MkBL1SlbP2wPyaOgqruep
GyZeRoKd2gvTeacO+/SzL1mD+5c+0oQ/dfwV8PCBtkl9yyShy1UEGFlSj0HxchDQYMdJO4kd1hWM
XhNb0nf/deZO0iKWslvtmwfZVi39VBlGb5GtUPNv2Npc0rwIKMKCOW2BvC0VGsYBVuFf2bF7R89/
amE1c21wH3RAUrROc40v2pFLWMgMw3lj80kljZX7FJloKtiPzrr9nWYTVhjAbm1qFubkuJ4gQ1lg
xlKO/d0tlCIYvWpo7XtkOChsXUoa3/WLQeQSCrypgdXWB4FxraQXGyCIxKOz8Nj5RudO7xLGHVVI
aaNXjjmFZm1x8OeWEgbD2S4hIemIp1uZpGT/yMMk6cCXLcK5tbhOXA1m5tDASlwhkE70RbA95A01
TZA2qMZt1JpHQuTiUKuH1p0lnEaeRtmyZwt4mdZTnJzp7TAidKyJYmELWRvZB/t2SL/HsS/+d9bz
QgIlHAuxBLMI+KMFkiqPuFi+d5ZCyh/H3o2rQLLxq1p5TDNs6HA/Cnaiftxjqo4VVyO+//8gK/z1
7MsEEyRnk6DdZM6CTU5MHWd7DcvTsFw2VBvJrwW/9mmmlMnOJ26tSGzRTbLl6sZ9a4WaSLQD2DPL
GjXJLcmss5hJWkG0hw9Q+c8u/RhR9mNzX6WwfhlAmnrvDTwEXMIqQRSQASlhs9aDxsf1x4cWnmRq
Noe5EbHgA27WeJD3V4eZy8Hm/k32u0MvnWvWB7RlUcw1OGr8+aLpcu2u+1P1jbYT6l7GTtn0KX9f
7Klkw0n6Q1llSVQd4eCEzql+Hu7ft98E/i9Fieg2R0OzgMyfg9R5UevZgo65fOrwbAue1pq7h3KK
S61PMEgvl8tnf6Z3+K7M0CcHsnhf5GInhXHPdnXcbK7QhDwt7zarGN4q7u/icTte9m7xHFYhzzgo
6QAEa93GEdPPvASS0NLAaHkKh/BnnJIiKs0zYOZ3A9xAyylQ2Zoba599rRp+/OehGsVO+EC8ycG3
oRRf7nEORcxrOg/r0/UR33aDNVFUxLOvPeH703BZ6iIPxevyxL/2TQ6+M6QLtJSpzX29gRDXyu35
+eiDxKqwBUFBJDfxmU2o0QZYmwYEzo6nik/5yhdmTM/c+TMD0VlMnsNdRKOfk9o9r3pxrmuWpsUL
3LoPZd0tAoZeaQH5pLZ8ahZ2hKD+l08fIl8Y2ESPmwVyA/3ykYxRau45kJu/eblHnQBE2wqg1ZoS
Rx05C9xDNGXAMfCnJEfXAMs6s+ls6iv/DRBLJmDimPqgsRPdK4vwxIXW3nwQhynggd8uBrNZ+1Nv
fbAvNZt2DYH/vsP+hlEjUybIbzsqAfa+VdABmEEgezPXzai+oi75xL7fMaF5R/FBN6fX+rBXxHdy
4nlTOwFiFbsWnDOwlhgvWS84CFJAW09mkOiTJ7LlF76nlv5UiUTERvgp0ljEfh+yTCBgBKIHg0T2
Rk2gOSj3UoHLOkD6LZbIVXkSvuBZtKafcX3CfDbFcerHB4Lu22D2/MBQ0zrp55G0W642dpqv2byR
LHAFVn9R1sXwZnkrnQQAqvn2rVt3akdntWzfAiVPEVuPAjP3bKu4ZFJzHkIQ4rW3XDByCV56TWyP
ir38xeRqOEDjzCibY0efcaYLHOr8FS4kicAcZ3UpZp/SQdEippXjFGZ7CeHr1oia77lfxYR478A4
QrZ764HyWwBDKcIFqs3NUNxEOr8XsGMJ9xIsxRFVt/tRFR8eQvHHjrwujSS4WPrsM0Xo4OITvWRb
jv68UxidMj5mO8uzra1jiVv/rwBy7xlBgPe8SsnRO/6QWgqDP7+gXOCU1XAC7l+a0jXJSZtLZBvE
uCUrt3Gas0lUxaepNZsnzzbex8WXNkzb4+RsmGRT8LKIWKnTmTyUIklAGBTR6D4jfjg+IYxwMzUU
k0pk6DOctGpaqptq3meNaFFJSgRtnX/59kqCH4VmHll7bHg3+nJSNXRay424mnqFp1GyngROzxYg
ODbQyIvPdwU8qOy0Q/yvTP9QKxND2f9RgMrXcMhIVizqF7OjIxYE/JRPFReXNe0/QKOfMGioC7+Q
NmlTDXB+SptTVPPsrGqdTITufLHRZVhGh+jNRECPsNUEkUChb07LCcSvIRXjT0Kkqxng4AaRISZL
RoWicCA82swSl1nE4eioOzX5jzM4f/dioep2EDC6wgI0tzHHEN7UcwNItmhbjfwXyfhWhbg6v6OE
3MoVRRYYlCo2/IoLQpLh1zkDhYOVgsS7Yj8Jmb5eMDS/hzEA61sIoZqbZkif0gziqQ/lbLNjf6H6
rHoGKiG47oECnBj5k4kYMpCkP9vEyYW1b1U6vyOnoFuf9fCZL51GdEswFwEIfwL1oXALeNIv7Vb/
0CZ0nYwoI81tLqdNF5fgyF76+LpK0m1q6qEr68F1x6aurvBgJNovYbjNhVpImfpMyBhCcMvrcoqa
V9TbqFWqn+lZh4JyxGk3wazVIFeGGIKM0S7Y4WPbiG+v5kMOm3nxNToqhvXN9jS69jFpE9JmfMto
g4NQ0YCBefG/CIZOTiDiqtW9zBQCrNyTV++213ToBsW6OrDF/s/jyyC1a6Y7LwTxP8pddecpyRyU
TTWHqpepVo/mQL49FTJMAQVhYxj7f8DU7HGgg235yAt6xgXEOIoAO+vUk7/CZarNu6eJHAFqxtgD
3EHCfZccy/Nk2wg54eKUjdkBD4401f/Z17d20rw8Fs6eehVzDCQbH/om0vQO43sfJhKUhubj0X6i
zY578I2p12ih4HDkgVeJXmRMeHTf/hZY/A/dUzwAgCHZ69a2yu/w5foUU+4QhOk1s/M7S3YSwe2G
qehxuuAcjuSMepmUc7H5j/MP0tZOe60K3IHp3X7etf+IU96PJP4JEZUBiRldDkpQfPho83P77U7U
q2D3H51G43qvLqcLy3uNQ9ph+nFHieIpzDQUClTexP/yJMWoI2dNoUXSYeDDTASyRcmLdEkGFN00
YgJkUVjipLPoOGSjuLbKmBmZInKBRh8lw5RARXY2VpKUwOR6kpnB8MQ5BMp0BNeqo6hYaXKdjiTT
iIAXiAHYH0npgS/c1dCYXeg27hSlR6NddDbDtTpsiVP5SZ/qwrmRSLC479Vdy/CT3dXhy5g+yXkM
hOIekGcyOGYASYsr2oCqBiBWmbZBYRrvOLa0HdcBR+DksPhLE8ViLjN0Ee5vlSu57lNuNADHykkY
6MP22KBcKp3Uo8TX77sazSnG8IwtH8dFOeDIlI5bn1A9xptvHAt1rmk4nQGsqKNtRkaP1zxB6E/l
nxiDTqIvXKEPEeQIZZDJLhTbn7Tva8Kv9UoiAYhvpQpci9GpdVoY9a5Q+j2Mgziv6GqPOy8g/JEf
8d9jJRR3kB2sh5FRmqprIfUhBZP6GJFOSAwTNO/9BRaShbFe6tXfBiAZ8jQW3AHjXkl0aXtbvMot
hH1HOD4T+1ToFtAyuf/PGK35S/5v+UqaWT6VCc3kEsmNSko5mIvANDtJfDTBr7+JXziMbDVXMtJ6
fw24KlTTfapaQq6DPoA4aGbT0EkfPK1ggZ3SrKiMrwGLVWhDTqTDPETuWpDEoAWi68AGKDx1t8WK
yom24lRHhsIbbfcc6Shb4ftt2UhHZ4smxdGnfVEIlledCIvjH4GzjkranwPZf2p4DwuW8W1FBcq4
z1lATLZ1ZKvMIu5zAZWctqx0NgJVTCBNv5Us6MCnZUcdZqnZCMIRMZz6Qa5/7WOXpOaNmApRwVl5
WQ7q6dvOM1VGvNQekb4B7AJ8lOLDogcrTpJPjYKcOO1ZNgpfLmSsA7ELcZtquOQ421B1ZVpjtKdu
nMwkrseElDaPxa1rNF6LO7jrFwssCeJrR5wWqV5BOK2HY8G3/AURCrYD4D7gPdxrsvJSJgIOaUBs
C0K0xHlIc9QcOo92uVe6Ow8sYYmMf+Nf9KToolRhL7NkUbrsu/8pzabZtYKnnGvgKeqms4Fjh8eV
dUSEZ3AjzRdCLiP/SvDxrYRfcOd6/uYlRqTpvjVN72bMwEdl+CjJTrakW70Ura/YG52G1VXgcree
ruUE6rC9dF9bRLaYgQfJKvGYPr7c/B1us3hD91AKxuvRklMeYuxf0s5PZpeHvDs5fi0mh1eywtZ/
U7hFd4Do4zMeQN+RlUJTiS884eTzHAuliBtJQ9wsnBuWuYDpB8pjfZkMh5lDDSIqGb8Axo8+rqMT
bwPbxW5vidRXePo364EJUCBZOdfBiL3yPHvy0y4qOctcibfE3bgOW3J7k+BB6pWZAXjM0iyYCy31
QsxIosKJaRjKIN8+PrODQhJtYP2CGtFfZe2uKGG0moeDCBgkLEoC/aI+u3MGeyc8S0Bi8ViCpPC/
Jnd6q3daSuxvgmLmFr8ifCB+FUx7M2Ozmu5C+u7TIGP1RdeSGyWDbx00CT7eD/OsLnH9oJdxtskA
9FYsjo46FpIrbBI5J4/tWFNmwHe3TG3KDBbVLk3nqa0VIdhWZpdrujo0uasGX1ehQVFsSIZTuBHN
F9GHqGSK+Pq93peFXYZwpRbvUlWeMw0g3s6Xhx0t0zsJJkC71Ov4gsXjdwoNUZ8XwevJa9M3QIlo
CU8Oqpd+5zdGjGu3Ii/cEgWkXI8ssW6LC/RYaDd/0KmczXV+jZdX4w2vCG6iPZKx1GTEH2hPsaU3
gd775va8JPJ40FJTcTPevtclt3y0DW/j+TZ9K743weGBReg7BfYp+1HARSqhPFai5CBIjjH9T54t
J2yXO1J4kgLKrYk4uvwYqZ8RwkcuIRDM4aanIBbKOGHyixKVJiggIm8BM2e5JrraOUQvClpZUWN8
JoxhFUtorawNq0cZ6jVGdNrUvE3xWcA/+jZI35SMXQSIXZ11DHzEE26JMkbMZmJ8G3oLprrz/3rD
AX8nGXBQi1aIVoxjwzu28n5pDpwFGdvDCR/6racSiQuHEKgncQ1iQKVUqMZ4m3Qu1rnLqKHkfhDH
Kq5/BjDyTKqbay43leditiAbn5POt63Ga4n46dLP1G6XikeZgLTVxSH2nuL9sJLIIP1WtVRZx/1Q
BXj5ipJ9go1gl5n1VpzpkVKLKPbnNuw4jDuvkQxHOl0PRl4fN0z2d91AA3TNEzw1Vh2VlpdsK9Iw
S3vXqbYQsJ9bgPs0jxXcXedBlxkF+Uyna8RR/rEySOwt75Nz1thp6dvFauyy3nuSTRaNdld0EFOU
JwH28I4oPYhk693FFbvZkO7+Fz/FDcYPl4yYZ5CL2hS293PwDXvY5ZTc843GfjFF3DEZILDM3/S4
DQOiwp/jZm57Td77uFeT2RmkN5QSKwpzC9Cb2eTfXXdnkCkkxwWP034oizU5Tpx6T/dlrqwBu2L5
Y8edjJmf9nvRIueKJflK3p5LnZPNRgg0b90DBGZIOJTv4Qo6SRa2RNhfDw9XN3icnQTXvgqT7H1y
GMJySrj6EwCArovo47u6Am/ySmRROH0J+mzBEdpUy3QptqInSKdBQHXZGy9AODuvraA9sEDXP8iN
B0vFPEKXLZMo3rHgaZMzYgFFB60h4R8gohf74aPBrWlTK3/dKbE1kptvJfM1QRs68eJAyMK482Bm
RUppQjIGw7NXkO0TDSaYWC4djma/5aHXUXBs+3q6mXBce32E+qOHwbCvryofYSaNjLisMrwlYG0K
c3lYZ+5T23cCaZ8GTa10kKth7aocbzRjq1+n0nG1eWYudMIJUeQyrgT6siGpOvo8pbKcAvJaxRt+
MmaCc6+8qndGxi8idwvELasu1SpQh2eZfLV1j0nywEB2MhLCP86vty27/F6PT+DKWgwETWd8wXLi
MQXRxfTrSy6jpiDI8InkcttgZGLElqcW9pNGCJIdlihkA1Gtct2v3XoYsHUcINRaIJwQsslUd+LE
FvnypH41AKIfjZFoFoIW5UqVsujyFvYWtNDLTji/1itry8P8srvcOokhlNx+Q9xvTivbBmTGGqZg
X5vLM1NUga4nr6ZPN9dNM9LhD+W90wBU2lxEwUItJcG8/q24SlQEOHfAGX+Kz67TPKeMT7oGYSiN
t9hQxfE1aKKq45Io6RzObi1jtgSNic/RRuudRDB2R1UpZOiL0hUSpcCo8MPFEhLwjSTRCZX2KXSE
BhqCSyVj8IU4hDUKuR9MoQhJSwTDDcK63IxS+tubvBNK2AJ4+YwXG7xYoqZsg04+GgpJpkhzxc1f
ItEQhtAOS/eHuYkRoRS4A+o8AAovdA2FA+X84LK8ynEqcQClsLl5EV0AAIQnrqZOi/oIu8DaWuo7
nUKDIHLBXAATZviksmrPiUdU3BNIxtHNLWixapsFdsM6PTOaW6k53YvK/QlPYGD/bWiAJTWe2lLa
I1BWFQKq5yTNoR/Oqkvk2DOfhkVWli3Ypw+9DGlQ+Vs1nicepV1Ebjrw+BNWhN8buzBIwJffvEim
FqKhAtww/przqG9LHh8OgFOzqcFC4hBCgtN2aEoOduufCxMcuu8uhXcxntU/4BEZVM516pAxNsFh
MSKvI6BWpDJnBeVVy3PCCFZDQUO61Xxo1QYZEzo5W2CnqIpyxRLKcYgv5HfyU3mWLiKO4MD/y/JE
W0iJyTp/8ly2N8ocVF2qfA8f6fK6QQfBuDaEJ5MB7q1Qp1PS4KWfsUg98cVxRYmDf8Dm3LVdkm+Z
3kHAjeWPfapX3nWR1NMeHNfyFAL18yXHh0fxGwRNGTRY3sWZV4qDTIHtJAr6+CvqdM1Tvd7r15ln
/q5sa6Gpf8xyNTbrvrk/cDQx6Pt7lBG221Qnda21C46sLrdHZmYxVoUjfhyCdc12ZcOmUEAjtYOL
T55uuv9U0lpiPTbXtyDqEGqio3sa0E1UazwrACNrFePJJKYTYw/v/TG/el7I5A+aAOmxR45odFCB
vy2Nnj2x9hdKDA53OWn2gXOKJHiXZiFRHHWnatuIPxzoC4BOSbWRAutXla327H9Mnr/ZYSwO4wlE
0pxGuCLLqiSQphBguW8/tXcP1buP3h11KZqUzenXobnvyGmf90Dlh59zlyhtyHr6CuVOYYrJ0g+O
tr6NUpIPwJFmQlXwhHHhJzkMrfNSEZYb6JGLBrnVhGDj8Wd/l1olHjG4ACEs3besm21kjm45RO84
CficlNxhgfS7rQBQP4rm2pwB+eyY/zLFo0F/zqYhSqkO27vFgwlMXK6CpD1ffBOFArfFB0TTgVEq
9li5B2K+3wuMZy2UlEKJ/o1RXsuk84dsIB6skpZcei5JjPcuJaE4DsdZ4QjyRHOe7dhuXgcn9sN1
wdSKSWU43o/Qm+6st7C5+Zfwaxs8Ifo5ZIehat4AcnYHGIR74nXXc/PSQMF7lm1wN22sOoKGx+97
51keSQLDV9murc/9XPJ0ek9ududUpeVUBsEDH/O3bqOHV5q9C+945kPoYYkfvLeyZ1F6Yp6n3Ioo
NBgdBpLkywe7OUVEOqKjdi7KDfHOZhvHjfuA5NoOIKjpWwVrtcX9r9dgvee25C/0H6lQ+NhzHHXd
l8FCLpDPR+P1nXU7uuD45Ns6gLIkfN6A5y/tIFesnA5mFQN/T7ZmmFQD1FueArwqbau5xZq8L4Xa
A6IfQ9GNbKC4aj3nyF/f3FCoTkBGyOtSDT14TQohkDRNoQHgyDTunbdbOkhPtG3Z9QLu+m5I1K6m
9G0kBYWO8paPkk/6v7ErXOz7ycknAGbet7h/Y4TGqWN8yA7Kjfwv0bnEXYn9/U/WjXqcM+VKspBx
BKxvJ/KixOjkrby1CpYCkFqfgqIO6VnyKoJAfSz233v6WplDFKar7uCyTXi5X7cN+fDe1UXNii+s
lNimqeXyGqyjQMSfWLd7kBxqeRFrVTzCdlFQH7VdY0FzJaVrYM1K7M+H2vzDqmGdeisXA7elYvi2
RnmFY3+kptFsDx4d41ZjO7sxAjByl/1ifRdruM27EtumYXQ6Q+4MJK0/wcjqopK1jR3tipAVj5VX
ydYNKV1q9KfZnj/EXI20OVPYk374si1NWoWKEpQlutDPmrNjv1KrNqXnsCm1kPOcAea9CWwarywV
nvlhWJWuCYurnSJeSaF4/gt0e6bvA/sX2VAg9vumxvWYSuG7Xd1xORFzDqUy+PiI9pbPEQ9qTYYK
zVpyEWVWtHC+Fi92x+Gow4pJQfl6X1QloPvaUyey7Zgdf9jh7w4IgD0+DZXd1GZQFFzQhugWkeyt
niI6qCZmD7ZdmmkVgAIlS/E32l0kLYZKHj2otYuDh/S/G+GqHxSkwIks2F+WoLxrRU6tqFpJmev8
miOBL3SG5eXSOw1F0wVaAcuyragBYzSjDB41TUa9nNP19sZc2EmcGqvxCW0jaxQuJtSBZ0sFIFMw
0GdyAXXmR1Kx1ZERJlj4BMWIE5zYXzGHMklzZwETpm+x78e5cURWXBa3VmLLDAM7eUHFjjq14wH5
rs3xQvkd3wrWPwQ7vKVSNpNXvXoG8aW+RmYmNj6eA33UbBva/m+tGOCUwOUtwCVCUrKu9cNQu52P
offBSddNWNnJY6IaltWqb2Q/ufMVeY++lsdDwrSqdlY8hcD8F7zTP6nugNUaos0XDSVuCe5PRDu9
ZvqMv4wq3w+7mBSOI8jIzpiBVEKj3Bd0tA98UpbHb4sognvQIx29hZ3STJmeyMBHjgIMoYWC0Kom
HIytUrD0pOnNamCbd2xWcHUh62C2tmEQ3gjUaRaGS1OvBZpBi1YKILuo3U91kmM+JT9qYlD31e96
WcdhnKJTg2gt82j0tbYazDqt20VJkRPoxejIaN6A9vp52n2EU3ajt8DOwRGqi40G12OcqupnqxGe
EFQ8jIVvddqCGb+7E+Bhgbl0ZR9rg2euJb3pn6ZZS2gCkoysI264LQ21pbcE8VUKCnx6PaSpWt8r
bcgXT8fB605UmsvcFQ34L0LDofI2aFLDBcd0EA2su3QK3QLKd2/F9R3eiA7sOMqas4SAa52B/nRs
rrkdW59Oej627mv7uKXcWTKx0kSuhvqH2fpsBdsblkLV4m18HrH+J589+mvYI79mYjRcmzLjoB5r
/aPqH2/8BELjjfDixfsOd3Yjnp/QsSNPEpjo6HZXZCm05FzZeRZCTVC98w+i1pe5+y8FtBGUEraf
o4jwJDJBMPugqHgmo3bn+AqafKe2OWVaQ01jA/ke4Jj1QDNy/yqFvz363O3ML8ZA8b6e8HATFGps
8vS9UdHXWcBrxGtb9iMvC8Z8vFNvjChmWKVMb2jUvbJkF+6J1QbFquPPkVZA7s7YCxj2D1Pi4xY3
kup5DD4ueV78OrGxfrz/Cf2LysHgUxev7caYlP1ysjO4jXLlqYinvt/QY4xZFeR6ndNOgXWeecpl
O4B90xMgleOF3WX6gY0std8r618gMrs/KycFtqQJujyQ8yaB2Y+2ggFnCTWOczBgRctgGcad36NM
61T52visKwk7y3a7Y8teEXHnl+2LNlBgnjNbcABq0I5X5Y1tMyazNE1hOgBb1IL8Kuk2XPkmx9eA
0EYBftrdY0WMzJyzgeS77MFSYom2Ec9WdVavD6VLlNcxP55r9Nj3lFRmAOaK0quU5Js4wRTg/7st
2Se5XLuF+5AU0rttrSVusUfx5wwWIQOghMsZTSmfGoHASYXuR41cteInwIrtrVc1jT0JzrTi1VcR
kHPKwQb4W406NeJIadgbRhUZqbMIwMhd38Q80yN/s8s8e9uZbnzIpdQQSwBJ7EzY1Qju2zhk+rib
/xbwGGqCZfJxn5fLQs9o+QH+TvvOr7D6El3JBwnPoacuRCDJC2NcYQnwjAxgOFV1wK3wfL8QPO2W
qiy8j9ALwSKg8LnsvbjaC9FvVVguXJLBnmSL7tl7Idg9+8+97kJyagmS9QAbq0cqNXF+Q42+YcZ9
ZTenwje7z6aadp7MRMbnMe3MhDO3IhbUzcETw0xx8wbgGLHX8uTmhn8ZW9DQyB50/7IFrEs5KZkv
pNknEHnDvHfZGJneSYvIcFb/B5WIXZ+LxxDsP81oHFsAqZnTe9s0BqohkP9f3wZxgQ0VTaqfhp6j
E8JQ9U+bYII3vsNTJmlxjmrWe8kd96EtHqzBfsY6SBz8XRktCV9HaM9kUyJv2EjB1hRYcKo4e613
c2weZGffJS/ESfJUDt/TJWDv77/Ja7ncM36zkUu6qMDlNWO7CKW8FfoLbAyFluUz1S/sWrqMBmA8
2i2A8PQ0qbjNniALasv5I0B9gZGr/4T71zRQo2ZTEgjr4uABfC37SLZNxfKSkXRHago0KkhgW4nw
+YTCndivHJbt8r3p/szBlX81hz4b9w+HCi/dutFjz7bOMn3DvQTDf9WVLzAkD9n373qtt/gv4JlG
EH7pw+j/pkcuGD2CdnEH9KjyxHlWbF05RcIUEdrqVje27YT4VFUWVRJ9zLA+6JcJ5ng/RyPxOe5G
VoOhbV37ZVuEB9L3/m5IsqfJpgySTY1xXMGj6pDBzoOfm5RjzoJqpnNVtct62lHgkyBhS5u4D4bh
RMpRraGcyxCUiJe452Q/KnysWrPdLqdodbGMDW2oH7BKpeLb8X9LCm1mVIfnTMeCw5vazD98rKA6
dkEmRUW38ApoY2icrWNtOiT4zlAzxNVrYs62iEra1+qjBX2nyf+qBTkqutS7NuwFmvvcgb0WLfWi
gNEeL9Z5ETqhRCCF4bObLjTBEAGt9QbRLHtz2tbFMKA50ewkNMn3TezuKPKDBMb0aiJyyqoqWx22
NTzxC8FIZpc73kgU0u8uVx4pICdNBa8AOmiF5n8wxsaTD7PIfgYfylo8Ec7hX/eTNc4CM18Y4zzO
KaleYFMqpr4foGZCgzarE2onfetmyYDvSvP6EcWMOt3FjNEYP+tUzPCbx0SDCasu+FrnEU/SKmws
wtBlBu9HWwd0RryXHBWrbsI+a63nife9PXUxwlUW3/ALxvj/U1pEEVy2XU0i74SUTwElschVhigV
JQ+feSzmJDhFKmrpFA7sqdQ6pyrbQXN0MraOJbWXIEGk1kKsPDB7Tq/tXmHLdxKW7y4w2uCubasH
XIy3viWfi4Zyp4Ou4vfxaoetQjErFeYStFN62ueEDvsovjhzrDc5k6uC05laTBly8quh+ahFyVLt
kUz8SqTqmEIorNW9YtcgyyY3a0A5jYUs/xQ6qnGDkF/zLjeGZNUDMrlKtKPLnFRoqa2vQwoP+yU/
NpC41MLifblwvcWaGo2+dr4YMd0dsfU504gC9TlWkiMMeMDAjGqNkyX7rvwMlm6NqTbpImvH0+e6
byeGeEonK3gurhB6hGuTzMaMpnsiwiRY2H/1eOTCog0+gugG60e/kCVCdTiarg8S2UlpCbDkUCtI
bV13GnJL00CuVlNJWAHPfYH3qRQ6RmgkiYsXklx3VuqU+A5kxzgkg5VfwB2FrjCqhD8vD12SJCTE
jZt4FrnfgvXbS8i6Dob0ODJAnYvJpUGmY/4YZz9qk6imlOzDiQy9HQs/TaWavlSu/pFyC7Wg/LDP
LG16fmnj7BLpjUWSaGBWfC5c85dhczp3iyv6mWOj18eUbMERBVgUMKB2Sc6x4neazbEh/4Nudw6w
6wzV8O5tS4KtNqWM7o6TZEAjKRkwIkmGtjA1N199GUhXr+4HWIpPssyJROj6iKC/fos7OTe/7u8p
m85ixHEmk7kh7G8T928Y2RwcQnurs5rOf6SKEHG3/qAcwvSmt2MWdlQ3dan8q8InO2l5jNfv+mKP
gLwe9J7WzUxOTvXXQNlB+XSruRhoE/U5d+u91Lq/n6jeFgOItOoWLE3usiSmD8eHWdFay2bLmcP1
wfYZyPMIhIsAmUp7ciJvgOZKrIhR1qd0tGdqh8RSbsgIQO+9BLYaQcaWCEUlQTPw0Mc7JVa4B+t1
zGQ99TTnXdJtW3XuFDw0OplMFNrq1dPbiaf1ISVTaT7smCzwdFYXjYi5457LQK2T/wcsQdbk5j2o
ZHDRSPHTRLUh9stdUJv6tc81F0COe6sNgXPmv5PI9c+cmuIRplSrFH1JrwAsfAO0zYCoR9g7G0h+
9QSWRcqOKD5YQR4XA78u+/P7ZMAH0kHW7dKmbLuoe1ZN9StKn3CNH9TZS9G71dSqu2d9KBoejXdT
Inuq4Yz8bP0BoiSJ8vghth2cQ9Gu+oAMXWTOzpfaHQFTq8vxB/8oRkgAL6ykix88S0hTfzwpF68/
ZNY6ZG61oddDIwZTanSXokWMQDlV4gv2j1wpUBcwTmhqASzKMKTsGELuvnSQWoz9WhE8ntf7h5s2
SVfukeaTAuJNZ5zYRevfIb6/P9ttVQRytWKC06fenS694gv9K+Sz6L3xoZOOZywpHaLTpqs+BohM
dVsDW40b6qgk33PBIq+8BShv3cHBuhQhJmfMsVJWRKFztiyrk4S8Mp5PAIU0pBLCWkALv33aLwU1
eDf6nMrH61iomp9DeDDctN4q5FvB/XHoeDikuWXiLSqY6aPWG39Xvxb7a4Kizy0PEwmCRFDfAmBj
k9pkJJuMyuwyGOiBscMWkuXJacTxeNACaqNBjpm6CPmyHdeV3hY6Gm2yS1BJlvmOhU8uQgxW8loZ
Sa84e1U8a514v/N6cXwdVDdiavtNG79B2c8VATyjw0nCb09xGzz7Oo2enP6DBZ9D6LNv2Ne+zi2V
u+HNirYXfBiA121zZfNJdYGMWnihVXn1kKxKQ9E9NCAhF/yACqnp9E8wJ5LKEvyPKLSj2QVQitxp
esGCgmMnY2VxwPJxXINx6aB/PFLaPG4y/Sck1kWxCN/CotBUsxJlFYk+RWEBgMdFvvGQJGjxYx2f
fYm4JuWEeuibgl2Vba/wSbZu3UbyOMVyFwiIfxEMOvR+RhVRV7cOKBolwsJgKTtf122cesh5oDCc
wFFqkMIR/bGDU1RSDBXsowTxEES2ka46HUTghLv9pCUyuDxT64oIwJ83ShRLt3v1wHX8HQzopeH9
Jga9lP5T8WLm4wf+8KO7vM5ZMlearW9JNsDfaoGHj/bcyWL39rgm/fLyIBgAOoIChOhylfiNm9KU
hA/Fc7ephh5ELEvaHLH3zTznh+zGkV3B7e6iB9KpdxilmEb6MQNuuLkGnDnC+Ebs9iG3xyMevnRr
IIf/P9e2n2+iFJbjfaPB1hhSjUoPrRcVfiFQlM/Vrm6LTwgSmJ2EQnf6V+WjNrwsbn3d8TqQ7Bwj
k2kqw/MFI6QEdY7q5s2M/VvtQNm2dlIhFiZk3mzffqF++UTjzyGxSbxUqZuQmp2kT03ZGt+dWV20
+0jQNxn0AETyhI4xU++rO2ZoJgwRKP7jVa7qD8mkIchiBj+EhFcSAk74Uy1NLDUgDrMJG0GW2BEZ
xJmPug9ZnOzGsTAB5SPgDXxJWp+pnOHDp2HqplX9VDNXDjLjUQmApc0EqNXeyoqyG3yZwlHQZ15a
gQF4624kQu3inhvkGmDl8VheBhN3mL3a4odQBIQCsXoFFvpX4iUDiibVPD09zMqz7kFlyiO6h4LB
BTuU6CnBw1PI5LjPYMD+qUOdXteUzP5ACdEzAft0pETdx3NwVMXQW8uJXsQS6DURWrHVqXVvi60X
HawUzcuxMquAX45gWARHKyIM8/T9EAqzNBa0bbegKgXZ/hRXcpoCXqQT6bkQxwF+StCD8TNhUwJ5
ikcS4j5/9GxLSQCf9BOI7Z316iNhDGWp5C88EVx+AYOMtA9dBkdNQ5geXa7Kk5O9V0xefGy9NaUX
aWFOuoktWttG6zVHRPHsD6OoxDurE3XS09RgmG3H2gMMudy+Lls0OvbBZuOjTh7b+n0mVWe+kAtX
HA5Y25Xn2RgfpI6NgfWJEsvuHwPGAqH8Xb39OnPeu5n+7oYPv2km76Locx6vPLao+WPuozmP7Eb4
ocSRkwy6l3IWvD0im9Qkp9wik5LpNdYCUNTBSCmEH06i9dpLoVlxqRZaE7gb71Y/zLU0y0fpeCRO
OMtowcPU2dzITqIfgCLV9coNcYmwObYAxDJPRHybr1tG44qTFbcaB4iHGpeBUuaFrN5lW49C3xdE
xAfHOfFhfy/XRM965B9bUoE1ag6l8tjRw+Vstn2iyGKU+w/ksLdvb5STNY1eEbaDia7QO+BpsiiC
kxuJBDZQrRSSRe7uQaJNRHm7YSh6+RPaZ9bo26wSTYbZeB2YuDREjo1n086QA77a1iNYEOVyGywt
MRekhXt88B9HP+cQVcBZygL4aIlJy1KkZtRIzqOjkoNIkV+LwMyIA2GXX5m07GzapRf1T2ZBC3KC
dybcXLX0dytI3X9CEAxZGfAsA1i7qrGkZydd4plzIDMH+PnczV4WMoR6fxgVPQmYaK59dCbzAYiP
7r0fV2aVPJliC3oLpYp2Ormf41I3mDVMDv/nFmNKKSPNn5LGcqfmwIGh3aKhnIL+HE5vHnv3vMpd
+fbsyq9675baK5/eSN/la5aOCulhbGzLAS7WHvvPMMm6f4I0SzA7XLu5tinXeR/etlJnizXf11Xl
3Y5XLriIptDEkv880NWVfnfTmpWkaanVRezeg2GUD5UDdOpUaA5gPDs2OLhFDGEl42uW2Y/MWUDo
wu6gDEKfgMZ1GoNJOSTLdK91DJbNRSi8uylx25oCsOG675ABppVNuFSeoDicE1eNiyNfd6kn+JMq
H4ABOfXxMgyaDo5Ac8S7KIUngOnY/TjY/gteZGQPRfFutn7GFPWlbU8GlI++p4aA5r33yJn3mOL8
S9HH9u9GqMApNDaunZxLUatvyySZUO7vyZvSpzrLE64vZQeo6KW57WFI75lYZ7eSGKPZSPLcisaS
EJIVcHhmhqeAxYn9KSyQ+j/LWqM3UOM8X5k9Pha2lrZnlh8ARVmBZZ70NjUXE+gOu8AlsDHAOHmy
XjFfD9rSXg347rePbBLyNiozGL/n8z7Mx/I88WePSs6sP03o3C91XEz86XACvSkJ4x8KJYhSwjty
bdlgxv3IbwzStRDXgSxkHxHJpLlARgoITfbhvU3SEbGUXV8U49bkWEHUn6tB3B+i+qOOzf/riRHZ
+E1PAGOgwcUBMwifA1mY9jzy7hozYQanRMkvjDMU1jaU4WvlFwo7QYJHGONp6dtOgAkmV9QwjTjt
q+3izI5asKvxqzabhINrQBcXME36D8QjDVenUp7z+00E3y3ScYJy/HYebPhrOMZNqtfo0j7j4Pcg
BjeW9qhhH9vYvutNetMtKnaa3Tl3WPaO+5Fw6uUkCAzmjpaSzBErIJqhaiDk9uBovLCYEyONQIsg
4DAa6ogLVtmLy7cqbSXPEW6Wq0Fbi7wRUMM7ib/kUNHvzluptQ3S/9TiVlGg2a3448XcFwUYT119
CUqV3NhR1Pahvpf7jVyB0vLJY1n8a2NaH1KzxhSdxluMJrd7O3S4tcd6Xt2XUe+hAKXPS3Nho0ld
3Pp1FdAmWLra7R3XBsI3WvoTA9aaer5kti6Sb+t2dLUnBxgV1j/ePX7alin0f9vDYlX5hXijysQ2
1bdZRN523oxvcWZPEo2R7NVIsuRn6rXzsnqsoWYDem92lf9Matk4DhpTV5NBZQkXWmeve4Ps7u0k
zyPS/jnfLsLLa8qXvs8U5kROZbN+uhMaPVSQ5vXJ+R2pMhwXDl8bxwYEwsp31WSCc27fj4p1FPZ1
kkUXdLHJKzVJH+a/nzxETbiuaz3I8McxJQWoOZ7qL4FBUbMOiYM3On/aDtTjTSVKu8Q+eMFFB1d1
3Nx7HQ23BKp9VwZP5WcboouJTrJc2I7EqRBKHBH18F6fiWmbpsjuy4xv1l706fXSjteLxcmm6T0G
ZTlIYthzV4sSEWHNsQOdLUdmu+baB7X1rAdrh4WxsullLw9bySQC9ft3WPjaW1lJiOf5MsLVOGnC
9YzFdWCbQsyO5sBIg20RI2OvLetp8kdH6W+C3PH7AR8KOgjzJkWCyfaBKOwI3xgIPZskDVnP9OBY
w8r82Cz4JtRWdaL6U8zS0QdfEVDNcuDzNF3UfBNn+V8rij/L0Fjrs0+kMeRjQ+NVrP4EFBktWLPg
lHKXPYKrkjNknvWXbp9890XUmLRWYEZYGV4TmO8JX0hhBMMlN4607BfnjmxJC0E1DH/TDSIywzP4
hTWDgWh8qlY+3KYXRXVAirUcT20zmh35yhEglttybWoYMPhCrfXXLlViq1xjkX7yK41msWfDl6qk
gLWPceP1hrwZrVLbc6hqgVGQXcNuUUWOjYltQuk5ggAnbGB+lxwqX1JOaGQIPdL1M9dS3gx1YBF0
aRF3AEEWPNXcKDVcs4nOtL7UbdQ7kufjYVcqWsuhGW74hUNyAdmQBXCNXyKEEX4DVnHkJo4CnJdL
sdboeMLO60TWd6WUVdy6Kl05JBF1EFp0RukMQJqovUdSQwOW+zLFVdscqWoMXzMH42LH5Jk9zXGN
oR2ynUDdmE6ohIGVeW3yzNV91O07EbqrfAFAeiJSUUuHhF4Jakf/7xDz/QE/HvArO64YpmQB7EqD
3XFNl5WYH/a/2zPL3TH7nhfIgYx3D46Pl2sej7TyC3p/5kk8eDCbKCOjnUw4z9UbvLR5sVfwdqeV
ITUAF4CdZRGg9cCDgKM7pS0vcSiE1dzWODnTo6CI0d3U4ZixqalTBwllbUZyBIGktsOJEahUWQBJ
mgey8XKGxpBTtOS/b03ymSrNWdlmQnRdsd65ICabi4iCb9dNyl4LP0gRGKLbfq/cXh2qp6IqHG3I
3SvhtbFqIzpUnX72OAlk1+JUdOrVEmgBqu7jvOiBtOiHQ1fmd9PPPDLlReGk1NJozcYu4D6FYjN9
5BlCTQLyjAvxS6UBuzgRAPeU87mWQ5aqElteMrg7djZ4RsQ8cTvH4DsNw41bCI2t/RL+JniuK/iE
fn2YVpudwCFuQEC5Su4CJ0gYzvHCHp6ZPWkvDnSP+2ztNSpuhSgEo/82AaaJh0QQYPGGmsniGxwc
pLzFzuNtH72LjOO4fuJJy0AVpnbbZLPOXOnby6L5BWXPptp9NxXyR/hU5s5/lKC2kHDn2DfpvoBg
5Xql4zCcDfe+hjgYVfC9AgxxQnDBBGXEvvcigpobfo9iAILAiMS/W3RA6FyUUWNqiIcROetO55sY
7VTRUw1KSgbhWBl96SudX65Ys7Z849ExZrIgw83OznXiV456O8VEyeOHtocRSVoXwAbL+00OpepQ
8V3JRVF+EfU5Jf/ZcHNDdRCOxonxNsKJHNBTmcpeYJCh+rQnfu8X2+pXP6LfitgDtVV6+dnEmjqr
r6rCQsdHWgawIr8+RBOeUDpfdQvHjVP7nSUXWUWNDJU2tdzDaDIFjvDYCj3+yI5fQnkwzNE3eYrQ
8olHoKwsKvVAYsRV+d7GIhAwysCq8T6YUG856ICqnHv1nNhcU6MH42rMjitSP/1IpXO6DBPm5O4h
Bx9HuW7fjPqkf4baymX9n+PmQ5JL4zFhfbZVjTeR1fIEv/mKEYFOH58SGEar6sTw3hL43mVQfZ1X
XYW05wRVAh8hiRgBW0Rv6Fcss+Hno+4XxcBYO92G7BXvJtZUQIZ8noEbCx8KNcdfcgDep7oVMR4D
br7aofTqpmj03UrmJDrSNSBZmeG8yRnin+29sZy0w7uFRO7+cNijOXE7rOFskFK7zH0mCX5CJfp2
ssNMSl/2i4MVzPDd6Y3J4rWzyVFkLehMUUN86MU7DKrojm6tYRRqaOUOJHd505mwg49bW5voI30p
hsswfIVR4hhQjbP9jkhEpzmxb6PXxulyNoGdYzIsgkIK8EHOtiD58mJvP4QKqTrSD8CaYkITNcMK
sRbj/cZQChgvHGillhlqWLuRukIHquZcW7zsMJzqc+j8odszC0UMLboOFjaoQCCxAsE0Xja47SV8
XRKEGywsVm5REgKewmf7jU8gITVcUZQsxj4OatvhBOsCDocSYG+9QIFG8Eq8+C6zpY3yVu+NupIv
iLBOVZvXCp54TywV6bbOuTWvfy+YazO4UmQ2353BjA7j5pnAIoM9Bf7C6pb9txHdFKdWvVKsVTJi
So2EyolTb2YVbji1US6AsWJxrs2tz9XnfGqntdsCvvEqsn2bgtu9DENgWmXXHW0hTb0EVT+6VUJ8
BqaH5noweTw9sv2Up9pYnRctp5jRibGsJG+Boy03Xya3urjs2OKUIuvPFkUc+/C14AaeI5gd+Tvw
Q7lh/whOFmv/hWI450PMv37NqGLoUgyZkRSBsKx6O0+uuOYaPNL8i0Tktd1k5eEjm5E6OKrHUFhr
N3ZQwaT1r+XGhktFy498i5URHOWbp1Yk0H8uDE127tODXbBuUsCaBiC3X8R06Q6o7YGnpR1UlzDs
42EEoMhpxeZZE+wRF+k6sfEW9OuTsfaFN+nVoVgJYuuk37lhmZCtKLVgLiIaDu8SiahMoo8JPx6Q
YlOHv0W+iUSImud2snuXBN/TXq4qpP7E2QGkkUace526zke3M9FQMacm9ge3hmZyYZp5xh9irdc8
IJNypfbzxCfrKONM8IGvjjcvy77A6TosMPGV9RoPRGBleTjdIrWbCkSyPfg7qoISUY60hKbYtcW5
+ebjJiskQ7ep5eu0Nql1zC49Itp7otPyYLXyZlxz9s4KRzIYaDlmkY6A9PN2FJBMGGPsjLaZfMXL
UHnrs8mx4zXWvmhWN626DbdLifXcyciZU1ckBxNaajbLZcXs5036xRzfUI1UY5P8qc15DxReujr3
AcsJH3rbz1GV7cdmRJKlPPAz1+lkM5ptZcrHrGNoKs0dCGqpRUkerisaX+SDujoMXDeExZZp0vv4
/YgrSuoHJsaMklYxPDa5mvB57yD0k3xKqRk/lYabF5bYbSluoP54uz2ZH3rBqFcBuERS/fj/GqwZ
9IuaFaRcM/3lcj6RsS/9zOTsgP99hA2MHxOuCc9kUcOa5U0GMIcWFJTZRWm704wtS6f0/pyBwSNf
vLPPn/XN8dTr8TC9T61G8kcVRZeKA35Jf4U5H17gOW4nOWBQv+7Qv8EEZL4sFs/1plXAzBT7ITDE
rj32upKzeKqx7ubaQEWk8G9RwB7uRAeXspjllTkhQZDJlxkEEkqUxMSnRNXvw7T4C4Rak+4ZoxHZ
D+r6ITeOtvRB8eI6rIAZG6mZHzw+1cKM1/PeKWqILJZuWYI2fjZZuQNsWmZIA7mtkTqdbmBz2ckR
w6P/Cz7DpbzoQ5w38c+xpXCFAVBlKUu9mvk19z7c3eetTDopDLyiZWApmI4O2uKZnwaMy3NPRgG3
Zjv4dNI56t6EZLDJkF3frmOQCyF42CDdc/FtOiMNPsJk5SaNRuuqGhWCtRvDHhVS+pLF6j3ouf+w
1dIvFbMBLYzoFqF5oO9spSwzzF4MZhC5dN3rRXpKu2qsph0I17Qio3hQNOq3C5BpSRi8GveIQG8w
dWxqUouZ3rGeI35/O0VpuEicCoouz1rqGBBwZ++VQrIm3g38ajdmcY3fB2Agn6tm5ghzBxcjAewB
z6n4godx+MCH5liTxio7W2oCiTtxeuCsLtQTMYMIt6jUjDIGra5FWNm7vrcZVb9HMNmne31KnwmN
UVjSvMWRB5YkEhcBtSiN+u8jsNbc0rIhqnDIe7uYM0vsFzr85bSiH+T68aTZA8aXlcheqGg5pQp7
B5Xpb9N/zdEhesZBZjhyhx8BHfyp6UZCuw9N6IX4hTZzD1J6SIx/pNSVBK+10dWA2bWVX/KbjU4E
CNtX/RPE3AdxB+J/oBat/Y5A06VwTCP5IK5zppPvWjD2qE4D87hr4M2X5rbv3sPW6wLAzog6mpHM
eoKP2FORqDrNpp/9HGj7PYYKAwgo6D5IRiKhPC1f5zPuG03rdU+DKUiF/1c7LvanF9VI6HkOzYrF
0bGUMnYkz5Qm7/hNll4J4dS1bOtZZP87OgoFPUF7wVQ1hbbLtB5vapw65qX9dzhIG4ELlTpbiVLG
xTGRy+ijw3XKwtCDm/FzU2Vhm5QSBRxm/w2YRQQwm47kKvoP/eusLEUM5USUApHTpS0okRQ3L9kM
cnG7rS/5zTNO51ljFl6eGQ1j5J4lipCveYOx3afwSDqmA3s2V9yErQ+t8Yj5C7GTbrdxNMRfKub4
ptq3AAsDeJMQQgREw4B2CVDA8lCD5ZDdWoQeeYTLr/h0KLV1WaR8HWDNw5Qpp/U3gPlsiV0wPFn+
7ci1Hv16uMbDzHlDGUCqjA8HCZXi1qhSB0e3qzHFvjgWsCzrYjg8pgIyFd/nKWPnBa4EckmmfPKL
Hvrqw5Db14/hwvwpzETDQNmfUPund4uQgyHcJtegBTIsW8NMlBEOGVfHFQFQwHI3QWgERMzBaFHV
773NjN2C1GhfMgrRnsk02Zu09SspvSdPM5zhIxYaKOKVXQjdZ8p5gD2ych/s/h+w280O0Pg250AW
By3vEAJXV9VFz2JYPL+0XVVCuBS3IQJUyNPybQF6t9poBMFoKvr+wdvxklCrEnT1G07ynkdOysYh
QhRp9Hmrz7vqNLamTn3kfcySB71Hn69R6rJUcG89KZZfdDs0/WbAoyOZZk/zkEsAkhpxNeqOv37G
dLjphWPUZ6fD46K9zrw3lOUiGenpg6llXGM4LrwwSwvJdtHzn/bdaEV9VbjnQPmiY995d7JbZgBu
U7Mi79R5hnTJ1lj7D1+rnLvEl+KnOZsAiJlUwDA6VOWpadvk+Hx6c9xjoqY4aTplCmSq0PAMZ8L4
VBXwRg+5nUnNgMX6xRFH2mqZpkBlypo0bdd8+KTnwjax+3G3sGAa6rFeK/tXHFbnv+xotKoLai5P
A9wS7iH2txU0E2UtUiHwGXOAFA4TNYF8HFddkVfHBJvZNBJnTkfqq0/AxOEbItKcujUrdN5sIy+k
RnMY96dpBB5d0hviRxKMMT60xcDL+eQO/YSG0KprmocLwjj0LlfkFwuzGdGJEwhxC/dhQQi8Aagz
V6OmO/YcoBhoDnIp82xLJO1eLBqMg6wOg8ZL5+BL+Xu/4Idr282xwg95wUlZyxpV/GkoomJt/k1J
DzBClROtGM2u0rAIi/H9Gj+cz8SJtx4YDX3XNTyWyiui9Ss2AU2CSMsxpdLzjEHDr9F0BsXmqDWY
jIhcJ2iVfLHbC2Hm4fv49w9rvONYyfJyWPxNfta3+nP1YRGSJLPe1ljjkouodxRV7efEjOeUOv0e
ECW1D7paQ33aJ6lRUbdt+E+CDCINWSUMaOLAbLiFXEjHGAVodpZEfrHe7C2TuahrUIbQvkTQ72D7
sesCV83BL0GuBb01+c+cjCkBUzUn1m+7z2A/XtvrP2opNE3LtW4By6ADixpsi2eTaqeHG09rLUTp
1urrjwMb03rd1yf3FGCOzd6CVfWFDZISfvoxDw9vaRk8TmV2+YUJFm2+MVlaMln46td1a2JaYZZl
1ZIF+xhRQaRPIJvOsDhaEKNxh08s3yp8Xu8p4h6CTJ9RV1gjqNyD/Q9SKeKCPnb/cHjqn+o7xrn0
J3bnJ8xwgt4Iyr4GsUhr5mRI5MUOuMV/WxhZPm8Vh0NCbhGHzRt/tKtIsgqW4JLEV+nXMIhkBa78
za9rEDbQAOsT+ZCNEm+ZYqdHBzSPkbI4u55G+m9nqbJWKsxOM7c+sAmbfVpsSiS6GdMlIXhYT4lS
ykTQ2yP+v9Tqp4yAWuwFDyZx+oPQGnZ0Uk3LLuqVuy7KVtFrcjeDeSibaOEsVLc6f2G+6g/gdNLB
duZNRMUkTKdi3qeEbFpXOF7Uegy+s7q6F6tu229ct7GtIBc68BO5+eFQ3i8nVJnYrBsO+qLjfFNG
nWpLmKb5mNyMgsQht0d9cdb6O3Q1cM6jGEj2f9N9xWokQQiF7TdSnliuQp1HKWpqmSPSaCCgQrWU
SHbWpxKnGVO3aWqLdQuVYrVqeJusdnAwqorOR0MZcR/lyjiJcLcFGBQu4XzDu4WLMjvcfBwWTISc
pDXvV4Z/13pCDGWiNlweOSAJ4MzWRjqAW+lLGOQMpRNq2WbTMddvUHmUJDjeJ9JlBvn1IcS+XdFP
uvmwFyoxojSgzh/jsHOBrJgxA28XOfFtQ6uJ/dcrchtXqXqe7kZHPwluWFgQKy5iZj0L3eQecER2
pzr2M/NFOXXAYtnSoSVlb9/JnRc5FDvueB9ejhVM4xP1tV32uZQ2O4PjKtIMvC+Sb1lWnbPNEhx0
etpcwGHuFYyP6w7Sbsf7JUg2CQE1wHcx5r5ls988btcKMubQCDOvKaX5od2BkG+cCS1nklQiPm7l
FQh1EA6CYkG+tmAl+I0QA5D6+LAFWY4Dy8x5kJXjmkMT37vGPY1okpF4jaV/hDuOar5YZ97dBybZ
1k7+YC8Q5N1M8J+rzUSbl7T2TcZcCnnN8EekM1ZfUNbuhB/3FzqycnTY66fLbqcR54RfkQg1duab
k0xUP5M8VRIXBYG4g9LVb5qPKcNQXih6Y7FG5djMC6mqCTZhuykaeNb3WMTdX4lORACMRHSYwGTA
tLnAzkUC3sZJZV6KXJkWUOv6TJIcO6ftsC8o6vFXdRyGtsPdR1hSPDVWVOysJp8+5oyTyM/3I2+W
4u2j2ViUkrXt+vhzP7DoY0r4jghdlBidwzFjJQ+xx5tf60gA35Rqrgm3GukZ584nU3APHgaGTqxL
PZGgHQKckXAs0xg22yqqUXnlVQGtOfSoCT/sdh7uee1u9PGnoCJcukol8jEXPviDyQxJ7wjGqINQ
XkYYjLAtcNLekbTi1xeOTBmYSHfZAduxFaz3iM6yKq9hgxhUs2V8vrPjBAcaa6tL+vNSOXU3hJLZ
6tulUrGqbt3v38nlawuZhMsAmBo36NxN/7uTT1JMKoEzj1l5RTHC9aQGwIvrK/oPYvKxA7lFNik4
h+1jnmNWaYOiMFc9ZylY3F8/xePKiMveDNeRHj3icHZodUQz9p8adAui5nIyFfQG7fznPspBY4IH
D2n0Vt4EkATU42CR+nZf8VoWoHbJ9E/NGrFMsRdBTlM2OB5P8Qt/QTleKZH2MLIC8p6UnJ6UM9JC
VNUttpVxO0s+48w8+KQPPTOcdMr/MvN5YltNl9dVUkHJudhJUCZOdPJjse5qMA5HDsf8WFh/1q03
nMjYbGu3KJl3OKYQNZGIiBkbWj26hO/SvDhkHEiN+BRCmvzSNop7jf/A0/Co5fYUmdRE0v5e1Pxh
gKn9bylW1mVazmB23BkeSu6PHSw69lQC5yBFOZBmUEXef3RxjqbdilKxqbM3ai+hH5pPR/SU3cGl
fkzTXXEPnttLqhcAMNzuW+r5EuGvunTtepjGDpdOt8dTuBDH1sGPquzSIZLvtVnpe9boe19eVW48
aVfsDYFOUElh5EdTad2o3Vw+y3NmkSt8RbvD2028Kvj+UsddpGWa7TRhgwCB1HmPyvoBj+xp8c6k
HrZaoKgCBB/PsyhrurLw+H4fVcDqa9I5nC4O7gScthh5bf+YhsycbbMmXsWIwQsp2lKZPsVtG4mP
KeST98w+kHamjIf8AD8tKo8jRkZCZxdjTIBIwKF13HyX0CYkAh/Ngt92WYRdwii9nJXI8SbhGKO6
HLAoobh/LZHF3Rl+Jp4yvDL+paUzMWdUP/NRkzDA0Tig3lqvhmDC2EHh7x7odPzWnYB2P9kXh1kH
TMUT8vV0/EjYzXMhD3CEkEXXfjbBA2OpO0IN3RYv+HiR/PATsB/2qK44+UMHyz/XmGimK8AcUfHy
CC94aLbBLCHegxcoXlzqCtnKJ6Hx33nc6buDG6QQPUXy0LcgHRfoPDoB0G1TcOAHjHMmBsyVqd8m
L52hvtLfUO4POTR3FyfU+NDLyrb88GAOpfym4NHzyPgdSL3lmk/7xq9dAPI665p3Z+CyOU48SKl+
XRkrVCCD8XBm60DxTmEAmL7YptfnvLUrBC7eYdCZLjGABs2y95vsJ0rC+WLusd+R/PX2keNlUBQy
WtkOvizKDqRc2Xq3n68N8vedr5ezwxsU9kvJnoSigU9ThIe3cLlbmcNwvVNwL3oaQkStXGqR8/Mc
aAwUk6j37yFiso/zAZSbIDWc/YXHlQqGtrv2O6rXZi04q8FJ8/gnOwHuQ97bP6rBO8jvBex3wRU3
5ePMVMl6LP/ulTWTla3oWQzqSchnelMwZFPPvwLZhGDzdC33fYbYmsYi8ZLLtDe5HLYX/hjc67Kx
sfYkjUoE10w6YIwzX1N5Rg2CEI1J94iKeH8BRkxgU5/iz2v7vLeDegMbYYPa3FlqM7ztctUh7g0r
npCkQI/zA8eikOF5SlkvTEIPi3xwdC930cw2muB3pS0xtxC7RT4dvIcEz3ozM2juSw4WA5+pkCus
pBc2WLNcf6ZeNsaTpBzwLZpSVzIZcPZ6ujYiDcKRaetbEv7R0yrFfz2abFk0ZCglZ8EpwgG34b1O
kF2Xt5h1RMAKZtNzBoWGxeM2bKPzZIemKSyPhzxp/N8j7gp081Ua4NgNZAnjbhv8a9hI6rDjcbTa
AYaw40I0LsniZSh1IKGWz7oGXwHsbnDwmSAb16SuB2V0eco3JNFNtauZG0o8vy4KGax5wsT1iMJ6
YTV5F9oJn3SxgGpp6QV9kouOyiVNa/aEW4OEuHeX87zumnfttAY+Yqp+fPTnLWJTu/Xh40NVHC81
v4TDUkHMm7dJQejkn6n/48p5SGVYj9gmikGXiABHvUCQaN3JtUf/4VxfgpuMPNwwJDhbXxn0ErTC
cKW3nbCU+rEn23af7baErmp8qGsmvz3LcJXwgHgVML6oMX6m/FeeYgzQF/86JxltSS7eKlwwxFgv
6staAP6UEQjMcOEWTSpm2OYTMZ4sCf8j7FjyDDj4P33cvQCEgoiyA4gY2LAxjzoyTjzPUB6OuRJ/
ALK+hwn+MzDmiNV1uaUlX9Ip+PzP4br2r3PmuTk5mGt0DPpBZpOwM3M3SB+cMS332UscQ2jsEKGW
KRncHnHF9NhTjjvDjDCSlS/px9C4C/7DJkV0JR/fDa+sYS4tmP1UD3VWMxLcz3Lw6eqmHRvzfVIp
Yo8T6Mo9YBFHZrqWnapFi0RT5Fj8In2d43PgZp1PM3s14nGFSo2L1nsLv+FeOmJBbADWImM43zJu
u8POgXG7S2XuvuCgI4Mp92uFwprc5gpBaZwz872ivAPLia79QgV0gZWwAHmKo71cMOqquEPZ9OER
qh1U/tc+C99nOqcXyWSNWvBknFDc1XfRSa0kDeBDam65dHXK6FTs01z1y7RKxGv8bthTIdOf3sPf
GkVUaxzjkdfcf2kN2GZRaeELKpENnZgZd4xr3XMe9YdlGMv620SU7kGenA5A8x9xk5UVz7euXK9J
VhGFJQd985k0neJeCcY+GP98QtnWBYbDEY7H6T7jAt7tzoh/JhYgmSsGLpJ5Tnvb7bMzMSkGZNpS
FVc3yyhYQDxdOkrGSjU6ALh6TuRN6eJqpsvmif3lN+Tdc6OZBnvbKj5ICHs0zccj/2Q2v6Iz7upU
d0I56Pqr6+nCcl+/r1axxn8GBcjMWXuZ543Ha0oK+JbhRzm4uGnu2x8w0mROdkBWhVbVNgSOJoY5
VK7Zi56zyXxtLUaqMy4f49WDWcSjbweyOhFY8cY5dhDyCl0UnekvlihVnzCJCPvnFMV9ISxK2bxK
NaVRqSdYg5NkXlja+LlRdI3cfiQhWQLi5e6iYfR6RhLJ5H8A00ckSofU1y54F9t7LGVqbyv8MnBm
Jq08P8+OmjQufHGzxzoe5vKJU+5nNu3sk6h6Y/dOiexdSGtvMZ4v0tO7pag61dtr5iizR1A6Zj97
Y2Vwq8tjL/gmTane1hKMgCRkgR2OVQpeQMoCfITBE2LSM1iqdr830+cdcxY+zLg+0Zfh3hO4pO2C
n9AyxwaiqqF6I1q50kpRtsx7LvF1tdcGUTwWYBQIVIRdviFtH0MJaUOteJcOl5Sl1rBP8wIVVY0C
E1pOcTRMV0L7bhqhE3jCuVcHkuQ2442fE6XMj3fN3YakEQHP6hpo77+S9FOcHdJAR8xBuwhJHT4T
jOZF6pJMEWXmRtES8FoaYmKsPmWIRVNUu3UZoR8X/mgTOeg19qW3zIClUEKlvm8WSo+ppTtRG/Uq
YkZqZ4un++MPjkF/qgoUlqtv/nsGhhIOsFgNRikG9+wblgw7hkxHrHRxPZDutmpnPsHA+OQoDg4F
dajYoiz7XTiWdTolvh1FZlNxYt3sA4TDs6zMZ5vNTJsLqD794rekf7GrlYIG3jdCSuWYpSwobo7V
WE1gmjI8hCfg0P4ra46FzIOFnMKoi0uGyDH8YjpERCcKccpO1YUrQf1Ozx0hd6rIVAWxl9aOaySP
rZIC2u/hxe1CxGLyKrixum6bp4iZYEVrK6NLLfVQ9H+3ZBNXwYnMfWkihj75U+k4muA8tPBMUGLx
T/XnfQEdjlX+me7VkFc4o/cBz99b92rI/Eg5hZ5w9cOEL45z3UmVJI4CT4RVhJPd73UjRwuVop9n
9jBabDqox60JkxzQKdJIdtougCXPjevzFSNqOKV9zlmX/NxcjIxQJux05zG8e5FLA0yevJl3fN19
8cBV+GoeYrTd4mF971/aUveUOhkdyIc2FI/hJsmnst778FevrbcCXwoPA1R/cfZBCHPKSiXcAMlv
vT5+VOnSOzJ0ZmhbpqZR6wXfFJ/zBHmgWUw5KturnU7OiWk5AilEtTpnENtlVRyif0+hnG8Y6Awo
o6GfQ9W3qF2k4PU1r8IoAzW8cfwLavqB6LBk2Z2gxFzpRL9QZqoHevI1yvMR5FhIpIf60iO9gGOz
TN91y80MUhsA3/coaFZkH+HhFs7RbP/Ib+J/ITbNXxYoqdTb4fEdzyS4eRrf4mtQlNCQqvpjwH+m
XbDAwWM0RyAQcoovMD/FiqzW1PKKUSQUKMkkEY2INOCNa7OJjpu31qZTRJyrOyaKPz0+hkWZfMd7
1RUk824kXo4bVqfG5iEYMaHUPhzMyFIhfDOBNcb0K6PZ9hdyb4cWzjYs55I6QQMiz4fbJfokFdL0
CPReGN5n2tCX1VBa9WZYCbWBJ5PJLpGAHnG6raGVHmXplkdLZm0CtQIw6OG5OIeuyxPt8ENk/et9
ffdtyh+aaBdykJpOgwrMTDaWTPWCxZ5l6fXMUNl+v+48SbbUc495mktKfWkoXcKVv12gyax2dE++
1s/4iO8PGjkaEzds34y/CQo6N9D1YVIA+LnFQbT47yty64z9iHHmrFv3zaRvlqxYtwppR01+pbZ7
v7iyr8TkMSzElnr3Eg4mwnu5JJxkJeGtq8uWpK4/uJ1nStyI9ZCp83aISkfd+YPDCYnT8jEfDTwv
Mlr8nMKpI/gj5GJfj2fCr24c61tQ2LoR7ojIusZRDY2Oy62oYiKtDAeLCWZiAWA5bOiH/bInkUxN
KGX2hNRmJy8ZrlLTXfOMlABtyWJwFM8IwfL9DmJXQgHU0khT6zm9av7g6r/2+uOXm8Z1nkplsajI
s7iCkK0v2bZfcrWMyLP/seAptP54dXDg82LMTb9VMQipiTB6p8Z8icEr36ipso7wL2B5RQkzcDU2
mtFZCIXAJO7vXMnYz3YhTpnINOAL434+awws1rNQ21LB4gpUpUoizx/3rx2UaHx2vmtvAoOJMIE6
xOcAqTzIO9gKLd9glhedb0v/Q4cKyMSn6xshW0ZBdRSWRyVWFQgSDrim1tcprQZ2l2cmNo7ymSip
iQt3mppaXnpve/Mx3p6mIKQ3O8uSsfhiXSYHS3eiobQLqIHq7vkJQ9TZzKGpf6YzKuehrF4OcRy0
DQ5YGwsYOOhHJIT+lEoaC4Q2r+SgxXlfCDGqWbliMcX+N2/kmN/qHiONHZ3Gmse6IdZODoZOQkbF
hg870KaAPG+jph56O16R/DT7aSTcuiCXwqkg9vk6ohYyeeqPgnwpOL3G9kS0EMMDJUcjUAwjiSMl
RUZqann1+Ox62JsONNSVZxtEDITcaeJO2/gP0dicv3b3SWMDzBTcbierkcYbFNux/R2djTnzSNAZ
YJOEzLEEaiqraWe2G6TIShxH6nsTJVx4Ol1CqHmnBuHTLuc2kVp9t5EE14jTqgIp8l4otA/R69B8
G/UyJE+uPK9XoBY+HtmiRyBlmHrTXm+ZGnCo7mYMeQnfFNuj9Uq+48ies3zTSP6TGmUQ+TU8aabT
9e3viBljnPJnZ4DYt6RkebchR2jaWQhfQTHdjfCaBnRy3+LpsjYuAbizALwMwV7nvgkMwWuf5sO6
4ZJufNymOM3Qk5Zh1zHLtl+0KZXus7UvrBBlziFMSInbdA2VknqALUwdGw4qnjQIuOeqY1iuZTeP
wDWPpkgYBNPxnkcXg9nblku4f2efEtZMCqpolu7XEDU1hUZz6kJoc3Ue0XdCHgUz2DH9gzlD9J3y
vhJ8V4W2Inaofz4aH1YvK6KuKwv3gmHp33YchXv3tB3iE169c0Q48KqKwkUMdIokHmDyoEBAoWmq
6Ru30JGaNC0GLf/b/LQHDTkeqM4rJzZB9m6Fuo+MSV5Q6eOu/JnM3CmvTkvCENkVVZhVlTMlXIdn
hs9yyxm268/v96tFosWSbitTa1wekaE1rAQg7+W5a+bWBxYA2ELeYun1jq9Bc9l66xDLpvznLIZm
XOCXnm2dn3xQrNawfo8KL/k39TJ4HSgIczJsKNlOzl/DOm62PeHcrBWurq0dDhTRBU+RpL/RP7sL
Jz4pogOiKLyESRTgXCcPyVnLMJT6NA8/El8eMsxRdwCZJbIFg8PvfHSYX+hzT7MY7eyPebge/x5P
lN2YsuDLDmbxdsoXj5jGsuBhcn3rGvqPZsL25KS33urg2fFRyTPt5qlqOaDCqnH/VDTKIvKWKCwm
7SRBwOcFCsj7YcLeN1xCVN7I9X6rNF2ena/CTw0Q+mCgVMGpW2kburmzGtAbpLpp9rgRjMqA+BDU
Wbh70PDiQURGxWvxt9rKej8h70Ej4dJR5YXaqXNnOOHBvf/X0SK+bbogOXoscfcDJxcSx5gRb7Me
iJvi39wO1r7dZokCPvG6bCyAAtuJxh/rIE0W1nhvcHDD8VTLAg7g4aakefKcIbWykLtoYG6xX0ic
ouY/cv7X59/Hl2G7/Dqjd+ypRmxVK/ysFhI9xrWB8M0f3Lbr89NuMtrccLfwayVL/hRXqsMfBAnR
/iXt2HlGrK/X/G+G1hG0e18E9sfjbL2NrLk8qV4vyQvFvJooiTp1+7E0uRQq1a/ufhYoK8C/wBM6
HnO7pvd6JiiBRbMHb047OTr2B/nw8cAYeBe5Wt6ujDF7xCsxhTpuYk9W+dZVBHcMyn1d1cZdiCGs
qbqyInZMioxBNhWTTFqiqn5P1qRBGphWkU/qUfp/ziGf5EFDYjGkkS8z0ho347213UCfg1wHBUkT
bGeMLhJB9SlYs1Rtq/oAlDkxl5gB8JOhY+zx7Am5NGfTLrtmFan7QySmY+oB7blMcSKFmN1T63xN
2p1QLTTQ/sVSxRvuSNE41NInmyYxEwvsBuN2vWvLI/kDEOgQpzTfVSrF91X9Kem3D7gDIhVER4Yv
yii0BoXIOmsQiHvqziDa/uIJ5z8vI8fz1cAGIBVM5HIVDAJF7dyuF8dnBNwGajypt83DZmN2iXx9
S4k6C6OHPykAsB8roZXwpVue5aEcPh5Wkp4y3gslu6ErOqMF9t6jJkLM4FWhhNlF+VDNAfn9y5s1
roHoAgJRDy5Yofu5qvzmWtCwXBrovqUzBKqPl/NDbk10wiK2Uu61oV+I+yu2znbMGYQ55va3cY3E
TQND89NPcTBu+CdJFuqjFv0KgMoyxWqgp/KZIdv/Dpkx0CjKjxu+e5aRBph5k0lhpjrVZM3YwK4B
C7jJJashzr8wXDOh570CqRjdF+j1enUcKeclYA+Il+Ei1jnDjvkGEmv3rE+d+elCgK7ThKhFgY0X
dX4PztnklUAzbQfpZnv367QOCk1xMAVmDweiMQwRCthApfGLq/UYJktH8fAcVfRty0zUIsLNKHB4
M4PpFy9TxH9BYqi6uhSP0HWum53AN4AbiGnahHe9fEqEDVIzP4Ksi1++EfKYbmrW+U6lwtb3ypcE
2S0I2+L0Tm0xpKYl3T+dJ6D1x+4L9IbonEVrVPhBVCtxCGJjNU3z0ojanFMl7Fi0K8YqvVFnMzq/
euIlfSi9yF23sbYGN5o/2kcJWBh+fTOgQda2HI3DzRMpukPK/Om6oD3qPAsY2RT4Dcfg+zQMS6XI
y6RqhONx8iDN9kHfv1tr4YLytj5jSB+AlIFhp82QiWEQcgjE/8SALm+aWMQtAMgETksMFaENK3z2
sIioB9yepI5SfGTGW9N9d7ynTD4xEu6XF81+q7KTLQYzTMxoiJF/L2ouaNlXiLWO5TqPS/0IvlYr
+PfL7jzFFd5lv+cOIH5gYLWKcEY2ocJWee/tA9KW8R7sLdik4iolM2qGPnX9d5WwkoiNLHbN/0pl
0TZFsGosS5AfGxeV4ybNcMEMbOAIsw5V7JB1cWv7IJKVcJDiWS2Gy66BXilDMqLogpCyH9/JfvIU
2z9NmCN2bD05DlQrgoJgToTmEREpYUCktw5XdZP7Qx9D+mH2ZafirQKXR9UfiXAjVEY5jZVLoTi5
o+4h/9wh9n0mGDPv5BCZxDdCVr09O0hjCyUg5sF7aljyOfUBg2QgxdvJNMAN5kxnP0f3yrQiwElV
rXXHChD0qgv5TtgmhOo1n4pZ9sYNR5A/iNQw6EreU6sQQPnhkujmzqYK0gruzgAgIGLHua+SAJK4
3ugdEUNV8Ts4EZAKmAkr2odvrRY1zHw5Tmk10S0wDqq7Z8YV0i8m698RN5+ld7Zgj41kXeR2PgTf
6r7M65PajCzvvBa+3yG6RtlcsS0cu4KW4HTWF/YRinjUz00CNsoaDJcroqegDgzQ1TSNyjSc7bMo
mEh3VdZlp6waTupIb3CNSNj0YAb61Uu+khYuzYsfBl2m5lX8kzWmvC+K7q/AYoFPMTYAWyZK8Wtq
/2xlxNRpmbRNIIeyIItko2xb5su6lM+E5jjwOXJD2+F7VzU7N9rCYY/pG7BuHveoz2CqyDek+klH
d4cfJNCrX/vMnboNEHVMAFJ4TiWXruDU6Q7oLv+irkYCv/5XvyTaqOPTCqg9IpjUA+hxrL17KHS/
0aFgKj1vUJ/ka90uK52x+EL3ac4zA2+rVX53udcsN6TMvpGWKXpaPZpXd2oGtrcOKB54bgoE+KGH
+0WDk7BigemaEVBqZZUtKkK5XKBHj3RrWAjfalaY+zGDF1AlaqBcPgIZigH8wqK93BjBwxdrPJJd
8z30m+DVn/z4Ns4AZuJ1lgEVYZH6uv8FkVDnlDZR610X2Rvy8w9LRS5HHUAqbaGzZx1zOYDSWFMR
WLaRvyBxkbgdHFCEjyx3sD1jB11Uu/oDlbBSuQsFGGBium0FDLQ3Z5R2Nd8oMxqnccDMPGzCH8pX
iqff2HjWp0/XgReu3GO1+EIhGnm5LvyJF9E7w37GGE8xFKGkrJasYj3S0CnPqZX0TTXC6XbeyViH
zNCpIOPQfIg9kEIu4/CkumLRos8v9Z7jIXjyrPyJXQ6s3/xk6rYlRSa6o2OEw/Rs23pO57xJffXV
8Y+8aRc41ODr4344IZ2gSKYVx5qOhLxC9hgeZOor7NkFRloep96PN0DY5eX56LBMF3LAJg/u45zn
FiTRnFymQ8n+f5aLaollMMlSUVDQPNb8FoSa2tndUUvhhn3R4llaUu2no+dEET/y3MQjX3+e1t3Z
3EmVU1l2oSku0bxDTrJXxlF9BztswrIePpQD/dqDaHUnkL4c3wVRUuN1JbcqbkKZG/yC8IP+pC+q
/4Pe8aXZTEHmErg5wbr+ucNYUD0Fcx6yV47PvG8yvama5dbENIlpNBFuCetnj7m5EHiMsAmyWGkP
NQ2JUq15HIRX6xMMLQhzSv4wdLh4cxQChFlrU3TcKBcANWHFJkBzWfiHqo4bqXSd4TBFnQ/qbJZf
VlqGM3SoVI+vUXuf+Rq+NO0PL3zoMmaovcarTecz8kLThCBl3E3pFXRP3lA92l2yxKLZD3gawoT/
WgA0orQcSbaCHloDRi81FahIy6PAsHvv8NfF68g/+DWjIWPJjjMK+42qix+14Hu5+/9rf0gn+if2
OB/PKLfhSagZ6brgltLl13Hyp+tk5njvC/3f8vLtthj67kSW4CEG4w7V5qASz9uDNmgUvmd+ZpwN
HM8uFrL2dmTUVigiCgJR6Jr+6lMrWcVGvDTNsRNo4YB5ZXY+5zz8RbswW2tWSq4YlJuMSGWCnu62
ZEBqCahWQbh4gUTUXqtRWyBPL7Rvcnkcwl+LZLSLCzn7Ib5gc8/fyqCbNTwr4D7oL/g2GeacEbc7
nsIvU3BVsIcTrHv8VvHTEDvoxnHZD8erwMFbCxZVX4sX9muKUVvP+grqwx8i9+tWr8GDU4io2ifo
C5PFdsNhogBajFRWrgJ4eH6qJc74bQLxXJKnVCztSRFlev503ATR2HWGYdILf4SRETANgYUJjekl
7lgWyuI31EAnOYjxMzTN4LpFvgLQtPhWsG5acYwS9/SBSHoHI03dwdg37ZiTih9ywW5xbFqBIzAu
D+FEbd+ktzIA0lcYVxFiFClP72ew3Ksxcw1Z/Ic4Cr9Gm+vN2ySDctQc2QjQPG+/arJ+bGM8Y/gy
RrVwugGc1cU7682bHgxEbETk3VNNmFpBrC+Q2YZlAaJM2w7HopH3sF0vzyHaWxc8fha7HG6/SH52
sIe5FNeeLlb9ZpJ4/eU5+N7IxXHMWCzYZHq9iyZS8Jiw1gzzI6QXpZYOyaWm5COv9xY+2sMEaoqR
OjtkfhpZeNaMyJ9p1prhdzBnQizwD9RquTc+PzE17EDxGqi8VcsABS5r2vFozouZc9//lFQ9rqO8
h90+EX1DwzlU95XKs2leo8yvW4LtEI9EHXHkqGdxObyepYn8Fl5q0ucgxIBotB5x3S+OTQwLUzdC
OOZ+5eHGY2bP0mIeMUuOvARKDDPtuLmK3PTLdtdZWLXnXRgtQQD9gqksLti/X2BL0JexS0FJOCK2
PugBdZi8109eHSKzgALvtRdQVPVa9SdHRC2oG1GSAMd1mn4cpjkqiNdIO/5JkaVOofNPWHUvmAtK
7WRR7brLYeItdRwRIS+KmnhMnuTXH3jgAPxhhxHrCKsbZ3eGuiwTQDEnRW0Fmkn2Y8ce85MFWFZr
9F8jb4Qoo1YpmVw75DW7t71woVVf4HSJQCPZAy95n9KYF+Uz6xC3nhEg6E0lIkL5PyVE+eb52sxq
8fFEHQ0dX6ItjdxPLBauVUG4rc+4c5FsGYG3a5VPDKM8weFu3UJhTCMnd2kvqDUtklB6/tTB7uXe
iI5pSZVQGN3iPZhHLl57PGnRWNs+RLx543Nq+SrJQNVkVlyrJXaH5PJku90dBKRaJQGUI49ZHtdY
YS5S83tBJ9NyWjUHWdlHabhYbLBtfM7fxs/3rdvHlYcfLmyxC0Z9gPAgwFv6JDXhqwNcYmRsSZfe
Rn9Q9Gf0PqKxA2alBqUXd12/mb4wrF03GEeUIskvd5x0q6ccXZDsi5t95fknFhL+IlbIWesBizsF
iVllHQcRRSTJ+r1rofusO2iWjToNmlz2FUp35S+C7S1dWaJX0vWRt4ycPFmHEUAqw2SzJZhChGmY
UhnnhdqtckfVirB9o6Rm7XhxeeXzjv8G9y85Ud+GbuL2LNc4afgLPUeUYTzuiBWyVue/hm01OCL2
bcF19tHP4XTn5EPtw+1M9ra/O1TpgcXv4REgWS4I/h1RX3Xdxq/MHj/K2wGp2XFfGhzMVwSR3jNj
O05g4RDuW4l8Px+m6bgELOnmXeVoWqHCQtnrBjFYsXfPHlfaQVUp3lq18NxKmf6UdQfeN7IWaoLG
a2NwmDBGsV42Pp8PnXjBZCRTww3+JXQKdBKshvPGJ3zYursdswH62VmGGZ6eNt8ugTK0q4ajB3pm
smxTUvBcRlIkIfV74FqIVG279XtgWzk0cCJxRiMVx5NLKlRFXmIDl+DLtJ+oCLxnc+xrI2qo1nkG
+gAtiJMxMNaxZduEVlEkOt/ma0yUuOzJkmfYRxE0osDdCqaBpp+pkUpf8A8ib7WKku5SMmitgT5P
4KsL4Sb7golirnxQh1bicd5YPKEmppn6blhQhaongXNzFwesiZsGdJrusmjH7ovc6Y+0F2F+3j0w
WU+PdTI4w7hBbHET9tnJQw5O0FolEm5St5sYgXlj4NJzCBYaqcln/HOfHUglfVNhtd3a2ljIy6xZ
w9VexcLpCMQfrIocPhcOmr/vAYFzrWri0nznB+/yPc65RWun7BHSlKZzGtmPRDAW8sLPn2bNiXD7
EqqmQMXpUojNsIeemZwP1haUVxR9sNtgBSQEchGj7wD4LxS4y1Dw83RX5bXZ2inJI90kJGghAXak
wgbouVoPzFpD1/fVyc+KQW+lKuugK3EE5qfAzuegZhk9aKrEMhL35u/RgyIJrzWnTsWDsa9zvx9R
h7YXzuzG9L0/KJzwAjKBcT6aXisaSdDKdLlew/WwuRj8RjD8Tyvn+cb/hyrHPLOCQBk1T+l5RHB7
5/4g+j2KRIAmK6UoSjwKkLpWS/PXs8OQ4fMofw8numzCAhhAlYmls/nKasRFZJg+024MrTa/rKgo
9lvRNtdlVR3nA6oRZ1k3b4dWiiQA4kf8+cZyXdTI3b9buPen26a6yWR+t2VkEcL91SYrYbQX0hp7
DvYYcqsFU2xSyhmse39Ik7/NKMHJP+dy6FbXwB6LW9m7XIAppsh99oTd3uNjSEyLZmtGakhBmjrk
48RoIZdpxvFYiPrUE3yZ0JZCGnUM7ZfLQJt5/vg7B2wvWhA2DCwJhQBoW6zl0NNnmWLc6X7Tkm8b
YUuB6JXUHE16gAdLcwI8D1NNO9tqWiAhunBg3gzB8wGPY7fTPENYL/liSl8Kmjv72heBlG2yjPXr
cFuSitEp5FpH7KPpf2Hv6nmzgG0CFg4xfmRGkZD4d0SsCc1OIhMyr1+FXceVjf6LRzfTSw0Ftyhl
0vC19nGYhKTN95zzuc7rscUE/FDh8EtaXChIx1NCs8Q8an9908nie8b366OiIkRHHn1hkdSxXhCR
meZeKXv0sO9k+f3rCZhPBjN0MeCDbOiShWwRPtoFRFoZwaspiinX0ZoX8GTO8QE8DuqIffeuUmMH
RcYKLau/NXw7kMomRy5lB9vH8mLg445kIIcZyhP/5vTDeKYlIbIDB5WZKFL3pyz8vxEcv2aXQx4y
oRrCKbxT8IJ7qETUF1vL/sYD2VsKAkKHR8vOU26hTZVeE4BquUj7bz6s9L2JUE+QJb6brRYmqCyW
1+nNO17CkxKBhAiirvod1VNwxfB5DEr/sBi0STFxUfrQZXubqm6LKTi2o7pp8jrgO6TAPJlwdK1I
9WkkOPdabQSzbfcG3g8puDj/kZ4q6V6tVqhG+GXOQH42pHqILvhG1YoTQfJuZYMOBvKO4HpY5HZ3
3M248XsCHrqIhUEvdmmcjGW1/IniNAdPd2Gx31a8+0ULugvfivy2q/myB2FVSJLY+GcSXMHQLOl3
M3vgf1sDWH++9ShfxR5vNXFi8i9xFp0klSHBUVAEag4GRzFKhAWxv/rjR27LYQEv9b4gNXV2VzyO
SdrxwzFq8nwcFeC73rkrP7G5OaZTWW9yTFdWlwPp2b1ZVsHSYvcFKOj64zJaY1G2ggN86FuqDIkM
NHf1NY4lGGzMdy1oLMYOcapSkzmKF12jhTQplTjva7hdrT10aEa3yPQMYWqlQR+lAf+zuYXp+nJy
/wjTBCyqoQEfqKjPHR7sfrb1dfHnJsPuHPSABj1nxDCm5IHmK3DOhqdBsijX+akPk6dFaRRCnjkF
TCIq16qDc3gNHSKfTpwQQMF4LqNthaHfCg0uXMLM0tjy/M33QRdno4oR4vdBHy5rpwXc94hczJEt
ibtjA842kzTM2iOz3Z4o5uV1WyGDhXeAmimB7nCTSde4tnwLZCAbFZZUiQKy307750FIH0+XW9qz
1raa+5RrjG0XcBOo81cy8CpJrKXdOysdSvxG3MLB7SBFF09dHiW6iW4HPw0J6rhEkknx8urSL7cT
lEqMv9R8BG/4ZTFdIyX/DvS9vG8Eqv7Qo+zmT1wgWUxrVXnlht6h5CRT6IzeKHPFyefilbE2kHbN
kliZt7qGCjqqg875J5uDn9OnsNw3p3HTU/VW8Huf2mpZeQ/u9uCMg+O7J2GssWn9jnSuE0zC5Duj
BOBf6LBoNacM8zTbTzefRnsf+lu2rlBpbMCqwnHXDpvannl34/phGIjaktkWzabalwEOs0sjo8Tr
ugQjQVuiJcbkNWQbo5u/UM9VpbLObo+oSO+dxFCBufq+xXk67UbDFnK9FfPMLwrjIrOiINCgCHg5
xJ9ZyevAqy2JAn5yuiBcVqOdbyDBm8tu+rZnv2vV1AzYhVSR870YWnNLXphGhDi4zLAoJnhW17ZN
A8O1egla8mUxWWVN/VO/G19jCnvcqhCV2j6/zMlXc6VuGDSu7Hq4DYZodCoIib/Defx4HPGxUtC9
i405s07pgtyy+w4dIbpaCIBF0zJcqJvHgxZb/3TCe+glWYkHY2iEbY6MBHyvla82S7cWs5eOfD5K
84bjmbXYFBo+Nu1M3U97inbjkJUroakmKceqZ821UgC9EsljihwscXbeRkARoPCKSqXXKd2WK4kv
T1FGfHGmdGDE1zaBPSSSR70GeF43CC75MhiccJsz5U1LdACl4WcM+BQPAWzmPnvbNbQZ6MvCCE7j
aDqNYukdpvvZ71yVgvMZAbjGfA/dZwEqSBS+coQRUKhjYh5CvjaPSp0Eo6nmIcIcdSgxlTOGRsQA
uvHSBXkgWjzX3a1TbE+J3oztforVdCp++RXpBDp7rWDuaHaoPZIhR9cW4HJue6IHLAeAsr+omOc4
O/85iFuNRsKHwvVSdKkDkJ8BQ4kLyB3V+RRPQgK4bFWYF1xVYBWoxZljktp2FdnnwFGKRvj6VOnI
s3gGiQKOxUEpBSSuo3grQrb5cv970+sbI0EGIULDWFK6DKr1bFF0GigwgnncnUiZJHWftaAQtwAA
Rbi/QMuXX7I7cvEt+feJm7li7IhloWCX/DhdYXtbTPa4Km04I+VanFM9ziwukg+MWxAC25UEXDIX
5BqnMaKcAy7hY0mWjVAIHuBQnbADrpiGN34BSFpRnmjJpvl75gW8/lil9G2ViXuUhqkzjBDM59fN
IpJFhegxerH7N53nvkA6/esHMCYu/3H9haOwBltJXNp+PeBVVhSqCFJQbtdSACgoBgeGiFdk5WaC
sP9y0Wx6uQbgbSxkzMCQXiFwHCm0i/e9Dst4CaibuE1TWX59kzGwm3REzsItb83n1Qa1dkStbCYU
8NEIuMs+bOksRM15Wd/v9+1FVtAXyq0YMSMCc9l5vb2VrX5+pE9iTRXWbOSBfFCCkCzRM8vkSFCY
sfxHTyD7kWbVxRKtliLk3snl4QqBQtyTVGyNzwOn1uDHFN6JlFO2oZcgdvzyq+/6dI3AFSxhq2zE
RV5HeBz1gYo4I1LP4fVCMiqA3CU1yjShFSAmS8rhAz/GWE+u31pNPuyanTRFDe3CQKqkHob9OLQY
O8nbO5af5shIcu/xXIjC7ys8veQU80BeNE+ByZova5sgTegg7HIzf6HfZJUhNKax8Dl1m6/+pswH
WpA5BqQ2C8mswb38a65o0awWuU/G4GerfWpBqxkzdderfztz62+c9++uPVylwcQeqAQ0CvV0gyHj
p6lHkArtYx+niK4HPDI6btmL5z24PJEn2cxkZcym0WtUsTrbcqfHXPHISiY4c+eBl2R4CXot9zHT
pBA147sD1yNAZSsojGeLw2zj6DqxPtN/tt34xHRDjwkxYiHjZBn2Whji4wtv/NhSuSP3GjyUGuMw
geXNG3BVohCym31fNpW+FzSh0wbk83Qki59ZGu4cCqB6vGl/iZkN58ztSLHP4quLx5HJ2kWG1Ulk
CHi6PQ75/aP+jMp4ivxoDE5+TLn19AyMQ8xU/oSBbb9tdEd8TOadBRavAvWR1ZMhAtF7u7Q3XANP
XPTNl93tEHr3wcf2rt4C0xq/EEfOrvT0ENHU7flUI9Zq5zpHKi6DdeUxFN27w+hfI9UiMuxnhe4k
HVSLt62potYklkAiuVVXwysaakV8tpAAOyq/pqNDtweBQxwxvJygjHOnKOiVGRdfyGl1rHiozh2n
4Ahpit8LHhOFIBadhK4TjrQSAGQAvxbE3+f8W21ZoEXec3/equ0h4bElwVXOucw3uQUGTfPnYfRs
yNnzSX+QCYXG0stg3bCBb5QpNd8GSFSABUust/itsOzk2NhYrFb45GaSLYjSu0hgC+pkBd2mQJN/
cNkNdilwlfFH3Pb7iLXzQ7/Nbr4atJbASv0dK3pHzr4j/DkVIon3cMxQrDwCqPd1OJ3rR3pc+Yyn
IpSLOdaJWq+YNH546AzQfLKWbJ0XHbQ//s9WxbOEuMhZbk567yZQZV6x7BPEUu2P8WrkstFG0+om
ZP1EVM+dWx3vVK1zlw5gyXWBnjCH6DAFm0sowveu0ni85HN6yBRoRYYMyvzBR57dy31ksdYdz9Dv
hXeB9khOXaj2YlzsLNr5hyw/uAwu1Ygr6N9HzcZCzeJCUpMKGqAZvz8w9GzCEMqChjzFol2btOf6
UHfh4/P0Qzqu4+AY608+Kg88ikH0gz0edJRxcPukldZG1kTyQFcOE6MTuI6IgPm646vP0vYFjmWX
F4DGIebbA/GmhSFY+3OTPP+HiyI8YaNgMWVk3PlwzoxmGFhARIB2GFSR7se5zjEJTP9n3ExGmLF5
VuRH6HFD1CBO+RiwkQI4qbardsgY+ubWDhy9WRZW50V+4okxUtYEObA7jqfMSFBQBzhQGkhHo4W2
PKIPM/3oriAYM6xpNXX+2+Hmet4CZJv0Hhooe591kK+7YrVvVjVSkxkJ2Mi+uXDHx1PVM0haS4BZ
lL/A3EWGl6NeSMdaLUxe/vtyG7lYJAQ5yL5LGRLDEmnwUilbFuoe9jBSGVbfBbaKiEkzwazD8035
MiwQCsdwmiBb4w7DJmKiBHOCheVLSVcRcxjct/pBBJwUZh3b2QCvA9vujhEbckzUOJH63U6QxG9q
kbquwG+TkEIqBVc80bSilGi4z6jGS/BYDFj04o347y1oC6YbeweeFkK5zCwl+AUFSt2ildYrUPmw
0ddWFInwvgJJC3Uqfehr9Gn9SdxOfXPn12Hnw7mOWmPwkACGTzhp9vy23k2h89gL4WZDwGrv8/+I
F4pzITunrSA+bfY7daK0BiWApP3p3VFTb/A3TKn+KFcq/oI6arvu17G/lDhdz/QBjU66//tuMGJy
QxH0GIj8gM9tI5NQrWMFsos5K45RQjeesCkgSEzD7gEix7wZVQ4QCSjneVVEp9DBk5JzD3rESs/w
2R6LrWp03Fj23w49ve69N4mq6pYfcAkrMmTkIefcXXpchduYyxS0t0etlo0mJnLOmD9VcW/ICKRH
4ajaNRYrf1J86OqJm2BRCZkqG/w/yhg4dO0s/URS3gv0gl/9dsH7CI4He4Q4EtFwtszMI+S/eDd2
NKeXXpUlON4e6OB9zdSdaD+VR48aGcCFCxLMWP3bJjDc6bL0NMCGq7J2SxmzmC+xFwzOPuzQQb9I
0+jcjTTUeXcGGF85yUEaSUgPYdQr168ELfZK9pRFZQBt4ASzkzf2JGv5phYJQaBuBhBtQCdPtsP5
/ToJzBqf+gQMvRd584E3J7OkOj2+TCAmGGCOJyIayNFNVNkcjLCFS5t8BvGUDSWex2uDG6mfp/w0
E/dy9D+y8dDr97en/VzkxjmXGJoqpCjShxglGXXOn4RnF67alisBua56xIJtkazCBTKYo6Z7TfxD
7OR1ridWxPSe2N3Yt3AeXmlAiQLzG4LFOZfVhmOzloSp1ZJrrXsx15GFJ+0/p+wQD5EqnGKnKbmH
M5MJPNC6M3+bVLglUvdl06CsbAuUNDTFvYR7QyY2p2IzqzGB3KtS7IdlOD4/1Qhg3NpjGD6adorp
cjJP7qeJq8Feg53fQYcq2rb21WmhKOJTZ086ClpHfL1kFHi/0Oa4MWnY09DgSTHNxTTsuZuKYKK4
awqSKsS46kz0gVZBZJRIkkXZ9EJepon/tC4+OUVtfuhLVaBcwvSObISkrX2HUCFVTtc0FQ5LaCbt
M8mhcxp1UrjxJbb7BrQT10DSIKQOCJ38vi1Lml2YKQbEHG8WswN2yCtHhCe+vOsdEoyjsE5loiD/
W6BIKGSmiUH5zlZoA6x9nXt8jUiwil4wca/PQ4+GpJR7mL2H7cm9Ty2td6+0Dhb4QWOJ3HgI9Ffe
J8MGbNThrXVxYTB/DdcjrYbPK3VK251f1U4BsWucqsQexB/a7eM0y+gr2T/k0EeE8Ep+oSjHz0gR
qMNkWOfwXwYytfGIBG9dUIz0m5IOoTP+Netq/mgaZeNXjLPsyOKjVpZJQyf5YcQILfA2WpJ3GoaR
7tzE3iYlKe92Vjud/c2OCIPlQjF9Nj0j4plCVwWJ1qcgrsXvgz60zCrZkyRu9Copp4Wv1cP4sfZV
EmPXR5IHkXNReh75tz22Hacc5p3OA/1fEYRZBwDFM5p9AHg1EOuufRM+J/9TKikmPHIsQ57znuNg
ON8/q4X4T/S9rBoz3GL/tIEC78JJnF489pGN32q3TyCzEUFfzOPW/Ui7oPfFbqylnQ3P5S8D2arK
R4qAA7jKBWAXdB1eqQ3XNJ14Z2bx/V4od3RJVVR/bYSKehH1IxyjfK+43OhTVOhiEu3CsteZ9ery
HDhcX2LWdfVaAOxwrCoDpdPar5cd0OQIxEpw/qrlMgtb7Ne5/i5XHFDkhiyK3Dp1zwASuMDanRcX
CMu+HQQG+W/DGlP4UUYL5Pf5fRpwQqcufq6hEbP/pwLQZLhPJc+6RactZipOSkc005pFS8Vn/rG/
DjljCt0EzljgNoNZjxGruQTsTR9DVk4/okQHl4vF+1iuFDW49UDgDfbdthk7xVPNn4ilCfl4rIxH
N7RrPx3erCLE6rOeDv4B/rthx/8JTWdOztRuAlTPjcizNRco0wMGGZ0YADa+K++cqLyNuxqfEB8C
JsR389LBC2+66w89P86RdABCcUdNSEhHXLBfX7kah/C3oOsvWxNdSDA0dEW83aUa4SqtDp9vvTxn
XBmTWPm3Dp2ogHKTZE3afB1UDvON6HtlPz62EAwudPzr73yhdBAZ9bSJ9XKvQ6IBhhS4VnWj1EQC
MjSkcM9mDJYMN1A4eLNOUMcLGb3uawL2Tgnm7GFlLomaF0RQ00ch67msX4YIFRXimd2g/uZObn8p
rIQ06rC8EggqX7OD0Kmel2X/5wFQVM4x4DbRBa6wAlXp/68uXNh7AtyykIJJfSCBbvgGo8CE1nLj
hJp+WCAM+4A44+qpEnn6NUbs5SZruA+yZo3xw+GKhFDPIZSM6tmTlBdLsVvMAKnT6Z79nahmIkSI
FFPMphGjb9fj1eBTE2DDk/MpgbKAB2VO+i+LXg8rFvYCz8V0c6LaFtvgL4tF+Swe3vj25Shpvjgy
RleiitS/ahxK82eRvPJe0NsPSlvjiH6eCjIVSuZh6NSegyi18mrPVyrQClS0O78WpwYVeaL0Bo5o
Hq93RNgvhegsJxKggYvSZRM2YAjdgeMV1/xYJZUV5+Uiy3ljwh+OU1fFMT0KBCdugLMSJKQniui0
kwrhuD28G7XmkGnzvRSJ4RzTxMT0pltlFRqk4ImQb1ETL+wKaDLYhewBhj4tvrGoVkSIfwNwrKGq
7nWtcYJnkSduVtSvhIdRF0hHSoCMOTOEx+Rc2IZnEitlps8wXgdSYLpXPK+GJxYOY2xfTVCqowNB
iVyqVbZ4OeRtrsGF0hMuy8hMlFOt632XJdCtWORu4GwB1VnqYLMZ5iB7sB85uN+ft4OsELG5zT3E
sPG09OxT2I8vMW/8qeiaiEXuFVlrHGFczQJWtv1oSvZ++/T7cwOuw6yQMFb+LX3i13EszRbMFc+O
+uicwOPXtMsHBodEidkcDAMxP2N5qpJhnYiTHzJdiGQ5OzrNL1cVh12rxxrXhRjx1V3hUmbUddGE
vxRQEYpZsWcCaw3yeJSwxxhlu8QMMRtu9pp3lepphIqptTSVSVj3ihu5jaQyJYwrdiIVkxO3HDVq
LdRc6Tx+1S/puyxqAfvcpEYlX1er4r31VFAlS9ociPt8F/Of6YvAaLpSJHQyE8yH4jqBcFkwQ5FY
fHtdu9ignTukVbFqA0q1SPbY2uL5LKwz4KL1Wg6CZyztJzgQtBWxZeXhTiChm6fcRU8v+BKjsMVs
JgO2fbSU31TABjCITJh9BIpVChXdfHybXUikmXLlWRuerxdw5JyUzYCo+cu1yKWYmePSDD1v10cM
Hu/fCE31kT1YPjGRZVblzHwluregTwah+azP75wfU8JfvdvBR4n0Gev3zTYxFQhs2xdZJPbkpai1
2s3OXy1YoCFUtX7EyKnJUNMcgUtbHOKNldV7HPHc/WMbPYNYvSBlS8WsLckI2Jt9ek4geiPc65Tz
yDulyYiE8T4rXQWdkv+COepS4V90qG/rdBtZvSSsjC/7HFL/Z2ukhdR6RnmpGrAPVmC9cQTyO80F
iNQ246cU3JiV5kn3ex7r8RUp2YK5y+mq8Y/HVpjfqHJwwFZ4wLfWRe1IiueHsaGJRtMykGat6Sw1
QciHfgyx1V24jfJ/e12lzz89uODGG9nHi4DQGo3vT1L7C5KU0DvCI0vU5u/3NUMIezXZBf4U3Ll8
UgKskeHSQplv2ED2DP26abdKQKc27/CVEuE3NAW9gqKWetNUQ0o7yGFBtyxtnGvVo9/WpKNcGFgD
ZAWxrCQ4Kk+vPbMoxqa/vFU/PaqyNCGhUTWLZ5CWrYz3BuF0tOXuNYOhAabx+tV1WW+gfV+dGXLi
SeokciNuUcri6cOrKsCHkgFYK0ipfEAX0/j6hTZsZz+eZvnYH/tn6PtW1+LLtdMwjdkloW3GnfuC
Hqr7lau1Kn7DNtS8s+X2Pj8h1XI0b4UdvPAmZigRT932GjToZdAn6W9uKIqtWhQvBL0hErgFr0QS
TdQDnKEfzD6fn1mzlIkSI0N5OdGmpKVlu4GXlxsw6ES6T/m7dKjmJqBfXLjVceknVNEQLLGJk2cG
CyumgRw3ROYDoCr1sqVfKu5QB7jFlyJ1I9lMvHCVi/FP33Jg9Lx/3FlRiTBDtXouk41bn+ckhP9u
p5MutW1bfXUauql1OmuY9bReM5BOqlTiUiWlxW6n1+pyR/r6RJ+N3kkQHzqzJZUU6taPazJdAPIz
nnfq1MK3dpy85Vx8pz4fRbeUgLpV1PzbMOboChSyfVw6EUmeMFuSYCdoc3A/9pFWFicOAxr8pBvI
cId3e/auollp2gFX0bstFW2FTESST5RVQNJJntS6xz5cC8drcvHlZIjWrKcCWvh7fUjjNXOb9u88
dFQ/a//nCfDjj2aUdeLK//C5YW9G7EM+Zz2/Aed6YZWbovn4Mx7sLSlKfh/1SBBL/rJsinXtFTV6
n4pKrtEnqNZslEN9EzzbRM0kZCiw7Jt9XVPRmRyPBEISgJGxHw5S6HiU0uFuCtluhhbcwPC8XdPh
rIsOmSDhnHtSThdA/XrNHw49ODRUVTs2q2k53eQgWA/SirHRlBi6LT6J+5IClocO9eBWyLLUtCsw
hVEr8LWgFeNcVR00fsRPpYvinrNflnaFvXo4SeEgYDbLQ2YzyArpXQMeymA4GSwJq5m6l5KFlCE7
SuQZvwz0AnCRSjQV7hHg14C300FkDLwQZVM7zsbsVjQspE2qNKmtWrwAUtXL/n6An31cJHt0S0U4
1kk9tT86Ozx6VCSbJyJa1P9FEpfqNxpuacwONFY8YE+BPyz+P3bsylUtcY4gRo204YUmvSAED0eB
+tRrrrOj/3AtedVLIsrgphrJfx/+LPm+4+iFCzqHPfJt9klNdrboezWtwL1PGQo45MVNy9Qqhi38
aPziCEU6DHRHARKdLewmZ0wABONtOL8zxoyO9usJiav2EgtMc5xhLR+6XOXtfeO5sJk/xIvM/+Vk
TXnpCwD7OzLiDzQjE8/bAHQpniOc2Y+m+kWNPnsRrogdLu/G1fT8a+7rD6WJucGg2KwNYF2YqvUL
ZrsUml0Hsk/Q9AYMN52Ygy6shk/ErQeS/HZY04rep5jqTX9+hCBHdDAuubHGrCgDH/LDBd/Z+qj3
MED3nW+FkeYFZzFPAOBv01xDoQhMha9SGO99tBM+AxIW8oqayb1kDOXvd0l/GMgPKWe2oLN3JvWl
fAvhY9jgkCLm9zLjDInyncfgR9EEBNRrJAJTrYabwjAQw9SSfscvZZXFtR6oiWjHC73M5WSWUBau
WTG7/sup0xLxbTDuCjoEv32fHihb4nrB00/bQLEFThXdu+PXxb2eyKp7rkf2OSsB630T2YCr5Dbi
xM1KO7UsDD4nDPr05Zfd2xiXxk+tTSbvwb582s5BpMjFitNLyLJxZH+7wc3OE07jOZ3w2EIbWi5r
DwKQARunoQ3RL+5rOH5rjtUuBCuWFj1467O/+VO20rKcjnd8lKNFpmPSl5KH/RVXzkuxmbEYl/fw
mAPgFcyzva28ccSeaxFnXacC5JXf7LH7qIWMoa13uz477jT+D2SQs7g2SDAiL/1uTrOQG4lzC32J
zizjwRnXivlSFeCuzEdGsASsCDPQitlDnIYEs7r6Y+kuo65PcuvUvHisplzezdHyQgJdFwYKPEEN
Ssg/JGEQdiYu9HftkSQFQCVO0zlDCg6wIUdZ3sRODFn9Ga3D0tZ2vumePlZDX9hFDwx46fEdNNIm
Qd+ASkFBZPfhfmOdSqQ6w70miAJKRxbsWSEKxVH5OhSujvkcB3mPzphaGSfclT2hfijpL55ckjNG
2I0zTq+7pJN99GzSOO4y9uxHOHY16MlhMCxtOzuH9xRaRpYGj4K0BjgjdhOmBvTOkkHZ4fzFZ0x7
smqCmijtf35JphEWpEnyew/ECWnvcI3ipGjinF0toMHNPdG6tb1gYlFugcgyzNVnFVZi7ZCViukW
EsTheIHs5bSI21/1PgZ4Af8nnvKMKXmJVSxXfqyEex/ys7jkbDiwR8fIOFIH+/966yjAQNRsFpuR
FojWgefQ8dmcJdd42g02t/x62vTEtZ/6Gbnb9dX5ylVlwibovq+zQ3w0O2VphU0if/ysPN0rkY7z
Jm7jEHit24SBOZUoM4TSfL4xWvEqRjffZ2gN1MIa1mSeaCb4zU7HsgJFpQrC10sOYMP0VUIaKwfM
A2m6hRTNfGLin7V429NKJWnlro8CNfpdYUo+HGNAecxVcWzzmXqTXzm/JBMuuLjpNeDpcUSHZMoT
6RxOnFN/7G/w3XVLMj8oTaS026IXase1x2bRjIo/JXGOgLZi1AQidSg1TBnD00gKGRl+aD2eGC1j
sd9r0lZ6uOhhjpDaEMcFMAXKWVo6hYdwPV4omgnxoitEzYGDohTx8O4IGSa4n74epN0o4fRhzsZ5
HDP7hO03gw8C3X92IAOW2m78U28YJmzHDnnlTKLN3AgPLgEzs7YMpKTkIw/+6bs+Ves+m9K1Igdm
j1/oDIdOQwHpgEyyB09V54MQOm5Xs6wrcRrXAsL0FcAufh/7UkGc2dsijBzc7bBuyN+cz2HQMlri
CP4GJGTSi048KBW4uo+7QRhZyCzTSUR4x/s72TD1doGGObCJs6sqKJ29Ez2heEJrXglDtLz6dptJ
3DNSEAmZjvRbWG1E7W1sOficVx3A35q87kPkTiZ4lteYyiC84VJ5ZDAdDAZ2jZCMNCMDQgU8px22
BS/V6EXC8FWKyHJIg/h5tMrYPQrQk1qC41o4+ilL6iTySsSU2PvL8PjWP6pvMljRGRGWv+4qODwk
WyNIw14XPWY4lwMzVT1Ymvpc6WYrQQTZ7kqKkgG+hQOXoOXY+VnOXM7kJAqmbGFU242akwGu/iKi
gyDuuHxVk/UXD3bx1VfShtCbXPLe3tPv7mQfnpwtaWPK6bxBrK6tlHW4hooX62H4rYOq5/cJmTAc
YJdifD/dehG47SvYuaxSRdPOm5gJA9CgZImV60XFbLvRYtYGm+gZzLllHfc3mYjDx5XE0uyI25wi
Pg5zunFg9iuw2b0D8vNsBFc8S1z2Ywr7LaasOAwVaBAY74etyutkpQhALrP7ZRu7IMIXb3GaFVeN
LzRw4M5qP3jKgSGVro8+NxS9AuPqaJ1YHA/kQALW9c8UZO5d8S5mHru6wXpu9rXQ3vLS+VfbUdEJ
SUII43tvX8/g2QFKhwxWw+pNbc9DV9476gHSoBi/qwoX0FjVUn9NxKTXUKlluX5BuVYjj754Xfe5
h/9W4zuGf7gh5KK36We3+pzZ4DVn18IEoYu/hMDtrWgR9wLivYZ/mFsSOyjdMgvTM1tAQtCSSbAJ
hlXqlTLRWGnlDGBeU4odWVmBNTYzQ+pNrjiHvXHW6cPscsQJWcVgILT1RpXOM4piM+WlN6PlBKrF
kQZCvnbW0auJdBICJOufw76X1ylKRadQxxzovAkEmw4nSPs12DCNg3iFKxVdZn/6shT7ac91N8Y6
tAy8nwnZEX4RvVzMt7OWATEODTCIDAI4nYMdZY80a3lVX58EvEGlySx0lQvmtCWBDLvGW1TE+FpU
WL9co37F3Y5XvyRdpoKwhYpU4aWgTn5QhFjG7rTOsdWrw4qjLogdRKliaAiFc5hpZd287gEE7vV0
j3pRqZUlI8V9mEFgbseWyxLwjBQFBU4ALD6tnvsV9MJxCde+hzmlQr7j9iZ93hZxLGk947CdmpX/
Jn7nS/j+LlgiwRXT5G2c7M6lh5OJQq2zRdz43buKWLR8X74bzNt5qtOEmmKhPuykUFocp8Nk3MG7
kN9A8dxHl/l6aIZxtUy6zd8RRzM+sk3llz39GJEa7sbnji21dDBsczVvest1Xvmom2JsCN/Y90e3
zQkJZR1fiycLBbMGWT8mj5SDKP+ByaS0lsoCU1iFCjiuMVdCSKsdMEAQ5CkRg0sNkrJLAOYocigR
v08QBtNxy1JlKhxEGsmb8nkNVcfN10pgxwwPfcOw2Hj0Tc0YprG0qJCRzcTTN73Km89QiU7BfCj4
C/fEPEu+dr6Dc9QzUuCeP6ovvZUUlEmsCJ2A5uz957kOQ+HKguTA2LPTLtnryOXVqxDX8MeAYUtT
nGWLlqW8UUI+kXJ12SwtYNcOjDK+QDPe3WyeQ2XQZB8dmDx1fYtb70IQlbxEVL0Rc5W7z/8tAWyX
EML/bJC+W56TiahRfnwosK5wh7arj+5V5UjK+5YGS6+uv0kFFcr6e9gh7h4k+25xmCzmhB2Z8IsA
j2chhxH2c+U814QbRyD4lseIP/1sBOYEBdfjK82W9G9GZm4MtHznkS1kNrSVPR0lpkohMJZGD/ka
CFYOtsLQ5kSxUtVHO8ubLrci87m/76dQJt6LYXRwgz/SXdFQep1iha1TOz6T2MzNNop+E9xyFM2a
6Fzqla6of4YbDCco3bNJTsF4Jdgd5GgAgQGCAxuuXof5Slaopwwiz34nJeTlpTbDqJvKhR35v+xQ
+o6c76IFyL50W21l5+S75FU+FVidVw9bB6MIjXG+lvK18H1k6GdYfyzKZy7bPH9D8O8XScM0K1fl
r7++LRPEnT3iD+n9D5V+gsuaymL5Z5kYQYaTApwPyE2aLK6T6Ep6cXzvblJP7LIQd2WkFdEUavyz
5DUp6Nvi4VrNB0f4VcFmPZTmys6+Y9ViZ+kK0S0Yt+3S9Bt82BIfhe51aFAzvX5+s4vDPkzKxuus
alB9wLstGHgxh6Q9hCsYI/ukdbaSn7vHCNWgodmTcmGXyF47E2wbKH+c7+a01hXMKUUGD7guOOey
hhMGWyLdFBxNL3sGl3qQm4vq4t1nrDp6q6719JKeuaKxn0dLXY9d7UamVC1DFS2Od+DP5CefznUi
LV+tzcTBUZIBpxpv8gYitskhVWheRsZDYMBsGZDnE55t0siNaWsOh/HS22mYSTwoo84z5LPgAFVo
KunEOVUfTYDW+HryI5R1sorZTGjL7xN+omCN/xMJAvAp54YO9crBxJyq96mdrYyASaAC4ZZDMMHt
CFLgf076ZHt3J03fJP07TKABKYQigpeXpSfdAhhXSccP6yFioK2EibOb7ygEDII5I4I2nFCSH+U+
aSUGJNDWHT4+wpq8ujO7QamIaGyXXeJvDFQFuXIiV86/QssYKHqXWKJwroR4Y3ScxLhSB7xb/Mxl
CBW7uQxtU4n3+15DsQpkZz2S5eElsjXtjzCNlXuTUC3ve8KSYKDGuSohPshC4db25y6lMK4nEcZG
jwKEnG7Di3XSv6r/ADtl7lD58RYVLPnSexAoBbeNAEADqe3/ebroa2xrnGgLEdbChWcCJuDN9Rfd
NTEn4OsRfH+7GCOFsxilDU2GLoyWYYTwFX3jvQmgg86Lxn8HLPVQxCyjKqE+99/CGPjSkETfA+yw
hvLl5p0x9OUsjAll2Fil2nQuZiF8+hW9Thk9Mj7LzLbHpjz62mU6+baMfX7CFmDGZYrUrYp4uoBD
ZwgkzT7BQB+XMrWGs+3isPi6ImpSSoVWf9tQgFvyA2UHFsBjnGWVQlzNOPR0Qdu4pzMU2d5yW09B
4NFWU02TMjI4zUdarK1XNuFkLsOxsnGcz4eSgTYIkzyF84Y1SXnub7/gCeconK9bK8l/XcCjpVc5
OI2MOnGpTKeYxxSWagc/ZaCCBEH4NK6yqxyETHmxJz2zFHDixjqbEBNVqVJ/zPJOR5Ed8TRihLW0
rlvtz0ePlcz7xWW8XG4ogqdvGxk1YFN7G+OoN/U0Z8sjDhvWQoG0uOB2ixuNmgUC/kwipYSTeAgO
F20Vlzseht+1xyNNbU4zKwl3d99jdJy13+Fijlg9lb1YYBERZVR+7Z7TwPADK4EY+WP3JogG5/X8
Q4Yuz0lmbsWRmCcOXrPSNNbAI6FTN/Pk59+BMiiLePpw+Wh2y5P3rvqrkm0t1M8MFqp3X4J8Jc2c
BI7BsGW1EvPf6HhygO47ysskzIGEizlqF3ruKrRjJfbgOnTJfbKN5Oq8F2422+pbSJlJIEgiexQO
uGwhGhmu0r8z+P12tOg3r8lMV4KNvVV3cOApOhNL9JGuuWQAY4IQojX2MLLhPPDtpeLP7C8R2kIa
f7hOzJGgxmKGiFyqigaJ2CQHk6eHIT7WmW8myh8kBcs1bhY1h4Qwd7S2fLEXlkpeE1lA27uXw5V+
Q8xL0PHloNQGzHizG7svScE+yHXsE7acAnyO0quI7H4DxyRDm4rS01Jan2Bs+axAfs0OyFDU4NP0
7KJNJVvk6FaqiBZsZ2v+vzxLEvBv89ICn14/rvVl44+uS/V5659pE5Rt3Ny9Srhgko7UIIp6l8OC
pLt0pGmWc4qpDkjIdxPWVSAFVeUms6zWoWQatQzo6HZEgKRbrgpzU9WX079D4GHeT+eiIeWrXhWu
tUraXPFOmmCNkm5P0ApNcftYMmtYbYdOIzNRuMs0bPU9eOfsyQtd6xIiPYApv7o6bWJycMLHP83r
f7jLi9ioND4Q9LpJd0UnE0oieMHv3aCA2tJAJAl4Ek8XFzDZExkn2zXRteVKtj6/QQeUabd/854i
eINsSWWaFv4W2s8pOYri4hIdZsNsQqlqe58ui3Eh8DH7a5fWuS1yq2CZwethM8DGJ8hvsNPulU6w
Sd3t+SefinYwzhkwW67ClCe2VqOSLZX+ai9du7EOmSMXSt1IdzoQZlkoXodbxKv0sbLFFmOkKcbB
PWuBolXiN2GL8wuTGkrnPr5K2T6WDpBqg0l/+E147DB+zJhyyCxuaCnDqUDC61chpKeQHdujozNs
TyDYZwunnUvFaPBgGSKLtHnf6UQRSn6Fw5CRt3+FzqL3HUehPtbASJ/QuuQQOHGS5ESSp6e37T+p
ST7Cy6WrGCzXNm/accRgtrSdUS88WBDMIn+voI6fLvReXZk7Hnr5/uWZP0Xfbdimf/KfYJ2Q3u8U
hGkwJD2mw8ZRYHG5BSw05ufIXJ385h+N2DcXVJE23SU1NB06xVE3BB+VIoJLMX7lTUhByTfxzvs1
XG5+mqA53J66PTBco+J3luHuu+QDtUoPTd3wE6q39pZYjpx4k9am15qhvlTPQB3nIZQdQx/emchg
9c5Hef7u1GFp4GiqpKazpyCWoBVws0eYePoBiml8PWyNyVt9eBKF7IvGxmSBKMqMYkFb8dqfC/xk
r+sI5PpbYmMWPF4NedesfVOQOQqIZINaShGlrtUvXBEZ3hPOl+ASouXtPWQwlhD3N1WP3of2M6nB
qlytFei2hfyrWggQ5Ho8KjGaQgru+txqXdaG/iA9dg6TSmwgtoO0Y8HAfgsDzD79EYkjHGq3yYg3
TuFGmMn2SVAVfoEgHTDz4ivvHKwq3K87mDo/Phrrml0xlnq6+e6NpsLK114wiSXDyeRsZd7dID9t
8b/4GpzwmcV/uBdkWd+XBMER8nGtFxtTxPICwTaiEer9Huseg4tHWxqlNbp0q/lnUkb/ojIbG1Sn
5vTr62TstAC/x65YGFCObI+iyjWT1T6HcLLCHOUB+Y+x+35gfcPALevVTYMVOdRP98WQZxFuoW7N
DKX76425VbnvmfrFbbkA2vX+G37kOj4Y8iL7UpIqNniQOvw4k6c5QQBpcPJ7fdHmBopLjzwniTWe
4Kes6SLrRuTqrgNpXNQ6coKbTfMe6ncoBrN3F1WXh1wex1iXFKl6r7RLobTs6WWXrRMAeiiT8hIB
p1ljq1eiZPuzCHTuahiKgPtWbZVdo0Vousf1yNND16z6WqTkTgDFhsQBbJKrbmahYJPWFlPINoyP
FcGBpirzjKV5/oRU0TbuZVSqJ0SUYVQFZyiSxtLMonqZ0p/bXTEI6SmsF1VZxFfOFFBlM+H3nZOj
38EhWfQa7CXIvq0he5yIGcXOMiOPqzbhx/0BGZI2PTNw/T7AQr1k8MM6IXWd80G0lSiidZR9F2O4
mYpm7ZXSfs/XyKkhIRVHmdNO8nT4Qu0Hd8iWxjljC5vqv7PVlyS+X0l3onGkZYGQjqpPU61C5HcN
jljNGF0wNa7VpiJXY+S63/FeSar8IM1cX8G/TfZAcbK+urn+w0nF9/t9IHVdDxkaD4Rdy47PhPJ2
S4TTz9sx28sivn7YQB1UFGbAxOM4EvlwzQT/VG1ajWZ0lQqPI00lghELNlxSi2UGnUnXuTesa16Q
jrilA+IAm61xPzqOQAWyb2SQAddSQ4Wpwmxi52vQ4ZZyNUD5AXed3zcepG08lPdPPhlp69Oh/cBo
kOEs/NMHHchdCJO9ETU31jvZ1AS1v4xOoHgIITLZcBExgbVzPLT8YRAymUmsYUcTJxBdDEFqQnTO
wlhrSZ9/VSHBGSk4bhLzvoAVyCCxLCicuN0IiFhS0SOXdtpHj0N53hr807kzS6+06ZK69Aak+1y6
PjzDgS5PDawhtlv7j2j8d3/bPC99ZscYRMQZetqouYjaXWwR+M0XOjhHCz0hZ5BlyoGtRn+SGaW7
CcWFdghS4Q4oO0hiun/7veAbeiuta4Xo6wPboJEXgxddvJWtLWNVX8JEP7waKpXaX7wttCAmZgYJ
qxRaGDhkAdm+dOwCawLdRgxm6bAbps/JuXk/qchJfrOXm7l6ErWI440f9ebAXIcP9A7n4lgnryQV
LFqN5B3MXsFfCO7k2/g+FsVqmS1MSdqYIUDgoXgZawr3eXb4OwZPEi8ShX5v0rQRoLQE2xvyyFPK
n4UjPLRpI3rmw4O96F+RSEAFiMcfM/kxi47hWIi7PmPdNV33YrF5BvJqU2HUCkU4yNo4XY2ESSlc
9n1OXSTJoSXsoYLYHqLZsHnQqg8FQcvZpwSAcB8yznN5kXvRTy1EWYjp7CHhPNYHy0NKKNMfLiSl
c2J3wD1n5ZB0AXwKSym+2Fy/Lrjz55ihL0BOKDJzwqbOgSEHraPyD6owhdhd85NAfJunGokc0rKh
AWsjCAIK6/3o5gemNM2LtZqwUsid/2cH30jAs9bqNeO6TiMBOwqToQfDECl60kdOa/TJlumE95AR
7ptp0d6hRB48/5iQLdsWR6nQZ1DxovQ8lZDULQg3qDtTJsXn+fn4UBBVMAw947nhvDsDq2M4hCes
LBgU8u/A58Jc13OGIqsBDtBDd5uhJ7+ZlKM4JVieCYDGonkZdXnSCQQb/QK83uX8+ENR7XInOgT6
glLt/B7qRECnbHHBfxECOc0OfddKhEtYIWKWviB6u3xsIVy71rtTvaHRUPOE08xFC2BrsBQjH3V0
7iclEec7f4mJISw+3gVChBMIRc1gdxnTl3dnuAJroYCOMVjjcYVb5RS8xL4CpphX20mU/PBv63N2
tCjTDlaUaQhiHuS+vtvgoWLO+UsAZA5iBUxey7HefFQOkHxVBJh6hQ0n+NB3p/IWvkkBy1Wphvdy
9cq5zLF1GCcKeQ+so6ViyqeyE8LQ28SwVHzNtimzrYj7a9iP/DtNP5R224zVBwitbTmFWOQNlwBN
ZX3wtNhTye3w9tHaCuRdrfq5JZptwywvyop/MN0r9YVpKfsEL+SiQ9h2LYBIdAO/+xF7e9zWSFQa
RXxB+Oj1rUjIV3Z9HJpYEv6dkfg8GIHpq0bcYaRbi4ZudtPHpzo7aAZip2iAfAvIM+vUzy56CaA9
vQ7bi8acdQsvXhbZhV1NpqPKrFCBMZDoHgxmbaZ9dkLUBATGnGXnPLjxqF+OE9dQrvq0KtjD8Cod
M1I7YW+bHk6P99McfQMxREqIO/ncUiT9sqZ4lThDjnbcrWZH4YQvVhuaN+dZJuU7maCoooOLJgyc
mVyD3eLL9R0Y6Mo1TwdqToqehoRQeRuToL0Q6Obu3tbH5Uj8B3GsaIDXlQYPs/9xgjuN/W0ikUYA
WZ97Me+XLOF8VmS1PqR2wMan9qgHEIkRqNUPu1tD589OlYHYYxhrzwtM33VvXiCsgS5IpE2+2lDi
mCyxC9Jn3uDrkiHTpuZJNSJTERECzEcLBbWHDI59T/eVWJU9SsC/IZYZ33xakGwrBZZkwSklYaCh
SxdHhdQzdKd5RchJAuC+IMiH1OigwI9hTK1Lkrz9eqByooHRGQUJ8uiam5t6WNi4VyirHKytV4Tr
ZcGdoM+jBr5qHDV8RxWLMLsJJrw2lMAN9BzrB9iNdTJaMLWm3cMV+DiT95JVcWtbxl8NuxlH+IO5
ZhoPlDVZxKhZrisXAQvXZjbvQ8LxLRpndzLHbLQPg62cmdX9wQQQsHrUq+iuuDDVAbvKjB67K0ii
yb/1Tiw6pbq0jxwtdqvKm+mXIQsm0vdbanNOPJZ8trhPXtjq/ofZUs+BOMnM0ErKG3YlYSw7Ah7P
YMauYHQUTZi55jZ+Ih+IoyPJTXMog3JYemeIAC463XJ50syjMgj7ullUUTyl2uRuGR7I+V46hDQb
U058TsHIaoV7goTh3qdG6rbQ7UqHyMAxmhT3urTWxRn0j6xFsEdllt4sxPQAvrm05dCskPY1n4bm
hemUlhAAZ/xspzSQevKmIYrCxikUYwkuFTNW1dEdGoAGATrFjFGmeV2j0qqJ1PZiIVYkadPGRoIb
WtFg3H8/Ga0pLHeEB4iQmYtS3mowKpF/i20gWSItZ4KeR6/XJeThdn5heTBcpeFDAKMEdJ9DU0tP
eS0LszvvgJjIBaaZBwpm/RPsHXgOTg2RELn1jucYiTqlj4c7ekCxzdKKAhInoy5jPVJR0jmS8tCR
CP5GU2SS5a+SdqnQt6D1TUDIRTbKct1gC5y/xEyauyicSK2ftGs8Ji15mKTVG0QjKkWjIQohuR85
GIAZZNKcgn3IIP3qWLOGgCJctJrc4zmHFz2HhfwoCMtoedKJm4E6lSiO26j1lRPjjt/itBiq5Jn0
J5AiOf6zQOYcs+hsC/LfpsEP63rRqx9GnBrPr6AtiAjK+peHvTj+Wa8Vwqu7iuscGScLpstpLxiu
XJrVLe6EJnE1IFyXyn/HRvxGFGUqgoMIAB4HNAaz7cs5bfVZUuFJUsN7aYtygQAO5OhkuTas0iEv
gHeIZtCEmts/qeCa4ar05DEKe+AeZzBFOE5/ocynpDaHT2ROEzsBzAxmwahFFG0Zz81g3trpmzjV
hfTDd2mNkt5O8DP0v2HnGAH78fahqw4ZrCutb9fRDD5tG8BRRWketJ3t3r8qatR/w12CvcbSw0gp
Knt05f/7yovPv3h3Vmvi75RFNPZCG9teyMfZW/b/JEHVZeutI0vnunw3nwGivVWwz8jEkYOEOOSK
9oTVzVC0/cCq98Vj0oMEV5aITAM5hYL5qMIqQXEHxeS1kE+LdMJZ9Uci24fBmgUl3VjEiQQckrsp
dSQsTHp8ac5Mq9EYRJW08ex6BGGa6y0Z99iBLlVl4hThRcikp0+I8SKiEs4sC/X9Ee23Rrpt0vBE
nh/TPy2zXGzvHT2zIb8OwobUbGtvPgt5/Wvj8edrfLS1Vh1zOW9sS9EDIbTxawsoxgfpi1zYgwdg
8eQS0+ipvcx+U8c2gVehjK2qrjDDZp8AOd60KzxMTtJpuwA1aRFARurzW8R/onbI5H/GoDi+I1+Y
TffAzCw+ayxprEbtSwY7IhouDjvTOsCwBRB/lh7xaxKFULSxNtwQXo5bdb5NC+d2ce2CZrNiVj59
UNtnppZtqQdxquCvnyYRKg4iisxcQR6C5ADPhttOYFHz9Rd7eMskFzV/O5lFIYZeWTwhTWoKKLC/
vLrKGUDgiFJ74OX5A29X2bkvjDQmmf2lvgtO5iA4C5q3E3Xca0rn8IK57RZMwiYtu5JduuWtuZnK
A1u7UMyZETK0Jf8gKx9hc0CZhZqGqBRfdoMmPT1NUJqOr7RcbIlay3eitrG6IClQsXW3Ara0Mjsq
oq8A6OFUNh3z5m3sL0QH5mCvMdPlM0oz06Imlov9VizP6RxiGRatH7UspBfAaXlkMqIwY+dCfniU
i5OgDMaTJIjzN9/OFIZF38QnXJuadOzHysL3yhUHlP1QzDIJrtegiyzR3toKwv/egYUvoq7v0KUl
7zI894uGGF4rxg97sVcH1zhXa9FTeDsbSvv8Oa5y6MP8+d4eA7sS17sww+m2CGwvmSHDMGo9Ixe9
5nTOOWVX/oKqz9sJOOkzBooCR3MO9fexXMiHwY3/LPnjVU8iueJ6PoXJeDHe68h9t81+fVJSq8jA
cCi2jn4IDK6gb89DAIzVM7Yzb7lC0agrpq0hPR73c/o0wqfXY5LGhVa7dBCygGE29jYOMZR2cLob
DwEyi9sOlRy3aINrfH/lNkPAnYMzS2kK26+5IcXvHNEOT4LzfJP4yMzUCqN/WiN++3Tr6yWVR+he
O0MtBpO9i1I+fd9UozqkFKEVOqHJTjbVz29vhL/DBrMUuzZrG9xxKKdn5CUHh01r6aks35nNq4WD
K2UZvRftoFvNB1KsGF7XcBqlo34fNw904Wy1ITBIKPQds3KGiQGRZ4su7KecLbFmiq+q8ydENwpS
lO/yjH2ocom87gXxVFe9RF+VjJtYuk1eHycoKLroIWHbdR796r2jL26lH+MT99lGV5h/rIZmWTQ7
DQxp8uCLdENPIJSEiJt7d0IP41QMb07NA1rkwzfvqjHavD0124IgrwaCwmNnUIaQFQbV+xBTi91V
NJ151nA763pU8eKcyrcmoN+hj8xR2YPDAnLZ+T2syPfFzv7Wd0fLVroVPONfFdGD0quIJKHSNIgo
zL8CZfSohLyDwoDi3keJNDjUKvAsDtkPi20UIqfEaGOGF48emBa/vC6QvI3j20/YNNeTjnGnSu0c
jVmudKhGf/kCIVyzH0NiNKxcnZifxJXzQCZ5LhFY4gTj3XFmOm3sqLIKR+BovXd1It1d4lRB8gQ5
+AXgCq/JbcU/eP+Bx2lGRtAIkeJGBYh6i5h8hw6eCF+gR1eUvmdqg/u/jDHQa5llE5L1Nn/GDA2B
+SbK/Zx+jbI/qUONXqDMxQ86SaBL0WZ5pyvlun/ORJeLtViNmuD57xOdAq5uYFkPCwG4BnMs3HZL
lTz2CclXS/NaDE2zFHp9oxul8E9P1d9fzcvYts6c8dndR6e47Y2dhYVjxVh3bX4gxKf+eTnWJ14x
Avg2rMYAzcJnDqj5FdJ0hxwp2N/WQiqhvxIkgWxjUbZ3Jn3cHrUoay9mizUcC+W2rWm5PpwUdZEI
7Y5tzcrDAdhByPctajFE4Vg/216sYt6qY1ZF7F2/EGWnefVynVz9/VDUsvNhJ2Vx+qNlGNXW8EDI
kHikrVyNDx88dArTJbNtj+DJYaeHkWJchVY3dP2c/p2WttWWmb/6QfQgV/+Lul73B0jRdaNTZfUH
grdIlnknMDDZJw2QDA8gKuuOFttL2alkYM5a9oIPtxw2+pfx4mDuQrcseLvnDajBPcHCdzhWePHm
Oer1ef6yT1Ip23Eh+kXcttiAhePLXuqUibja0eVTTnHtu7+JwOIPWpe/KF4Snuwcj04Y9BoNFEkS
a9Nw6JAS792YffG2w7wTWPDvBcacqrQQ6bG5CEHl82X/MOV7BshVavtzNZDuBd43O5UT39U4AM3J
1LGdvJemQwf8lcg8LfSdKhcFpPb14FEg9fCh0WCl6HyDeSdT6zaGJTIb+kSqJCQWdX9fLZJst2/L
sV9hybCEXlGdUupTZGhXp3dmczlWEdDrhrgBsqANdCvXUwvHFH77MOmlrhHsrveTDc7Xkb4Lu6SS
c4TOa1+s/Jhmjj3GoUiDhWGlSW0JQvO1Ga3xgmEGC3rfX7e4RscOrjh5TZjMmlzJAWdQqkOAcyWD
D51H2HP1PLAlF4yG6/HarXQZoT1DXriDHdZ1ejHRuc1Y9WjIJp5/pnYd5x0BotpNqNpTSYeU6tYm
QTR06X3SNJmKtdm9hFKfamslIt1ICKB2gWSLZHZfibRsNMbEOD3hwBjc4UV83ozE3FVR2ypv5Zi3
f7kQELUks7xi/SH69xIh1mHnIqYs5x4e6mgnzvWKCXoxfU37XQLkz+Vr/2VrHgmR8MByQyPB/U+Z
5XqJQU3pL+CvOQLyA6KsdOIoRYliDCHasnbBzDGFC+q9dTI3TQiN/3jHcD30eJbH+dlKq98uNnWK
vuYNDS+b4n1fXlmuyzeKCTlV2n8U5LrvirLhZhKxA/LyZ4PBE3ljcIxWlaSq+5Z3wcmPHp1Xv4/R
+Qc5bJBMVwubWqUnVKFa0rNiEqmYVXhuj92X/dZ+Bzfx60F4S+uPZpdLxL3nIHugig5wBoMc3ffY
mvl2fCjIgNwtKeESaWdPY5vbjJqq6Bn9pI4GoYLpP+rc8vOv+JiM5h3BvIZw0UkMGDV/Zz9uyBeu
SRmnG8I4QJHw7YsTK3BgG9dpaV6ouz1cO33olx7bhrGrAXo2OqZ77XY7AlFDAhQBjBSJ/5yUynNC
uGmNiC+/5kB7Q3jhBh70Rmg9l4U1xxAC6LRQsWfrBbbnPrSB6KhXmqJRGEq9E8FB+rRpkntAtIqX
EL0W1133qOWDIGNYhQlMISuRlMn1TtgYxY3Qa7SwJX+rzcqCt584gUJBOA/KwaKBOkqco6E+BX4F
dbYEkhnNkgBMZpt09AN7fGxut8CTz8T3lxXnGntjSLIyjVvNXDS8SJ3maHSIqmXRV4mFA8aAC8eq
FAd2Q/v5HCumDnk8BxM9musCux9K8qj+kzTNugpgZMNJvI2IoLxEuSZmoMwGLqUJz1wUekNU+ahq
6RttHCtGaqSu8629ap6uU6TW+kAnQTVg8VwPwh0FpzDKo59E/YIDyBSJr2jXlbkmYb7mwWIY84ph
IK6rkRuNDhvjiBhZXDC3plEIsIWFWW6CQtE5a0H6d8I0La/SDqaxPpCbOjabU8N7hcny53y5ZUr4
jbi1BNePuBWT9zitzChFcilOs2JtU1wsyyeL+GgpBksvzzmiCj3eYWJvSAhiNawBS/9OT/RRAn1q
GB+WGpNKriHpCqbTk5hlfNXWlv3Juqh/eEro9g3IYrvQ9x5sZH1ExNioA/FUg1kjWkA9Uwuoh0tz
/7uwbNYHqswBKV2fi+dO+1uCwhKzjiEgphzh7GVS5/1bikrF4DQlEebhRgJTZqtK33TMjjGyWHw4
TSpI00GyKBsOLtGunQ3KWV9oMuTUXswFqEOB2hcZDObK98O/PFI6Ep4Fbtnqedu4yh3QhVkebIMk
Lac+yESL4r9f+IGrFEC2keZTBzti97hfE7Zu3o0RKTC/gwoemrsvxza4z4YyMgW9QYPaq/ZuJfDY
IfFbOuNakiU0BAbuTCvEDYb+apu47WYLzGLOyVju7KPRt853daTB7C8l4Ku/njI5OBQeDiAvsaon
RM5V1GZE5oec6czzW6vSW6D/327X6uIh4Vk9F1fxiau0LYg7qv2psIIJIV+wi0AizHLHjArSb9DA
U3Vru0bpycGS3dFWGZNvjoT2qO6qwWvuOLdT/3prt/JLtmUCHkhgbTyeziQvLN2BM+viQiCDBNWZ
rh6bnRrC0AY5BAEeRIBbjA8ZvnMsWdLKN4s/kO7OkoqQf//8/fJ4ZqRv0ZDqp7c5W1wOV09CCSY7
wfSK5OrCbuOJWpeZOptnGEts2hFdCUj8YZ6oUBYWq1D0PVRharS1aT/ZnV/KhB7IjGTP2Jx3nNkJ
bQB3xwwff+K5eJ4Xb4QD6lUfUqqtUQbHa33wXJribxMqSeUs2yzO2LwOJTd3XpQm5DoO2N8Ty1+j
ReLVsygMjEEER4CNrC6OS8OIxZybz+LkVWNG0CDZrkEB4ycIK+aP0UYEXzlgr6o/WrVZQbMfR3P4
0d4rBr9hETBX4kLDHZ5NpArny9cG1jFZvq1Ab914TCIuIo+DiIYpblldW4qoXo8LNhrQTmUsTERl
7ULl4u9NrscEGXwiPEiexq5I2GZ4lgNIvuOzMNIzIm4oGAETGEN6EgnttbhvFm+R2nshwnSfU+W1
erh+UbU98jlkRLKQ7sbTNiAV13EJlbZzYbEJdvoRVf8zUvh69O1WoOunscBX/sIJo3xTXioUnPlz
9BxFWIEWJ/Pe4TuLT6AePwGLA7uoXBr041iBiBd43yo4yN8SXaa1M6Z1vx8yH6pyy2HyZl5WQFOu
HnC1qocb0K64+JRC+6RlwlCDSDhgn/jGVuTMmuio2IL5aEQSXNTISmB6rtwH/oX0HVAz3xQmDoVB
4BunsSNtALB8vJ8j5s33rfG44gPB68Kaufvc0h/+2SULn813FgAfa5VkUxwAEYsSO5S8RJJoItDj
enOyo25PPVMWduSOSVFLfpS9wMfrtSkZIcV08F5wHjWA1LDSHrvIrMqcORNeE7c634G0TXGAPW8D
5NA46btMvaeFO4eck1TxnY3eFro/FisndZVZrejZhQCG6rKLtiHCL6IlUWpGt7ESYJvCLR0eisqn
BcQfPhUdymR170bI018P/jGGXZZAGxNdXK+K+jG3yf1qmYcqA+0PS3IHf4TAlHTkKZjf6ft0NZtA
Ok+s1zBMsHbB8QkSDZWoOBN0KVWfyn3fBjGmXx63YMhSyqAbYYCdiSk1OCDl64sxbN5n3ULusbL4
/dVaKWCTwi/JKSAvdq2aVjt3mD5eOOJZIVXaJK3II9/TgnCqoihNWx6cAXaGQxAfKRlXZ4UX6XOe
Xs60KrneD41A57oV5UROyxatQqx23YdP76H3te70HqzP7L+gTmmdiSvUiN+CvNTV04dvsf+jFrre
V1N7xHD4dMLEEuBjxTuTntMHW6pCgcCkEARuzv0Qkj0uzib/YW4vCTjP+i8TsjfSrjZ95jOvFCid
MWxDPN30bVrZj+uRWKIsAOAe3fZ4khZP7L+/r8DjtJyEAmpMTXYlj5RbKnxCjIHN2ZCLnTT6DCcf
/fKQiYjjYL3sBFkUCxPKCOg4ad09ebp2B4CUhWMBOaiuAmGlZDnv55cHeULk/teX0CnvHNiIEiQt
7Tt4SNhph6XPZWrD+x5A61Pw3kK1RHEqjUIsoe9vzDTauEvb8tgv/HZQfme7fXL50oxeWXJMEdKD
57pqg9vJNjJZdKbQskSsss6Zf1yicLbA/Y5HUMtpxC+tEDjry8QvwI11gx2UHoHpRAY/nVi/DAeu
BAfTol9kuinQSd2xSHJpoFDMTVR3n5GEI7AR7Tk7yYxo5G+vEyNZlaoWAXYWbVOKKz6kPSpv0EfA
+4vERXm95IaYTptl30E2yFCf46r2Eop7bxvv4YEsn4xRax4641JZE7+upS2ECviBpqPl7fpHOAVF
OgTnFT1jth8OY2v1dsIpR9dCxr6GKEoa8pYe/ZRqVyfioiUtlWz40d1yJT4fSO885X2NlmnItaTq
Pf79ez95J72kusgDN8SAjeTyzYHd4heDI3JIq+oLjRg2HasxgOPZAs3paR8uCCrtN92pff71Kt/K
mmYdmReF5s3CFtX10QhRPiNl/ZMfc2xF51sYXPJ7+jlB7Pr39fVclkWqDYmtn1Bd4AhY2VKHufSt
L4rkBwr2iBCvrK8CFMPIGvtfYYevJUGLZNC7Ofy7DdjbQUXWS6DWlzH1fwcNgvOXJvmuy6u97Dhc
q98hkGvS/w4pdyBEcvSAPPDo/6fGOo/49CwEF0Va78YUZcrjd+61+aGbTIVmY2GGwk3v3GEmUnS9
bXeMFUX0cTjf6bxDKkqwXP8JdyoucHQiIrj2z8CPms/C/llaegBospuOVLDveT3YlBgby45Y7Z6O
KcJOPTsaTLaNjCoDyyCVb3uyOJWO0738pfmuVQifddOabebGpqe2cVPqp6FwA1aecT8NyEZQoTuT
BkBJ27j6bLl5ytGedRc7RyX3dxnY5VJwBmsl68nzK5gZRa7ZjrLjB557MLj/fJDcMd5GR1NKL1HE
ZQJUI7GgK3Shfo15w7hTCKzxH5627J7BHJlaAqoVHl+AHh8DQD/4YMHNhNKnFgH9/l/EKYg5uwOV
Dj7UDvgBthwps7ngwk21yKTi3QctSPmnfZZAE0vc9NNdge+33/3hyPQab5hSJkm3dYSPzBOAZc8g
+/V6fqw2lArywc8eQ3dGoylbLGpaolXUKajpmhAnE23FdTCwAQvPpWeMmw9di9pFBhryfBXOQlqy
4yQGYh+dY42o2ZTpRy9wOa31GezN77htQEpu4lOsVRBV2FjPg/NANcpc4wojG/h6fO7Abn7Bs/YN
OVNNZHxscT5KdAkD81AEbrByJSCsEuhp4uiwhk/mx0eZ7skGPR2BrgTOJyOi1JydFaWwB97QM+cH
5Px0xNScS4Jl8aRyR84ZOrAtMgX0inWnojQowz01bilNrjFcrFlTQNq8Yp5FCsRQ8TKQ1nXwDSVw
LF2B8wNjlec+HKxsEmsqmtAJLvJJUn8jWiRcFbozVGAXtq3ekv+0HGEd884oJKukScRXld/mMBzl
JEm0OStCQ5Vd7/7F+yZJnMFha5b+/GDrmXWlIJ1X6li8dEWXYUw7ccVamza4vfq385ggJC5jdCOC
8J79u3erPw67PnCIN1xfxyJb1gpMu3UaYyQxxPPZ0PfBVVndXPME1wvW974VsGFEtjp1fpeei5Ni
fyNVFQqnEwf7Bn/f2Lt2eic8EHFSXjKuLLJHc0RtEkBIuXT8XwVDHtCeNxlWmogQNQ79eJAdcqKN
Xu22KTeIMbvD1NUm6gyOG9WTjC20TL/fXbzjYrQ1Crp/2cj2CuM2opVZHDi7X/LTko9AN7iDcJXF
kkuuNuNAqILmqa8MfSBXAhntV5T0Kow7QngZMCc2eskrPei9GrpgSV2CwpkFbFk+FEnk+541ws45
Jzd+xoowRpZIq2xbjnD/BeEI+H+dkhdGqhFCyjchO/J98OlFBX6K++IK6XoeP5Kt8FR8YK6t4A21
cZz11qIgk6DBGOUVNm9gV3gu3qGnkURoxq+Nsj+swdLMj4ia2a+A2qGyVxuVUVDSDdnYFJ2YtJfY
PqZiNvGj7v7+ZYDWP0xvjGRkssbF1m8X0BqWNiQqceG9k0+huiQ4p82BNPcNWkY518dIvRlhhBg7
WqzPW0DfiubKTWMCIv+AkzlF2mtjBKfLTVQ0G3bBKX0WPeaiaRvrjyE0r+E7XeQDWF/+yrK1kGdK
qyhrZg/ZC6CzdHhLrm6N+XaZkyuvTRWSUxMb4P9+JQPimWgnW7EnPNcWEUr2d7jJRI6SPuE71SbI
AEYarpSaclg6YXYAi3RLo23yOtoGNvcGu4ZIOJA6sYgSdnQ9Qe/T7N0e0iZUtwWF2bO6qCNDtZZM
G4tzsl9tIMrouQ+wgWRvggNBqLEAVgI+/GRkQwqRxoZFkKbe34Ihs8pEk6CK9kiAAdWgJyQwNvHj
Xt1zeaDPE3Pv8wxoUz6CYQRO6cfG/EISbg4N9sMtXLwVXZYB6hxrPfrX5O4YZbUjSwm+gsFOXKtI
JcWKCzGmvMU3aDyarxTJUc1+zP+cJqNm/Y8qSUidFu/MNPDLhNwd02XS5Cvy/dASAiUQuPSkddHg
Ii0ePnMa4JVpBn4NA7N+Fqi3zxepqsiIRcwp+BcHSdoS4fi0kRCLOkBFFZk8yisGrlyKzohxFvAc
69mqD0tuI9VS7X9M3pusoP1h6Dy5mrflFRP1y/ve8NoUO9HMJ6wbxuygqI4v4/mTjnyL84EbNQw0
ampmnV2E1S1acOP85px9n16bhRsMv+J62WqzQJkQBGObWvKovjGptHMXFzktaQ/Oo4Ir3Cfoh8G0
gBelowNUiXdVYRmqNk/tsj5y2kBUul27acNC2nWHDnrQkPi4OEEVE+uxdI29hq9+gSWqRaDSHnmB
wBXD5tLCw/HTOirDtHrvNUG0HP6XsLRhDQp9vj78rjvGJgxUhwV/X36yJAJ0uH1W1LbWo9NLoF3J
iwLiiG71RjVu2HdEgeVaSViEVSoHxNjreXyXzJ05ZZdpnE0XmEW/11yl7c7RFic8Utt3Ymd+1kg5
KBCGnWJ9BwoGQVhKxzB7hsnZtR9qQqm3he+m1BYiwABp0TcHjfsUxQHK4qDZW+QIYY/E7ib2pjQ1
2sEkZlL8zXZByhJ2EhwkM3anFQd5he/CvcQIoIiWwr76j2GotJitgyRqWk5G8v3Pa/lvCoLoyhOT
a7QWaGYGTFKk7+RRRpZkimB4/iMR55FKONWLzvAf9UBRtVkNes9oA0hxJbWwkND7BncpBvlHbaZ7
zouB4JHc4wyi9FluNOyuT1VLVZ+fOpvkOgFdYU3BCO473LXq06XDvXmeGDdDMEWmvDgE0KduDrnj
zohLmGI8HR14+S3DEUtRTLof4dRKsXQC67IafD6gRdECklr8Iyro8cxUzUDFVuufhlm9Zc/5q48H
8/AMlV7OW9J4PWV7/Fx79HhpUDXCm3nmoBYdbgWDCDHWCc6j9ntR/A6iO1Auf90eUhIg8KEq2pkB
CGCNH0ez86y63XbyXJmcMOiF21/vZ/bhiWN2r3rhMF6dWJh+fGZ0I8usas0Y/eRpeKBdmrGlbRAd
lIeJ6+K7wmnqOUjXa/67ex8VHNxszBIkC1MeftpWteykGled4dZbNcpMeT1B8DR588uHpPHIqSeR
e/Soyt1am3YpZJHG40lUT5YtCEpFdCKzGf468+74A6KJJjfwIOhtcsn6ohHxplz5okwDwiLzNaDT
wd9yzAhk6FClHqK3JSQ1bAYLbg/2PD0RBh0RbPo3/VvgPg/RKv1GJLGO5/p5MT5UrPSemeieSYoq
Dz9VUNcr1Vqb95q1Aw607a/TVgCu8tmAW/OsCvixO7kiDhvma6sU7y9xB7NbWU/TyLme8989GLiE
4grVqBCps7lCqtYyLoItK9NX7aa8f4VevAf7EIvAHxL8kb0As4+Z/Dxkxkcf4/8gvFqRAoEwNVFQ
RPeVqjmxTw1w8rSkcOixvkS26Tam0FhlBzX3NCKSc0y3f7jcnCvqjBatDAdvNVx9AGCuHoiluLJR
30Z0/9/NfHQaz8bJ5+x2RxF7KV+qTj6wWNTVefJ/pqr6JeO1dQdf5IUOc3sZAyltb/le1bEpKo4b
MtLTCTuGMj6CqJGdEvhlxHeLnA+oPUk2rXBe32vFJikeCl0zL5nQJXL2pT1+gb7GZu2Stsk+TN+v
6qlz+3MTIMRQ3cZKWCG/Xr1FHViLFvzZ7RrXMjeHlRpvCFix/7zHjH1Y6i9RB9GElRye0ks4djU3
I7E+l15uhNqNrRaWEdXSKTZYMH0MEFdUSHFgBusrmuWgflkzfyLI/JwVa0RRLohNqniRTjK1mac2
MSjpHSL2Qf3q6lKVdAUd6SrGNbX+/MnK6TfB4+Gr0DRxVCKk6e5x/R7QWBAhgiA44WlbK4YW8Ejj
FQUPpzdDHKNRnyOMe6jFMSjW7dF3gMOa4+WXCQ/OxJ8yXvdtmnZr+BNxJiRajWUYdd9AD4pZhF4U
1zBM70C31Zo+dHAvL+U1Q/gDNF/5aBQ/584t/ZnfwvNGmPN7F7YrWu/72GvRqbtKvnvZ3anRReec
2LvOkD5tx/Vz+97hHWwcn9qIcuq3XgrO21kAT48TGBeTjRxHXJbI9C29VOXjlp+CEog9EcksLUyW
701ZxArWwBVoGyQ8Spmw0GQLQx6e2JSJbUdq4TSckf5Coc+fWiFLWRY21TxvVeQFaHdqioAg2i5F
pZemoBSk4Vgc+NWCX5m4vAlmcj0EiP0bLrUeY0eEWkmoD/CfCPjnJZX53oohWu1H6qCuN5ZaEdNC
2aN4xxwJ4ZJH3SPQLjOBREuvW6F3Pql54i1lphRKkLYr/s1xCrv3tuwUEquyn2WwqBM+8WUmefZX
hakjnJnjeGsJmjL2YUcxEwFlB9qLBgZq8cYnZLERZo3B8E9Vc39bM6ZO0FmU+/5XxdVH18rBc68b
4GFPzW9kZtWKBxzzk5hr3IKGTUYGuM5/Mqt678wrkQVW1AjjjPjugCOPFbjeUyAf6WaWdUH5spM5
zznqjIu8vbjLntM9JYA1Z7pL144bsDSjscEn7xsNrEY7YfFcuVO5+t0KxrYNKNmLQz34jAxYJIbZ
Dz6b/OSARAda/Sch3ggqUZE2e9suIOSc+xfbYGsts1VgtHl/rUu4myg/WyHQDQhllA+nH7aSEkYf
RhjJQFCpyjaqVnvCh7V0+YmXpis0h8oyc0M76jnyCLkpfS+Qz0ILqyA4PWS1bZgURM10c5CrHcmO
7TRgsIVLWfgqOi9IYpaRhamb1dlircV3LZy0Jeg3MsMKddF1LMeti2yvja7YM3xysySUOvEs74lG
1tWp4O6v5NNJFOaCQ5a+J5osTEZvXIqvrPT/BHTTRazXTQZZQ3n33TN01cZ7yhY33Gzv1exfIErv
Qs97H4Sxpx1eJU0cOoXqkr/rz0CgObXJdiD1MxQ4imFJ0NuN06AMDpMGzOp2OWAMBz/jDqLdL+f/
drdOJGWp4XAV4ylYO9owInA0JPcrilBtUIsHEw8yxd6r212nQWEWTobhqRND4feoO2PKlIoMSS7c
2N1ftsVUj0pDJR1c3LAqELih9y1IVxrQIoUt1ls0mMg1z2XYvSuJG7EoROTMFY9CvP57DbrxzZcQ
+bMusQTxUkOApQDjSIDGSCpH/mUBrDK8TTtuB+4FD6km9QKE6jCUk0yg586QE84HebaId0awhpKd
+S8YSmRX2iPkmpVsoKhrNexR4dio8lgRiKluVquQd4D7z6vY0LUlA3vTjrxdv7KYek2x8nLsvJ8R
0GTv8J1FG6hUoautnWDHtZYCNaGoxCLz1E4f1LeWOpo2cNquXBtkfDNou2xe27bsb/WKs4YejA4j
yn2A4JGKZRM6PSbDA1jgu4rkl+bSFcPwyUVVxk0xm8FG2CqTL+y6vLpZ+v4ECH04H0zG1OWf2yLY
CV5XI+WB38FJKDIEyhO/1rOyQP+MYCPhrevy2ffTOyoZ16+auuru83V+zpJjzDfI6hWFJKD/aKtV
9vDpAzm/UifTB0LcZs88j7zuJ4a9/992ZgYnaVhAB20omUpMLvM364fyxWSZAiBZD8SnFS/mnf3K
fg9rab1kDVW4MIYzqLgALU2SO8DePfAd2n54QSoWXSWJNWjn4z8aIWvVk/yHxHl+kSx5GsePItfN
Fp0ue74Ktu5Q5hcgVIXiN8VLxAMRRO/KB6g0zrTc+nVc9QXJmXNxNTIeCpAdGycb62zVMtsIFIVX
jKrO3XENxeeDt0CJ9eOAvlr28/mXWTbuz8Ce6KCO0ByJc07vd4RCichyMFTlh7HbTCxF8fwVJRdB
zDnU8Vh544BfBeyDGKUkb/l4yn8kdWjNFyQrxmy+MRjmyGj3+ua774ZNhcpq17V/bEpz/FJEGJqy
VTIdIo8ZkQhsQLAhxWmGJ6IvwO8b6mWkj1ti/CFJC1t9V4j+Tcqd4jCQujIMaHp+Ov2z4duBUl4x
L/gwhaYMrbMnkeQrsP84Ail3hIqb1QBnB9ibU9Sbb+bMyC26mc6hCt0KSb0GvRernyYdEAFKok/Y
KwByUVmV95QBymb8vyM6HiwgonmM9DPNmY7RrAajNHWMTB0fkPc+E/v7+MdixrMlbMSj0Ag7hHsq
odBiIFYzCTXZ2G/MYqrBv0IMqinL9aQ6p4e/7ChpVmSTTwiNZvPqMjLrXrKNcKAaQFrnnjNVEsi/
er8nSEp2vBVd3aqpBOqjkPJAnDqdV2NRu+Jx8+K5DrnxtnSMeJs/oFXWNViNvuFMjpi+rIqQFE5k
MEdDgm5BCGeofx86EsXB9iBELwTIYpZxbjlbifvdGhzluCwD8HSBFRkL7BnjUdBGP5qRdvkZZ+QI
YVhfjkuxGrDXPmQZPvEmMD9c2hVc7vr/vC0jXJQW1QKottDbblve5D5X6Db9hYY/KluCysyjy5Iw
39uWR9uNKCHtBlir330HA+Pr41Jzsz+P4b2WYKF4O4B/tEO2L/m0UWcpNV6ElwJgm2qnrDW1ZWiq
pg58Un8E9fswkWnIr20y0/mqVWu63mJplayC3YgAUF98Z8ftytiBf5QtrPGr/mmr2XVMcPmlRqR3
TB635Hd0QYQ8hOwHowpWJTh8saG0oOsqIcSMgs5zEI3EaxC/05H7gS21wJiPVqXN4JC7meYC6HUI
56WGypu1X1egGbDlwArnfKSSF3qHoaVeWtHJ5iVzNLoGGXZau0io0SKggmMPyCkM/KB3lvRYCGCM
4gnc3nxjq6mI6QKWgwcdTQ8xJBjU3f3SnM118BGvR8DNFWEBYNFBz+ktnBscK4RTVJfnLyIh+7GO
UviRGUkTlG+XjHNHKc53i2iFaRv5GmrK1TIG7HgpysutBoEejfJ8/WGLNimvv1OSk+FGCdWwxe3B
yY+WfA0ZMiAliwv3rRXo7muXVMi0lguRW5aRErd84ZGPKgNLxEnGcl6xETSArEQ/wQ36FmIcP76V
YvmGnuqF2v0IG/hEYb4slC1B3TGXPU8ATscAgsnA0UAJ4oesXPCwOTSvswmmho/QYIdyiwoet4vs
M7yIVrxOQB4sTgcfvohO3+i7d0OuBNSKwNfNM8SpN1pKSFFWqsopbFq46w67/6Ez63FXpLBv1ZV1
xSaTesC4FnvpW9+WbIHLuZ3wNfqt/3dks+Uedyg0SqtZYfHRGbkqz9BnvvonQ+Km3maTEFJJZKUX
hMLJGkrEsDo4PRogxtWFCHz4YRnMTZ/3+CLoS1kOt9cfR0JvsCe01aOTmt2xh6uJYfgf9fxDd8Vp
QhsEr4jrJ6K9SOXze66c46uflyL7+d53GTQm/bKQhguZH6eK9w/0zb0W0WxjQsb5DJl1YDljgSmu
y/6r6L/MzU+O2wIZOhuS3rgIQdJ4oVgLo72C6os/oUeYS1Gd/1em3MJALTaM41cAgN0LicPEQasQ
U1pvv3FkCgAI0RnLUnPZtDQFLB2zyAoklKJTfKz+1S8IbHwHMcM6b14j3L4DnkqyGgW+IydfPnnz
RKFAvjiHlv66Y1YWVBvaOsT7nZr5Hcko7JqQcKeXMVsedGGyBOq/nPmbr+/LKntyUt++RQZipmvA
8RIJQoilOUkNLySgR3gVmA7dwazB+zJIvWyuwYqJ0unSk0TyH2+WcIxzHxB0BZ/vt8EXBdynyCZr
J5AhB0Ht2tZR4Ugcb3tIOJTMWSNueTJAqeartoo6VoNsXuVNrL4DQJ5dmX8iZ5HGdRdw7K7P4SSk
15AfFNwj//yklFDg9t0Azu0mYOlevtPG+19o8EZS84ukJw3REIBqR96f06pOcbbesBdiOruJJoGK
O+mo7ld6aNdftLQZ9fqgPhZmfeKmJbbcLev3VxpFGjHsMKKIeiNjMPnpGg6YR6fWP0/R58R1c/Go
Js97RZPHxKEw5dvSSvzouGg6Qq/H0jOaxgtJbQgT9WHZco2Z7zHA/IpYKPdT6rzR17XXiMLAujmx
fH39YohA/xf8MkhJx7BLaCGN2UMSYiruuy83j6TLSvyQLY6Gr1ST9yrWlAG9as25ig56i25LN561
xFoGKOr13v5ARt3nDLO3zzRPJicg0FhAHaR5GgCHL9AeL2G2WM7W+EiQDdGgeY0wiO77N1/5DqmN
ZNml3A+lI+zcO/UeBh9b9ujNtHdRe+wg6Of/ZKgqNwSslQidSb18EH52xIXP4tSwuaYXxDSb2Iv4
1rAzhT+bw1nP+LXcxhAZw3G/PU3rbS+CDJPH8iIUvE2WkNaYPZP3dk3xeQUXpvK9zvdSo9cWyeam
IL+MmRabw5yXrRalYGAmzzAcT7tNYToD+6ovmCgapDjd1VZWU4+S6zZegVMY/+PIbbyS00Fd/rp+
/wRzKxHAeN7RKoklssKs/CVgG/u7UXaORN8XdXvNiVFwaX6IL+wlrPC8XPK6HT+lgz5jSC9i+8Ie
oxfWSlvFxC7fCGwGM5dBc26iMmPf/Bht6YN/DJkXlyowip8SH1D8CMg8j9xymEY76s6owyCsr8Qm
3pqDkHa0F6+ZZcK8+MurBNZqYFJ5yifOfzYbM3Erf4cc2m0/2rNofBpgapFKU1Gi4D1LJe/T9EYK
y8LKsqGr0+CwTJd25/YNNoUlz1xwqDLnn4heS9fKprx0N1KC/yxulAsLLBUeUEFIx1eMS9maeOjr
YnPw/KbfkYt1wSh3kpRGY/IOBNpNe8SR/UR6xNszDPoJLe1utbAxPbqHLzsh+l8XjVxLdMLeW1/J
qDX7cfJJ08W5kPzRasGNeLuyO+zolE/vQ/IBL4ehvnS7Uhg4Jn6sV9LqfFzEyFDeudAECaL0j/8I
fs4X3ogd8ysV1zOJhvkwvpwyVisrwUdOV8OoayvEZMfQuh6trMTDUl658fxukPsN0ramZmYf6Py6
XungxekIFqv5cE61u62X8X60402a0EkVy9yr0r9O7q5548FjyUhg2D1bU7SXGnjngIc49MEFTC50
ImPm+lOw17EnPcrgOztw4PreKU4AxrVpBJxzEpdv4oVvTDCidqQS9XBUvKaflJrOEVFUdloBlfIP
8szCR/Jzwj2TLO2KQbduwso/i3loJNNPCDqQTRAk4abZzZlPqWUk06a4O8f9HpVXKmbR4LuRBswY
2I8rV7PnNx5Vfvfht7Embf3CH0d98e5ayxD1VWkqu7bimsvraHaoUmTknFOPraMUGZrHuKvVVQjR
2ELnKF6neZc5vhXqw+2i547caWt9XpxCgnAQEJO7MDNhVv8YMqQjZaT5U4pjnxjVWrOjOfiXghCx
C/qSabMOnHpZjV54zB9WsXv9Ij8usOI+CXk3p958d/dnPbRXCO9jxzoewO1vzPXxbXajf44VESjJ
bAq2tvUqZUidA39iNYEOFcK2ayjCtBfBi2Gsmz8KYwiVFS0JQcHR3LT1FJl6MVVrZ3C87YkDvkGb
vHEkzJGpuAHcbalaKnX3vFpzAfVahMUmZ+msDLaLGqdmLdvQmaPESbhWD5uIIPmUz10xChzu5Gbi
cecjml44tVPQAOq7BqKvvNCi2SJw7SljD0JKXZh1J9MN32V9dQTUMOErb9WTsYM5kuRooBzhqRX0
REqT0kI66S+2q/iesg7nyu6VUgtRMuqUE2X2RixWfii8/Lct4VR+JkeP1YQh44816vPV50NxE6LE
UuerpDlcnLHgxp5SvpM/UGgJBJw1ZrVra8wzlvhxQHW/qXFHKg52MPy+x/mJgWJAbCKFw8UbsPiW
k4hXikxKRXjxjzM37iVknRd9OwgjP5OSqKy77iSOzf2cvl3AJLoiBsBVde6sqthdg11NMajskF3r
WOEAKhwWQRNN4FvxLArMJPA1h9aOk/MVBOqyV3OfluLSth8jTuCMOtG8+0FPrYls6upEnUqfzwh+
lhVBEY1YD2HSwElb71+3YTEZtAQ7YGq+So9wTAnIcKrGlxHjES9Ebp5iXGB54qHT6A5OSsvMGA1X
/e9iEvESzN+PYzzv8yKI3IGxK3cvfItfXwMd6y8sdcAinkVXGX5zPlCudOx9TR2BlvWdEeLqsUE4
aWgyGmyRNTN9HuhBpmkQoLXMIkiV21nukbRSWiS1/zxetd6rKZOZdU61i/QjsfgElt59Wa/MyC09
m5shJ7FLPRuwglvP9Q72hAOeuWp50KW3R9if4yOpUSnvd/4MHlVveIs7D376k6b/dcHBvkj9d9La
RteCPTuZ+CtGfa4pfNEsmorf1KRaVllNthUGl+tAyGY1QVW+wFLW95tq0YpkuiGxoYeA8AOwv2A0
p4wWGf34lTXDlDvoML9btqpLmuQoGcqmzF26CUZJHv+Z5w4GWyE2Sar5BUsF67xOIfAVNYUYkfg2
pmu2H1gkjCIYerEP2D/3QK+JW3t58GZEEIcN9GBK5J4AZpT4mkVUtHYp2eH4IGPOFYt1EwZmIems
3yw8mm1z4YI2GZRO4M9Ztcf+esI88tqS9W/AS6Mv4Acp/cPYJGr8gZtbZXVySaReDZ6NoeGtsq/L
W8YBBkPQnN1yguVESnlBJ137VVgmO18J8yhLPDE8YtDgz5KWQ62AUO/q1OgxUmN0U3eh91R9Pejb
9bj0olfbi+O9I1QkUXge1Dy4kBiBIVMQLnxxmdkn/P77yEQyUhniGJGp00Zflb4xD68aBnJcslAh
cX954pJGNZzQtQdWp/e0IoUp5yANr8yyFhT9wveugwAItPIjgz37vBCTG5cTawf20hWUnAKlzOc2
UV1vMLHDiw2X/FzFuByvaweH2w5m+ABd/fNE7f47ecL4qG5NT7BZRC7e3Ui7UewZVYICuVEhqcC5
YHZQULRBEhLXROqWevEwAT9k5CglFvMu0ro/rLLyVGCAT/liwYbdheBJWx23x682hDMSW3T95apY
NPupCOvHtPrz5vM0fSC5Tp8VWLQuh8WiwX/YgR3ekZ5iyk5bowE9Cyegxm+pWodGNQi5y4VKkoJ3
WUrpzqVInD/UezpIPHoAgh7bz0evGAQ8lk2TITOLFTvYhsplpCsuZaJ5C559OYhVH0IdLLCmINwG
K/tE6PWEozWUHX0qkPTOcOCuTIFwXM5J6rV08Ys2GmPwvtW39jv0IGksT65uWaoXJGW7M87tuL9H
BTYayxVKgm/ikHYFRo0iSGxs5UJ5mcnI3KV97PKUbxm+ZZKVe6SVqoZ5UTK6+3CW0oboIigY18Mq
rzw9ZoLbuXLT0ps4akTNzyTCMBDh27hp/ToB0lTkwVmIFC0jWqTqoedSH29uosC/NxdaF8ekEaP8
qbsCXkriu0rl21f/15cg0xPkvHAUt9ZyEUVkF1cYgAXLll3j9cnaz+zduN1/4d63bRvsQ3mI0QCR
crPMVos+jgdojjBDCQ0e6kMR049QfTFqVxay+XzjaySvs3kBLvG08zN3NCaJzDJKjSNFyUFRi8SF
Z1HNBZxoBzugoo7LZ47Gw1f6KQbyrgl68FK7ePy97vTVs495AMi4b2e7DjLchCOW/JLXvBUQfiSe
nr48FBTlgpyuIJzF99WjGdBnEhl24dAbV1lLEd732viAe4kG7ZrTR35rQb/zc/hP99LT7FEcb7cY
9Iz0nJgLLNzhb4xuma2E7bNB25kVS7+qasEKqyy5b8dVRAx13wsqmrjNpIlSR6BVx8LJ0PwoGOTo
RMUnNzKH5WCTgULEis53IAv8tlOlQC7u50VrF71M8f8Y9X/DhjK3CEGFmgCh3Nm2wL+xBbNUFZuU
x7qSZ01HFgszDjfofAJOVtAREeZj5RplF7XCmdSWwe+JOAXAAjY1pC+e1YxlRThSvpB6q8oNJFNg
KHeRkWgN30lrcqlmiWSdDjs8aceSip1kIh5CuQGT1RkSZN9b3ou6XVHOIRpvqcCD66yOqTKOXH7a
SkcJMqWA9Lp2ennYUb6+070JsfdNb5UC0t+K63vsBWD78w3QrtmUVE7QiQKWi1JpNeMocBGHDfCB
EPGnNCeaH9o4F8L4SrwXbbctEC/diKhj+hrzIPVZe+inuiOxmq+ZXdpiO9p0JaEGYqRFFZCSGhK6
WCut40nAmrVMhvK1kBN7AD42UA7qSIq33JtJhXzJZNCtWQTC0hxVGvkyNu0mFtKLZGMaqoz5Eh7J
RPshZaBrJ47YE/xwf2C/gZVuEzAeNb9e1OeJfkQw/VmeyzBqvf9J0xxrTmz/4h7njC6Hul2+uR+g
s3ZGMvZ78LbzH6yet0MeIWRDu5EX+CdGMhff+sBwr+grOwMzc6ZQhdNq6cHhWQ7zsbRil+u8PJvB
8AGX//t/TNCKQb0wbSjKNg8mGi7/ECVE8r3nIZADPdBDrf7VwmCGudWZf0JXOMSSsRU/rtC7iH3m
SHyGV49M0ETsqjt9yY4M75aZEbCRymFMME2f/fMWSLuC65E0xml0p3Z2VEqaQ6UsWS9Gh0rj82sj
FuublS7kLLmhMHDg+7XtAf0ln8abIepMhvDgU0ieIGYDVKvJ2E2ewIeYDyP9kpV1Q0gjeLrd/1DR
Te0ep/4kHQYBvFjl85PKVGP9tKrFavhl0FM6AXNoK/cMxoqkAnyxKMKzkj0s0xe+VMbZo8o5Z8kB
pKLRPXbd+IRpCCQNMTE2ZtQtCVpNiORt05IEbxSRclJKENpIquwPpL+YIa0LXfmDG7wgKPiOKXWK
20fB6ReDMQJ0KwLhzHsVvnIJZw0O2/bXUoXc4u0Cs+zQd0t1w+tkVZhLjQ6teNtMHw+Syh70lkHF
QurMCwkRVpIvZLOHGcN7E28jCxh6iC3KcphCYRmEIsSRf482lE62J/TTOLY9T5V2r7nd4JrzRLkK
Ckdpgk2MXdgfSuUSotD/mUHPypHPVbE24B9S/GO9TSsLNxtUK9FLJ7ArIXFFgMJBAmDvsZcKZjEG
rmVKQTe9DW5ywULeuSSlSTHb3H29mNgwEr3WVGwAJDCX5XXjusu6ByD2RXtZbEa2eWM60/E1Ia6N
JGyyRh3Re21uy3bMO/8/Ja0yVFOMisQL5AtV5bHIyqv/P7gMqDkJn/r0B5vHK0t0tUD1pkCsyBCq
OS8CZ7n+nzBi6pwBvQsddTFT25tSaSjws4BVOyfNp538U7mP31LgntrvyxKmmXgaLD539c1Zuq90
ZyBmUnD8strOhlTtNbjf7uf7SkMV9vtYlZe3J8XroV2quc/qO/Gh9CY7rM+4OJt/Ssd2PxPZrj8C
pnqXGiAshLGhF5Iw8/VwMMnkyGWWWDsPob8tGl3Mxdn2mZ3rSs7KHkYw/iCqn6NGYi67zZntSDCi
QSGkagK7D89FV1HCT7AVuY5Kb60BxB/qdyN1iQCh2TQ9xz6YkW28i/0SbopKV8Z2tjJNnoJowpVe
hH5vwMH9oX6YvjdbAT5BaCiH5XuSnUdlqNXSP1rv+fhGAtmokuBVOzMzupt/CCCIBxgg7F4WgR+J
t/lKuL1U6uWFyGjw+vV18W3ZNOVM87DA9GxDeFdGQID65gB+78lSqVXNLwFoJbvVgxNEDsCDc4+7
MkCt88C4dQMcBrF9D2LXk9cplW54lC1fxkFZOJmnz8PeHv3INmE1S6IFBr/txY1grjrPnpAoeDHH
u8zfPaYzGDcSRT/xnW/yVWlL6hcUo+Jy3xv01uXh8SucAzTlP0LiD+GORMoSstBiuu7tuyQvXiVB
yeTjhXjoqi/MKoNE48H3osRJM7uFYHqqRWLfZqGUrC54y28NnTpEFcugmsaNG5GbLmNbFKbVxHRR
ZD/U3KVhN4D+UntGDF+B0BFh6kFRYuu91JR5Sm2G8gzu/zgDI+P+erz/KtbGXYTddjiIujpOjoMp
MLTBYvN81SAVDXZCvHoWHEXA43QVSC6OX5nHCQ/3fRBHL67kld0BSDbIZjKdQjq59XIrbPBumCkS
VTiIAM24LK1sMTBd0pz2qqEMAg7uHPPiJofG1vwUawohT+sasarknR/HqvvEytN2z2cnvoVZoFZs
SuqDH9tl4QGxpyhhsrrFudE9IFAH6OdoYMFXMWFbahHYAFsO7rGUZUpM3UcD+WpmW66ir7Syufe5
YSZ/kSkw/vea7O6zJdj7LLLsef3r9gfVLqtF+VJm4chpkQQe8E6OjtmJf47eJ/gHiOgPA/M2vC0G
0wc6ixOj7KE1GdGGh7sqSaQUS34ef7bD31pRdXHe80VTYMFUhXANaLflfkBa5sk1Lrml8krRG2oV
iDM8I9lgIh5SWkpIJP8UCiTUF2xQKCGm2yr92ueikBPW4iUE2wnJ5an73J/0ZS2yEFTVWZfhzdyT
lGSgdYLIXOwFVGnUTbGJ7ovcwf8iXIqvyQPKi6Q7x9cyxZbq3VJnztStriFt4ZqVIc0aB0O+x6aY
2Dgz+GNvv5ePEOuzTFVmOl/wKzuL78EICR9bpPf11OrW+B0GK+Fv4JTwGA5dz/zUYSc8SGMhgrkd
wAW8P4/BotRNwb2YQLw1ycYsoRvBMFczl1jPnj4wceZG9uXoncGmOJsByCyE9tMr7+UHXyI7nIEK
renPTwxNehBUMrmSUWmVA/5ztjeqEGUF2cO/vx1lh7wLUMU01LQuSmh7yJuCwvxFkzKVwy1p24cg
4lfpuYHL5z0fQgnENV60H/RJglg6JsZzUjn9MB5m6V6UBu5o9hLHoX6e6L5H3I4col7C2kAd8xHt
pA2aTPjiZXUZF0iRwDyT1sH8V0HOOmifD0Fh5Rod8B5yNBOOo3qGaw8ySkhqQFqcuyQZU5ksrtOs
CfxEyzvd8ZoME0Qahq08xVllY67WOIwrjN3bvzYu2JUrgu42pLaHYyFeUKovkDMpXUiYV8PvTrI0
lhZ7+kR51Q5FOYNP2ME4bsJMeUY4e/K6lTJM3rA2qT2+ocli87r2Y1cmwMs9/b5Z86WcIQuceu13
HBwiu4a28YNpVo0cSMWUUoWuxlD76Ja4w1aI84Z8o6UEkpYqKUqMpEDyw0TE6f/tEitk/yZbao17
hDis1S5oCIJkfi6cL/RbPj0k2qgRxL+yqN6frbLH+lPliZr0CzGanB8otMC7XcyMwpKU92GRsBdx
x8qbb8b4B80bvDdUJuSrwz/IA+Fg0noFrmZJ6b5MHynH+YJaS/GLOTxIeg6U7ySMMyYoc4I3rV+E
oXi2n7kZ0WNu8JAS+pLGGtkOKc611VRFAqgirl+OAPqZGE559BHZFiWPtaUyuj6/vtmmftQegkxE
FojDoCZ4AF+dx44eP79BA83r0wWjTaEpTJv8VJ2eAnAE/Y7C9DRImmHMSdvI0NAIU2QPgQ4KxPkL
CYmDYQ28XZ1O3VmwmMrlqVOk4hd6gyLxUuQCy8aGsNyhqei0ieftsroLjoMbVGE6IOiQZsnd68j2
k0Jp5mwXOmiRjNl1p7EakWTT6Sk2bHsrdaIx9JH1i0KHr2CQhVz75AHk6a1uy6kD46v+Gf0e9hMk
1ayRaTCtmW2fufk1vDCJBEUdMwsUY8tjlrFz5PHF/sWxW2m9yZ/6nVNZhk9FHA570vZgX8o4obHn
bFG7axLqdjQQenDQ/G5+Kv7sPBx266kDEhUHwRDbpJS9kyuw9uDJBdoqG6o54PoEzCe0lV6WRD/x
IENyWeh46QkGZ8+I2XG4zebx2g1wco8VMziNgu1BLCirShtR7PdpJAwFE2olWQrg5D9CT+YZXhoh
zxxakLXIpjuux9fmzVCFQIdM3hixrJEnp0sK2vTv8nzWEPVUIQKL8YFN92xb7Ky956euWBhxZ6Qe
WJdIJDl0hf0gJFsgl0NGtpEsht/T2Vprsw+asFjSs8qoSKrchcdwYO7qEms9/V9mPXn1Lyw5ZpAb
DS+OUKysGMf1DLl028ik+QmoYOgdbkSuXHJpeDYxaOy+0MDjowDYAbBziGbLuOWrwjWHUOclinJE
OJDevxLmpMhXc6tNWz7zv63PPK35aV6JsxbiWJqt5vUZTGwNaRysNkeMM+8ljYaptgvIOJcFaZ5j
XBbeBVZCzfwoJUHpZGwa347oEh6AlaDB4eaF4TZTi3OR8xvyvukSqktDZJTI7ImiZtxjsnrcWArG
Qd+gzZyZJvXPc4b5E+f3GWRPEHeQNPAZaKDL0t9YMDtOllhpaPBImtP5Tiv70YrN05/NXVDWCYxH
hxpCuYIvNUQ5zVFwII47GkhrNunlJ3Y3ZfD+hPl44QV1VMBHD1IVX37+SuT+hdoHR0ECIC2TJQat
bGrKY+sA6IHVzexvwKS2ZzQA727ZmCrlEzSzIa1rN33C+sGhQ5Gu1Z/UogdXnumxngs+GuxFDbO5
SmMrk6pDsuPB6EuUOo/7c43dY3vb9uzm0Kfr9nPRcsjx4xmFxybe29/dYufBdbqTzIPrM5frzc73
99KGSIJwsbP6gZ+z3XRIqYaN6NvgQaJE80KfIjPJ4IGsROxnQQBoVDkG040d576sdlvu2yHXk6cn
rS+oktRBgUht8P2XAh6cwFOhBmqTfuW827JRJ+6PiM5Krxns8sAkdST2v1rCNC/7fs84W+MXCDEv
giW7NAs5u2J8/zJ6AD9GieCbK1xG89eeulfd0xjx5/2zEL9wK06PtK34qG4o32wyDpeeUt0ctb/u
tGwBqex9Vjei9pSr/3+3aozAJvozLNRAl4KF4F2ooMCJgQ04d0XxQipcT8NInOdkB7QmVl/qIQdo
ZnN24QcHgv43CpHW/HmgZ9wRQ43d3uO2CCQ0Z+mE08X7HpRIcrRQAF7rOhXVJWw68Of7nS5sqMWt
tkqi7e00fTzit69DY4CJ2oMb8d0+XQLxK6z7dHyFXB2aLKGsv2HyZj2MJ16LD2qifECB0MAm1Fjr
ZMBdR4/CAEnL1Vx2dCqY6PTXMVGOi2Gz942zzya8rQ2YkVpoYt/xM1Efa0TUpPBGSu9gwLGkL9uU
5N4u/y7ex63iSPbfl6k193HxSvwHM9d4UyB14BydmBoXps/hGL10gMrGOBKpQaE7rNHq5IgTx7vo
i2blB7l4NeXKKd58Xdpcmbxcgu6DwiOJMmN8MGHJh7B6j1xHf/QJyH80u/3deVAgwjEX4aT5BS0M
c00BIiDR8MmK7vgrjol4b7KUAHDR/xbzxZtoZ4lqvjJnUfiQ5ToAD5QQAShEk642rwmJ1Iiv0dDS
1BlCa+zd0f2/qpAOd4tMzovJX5LP9dIsb4T7SxwFW+7ZZjeeUA9mBh4E+Zsh6pLyS6sqdaCLvJIt
cenlYmSiiq+sXcpnKrCA4DLQUd5flmvHynxfIzqfKtdIFNAq5W8PIot3D94NfleCFrpFEwyw/sH1
m7LFwyjYzLH7fvNhwxcBTa4uQiiTRSvwPm28uNrGQibfulrnpRUgQzsX+gJqNNtzmc6BXffhFw27
X4/8bidBmweBotmO67TKc6aKO/J2JNdeb+TCjZc+xpunDZGPwGPz4Fv79o+slwNoN+WCqcdg1nOy
E3v89/N8q4b6S0h7rZkIcM9JmtY2aLVHPiEcsvW4buPH4HstwuILGucMH8u8NP5EgRTO8JDxFGtT
7y/Rcd+ciHTfxZh6a7wQ0KYY/Aeod1XIhowVq6ZKovSnF7Dgn+W2yapq2dBN0g/DlhAsEfgmzdaq
HKqDDJP3lrsbGaf2GqoQxl/DcPmyTAtjXiaJyJPC2OUNavOPgRTu39JiRgQVRCY+KOZMxXkelLYv
Mu4IG6k8aOgKy9alkXKqufJM0oI5vpO4TdveSQuq8r539P3DpB30eoJmIJuAM1s8LXl54mMCZVeh
Plsy4UtpyqUOw/hTSOC13U23UswHyvWmwhrTGulQqw3+GkLUzZ4PBiGKiHMBAI8U/Vd0xv4cgOtU
1QPx17D0yJlCjAI1Us42Qr1AvUSJi/zaNiEFTRU0TQcJSVlRTmlJl80ihJmSj1NezByOkGt5T2U7
f4c3MhkWEyMVcKampiT2OhTYIywLBGGu0eddnSqMBV2yH+FLz8nNzV6P0kKjGbmCCH4TVd1CRn3U
qs75ytBi47OMWFlGxqKtcaf4KVDO0KbAmkN9yxD35EMufd34repy37smcB82i+NwLk4TKXY01LLk
/SkYUI6bq7HUvELEnliNEXYzx0axhr6Mqm5oGzpvACRtQnBI2sP41k3RXWthtzm0cYiUGQcnsJjY
qXu+ysW+jDyOmSUMulmNqoPhJYkbCHinKQDkobp7r+5mqWdJFEEbkMEvF2RSzXVf2ganoH+/fgLZ
wB/wVVuL2VIMNiZU3HgmQxFiLZgxCtPPcbtmhOd40VuwI4h1n3OMQw0eO+BI8PquQqBzDulZe+Ps
zWSyshOzfwURvUlrt5xt+8KcTjSNTg30+P7tdpCKd2erciZUhRe2+dFbAdXBT5EWA6jxVvZwsdbq
vEWyrgEfm2pJ7LauiU82bTZ2cCk0YIGrQzSk9I3IDxbxMGsHX7Hhryb2UGRW/k67sabh6tEWCYbl
jToWby984SlRmZM9J7YP8sqxRcyuyDkI8fS+lgnTWy/aN2WBrzYSZahYtd6TnHa/DvbIgjlkilhS
BCF53xmS5mO1Pc7Khl9Z9hFrDO/cS34UhgQh1UV5ABSNIVQGIxKLaJzFaVSN+hd4HrC2b4hgC8Wx
Le1ddccdrnmqq36LFpiIXJf2aq3YLaI6V4its8upx67v5MzdDjWU7+EKnkg1B70McHGRuOOTrhOs
eszlLPgkZatIIf/GTBLvcg2DwRPQKIXHQ7WZw8fBaO2zoWiHOSozl9eaGQZNrKzzVfl+vkVh4aFu
wI4VCSw/+GPSbtTAYhnrZnFelbzFS8dmeimC/U1sHM3tAHDmf7qxH8GsK0s6pswNKcZ/RsUc9HyC
DyQr60N8LD+WaBVKpg0qzUd42H9Dn7ltSMZBRh5ZZe4yNA4WQ9vDm5BdpLJ8hkVO7THVPvTUJn1o
v1wftkmXLKw6JXGbBlSPJPxFrjClXpV+LQiPeEuh2w48SL1LJhLAdceEUJhjV0jdFQiRkuLoSUWO
uqCooR47+q5TrPY/QIEjoCMVPb2BRXrvBNFBmh6QJV4HXnHiEoEowPa51l4o7tGCnjRCxPpdE/sS
l0A+UbwF2tXj626dux+XGT19cJV4/ifGd/n++lL+ew++vgvDQ0JXWutlcY1l0DSDfOQaMKL+04CN
HhBLNlekoDd9SoK+E0rdIJpnqoLO8bQ3aMpywZWGhjNjCIFzlmpkNLfrtwD+WLYVzI8VUjg5kT2j
Mq22GSBQ3LyaVRTNPbdQ3xVoEYeU20Fl6mSlpexSbuxKH8oE2RNmQ5Fib/c4iYwGx6w3TsU+7yD+
hnRSPSI5A7ZjHBQLI/OmaloP3op+hO1xGLBMGkZfd51/Fk8avWf/vLCxdUOaVbUHxHCLSjhDj0qc
1rX51ipJxJy1hFSXkOrIvQzLMs0seFS4cgywJse+bcMYxjD1VWoTcvVS5vIah2W/19DScmeu7keI
p8SebdHr8Tjx8miVlrWNLpKHf/HzuSKcxb0spVCoDr+KzPvl4crmpj7RnBNNlSslc9Q67y8yIUdi
n1QWM2YjSOWGWBbBrCks0WymIlT9giGio1m5g8wRcF+gvJ01kcWt3rbAX/Hwkx1avZ9k/SVYBgSh
v3ZNC7bTs+2nHuXw4DjDkKkgp4y2033LX0XZKIoUl2TWvK9E5K/q3dW8+cSsgvs/bATNegdoY2Ee
BFMiqIQukS0jH6SRtQ90LxvPVALb35VQ80a7anisrSfJuK+LJj3w0wYCfJXFLrehuPtWv+qMiH6e
yDRfuy9NIDGTlEae71WOxkh4rgG+fC7lXuQpBECH0W4Z7RxVBpCz/GFSHEwMdONbs+mxU8juEFyg
TwSN8q65ExnYYpLMk34AjqD8Ui5LPj4KLSNOaz9KqAhAjoq6scZU/drc0YE9Dyl5eKYcbPerXzxi
Jy2IfJeh0jDIUqExJ5scfSoRLAUXeBwe6cNkvlRBHJAArAmA0P1YtyHx1d9pddPXYlA74esnJoDb
XzSWXc/1fYkDyEPhUK+n2X+kwurrM0Aqjh+5xqRGFxILAy7qv1AOrgeLTDZAYuOjLqn9S+X9tSA4
kEmPvrsatYD7WOAAaqhUBo++0UyB7me1Tya8NIOIDC5K1QrbMfZyy6nUI2jEIJx1Hcu7dJhTIc5P
7YKx7Tq/p2ybAxE/hdylxuP4056zNY4KbV6Tg7Udzn724MABsNNSJeupItuCzkP/dX19s9NgCYbN
4twKFf1jW8wqKsVEFjlDdKxzBld6R3sbyGPyt02Oe0090h3ThFQPPEsfZzULZW7e1cBzgLTB4C5j
zcCy9lRL/EH9EbWCTsNikSOT6KRZb76qFY/+vK6oRoknw5RMaeiFcqRSIY1cT/jRPNT9AUw9iUMi
ucBjewm7n7uTnpv6sx0o/Q/sXuUJCwc3s1s/cURid3N4iRtzsxG7GAN6v5dKFdCeJtbd2wB5JqsH
XggVj8OQ1wud9Wf6n4GPaz881/OzcBjAc3/4Jcfp8vkiA+ZMlEyi+sXNI0kSkrojxXklggJejzbO
VzedoCqdtBHeF24eEdnBaIK2kW1kxfNTxY+Mt4vPQ4IQslsKbv9QxmhZNOc5NK6lUPbZBq/+tByP
GPyrhxe6ayjVliGAcLKRnJiT2FdBSRXrBqqRTa1+IcbHSqlnMNSyMJfPz/tUXC1OyNvSN6JegubA
gMpKPM6t60TqqZH3RwIBTpExgLOmvtbRUpiBAflk0Q4aH2+lkKdzaIp/VplWVt7q4KhpZY8CsZka
O8BkHxIfpRTpLqmXbXOLSVjeKxrba30D4sFhzffv7eY4Zq/V6Dw2LfJpVMs/Pv13UyyQpW3OxLXa
f6HgC72PxGDUpHCHURBQoRtGVEZU4MGYChdwFe9YZUa5tWUsgbGS/peS9/wwuOgdokV9qzhE6wdu
U24Mnxir6VPYOIZ83RtvSlR32p9g7uhrZwOuenOJqYugIe2C09Vd+n6p5zyc81T/v0m3q1uL7gC0
rTONUZPnwqZwYoXzk/h8w6qFetjEZj4eAtrA4ptLePyV2Oy4Dt7jeuN3aMlJ5XPyVfb9PTI80wMU
VN6cEeZzZClxzpYRKMXX/aZDuvBUrvTvpls2Useuo6JFbciyowpwUebEGD9O8y1j5rjkVYX0afA4
0KmCT8EieJC87Sxt+CSb5/d5KZtxrQP4OL+YR03BOc0xoaXDBWf6LH6X3x0fl4GTQR/7qkNbPtKr
s5OF6IeAfJGbKRUc+Q7x8FFzEvxjymn4wjdgYC/CfU1CT0m54eq0XisMYYBKaki/iXQqhvE9cBI0
Ki5eEqhNKbSWD0uDoWAawOuXLePKqlCMqo0EToKlxA78HQKGABeSE+EBSq9/kgUufiGprCaQQpJW
BgLMqVNiM9XGXvswVA8W/rOeRQ7sikwefv4R//i+K9022gxwaOyY0PQnSK5fSUndIMJfTlYhbdkl
Dz23OVtZ4W2Y6UDN7qZ4VgaulQUZekC4ibTClc9Z2VBmADRO+XxzgUq1mrfkaqsQF6ME0CQsIHEQ
c0ovkzS0uQT/UkCe7Y68VorldFA/u1a1N6EsDfTGECyJLw9ibEiKpUzPqljsSWx0+PDK2VgFstzz
0q/P6KFegaWl8tZrPN/dFHgk5BF2sHDgtnmXBRIN1mfL0mua6LiKl6Rgfn3sHjqdCS2T02JkfX9/
YZHll2kPcgu4hO9LUJmVoEex1HtcA+l40OoxoDAFeuK9k8L/HFsj7vL8I0hk5dEh5PVAuYRZoTFG
6Hrs2yiqfMBmC7504+lBgZkcDGy2MK77Lj2yAOgCxcAAK7kjAk4SdorEke6Z5qIlPpWlexlNuQeH
cacmFOvccNq7qDucC51srAVC+knD92OT/UuRYnGo8Zl0VAsr1iQ6McffQSugpYvbZUE5CELkJZrn
d54NzqTf+iUbk714bg0Vf52dsNtFth+GO9eWYhOGRrdcDAd7CEShtmbnOhM91PVhJpaW9SGhmhE4
AUEx7tji9wPAzXrzW5ctziPIWYw7PIHuc3BM6IKkFDPttw65V5dngYKNZNXSbiJI1ZSxFZTMEPWg
bFmSbfCLuS0LxvgFfeIejwnBeqf3By0sjKtnSJJvF+3R6aopWY26tXf5mgDTtHA8ZVugwmo1CgAf
y7cn6cy35hxpeYzl4S7AabzzaJ8tA2cYXkewQ9A7In2DRB6cyitS/rP20jC94q+T1m4Dp4qnL/xV
QZtidchibuoo/TV0tM3oPCnbflguo61tpDvAJN3ZGBR9hee6jOnzF8AjhlwfvCK0B7AnxSqTophZ
pzW0eNjPrx3twoLRz8VzgHBem7BxG0b01qqYH6enNchVRsUjjHXL/uPeXV0EnDMyhDwwnG/4HepY
hsk7QnTFyLJwCMI7rqdrnl2SPilNJhGDsHALA1ZfBXdH4gRkBSDd8Suzb3/sgI6/e3JGOZPuurAA
KBXOmIDtmqzR+P2CDXz/xYQ21t/C1ij/4NhL8xaPss9X5Z/2onnl0gQN3DyUz8AeDjn4SoeiW7mO
H2YQMYFangcuxVUrWnsYQUmog+0MCSMbZJfMZiQ1qthHKu9iQGJ+eR73bLzM/irBh+Na+y9uruOA
smZRPOczJG7YbW5DU8ovKRwCWfaMccwJ91tcOpV6KngnMx/tX9jd4iPrEtYzIFffx2k9Y2t8uYCs
Yax1TTR1TeAnhEebPCUxarZ56dHuBOEFYHeYMccQvc6ZamjDvIavMkBHlyR+ZzUErupe+EmuxbNM
V7vYenpERd7Qf/fA2saAml9wo9wLwirLa0jJAOrJ86/GV/D+arwRq0JHnAtnJz9WhDOWhqL+inBa
g5m7KB5Sqv6LwEeK91qJVIyZhZqqYmU/sP95Qftlc6ElY2NE67w03Eh/P3awJWo8zzyINhPNlsb9
sBNEn4Suv04z7Au4l1axDohryWW2Q1HHL7FVsYYUSlUOFpOrX7nS+uD/xE5UTo74HhxRscnUtbjn
ufpkkkHlDUHLU26O7iMiELlmNmssHYG1ubax6+EXPR05SLURYdE/dn97GHb7tFoO9qojZFXEvDBU
MCr1kOA4ol3WVu+NRTsJggWc3xEwcb+7UzgapVKFkCdjtikKtlR/QVTas7bQiKhoHh/2MqQjmpiq
mpXsblg9tXRt/3Y5aS6BoGsUnnBDUy4nEM2uxiPjW04WIUcwTcw2us3jsTaY83HkoMBYx0CXy10n
vuJ7CaUnvIkmZ/5TusKPUlQpHSDEEYWTI70A6SwhF7u0feCWLC9XJdG/0dGn9EyO3J5fMfYQ4WO1
i9gc1dl4zOvNyaElkU+3bHGv9Zrnh/V5e/lJOnas69OoPtu4j6bTLbysy2M1ZFg/KTYcARRo3ilt
FIU+/s79nGXMu8EveeljVc8v7WGpNnMTIn6iw7x6nngjWU9w7jEtXS8IIT0l1QPz28XdKI1QTiOz
3yquo+YJ8Di/3RPV96FSUtCby7v/THGI0Bjw7o/SQhV3TaHGINXwiI80cmeGzQLy2A9v1IrOwtEn
7PlBg9AacrF9mPzPO3siYZIzsuaBKeqHGHJo05it6Ld1mSo/LTQi761P0S4PJmemEzT7obbfx304
SMd0lLXM/t0jQGOpHm28NBgTnfhRF5thQlIBS7OXv7ckXk2czM7xLEBez0TJotnmuD/m5zf8500v
bk/ulZY2/7OBkC6krftsnTC7LrzMfs+KRp4sSS/CjvZyr8Awy9YZggFdunuNPhRFRm+lxMI9n+t0
vLkxJmsLVNjiCK2eGtVkmF4xtQOVUPcMHSbtp5JKhvkYiwhRkf7o5OX4Nl4Yv2PZCIPAyuyjgdLo
UR3+ljjd15tIXyEDbAhm1bD+uJnJ1apLy4r7KrVgOSae5DpDFlXg3T9msTmf3QSQe8K+SyxFYFYj
l9K7bicGRiJgkfPrL/9GlDc1jXg+a3XCo9gToboaDOnCK3rH0xI7RQ/fxlCwtepgBoqWgtwXlR82
L7WIG3376GLRWbXNNLYAVA0vv+/djXr70I/Q6tVO7pL9GqrbzForPASdYZrWKdnZcKltMKt76UL4
/8Vzssl4oXM34lu7TrIS4hg390Hk2x6pyulEaey0sV7YChqJRANSUbEKUfXKEnOtxb2iB/FtItJg
iQvzeU2RIVnYZkZRg4z351m4niZRKDhPvBzLRbFpUHjMsnBlyGTtGYfcuNZefekeoIslLP2BWmCx
Su94fZNy8Gh48c7jHzBQTwPDmUbNxk9wxI7tlwXAvAQvyBhrxfKByuRMK/HC5u65KmcFehdS1XsQ
j1q2ylPLoql8rSRJEWLt3Skt8v70TCf2jYX4MG7dTzhxcZHgDekdrHZpW5NN8ghjgvkHyGNgbzgH
FOmLW8yl5CW02Aryr7/ZKYn0yeMoOEiru78Q0QWMe+tJY2FB3b4bsr1xq8A5RaGkOPLB7aM7pOmt
X6wZQxv3ZWPy/KWngwRS6thHeW8dKddhMwYBGunoFmrOzJzovUeGtuPHfzVHOJoeNNOz/iqHs6dM
UurjniLVJxNMKvOHORnCVbcvQ05QT/As0LmscDXRjp782aYCinS2T7RcBzxqQ44nQ4WsQQW10yA0
zeASJGchlyabg3riHxSDSEJfP+SuoR999HhEX3QIDmTTfiZRgGYTHF/xwJoEaoGCPhxtV2XQkhkS
SS9tiJc4G9nI0dF1xXYIyOEXD8r495qJxHRpAplo/dmCXxAwW0IEJBkrLSFggt+Q0OBT0BCgDu13
LlPqQ/TBU0Xe/ligafujmevJWdmyKd910boqg931sAxSs8f+sXq/zkFoHgTw3OkEkeSZPS+1OTZa
55RzjxjAoVXJQvHPLNI6En01f8Z3G8CxTnKy0Qt8i3psVAZBvY74M9SSVmWR2Ykr36f1yPyKbITQ
bSL4dMcuHBQz0gcgLFT9uDHRQmiVlGwKqgpPs5QI6/3FKwGDztx1PY4P41FOSHSiRNbncwtcWUKJ
JCa6VSUTnfZUbDtY5mrtJCRuRSsxho/oU+yyFaJNa3BYhHpVvVTeQX28Kwi3YKcYJsLcPZJbTGJv
kalNqM0Rd931M1nUk8QFqqZ35Ak3Jk3Zg+/0DtC1Z8maUcVlYtBz9ERAdnCAXPr4ytqE1kWjVG9f
OxP7nUBQtj2cquFlUnm34lwFUTP0nbFg/t4u1dWVvoo9fguYYQveYdNqLZo2MAirIBZg5b+hreZg
t0sATISImBQcK90L37aovP8NF0kuZ8XATExjn0KtwnAhDU5Xulsax0LSCZgKCCrpSRV66hOtVF55
oCMo0Qi62uUVoni/0hTMvdwcVwDPO6n5VbVTm4Hcrb3V52Jwgeahuo5fvPMoj2jJxiWzdSaRVKMi
zf1fSA2PUR1QFRa7vN4fa/Y4U2tdhqIbGXNi/4IVmcEPXA8NLPewmWROzyenCJ77BEFRjLQLnH/9
uNT0kSGzjWs5qA3l1w53vvSrMJMivGkzluPFJ9Y/UbNkwfCv8zO3lf2HKkmdD58LxDgBq9QY1IRT
7S8ULts7za1m5dtYnU+cl9gqVxvierbWuGBLlc9gVAWjSW9LdcLia2EqG0tIPD07VxlwtCxGV2C4
uuCJ9ScT3v/21afURLurDTGoa7Bj3QkMTfvw9G1WOt/wp4p+XiyNmIeFdZgoWPowxrSzMbq569Wl
0FEZP+/UGAd8KTe9LDYX2n7y6n5VHyueGStfGOITqNmmdM/ZS0iF0ywKZ/YSbzBPjqMExFIdhR0x
PetiwgTG/qFHRezknjDpZffzICC1gXLx7XShYNIAdpLDSye2GF/mTNZcCqBedmMwVFBzNiiI/gju
QqNmWZvszE508HVU3FuITkwuHES9An92tP4WhIwIYoZqkbLfdkLzEoj/ZEVR7As0R+cJEbAeymeN
gbcFXOLYA4rjy9gfDuU7aAnoZk7MCKZYKIiZu691Hr81Ylqw5ktCZ/HM928rqy3Cx3XJiXMBRRiz
Q0c5lz7efHkOXRdGaNEwedAnb7St9gWz42pQSFue9jH5uaC4rdJAzL9s3LB8QLk4rmtF7ing+dOW
DzwtWiXAWe31AXYEU/iPiQfO3begUR3mougbmKhXDgqmgu4pckDFALOkyvc8k2spTEww0+QyHTbu
mpARrBczMCgqAYY8TQHRJAxaqVuWcraqgiodATVXsRUolpn2LRdubQYepG7GEQgua7KlsqNyeDeH
d9Gf+F3JUjctPmB4cjG1XDcUj8P0InoH2t2miunw8hKcg4j53i+BtKvIaTDBXiFFWAoxWkWeTzig
Z6+4DmwDnIlNscuO23yF/zuF07NFythopbgxCRkwGNT+VSbNWJrvQ4AOlGp66/i9eakcT2h/oF/L
JvVRyvVv1YHDfW4pousa6TsbAV9FJd19gj1mxAVKMDrLg74ZdgErBEm/ra8t94RsxKZ0Y/ypUkLJ
edwQO1omP2OxgP2sDRA2s3O1dOopRT5GZp+rjaGR9rst4Adqo7uB9joxFZCP8Fem7U3EoFM6T125
WsWeZEoqxiUEm6NKgxdscd27V7UnkwjrZ2tOc1s8ktHtOOFW1ijl6ukaWmEmZmnMrrFsABnw2n5H
wD4QpTD3aEn8NhjkkE/cgoQIfkh0yjIlpZPlPI2NRwQcXiXNSFUTTl7fBLnx5MUyqJk63S7vWTYa
NkQjnSmfIw6qAWxA4/LpXydWg86hQ+6KPBpx5bH4fqgwO/V+fOYXPbtPvUsX5AY2SOR5FPFaLFv6
OvYvTV5cWgjrUYZ33iLmmd82p1yCkjApwUkItyXpiaqSdJBYa9SRz+ipvOOhYajC5JbxeiIog6pV
gKB3U3Qi9TJxllT2tu6NW7y7G3rr42DIpnT6qGEJs8GRkAowmk8Mbl7TkDzcH7oRyL+OXRYlrbyY
hQtnZnFl0BFEdA54Le7EDhMw8d1IFLku1ZIckR4VBHC6DnNyOhu/FayFh7PVPqV78dBAg+6FVONE
x0iamDnwj1taM6OERwFQGnkWb2QV+LPo7o8Wzolemoc0E2o5iYMWobiQa42w+WBsg3mfP5KbFLrf
bT8msYxql7bl4MFm6xhK1sDEPgruynrJ+8CP8+Zd12/3/J5HPhKdq2okQsxyEr7lpRex45NFgRO+
/zWGNqZ10hrTOnlN63yoeQH5f3Fh77lyNplEz3xC8UzmruuiHWSxjCNiED2hYnOXG3edoaKsXtHT
VK/zvgUj1nU9QnNTKNHGKX31svIXws6ZSEm/HjbKXpSCaGSmD7jZu6NDGkOFAra0gi0Zu6L2XoZG
EXLX7X8QjEICJO35BiIA2zfbXm9+Wg8ONGZ8usUKnQFL/KxTRLTwiOSRkfQkcgz0DRu3TMFxZHh1
lViYMc4wEjpwNYIGgjTxG1h26a3MSJqBrUx8ngw4ytu/bgb89YcUA2hsfUybqLGrmmFxWV0V49L4
Ow67B8rXGbMno9jNJ5ysfkDonUj/tj9j3JaoT+p8QaBQ8aMjyBkBSPflHldc3Tt28Xdp5YKV/02R
MBSx2W41HBM4DihQuuQiL2csUo05uUezLt4AfugM6j3S0crHFSaQeC4CT41G3wObAE0GfTM7XpEW
3HS9mNSmQszwEB+vrA6Oe2IVqWUH+xFXcfCZmA0Cspk/zLezpoQkO3TNMJGEdsIZ3Q6mz2RtlT+l
8v/tf4OXjnUK30jMmnBgjiBBwvOwwhCpWcHiTjpHQuQU4fV6Z03tI8IftjBhR7gMbwGZpgx1vE/W
xmzVAE6YT2vjiH/m11NP+TIYSQczBsa+H1zo8CACJitCo/4L7+p7JurCrRxoo21DTtvbeFddYjbn
kLz5/ViQRf6FnJEl53TMeAbn8xR7bCnOjKfi+JL9miLEJZ679JM0+pFDrRsmnQcMAphtWWNGX5r7
qRCLd8OiWSeQVm4IQZ0tItrR5XI05r1MY6H+R1URpOY5/mMR6XgtsnNSGl8nQaKh84ePJI8o1M5G
MmlnohkpX7bSOqD+MJeIXk6CXhxR+UL/Na4b/r6RrbVstdLctgCDUIXE7km/O4FxI4gmynhrbYrp
hwc46rEhRklxN3GoyHEc3Z2JpPGP6PNxo4AtOBGi1QZEQ1ysxDcivRRtCeGqmaoYcvhOq3rIU/9R
g+0xlxcWVkwouYKbjjzVtk8MepF4g3O37e9axWZ+74fRDS2Gmctekmmybql5Riy98AHnrpUlmItW
4UMP38ChRehnn4Lslc1y/xDcrspgJHsdXmogW46F8Zt62wW74DpIKd6iAbsV5iHOF3vDaBoc09ij
pC3foSenXN4TRGkzUvkNry2hXyMqKqxeERkpA+gN+NNIOc+6oO4uI7VpOJtaf0y2XctKxFDlSUSY
T9i/O7dfaOvWM2LvYSD0cpz1p9RV/LbPG26LyEDFawUwj5b+ZfVWB0IpiHUNQCxC8DV8AA9cZiIE
vfHMoYbFH6hWHV2Ut9Z4n9TJgCmChqA+l9qlearhj7pba3yOPbjoipVsm7ToGYY/pCqQ02WVYkCL
vsPGPK+rU1/h16dhERH17partdZyzjP1qL4acHaHUIDyuXGiBrnr3dQvQNPrhZvHBlqWehlXl5jM
XBjNFxTJYJISXkWTRCfpPpb82dZkC29y+QTDPVOnYH+7TNoYtNAJ3v3Y4bUkLYZw7BHDOh8rRvh/
ImeluseNX/fVcrGrGJULTLWAWLInYg/1iRky0xLKhboGM8/xkgLud4PebVZS+ESlpcsy8eaxMfWi
trQnbIquQhmCYl93zKYhPbNTvu9zzW/huAPQzPpOWgFCKaOhNRHY1VcijsnPGwew/WVg7kLDJ7QR
Yu7HLAgtpxxlL0ojBp4Dy0/FErjp+VdIN5PrAMDMC/akS6xGelV/eSQluY7A9wGdKJcreX0cID0+
0rs2c4nXknn+MvKr6R2E7EpAguYOWlUXcsy72/BuM3ZjB1VnZEPvaoVsmO6FrWmu79wArtcsqTaH
gSWcb5WBABuqr28aTovKq51r2DFVCIC5mSzyuPh5hElVVsTRPlSW2zFS7vM9otk5sC5hgBzEZFYy
FXvcFr/wZf+G5MEZNs9WXAOJcdjBxGhL3jXJz7IQarePnIkW1t9Nmhoj2BlqcVZgCaQQL4S7vaex
pmEbeLGkQreB5vuFUV8gGK1jhO6KM4u5j5/qDfEU33Azipf6bDnSC7yRzLkNV3STDHJDc28dhlGg
ZblEn1SzW4Lr1wCQSxKELFLf/6yRvSD6GJzxfhGjMaCGnzfTK6UvC5PfwT7cvLMcnik98ziz/yGM
YPVzLxlD4EwvJJbiXz4FtyI/SKFieHuAcm9YEawLOXzoRVztpBW0wnAB8thNZJIO8O48lQ0SAxg/
mV4zvyg5bP+u9DwmpUGhgWYC91IIfxFqOjjwGunCoHqocfXDgyoVFLU/L7Gc1nLfpSevq9hglSuX
yadwX6fV/KWVcc89F8uG8vhvVJIn864w7PzstAkAHE/fF+G6NJ0Bq7IVDO7D4Lp4jFi9tAOf4UQq
KU8KQrPgRTMJOhC+dBioN+fSJqh2kyRjHZZ2jlatLHPHZzNR57cg3O7RRIO0lFgFT2Yo6QRFFdiM
MsVwHJCJKgQocwH5lB3aS9mvtvwYFiO/WOm/wiTCUmeerhIA50M+pJTUhPGbfuGd84XjXWg/ysfo
8GOzCDJlbEfVhfiIczjxUya3eolpla+ScEgHDIVAfNBXpViTm0dSYffOl2zUBCpHIRmE8DbbILC5
FW46H+ebqhEqPbY0ZSsh1OvQkGdIaUcITxzIzfoYA62WJ4JuO22WNWrdbN1KkzOMo+n7IvJE2ABF
0QBtrW23yCWqTmgc6rVZ6j8p2qMcxeTjfwkjQzCxZF82tUShiW51GSyeAIOCzh/beyis0or4soVg
AJiBsyQxUAOILGyker415VWhiC0MMTgUtpz8TxIFP/vRsrYW0xsgi8X3342smVvJfd3lDzjNGxB6
fC/VHuD6YQEq4SKdjy6Bb/Ab5q8UklhOvuuQVJgxBiGB7LIMjGxihFbjUYbARFyEzqvhhop96v8t
1XIFrECYSVLQCT3qYZ/azb68+gAVnjXjdb5im8psmhAx2wv/MGP+8oqKi8hyY2T4MpQmJvzuWm0w
QPtnMRCvscXW0iRhjLn4HS1B01f+AazikqeeBHr6QcwT7JWZ5EQ7/JR2x0pBOorY3GLy3nm3XvMe
wQjc4cNL4i1kr4ZNYmE5LmjwoAQ25JSJO3fsGL6Nw+l1yv/oh7NQvTNf4CjPaQ7bjE1A3XUbrp/h
BN0Ff1uY7z7yfkKMqgz1NRBSSv7DLiERFi110y6M3LZThQwGURyG+EGw846mGtoPfbyaEZVRniha
DjHaWuXq5nQdhmMVDBReh7JedHP7p1ZnPO2wk+aWpo6mb005dXh3IH7b83p+2jogsw3xCJQSxbdK
DXkwsTmpl4r3+8n6pKgTQPapASLj4hMcwEc9OSDuU9cAEGn2hBYvnpBtG1TDDHCdRMaXKPZ7+71u
eEyPT5Th9EZiLJ19i9oFUMmTJWYZCHH9iXnoX+P/JjCUL17YzsKzDoALeTwg+PwwuKx6kHUUJJwb
nzQHAqqlUVtsSIcaR5LMWQkfJKGVsCzdNVD0xucmm+D+2qUhtRiaTRHnT31zwz+BywS3yrEsKYld
w+koAUuci8ZqTjNxI7olQuJOtHRW0ORlwvRToTBse1WaYXUqWqnqgByLeKI34wYqdt9WS80bbFoh
niD/I+r6j8RKyAgyZmEtwDkUrETqEF1xmkcYsjQ2D2impjZL2ey13vO/SjBYS2Ia5e7ut6Ews48T
sVikznIc3nDTklirJCm0gEda5lwvDVo77fTwclQ+Qf0mAeB7SuJpp1DcPpAnX+Jps75saNnOagT+
tjhCGZrC00tu4xbp6wEEYGogOAgpDUQBA62RnU3CAVKtZiFfBBGK5Kgk357F4RUSa2XP+ASsVgua
7qFiMk9jlxn463R2RLsrsJBNu6daa2atX/4c3cSVI3KN4gSdSO/99crP2Z5I22I5TuWm+aqx28wo
tjZAheN+P0wpmCTQGX/nDgFJe1YSdApDmE21XWQ2p5LKP8O+t7E9j5IX5afCJhQ7RmClUIZ6Drdc
4C6uJFKRaTqzrizVxKEKnslkPH37XqTN0OuEethr+XbhJneAF3dAAhfY/wdnVfFy5rrylgt2/XrN
CPmhtOS/SruojZvYH0uNkK4yP1cwaGsBqFmfP0N0huCtj0qSxntkZv763eQ3VSNznwo5X4/VbGND
2cPpUjCNStqPfrlWPLLpkKChQiobS0O/DTqj8EnQ9MYI+5R0ZGhZR+VfOPNOrtBEimkHxjIifWI6
H108JgLjjXdA5jdm4EbfXlrd4roBSF3P0LlDiJHacZqEtsHgMdyr4yct5qHxF2WmCFycGmTWdVwH
9yMGDb4vOkKyAo9MlKLFz/0u7gcVw8+RvEKW3C6ACqa/D3HHvPPVDKsTNGfss6W+NW2EBdC58qqY
hXcAbvB/JQEPedKjXJYgfiQoke77FoueS8BLyYwhby1Ncq7Bbs3GA1PP4+8ZeCgCw51BYcmcs3bF
xleiqsseFJqqfBzXgAWc/JHUJmXLW49yFqpXRyCMDGGW5+4S/hMq6pOtsUVlpoYyi6wRdOODS32x
L4j1cZqR2FT9qheW5i+Yj4l0qSKaRiDoS5YeLT+5f/P1FvZRY7WvRxyzF6X0csYiidjz2CesQgfk
tWvxPPxn0Nm+vKJTf6JdOZ2ryu6hWbePKo1RwsdrByAC6Xf3UPMvvTfE2UtBkBImJfZ5LFDfOLfY
sgyeogeGKKXl1Jqf+/8Y19+YCqOUDApTlxFe0F3AHYR1Cfmcdmmiv3RT2v4jiZLlXfjch68wE10H
R4XpzRlnffeQm9K4VfsTo/4FLRVMus8R9au3qM332tcB4f2rgcRfJ1EiF0QPXf56l39X80iyEcpf
CBpFUZg4bgQ9jwVh669xo+K30y/0KRbhOqs2haeqWfqY4Jsj7UweV91XGR5dojokEFdZASX6jdNu
Odop/LYa0/v8gHjTCVrsDUqeh9bXVxTUjJsgYvOMw4kclQF80ksQfz4b4hU09oF056Du5/pq9zvp
Wh+rx2n4qQ/BDdvT0NJRZvi9nB5XGDHip5+bJXMWB21Gky81weFT58cVLvWhfyhWT1lBHSuG8K/c
Y5jA2gu3WGmMKvtbEWlaazj4Vw4B7Zya3sNs1knuITZij507lTWHsUDJPQ6pnSjOICM4UHlNeEoN
6ZRYX/hL0OGLAa1EUMmvG307Aa2IyW66FztyBWi5iIMkdPO5xcEh/Pee/NpdaZprXOWXf1Dexq2c
FziB/FFcvpsxOZ2WVpKf9Ixiwohokzsw+MamSRipIXfpGeA6f9o9oeJKyPZ2w4k8rz9NRX/Q+0wh
t9s1+TePTQgWQcJ4OiQy0PUB9MaIsQabcrC4uDLNpFavdjrcw5kcuYBBNj6kxve/DyHhijGEy84x
X2fsmki6ZOSGZ45SLIxMbmS+YeD7zd9sq9HqwBDB/Q1moTSvELHYOdM69/OgFwIpSgCPKSM+ppxX
zOlAZV5E/0IrjlfRhb9pBfnnuzPkqAtg4XzGWZD2PIrRGACt4OiRQb6+sBpHziJauJgWACz0qpul
enm912Os8tTbKqxU8Qa+IJL0MtMNPFFMFgUOBXPoViCtdfsXxOMPRrFwwX4Vn/okmShs7626z4i4
65d25lkAtGss7kf9KanmA4uq0/e+otg3SOh4WWP36esPXnNhHyWv6hzK6iK7T7bPHNsEJg5Qh2Qc
Yc2JWGWiL1vmdvuuOCtGhhN59SDuFmsKMCZjDNSal2GrKLfkJ2esqhp25MW79HyA6Ry+YtpR+XIe
h4IHOcXeizWlpjaoZsfEmaxtLvcUECiIi2bcPu0ASIx9KJ/2kK86W19JMEjcgiM/vdbR6uzPTLTf
S4OhXymvpmZTiJ1I59Jnvie1BI6MeZEmdZXwYw8Ct7EeWG98scHaAKOfUe2gTQC4qpQeobNDlXpD
0AvcsyZVZhDJDOyzNl6okOtOWJ53xsvlvVz5yuHzlKe2pTZFHZbX/yUTBpEPt56WefRrFE6Iwwrk
H2PnYeM2Z1l2pc2vLWotV4EWe/YLF2PcOZSxAIwrQL9XPpPMmqkymJoCJp+H4WaM+ma6LFIT6nqZ
Xx0DHHlfuKK5/Fr8+H1Tg7cTMFBA0XfPVp62C3lyDzQJpdi8brzKp3bNlgh6kvY9cSYHT4gkqtBF
nr92balLMb0WfedMdFlPndGv3OscoGi7ms0BKnNxlO+FeGn3NXGZEUjZpGIzTobaMPj717uY5635
xrsaEqN6bZDTZYjxIBzAbFJW+5a8+TPAry3P/HZVLhtus+wXsA6dUcPxNyPFzmn+YWBndjWJJs1w
M8GyBKexWtQIFDPlKuvx6u5DlMS+v22DWxcu/KDfNSvbaoZAh2RmogpftWSxii1CjWzzV0ekj5SU
/ZuDH/DDon7cWmlNcVjabo6s/FvJ59lhXPozwWhtMbNbeN0I58036aRUIY8YJsvFaHJv6UUIttp7
WVdFX4CSduBxIWiVthYJDZX3IlH08xzJMSn+NK2NEXcrn9pUbsO8hoCl9BxtFWY3BSpB/UivYAHr
J8Lo38aF4lEZ/I+piANAKasMAYTa7vrluOwyzNsR5odYO+JsYGZ5FILdjNmHqUoOqbJQKgGimgZG
jCZn8RwwI0oUIgFZ1xomq/UBYy1+dcNoCFieHK0mbtwJvNLZv3P/mQD7X2s+5WELHohIozaUBtvp
4rd25BSrq/gDHJYPJtIRLHsm6L3DbeZ9P/zngFL8oZniPYU36bdpoCAHhHYm1Z2fElvGZnwX5EVU
wXUYQPvvdwZFxeTwGYqSx1HOhMjw8D8oekLlYOr0gEAto8gIW5RnY+q7Ri8Uhq6bv/C+Uv7VAzi1
KWfTTSGPyySHbNlVEu5GFFiaFpE8R1tICX8rXobsunNKvf+DJh2krPqDXqCNcE2TK8/ovOSktV8r
quL4ypC4ocmt1ehF1/5NdLl+uRLYyvp1jRsB/JIAGS9PIYgWIhXXNER+gIeTMwQ7b+zvvXCPxhRF
w/yH9pSnMmTLJ5XfgKvKUkSQ74d1LdamzRBdJjuyzF0/mIsAQuOhpYNpWTn8SAMLFmOqlPuhA2OI
dkyvMMoPXs+0GZESQgbeDANLbKUe0ZQU9KHXtBNa3hxVbAVuhnjUQz62HDhVzFFFaerbcjGeTG84
ulaINpw0PWGv8wY+Pohu3BAwTxLCs34IYhjWsWRQ2uwgKUnODx26nfuuriwFc0utX+VVSF+G7WP9
/Zm9X5AoYKerXDeK/pwB0Qp0vetbwrIZbqGFw3wPO0k+UknjXagw//6tmswhgCbRytjPjxMa2yP9
Jp8me+wtGmVoNg+Aq4MzZRUGdLGbzca+aVLeDBZR5pW01WLj/J0is2vGHJGsxTenk2qX8nlAFpZ8
o/36N0A6hHNzOw1CqNrhhhvrN77/7eFTi/SSnwUx3cl/TcBSh7d4OP2jhDzEhHbz98rGiw4jJKid
PdvCSZt278zgLkzJ92weF3EnaaPHuxjQP6DoD7nnTqq+ylXNVClbYPLbfeC9H3LzhtrXeDmYW1ao
E/ncBUnEvNIt1CcoR3gxeC3XC/cvrfgNAHr960zwm10AzB+SZuJ5xc3+Aeu80xN3WWxnjpdBIGxo
I8XoZQdPdXTKtknYQkUW5WchixZtJUoHs3jQ3wXmGjmPO0ykJNe4OuYHqQoPxVFk4Uer7aa8Qg9o
xwiQfcZWcdxP+x75K3+uYi3QhRGxWxTTY7GGLOnTAFmOZD5/uc9l3sAiPDonpUyUxYDK5DO/5mEX
Jk7I7kebgc9+bzawrOmgYniMeGb+F5KbFpnntSyXZc42moh/2BogEcFuPC5e/kg6YpLEsuJn1xFm
bxGWkVZdfN+9FTg8Tcjyb83sBdKcZrXGlVoRCQQ522l8anjT+xTrrJU60P9F5TTPukTpcYO6338L
CfFa7nTl6//ycm4ZWm3z5KY3soZ8tLIz2gjx1KdSSKirz1DEuCnXd0z4puVdRbEk98ZrWEwmyvbw
7b64bey4MyKfC6f9a8TYVc6jS1CnDQYJdOc51NoawYClWmfw9y6jexwC8ddHewOvCXynHpG00FU3
1UFvYbK58xG3/543l59rJ12/Tzfogx6YsKmedPWirkeHQvOV7o0KWeeVRScj4A/ow0qQQOS34F7y
8mtdpU3MbXFzOxup508QS3XJR824GNyjde83L0PYgC7QYknd3x8DZxq98p86AFdIgMg1uV/cD1Ko
5vo5wHFREGC2IIIdAFa19YaR7vixGucTXU4pZCXq2PYrbYJPy1fYSd1/oCbp6CDgiW946A5fiWVY
DXb+RJXgXmAqfEmcysgrqFzecs7Rf/ZdiMN+UL+LKLJRWHlutdJT6aW7POQBEGl9tE5XgP+a/J6J
ymhLD20xfk8gM887dEFG5xHQRLRErOFra18ppsJOW1eU975QFbrkvMZiwLXUM/Nb35CmHS2pETfl
kzOKRTNDSKdtnRwyqW8rorQygm9nPVY9mDyzEYHYbRWLSyMtO2h0NcDItlaH4/kw/D2jIYmlZ007
IhncQLk+F+8afJM/UvFxaq2r2MiK0r2iWzgRnujlpEiWAg+KZLy7+m6qVT5Rc7t9Tw80t5/hlRfk
MEHjRe1ASjn8rptP8GP9CW8JWcXR3dfelJXFgtEzxjrvt/4qc7KTawAxKwC5a7SgDKNkA7tIJzdF
SHrCLHNrXDincLkcN59KsacD5F+o/zVvilpgpx/uPJYAw74hDNMYHmdoR2am2Ho283wpilLvJy+I
tSl3hySIfLtNHk3GMvAd+DZZa/RdQFuikhz2VAF4hpFJcvkW++p9kUQpDesbJNuZagIBPvza5eqh
FjB79Y1M4y0EhJMpQmu/Zzbo6wAXChFvn0eh5Fn5DA75wTugSom5RDusYE/f5D60Ve/pdf4RVmKx
5NdpnAZOWs8fjC45VxkvftBJSvfkCICDnlaR+wmY+m5gboCdTrff9byZM88+qf7Hlwkh4lK6WTfu
CTQ4yDwmBC5oXclDjldc0MrJJ9Fh37gknzqchJ+XuuOgtixyZAaNmjLkdtqFBJXZfyNos+dQaEOr
fRTsEOha9Yw3qDIC831I36hGieyTr09tq6qUA7Ix3tp+wf5kJixmQHCHA6km4+i1mO+wONtEMFI5
AhGX4xgwxtfjK+v3gHNOFWisLGFp3PwExXDySASpiQ312zAueAXhtu95PRdevL4xhB6bmSi9Fizc
tD4MQPxdRDfGCLZey6wQoCXyEfFiBcxGs0NXKz+4oA7uQE6C6Wljo/apUGQS2c5aUEsKtToccKtB
l2n3kD76yCBbxYyEJpSl9irMKQILDBKIdOQvmh53G/fX4PK7sMkdD6rmO0VCMKoS2NZCkJuiRh5V
6GdIaQbBdvz/7p+5uadLeJH0ci94EE78NkdlayGv6/BHXOqlJEUX2rHJ52LEF4sV12qucwYQ/QtF
DJq/AGPkcNZjS1Qnfk2zZ4MtTVqltNppIogGlTuZzXj6S1NIJPxgVqPAXYwf34BBjZqnUI3wPApZ
6UCEuX0qy6LOh8ayMK+fKjk0N371Xid3nDrkRa2BQRx59te8XPHLSGQ960PVVjzEuLhxPkWogYiY
vKwzbAaf1bvcE9r98mkRCs91AXxwzqP5KPLs43p8QD92ROPHfi5RCkX3Ruw035zRMxCVXrJ1NjzR
uznxKvhe4EZLXgBE5Kq3EftxmLHaoYjYN2fpgS9JeLoSBxCK3OOyicgE27TRE3h+YgL4qP+0Uv/O
WxoFg3elN3zDajY8lScT9yw5RDl4+nWOg2FnvNfxWIZR0TxumkzqQV0yDSRjhIsIQl+evp8UGdLY
3CDHN2FYPnYlRKChd4UPj22f6Sl3QPia6COkbF3cCS2YvIJagg/2rOxcNjA0j2eZ6UH9khDoIKvX
0eH3OzbERCc+nD5lZePXI9S/o/4rScf8Op+OS3j3W32lvU+Jht8oQi6YCzAWu1O2oAINKXchduni
zQnm2Nz8rYtBtlUG/PHMb67LOPBoXxlHyH9iv6INzjo9Rfb8l40GkMJFh10DbfTs+VcCixCG75iO
yH8qPKYq8ZIGaJ34cUp7bUBGPi55io6f/3+THG7SfkzRqutpPRN4qzaRlvSXTL+s3ZClSmus3Agz
ogITpsFz1OdQQYySQdUjcrhaZRH0CkzEmrSL3FNHbymbiOkpuqs1fM5t3OCxH6SxYGKPmSRhsWwL
FSglkeNx44mbTTIRPJ8cgVVijq9wQ+hQPI3QLZAu3wZthRHDB2Ib2ZJ+oEGzBjbcviu75ilhksf2
xWxZLRqZRCDXiL/+tF2CyE8v3VyiLEStzdymX9TFk3yIirOiZOAUxYd/b5ncxZ5O6/9GY2XXvGkA
QN+Wd3z9gXMSh2iuzKIm3JIJAjGkc1nW1o6sJgp042awEmKtsKX5UqclFWeNgIgwG/jGbWJgxoNt
h9qlj/+Ygs06JghoIK4rLT4vR45TPV5uY+MTLU1kUnIiJjI6cYqLleyqtcUe0zcK2VDHwd77bp66
FQquzgCxodr/sCFKyxuZPHKiMO6V7xcYdIBrQ1iZaa3rJwBvob5du80fptBG9Bk5wemTvJSeCxtv
h+LQHwnA4OdQ9vgGAXZO7trF5F4tOA1JOhbhhSaHNTG23WRFzRbdSVvnEbx6exs2xmrLyiVvHo/S
V6eNNP1JHFwHmqOziSi61yGRoN8TXdLPGQ95/XvQmL8Q4n6OBTxC1dSgiUFeIRMxQoRO2Qpc8Nl2
h+Igq/RpGZjrvzDmOmjE4fjFoujAssSb+0xatPJs9N6im81Q6qhVaak/59nhnngj0h9zXywre2WR
O2VtfyaB8pjdXCwZWKUWPUkKQg7i/RPsa5ROa+4clXx09xYj75XNsLmDq8aWl8nRKFFA7SxWyZSj
3FVq5YD8Rcl+OEBzpTFMA86FiXW+sy8aDpfufUUfoqoJCxC2lh08x8t4ApU8k9CRCHVodzxZxQGM
YY9k4xjje8tQKCa458UcoU87DJAorWq52396VoQdEh0O/PbJOvESFY3LYLTimMAgOy/CSN5HdBBc
iYQbL26M00FNUykP/rLR6xkzoOvHzNoaeK9ilZSCQvatmG4ahqwF8Mbj+O0bKj+0y4oL4f58Kh9A
U9OMdxGsVwfzd4dbWWkxeqXSmQ9CpIUlZQhZMXCFxZ1+Kp9hpGnvvcN46aOubxVnfxUFoi/5beE7
79F6UcJBPg3xxo7dX30omzBAFVhQefZu9qNQVlOgC3T8QKZo4ctWrPaqKS5RlP7jTSzoLKaVrBjZ
45iJQzpRhAZ5rSEXYlA4Ksv4hrzfW9pXCoAvBG19AAIW9YhbzNKdRG1IYuK3Urk+X6o0YOZskz5t
xBNoj+xpG6GOOiCDtod8p39eF1ycEQq2dYYaKI/vI6rP8TIJBLzYIPnMOKp3EIJbuIT8yoRHy8bA
fOFQXaZMKwO7+c+LYXl751xZaSdgXs0Hznb0mYjTD8VAF6yiBF1dxWw+j5kz3azjJ3aJR1mpe3WS
7HV+JzwGKNV5eHeqljXuev3dJD1PKJI39zTzC+5vHeQuQmdluYOibhcrWYpLSHjvUYHrFTH8dNqw
6hOem2HQKvfglVQB4cSonrx2jLOfuNOADwszf/KvxDOZz2xja+IkiOAf9RklvEVN9oIkiL5u8OlE
jMe34sRfToCxtCFWb/w4Ielm1U+8Ua9H819e2ujmhFwOUcdkXVUzZAq2t1KcLonkT9XIHh2aRGGR
N9LhN5cC/M2yEbCmwsRJtVujE/LEbisvqZMAor4uNe6zo9H5nkNzOuP3nuLC28ISAm84zRobnAm/
jPkR0XMxc5u8CJuw19Dt4S6sK+w5ypGpobqBhO72IlgN7LpfqoQj3fcep9OQvm+VK96v6hJatI5U
RKhexMqzukhBrNr3lrSqlA9f+0kgMMOlgRB1hoQ25m6ZLC4yYQpA/D/ABjz1eLlMRcSZ+sy0vOtB
oT1/V8Bmxk32fxHYdpElQrg5zrlJad7xnBRm+k12+nXbnL62XOGRJ3IBOa2orbBI9hyUqjyFW/03
xRmB4ITVPGx5E9mVmMb2r7ME3kZeqMHiAaP+M4RluMc/iEOljmiqe8byezsJab7cCpIlon2eWgQG
MgM7VAyUmJjFJRRFOpfWA8shqK1vwWI06rHF+/y9SnnU7sFIC8i4aJUNZA6AVROnSEJWzz8KoRk7
N/AOcRMFgzYEq2G2S99M5BFpM/XM6AtY772ydSfQS2AynnSfT84Tas1/O74gB2JYPL3ejv+5864a
3dyFfzI5plIXGOC51vZE2o6MhMMNjLlRkAuNSY2W50e0GOb+KFOp47n+ezw7IqCJLiJZc0tfWir5
IAVeXgXlbvY01QD2AZxraWwjeSVyb2Iwr2szCUBgdswWOoj0JwRDBVr+5JvPzdPRWZGoabQI097O
o6O/iNjryjOzYzrcqxh0kw+s+TxxZwHeJvsEihqiLJ/gnpVoi/xXsuVJDPuwOYlO5vlg4FWQ1F19
ayFnandq5pRsPG6BbaGT0OTqdODO8LgbaO9XkOws/IYsurqnIioyLOinpHw65jQ8niTe/AlQ00/o
3QuQV8tqGJFsDJgJRT/3f3KUleh56DLetwQpvrl7FMPRPjZnwlOAACoUBSBHXPkA0cAn5jNU7h/X
9TEBcHUbY71laVARYA+ZuJmENUNzFZ/6PJ+eknc7Zc0Rmih1D8GKLw9QVmA4seFmIvbZAJ7LPBjA
djW1m7Sz8gtyuZHmgqwKffnG+Wis1J/5D2gjDA7GmzeZqBD97+swuND/AdkBgfsnkzWy2VYg1CB0
4Mtuzi2jGoS1lXrQmdIQFNhPEgDH671a66p0saoFV9pOhhNJ9w7dCgpXIVEKhZbQKrf+M+jqd14y
tWrGkAhDHWMu51ymdPpudTEWL8s6qDb9h7gAkgHAaBl81ljUX68FUGzPgGPcexqozIxFuS27KRo2
hLp4mjT4cV3IvF+EFLVxWIpxN0xxuXSeCffWMAc1TX6/gbjK2hJh6BX8IkIC1dWTohaZR8QhcWdB
2WUiQ/ejXZRKcCkAX9sLb63oSdtPbvqNPRWoUUPS4354vH+s/EmgDpTU0to79ZKLcK2Gz6lhutjY
5x66NkKa92euCxrT6VR2IjqhHv+HJS0ZrjFY1UjWRMNDZzViyox40Hi1bGJ3RnEle9DJPaZE63Tj
ThUJGDLpHngW2t/bD00eax9vCfaskKkvHJVTLo18iUwHpdNPURVqu10DdpkCvp77fmIJ9bD4gt7c
XR1TJh4CAz/2NtC6im5lTfLylj+JtpBp5ODCCnmSabwmRggQQPUFw7GFVL+mCJin0e6jRBfIGYP1
8c0fYlM+jcD/sE3xYDauHbWoQskK097Q4GQLzXhgxCiaAn1q8H24QQ04Nr379GoyL/YvVv0inJoE
yQjAc4wAewO1BHGaS1GFQIXZYvBG9sCuTGs14kA1fTdYJUQU+Wi2NidBLKulbCDQ6EH2gpCTrW9G
gAn2552B5C4QopskM4W5nfD4/GIzm9KHOGNbYagIn3sW2JLJAeJeYaW39ckacb4xMBUSbi1m7yGO
OiKtE38qjpkwmUESMxtIg3rHmhufCyfXY09XyslwEMXDdkQEL+w/+OpUlgxiCj7jXCzjEWObOJD6
7JCaiTAplQfYR+XD9lVH9yD68uTsFJwUy+f6Nr7vABPXxIG3MslGuaUciAAmvDCDa0IH30ok++NK
jfpy52vH8O2sLpHbnroHamLSQAW7FC0YQbL/w8iAs31JmnB8CqNLeQK/qnzzXCC28AnY+P7pC28c
soBKFsZhp4GbUgGIKEU5pqcg4IceS7OGkYOOuzt+sSu7il8taI7vTXByrlPprGf1+rODvPJHLT3B
9t2A9YJjz/IegpaVQPvLqVDAWHiA6QG1vzGx7i7boP1hTQjk6U7DfysoxCf8m9r+XDU0mlqFnWiC
8HCn9TBaHFa/afnFq6auFGNx5+NVB0a4zse3iyX7VhfknN/zaLFgj+maxuBxg2RJzA+R0CfLpmH7
e1MjyGLuYUVUhEqzmlD1iBAIiyruXl+r3RUahBEQjk5emT07klP8ZsynzSSvFXCKcyYxj6Al4Nc2
flBq89P8wBEf0yWXKchpb5fwJsDrJzIndHeexqx5rvDpd3uu6sz5LvdnKn7jlB1Ceai/HG96sGWs
xqr0L6D8YhYb8j8aU5UHXe81UD+0CT15bFcwBwrvfWAH/93NXsg5BkDHroF30rF32N3kOdTyuGVP
MYZFTS5h37fWl8OgQYk9ixji3oP1ptjudkcs/Kt9OMY0C1gH6XUsKj5U4O68ZLGKYLuq45FnsjXK
mxFAqtU+05TiWHZM7BAqN+nJmnAW6vZf6WSPN5tdEC7hN6PLLlLnLYnIrohzEUDUDcYTfAElpYKz
a5tWE4e3XESn/3k+9g6hPxw03NFelbp4jlkDOj/iWk7rAq32OeDkzj8OhPsrfMEy7hL9+b+a3nQF
qi8bWclWREI9Y8m78rjKhSxBm0zLbAY1+r3EtIP9O6pUDBhVIWrXS3BvxM0LH3ZW+qVeNxkIV4nb
AcFCc52LQc795KaECUMgCZarh7YYaDLldG9x5+lO+ukyY5XZweVAHA6gewylSo/y5h22quFqi3DP
gme090Z/wU79+n3HWH9M/Nrea9PYDavDw4pJYZitkRii67AMcdJy83JXafC+zd6CeqXtMyOpVHv8
1BAMf7x/rlIc1CQwpHNNJJZrurBefMDYKUepdF21gdQ+EWMJwObv1KanoTDo+GQlf08Ky6Mi2YOv
ppEYy8K0ys2Mh8KOmacjAa/+2TDQDgW9wdx9+PTAUIEsQ5HNks2gEXh++2+coEpuQuLD17Y+ZNff
4B3ep5wMC+TZtW0z3t0aVCZGtqH03qWUdB1GFAYOdGt7tGZNy9mKyePpYmBaRzgk9CfFUnV9OUm2
Y3BtEiHObcHgTzywfbEsVq3kC6cFeh0AkENaMkYcJd1JlkvMEgJnPzz98dFpKXgN4ZNhusIk6OeR
CZ1O5Q2OxrlUnmwDDnLcQT+CGrF0uwTUBCm/ZMXtaTzoleepwDUFKYfWfqj0ajn4wfHVn3o3xXGI
YTetb0qCJdvUNfpWIdSf/O9suwz7fgL9Kh+ziuJP91k5kLfijiITUtkgVJvJRe3W3ebyX8HBLUQj
aL5QFCtfP95laUVXWX4ycKsJO3N9JGbXTBbVAfh9CbJpeINYHvnAcPHPfno5p9sd/nkNyCwd4oBx
f8SA7PZ+cRp0x4iZFpNoxL9W3I+6xMeqN4/i+Li8hRo86eRUOMEkb12vgRuHntikUcOse360rZvV
Q7f32ss9l5GKjWOVHXbWD4vRfcmScojSQNOqn1MDwaKtuNkLZusnnb8vFFxzDJiNmj6OpdN51BHw
eEB+4XPMX8gGOTUK+Ydxewu2XD39x5zBIFYw+De6LNUsjYUFfp5jG7svnyQynH10WkE1groUVnPo
VPBkbZZXPk0Sok+3ztsdeYmJw2HxzSJDzu8qnmVVoNO/Nzca/M2JNZIUR3dYrICpjAawYgQQxTPo
oZ9XIwkitAcV/ofbymte1+BA3uac4pDoVoSBGU0Cpx/tC44KjBJ+5TXknrfJc3/9P94ngZQJYeDV
soEyuQTPlH12HZmRd93nYHuWjRmZBlL778CQ5ibaB2WhHGSsm2GGzv6AnasA10QYsFV6IjCTkAfY
UH4w9IsfbcUE7RpcOjPBChqpoQ4jNfVKAYPPc53dY0dVsniTKu1Ps9uBNoUAcEJCZzKDMeDvAhlh
GUfJ2sxZdIgqIkc88dAfnKwnRSMaIyUR4XUTonRuj4OTYuniQhyAqO47aBbow/ReGafyvZtROL12
aZc2Oe6rvoMDFdnWLqvvhiwVcVJguPPR+AC8kpxD2sD58pLhyWIG4AkUuujY0u8l+kWDVOMmfCQr
aokq3AR/yPzVGrELMQMCSvtd/MgIgqigyBj1ImBDUdEAtHrQXTRqjfBAPCGbJ4f7NA9sFhQBEBlT
lNTDqesJv92GK0rf/D032xK2lCOIx29wfQykV6Us2KFrhDP+XwEwzSJR+sESQBCSHTEMJZHgsMef
18iOWjLnqlQIRqJ+UhldcThgmRE5lSOO2Fczvc6M/hwdafEIG00h44HCRyU/yu3DvNhKibtWckVb
okNE8qQI26lD4cB8NC8SWY/SZe96FTM4XkQOgmtspksJT9dk5503z5LuYcRF9bLyvxjuEjbGzWm7
NpA7Bzeall+6AXsozmynLn7k9+e6JJQbZcigaz+tTaoVcAP2zAUZqKXV6V4vhbXIx882uO6RzMpY
9Y9K10C8C9qzl+K+TzIgV52xyk3p09ecttN3LLu/n8hwvGRPoXvWH807Q/JI3hJMGkZMI8oXBYgs
W+wrZI/uMUE0ytxDspY+s8A9s3PUH7yeYYrqMkDGA7z9wQts0UCVSL45F/8tZUY/U2wJ9nKPC7vU
HJDZwecXGw4FfiT8LN8/JG18DsBcde2QXBaoJNQcJ1MMMyH21dh/XKm9p8xyqAMgIGTaSKTZ+uPq
j1e+t1DYTiJMdczM8WqMmXQ6r5weo6iQTEgHRCW1JsCiTXCHaCjyZcWVFSAo78+S76ZJpKh8M+Z8
PQLXiCNmGKexaEb53WTrGhYQisWynVHaKsXOulQcvBo4thFAVbI0xoG28ljZyoFYngA8FWD/x4KU
QxAtTkiUw8+fDni76ASmnHdcu3KHA6GFhqdjH06bstRWvg7HXoxOUxXLVk5up0U0h+gTmquqQtPT
MBtthJrGiGe7XwTStUpjimsbHDODdum/gq+sp5QSUubIZdMTDN2j6oy1/zro37cB5zmmVbU1inaq
SohzMvcR4exWftb8ITGQz8/oO9zDbfoK6lvHUshYDQzDaSKtx5fV9u1ClLQ3Wja0ijGCXu5GkMEx
y/wntIL3lhtu5BDJP89DHmasCx6/TMznSYunI1mtI7i7C9+4sD6D0XckJaZ2QJ7ixRr2yh6V2kv2
jtftofeyI9gC/DH/Ai7aoWuhSQ927QselFDrl/QTB+8KsE03YfAN0aHW/mDPI4kFFiMAE62cmQpK
lcFfoJSdo4ZELbbOqU8ngky8hYcE9xAdSph0eV35s1kZLuZlSZWNEocObsoM5Eqj0Huuh+jkGcpi
bPserJ0UFkpkZ7nnUE4yxd8a5Hd29whVEq7rSnvhjh4biTfR2hDBXlKH8aEJKldS3JCkRgjMwgJH
j1kgp+HE+ik+kdTi/vkEagtg9AG57X3NcbL58zAtRgQ6I76TkcZZ+AKSYjA+kMAadm3OXVAW7oLr
qOCYmluiptGoL7ae/Q3l12AIm1+5ff3FAtePPA4XEyhnTHGy9jH6gE4rJfoQkZdw+z48ov+qRYGK
7tUJtTvDhxKX8efEAcb/SjVxfjSolBolkW8+NXlFJEjOd5mdnasPTsW7Bt2BCoL3Je3HEu5rXtIE
ZKj53T8teqZq+8RJVo485kaqkMePISVLpfv5TdIVK4tiDuEJXhe+XG8V6LyLTSm9WuNJlxsnoe1m
Wof2otALT6Qi7g+GuWI/fg6N9aM/Xoa3TVwqA72HasYdbwariPjyu6k9pWtfFEEctbBH3c7SlurS
MBTn4GG+hxLzeQDucxujcK691G4VqIDhuw61VSIj5DdfYjArkNVOa5ukGjsh07tfv1xVzuPWLrLj
rOUGheF47pm9r6RF+CL7dRBik8SRBD4dp27WbdMxK90a5TMalgr1WHQhhSyoC3oC0HhkIj3fQY/Q
YbiT/fpyd5kO0C1Eyy39f3tFiphlu2ayPL891ZExYTq9inrgwoq4OKrxJ7V9iDvm3JN9Px68bIIS
crsJumuhe/lCSJxYGzrMW7ZCOggqlOeE8bUDLW53e1pALu/hx7LDhHJJeb+xspH+rEjGiY0DSmJK
UCRhpQrEJRcO6xOKHYWMn3z8aci+Ije/Kv5D7goo19qZqnp0Yw8iES8KFqxJjH+yf3TcgHUb23yS
x+tdIgCwjU5Ovs8VgOHaVjgb7JZjIKMu/pvd2Z53Qbp+I/U5pnEDo2Y1u+5SRqOlvpwYYgtakeSv
JHQ8pRQF16XuT136EqYlksNHuPQNpzndD7Bj21Gn522LMRl053L3C5UIFu4IsJ1khzgP3p83KE6/
0zn5J3vZuZTNKKnIGTfoSvVdKjPzJnVxglA9KJFZdto/DDTWhg1BgnmKLTEIXxjOfgLLUqd03uvM
yr5vzNGME/b+xyyfP1sE1wBWHp+R1nhDvegkmJOmQHIG5+jRIXuhYBfdTotXHjn7JEo2+2LCcKU+
sanTBfz5tPGBi4IVrxT1GpK/Ma5ZK/gbfZZ1qVb/w6TASEZxhsA25J90dZUZ3u/4dOjJIlK+9wpx
E/o02BWPWv3AR+tQbw6GnnyRPbKREmXGUa2YDM4zQq6zQRZgpOGZN46fusXtX/fCC/NRcZ58X4ol
omqsXxIEaAFCGSS8S8M60uiGJWzKLeGlGA7unYXO9YQo8EXcoK4TN1YxZ3mw6Bj7MPKgVOjn9GUU
5t53JCewXUwnsRVxPNkAMQUBtU6GSawpE/SJknvsXgTtb/5+oVMd4lNrS10FqI3TGtrkOCsbF9ry
PNqi4ME3B6S8My2hiKbhpp8YXV+uA2PeVW13DFLjLDiHUE2tYwqGcWozPsm+Ux1+55rC85spl68f
edpRIMkmc3ehuRNIeayYWLCzHXgB5prWESlMwF9KaOpCdRtzUM/S99QykW7wTnikKzNrsZgc7U80
Nt3iR/q/JQH7gxKz/p/8uY51oFi4/1wBkwvsRr3m18y3mjlXiTn6/9AfBMoHY1AxOpGnrqSTS69b
baZz+tGG8FeTXbbWjzGm3kfA0uOZfTam9uqfbS78/X2LHC0z8v3ZPqjxGtjDcKlILMs9QmJQFhUi
rDoKkfZ9zzibcCrWKfl7thh2Br2hsec5xry/Yx7X9ek+Kf6R/ukrGz1V55PeQmzguGYRECkNTyOB
rRZ9ndB7t+ssRudp9dQ6/hkgUYbQC/4piCsx26rS3zK6PfGmGkvRLttSXPCPqb8A0ZknZqbFNmti
ZiV0WLq6Av3RH8KCmWfnksXMKiyYYJnoNniBl6rRwgkw84U/gQodJaNBz/ILtfLEqRg2AgULHRwO
WmbXevSdyX+n2AtqZRbvBBZRyphVT5Gr185U9EcSGG6pwMCK0CjjcLdiYA1mDyIO56ghdCSreVHR
IJZQx2Nvd2QZN17aaQq+pQQ4PGy3JbZ8XF/UYUAKr7ZLkdf2ZHhPEndrY7xyR/kpO0/JUotbX2zJ
XdnH0+fhGXGkahygyzInYlZIS+YRPK4c6BLG2a1L/NnhrECdtcv66IMONb7QLvT0eUsbEnX0o14t
bMb9YA2EXuVKUAsRCE8RRk0OslLW9he9TjTa6tOcDB2kFjpxQfbq/My+U52sBMSeKsCzSO0thakQ
vLJTtTJWQ3ECiJda689RZEY3ounnIdaELLM8SbH3l/LDEqCGMC9XtqYoubcrTV6A8JhuFfbqW2I9
NzJYJD6UL5IkxrPwqiwuUlJTHizZK/0o95hJAHLoUMSjpM8FlX+Lc8G7/jMdTSvOksfoQV4Z7KI/
z31g75NjCnUZ96qEBUhLMWztY1BAXAwcEYKo/T2vfn1dHPloreWAmHoVfAQKnSHlOcD0SSlgNwX/
EavE3fdwhzlzHImCtwmf50BTs6xBffEmzXjE0Jrhsz71vO0Z7TB+e9JTPGuf6MjY0wv8PKYdr4Je
wODA3x4s1HIZ8IOLwQskHNVJoUMRc4kyXZJae14u52MtTafWn5evoelqwTQ1mqezRT9w/5vbePbG
I2p80WdhFXNYCA41+/lmRN4kf2wscA5YGeILj5Wxf72vPEqKFWl62ra0ZTRCLCp5WitTPWzN22Wp
UCZvWire7Riqm/lClg8FnnP+uMb36ixk9wQmbTR/HRPYB+VTiKf1vUumGRjGye8x1KH9S81RS1aY
FhK9q+OZA86plMTM0RnpeoFXicQDmIHkK5ijvYBMImnNAXp+70xQ066CrszBqRpOa18g7ydxLHdb
V/P474KYORJOGZRiID/FQusL2QP1uo9h03mJ4IW6q/OmetuRCY0q35tZQrQZ/Sp1opf6EYKFl0Lr
muKP8nOEnm/LDQRg1Rnka+UA630ICNgGxQyu93mEalitCXpQWVcYvNfTRbFkjnyG/SgBO575HI3V
szA9W4WObHCNJX+ukWQggYnHysKSQu/KZgXulFeRS2Pf+jpiWCL38jQeQ8hc+0tii3ycWrypihdG
9VhUH5iZmP1SXDlYMMkWLXiOU3OH2ycAh/zl9CgdVtsMtghKPNupHonAFk1ZEXwTvPhCG9oeoJZu
PnKlNv5PAvee0D94jREeB7K4IVO6RTSImY4Hm70DdW1lhefloPNO9kMmmvylPDyLbYHzqfQVk4L9
X0xyalQf8n9FL5R7XWacVY5iFSr1hDogOBAwqgSu3yCQv0E2L/+L48NkS4+WxzJ0KePqcUpGUPJw
vCZelWModijalPZnlClq7anq42V74V4qd5yBO6uLZ/YM2QzX/M5o8ZItUP7p9294lxr/TOlEfIKN
9TLjLRbBrpGCYHP1FtLEtcKeJJg+IGhBmaqx5W7I5mp3ZCELgvlAm+K2KJQ5+0mNPGR4fGh/lPXc
4KvJilpbxI5fbyu0Bti+WhfPlIQuDkAncOElX2jTgAb9/4ksEwMT8qaMLdoerOnlN70ds88LmaAD
obUZE1kwrFwZjvA0zMr8zgS5FKZlbsuLncjfuk//RS4E5lcPqC9wOQYpH4vSSOuhIPHEr3on/mMb
CD1udk8ALKOVzO19++3HLiG9sqr/nOH9GGBvnfAB/iq4XPuXHnCo0RrW3gFY/lCqai9Gk5RLEBRL
C/rznAVsalpjbt4Vz5G4tJ1tuCecGdkKMEjQUSqcio079k3cHOj2djYNKz+sL8/dtAhD+Jpw7aXf
R1vCBFERvgG+pM1LdCRlabSCKzklGO4ReuCuveS6ixDL3J+wNDkkBTHM/jCyhc/90W+OZ2zdfZg5
R6ZjdPVPlbxYK8bTtbbya5RoYDMCJCf2WotSbnpvHnuErsZnpxQ6HlB3Arxs5uNgKDIs2r0ddGWY
wq+G/ZqcYe0x4F9NOW4ykErSuo03CqtvPVzvHuV95R5uh9x2VTaj4xqWc6Y/HCwBqoidhYp5do6O
tBsA7uMEdMtr/AH0LZkZl9i7i0Wjo0RhcApOm1JM91hoTBzH7yqwhu4rZhAkhc8/6S26b0pfs1ci
/oBNDmyHudbTZSLVb/00yBS6tVU54HUeYhlXZkrKrglI5t2P+ehVCIRRcFDS/WBUa19hdkqT2fJ0
H+YcQDlLa+QnVeLntyOYQp7EMxR5N9WwJW0+LZp3vVdqsKE8QURDT43RaBP92EVW7IN2oQ0FCspx
ug172oL7R47F/EYESBX20j0DkAQQBK0JtgrsqePbtR12wHYS9qbThk7VAQamruN6lCqxwjQTZItF
dZj8EHgXtp4WmzOT/jfIP/PKl/ibum9NtAHLBu/WOdItx61JiZ5qol4miAYUvX2byrqTSeyMztym
FkrTO+WkRxlVojIOcLrK6TLoTUDN/MCkQ0yPU5YwkEtsjy6DWB8koBADgo61FhLbvLV9n+a3u9M9
fm7VINgfs1iu+tIJcwEpa3vV0qfCMfg5QMjhdF/B/MiOhvgkxPbpCjQHOuo5+fufMcTqrSzIkdhX
b44UyA+Adj6AF0uJR3eULgojku2KFuqOi/EJnXZOmlYlnO52idn+ySMd3o5s40peEig/pQd4UlHH
BWoSl+Fax1rICdHTasA12FIi16aJtIw0e9oSq6/lZeB0WzoakbU/cFxndh45RuQarz2ljpp+SK0V
oDfE/LneMbd1PQNNrcghqZ/SyRrJJXlJEmf2uULXQ4xiHaQPdX6Zf5LmTOCFeiFth/PRByJNo1v6
vP+5SVEJD4kV7/PWJD+C79lPix+g7nK5YveT8qL677FC5zVkQSTxpg5e6thfQJXNG8/qYAu3bW9x
hJi/V9SOwb6fPQXidkDEOMMAOkxD3LbeEvTRc0hAQfP2i6stehpejRQP6DfxBnaVYX/kJKdR1e4P
AYO8NsN0Xt6JRk5HXi1OWnXPa4O79xOPQ22X+hu/X0RLHDZOjsKbKMGPU/hGq+Gu3Ay4Fjg/B6vy
mRseMEe20a/wY0fasZ91+Rxkp+3EigBdvpziRf2D7Ep3q7YiCXw96gckZt7MM79ukjSxS6aPFYtK
Y2JxZ4yYS8YuPrfW/su+ldbPo2qvOKpuoXZAOXgNxWa1W1c89oS29ef7VuzOqAv0HrxIZekHfD/n
nAvD/HDfonjsSTd3PKNmqheCwPIll+05sM8cuOfGbyb9da5yMkR47QJOE0nxowhFidpPephBncZy
OkFzQeqc5hSDeGE6+xNjFRH5HYp/JIPm0Ke8PqkDJmm7Q0Czq7W+gvXFWKI33UF5Y2rIvIXcE4my
CxUBTuAHxd1dvs4GzSwiNRRd2C5EU2Ku6pixlPPq+j/QSKsyk5xnLd4qlGINcqnTOhTOcv8xaOsF
ZE4qaGeIhGUPOykwG+l8rjb7GmICVgXpb5RA683EZUlDOivPBlj0rOqPBNoZLp/mfGlzTvOWDn7B
whOvwjG8Vt9Z54OxFVRlJBsAiWKjZQe+UUh8+kvRtLOdoTAC3nncg9Uo2geLkiQuetZEFpeYyr/U
6gq3QoMk6SuHv1HldhvISgCjxtZ1Rou0OKciyx3qbwkXEuYt/6qIbBne9EqRjLRMH/3SdvNrgWKN
ZtiSQIKtvuF9a/I5wOdsvaVjK4E/TiyY6zHmAHxRvTgkGe7xX0t+WBzjWr6br4vv4Qju6bhzdvCH
mOEwyBALiBsgCwfFhtH1R3xfW78comUplsMRavJog6oNn/DmznmN5JBTSNJ/PijXO0zNf9TL2X6n
WOdBC8VxX4pVdnXShdsRBUcOzy2vQa5JHZxkRUo4WfUUVJNiqObfHcAR1bw/6MEeqZ9ukWJAV1ka
twBiNi/iXKFXik+MgG365kD9lfCiheGxfaKa6GkjtN4RBthwZW4y1jkPfIwYTqfGoTG6fFqT7Pdq
1uMqev/cOrrJtAzOhl5GTXcv7+1RtYbI0JK1qEqqMVDsW6/JYMD+SicQu034Qzpg253685U3Qsno
/D+YCWHvBF0xhQkvKuFYNPEupqukPA0CzKRwR494jkkd1EVEkHOFQpU1ZDDsqq4+wlLE5A0rZ7Jj
7JbberNAIUWBU3PQBWMjBidZKWITL+WDrOZhL2J1PoFcKNSjSizZr2QsZAuWGmkartj5ssDpl+50
rnU4DvowYgamtk3K7eI3t2uD86baldag6MMfEHx2JV4iqR5PbQusA9iEeGMZMQGSMwkBAwKFQdae
0b4AH5WEqC13vL/cWgCYzHkpEsgmZppPvujGBd2yXVD9GE1bzqGKLnZRnAsVUp0BjZ5gfzsHxZX4
dVtGKGQ9J6QMO+P5Tnk6rWLUIZkfST+4ax8c8F8UzoFidsJ3++66PY1fQ6wQ8u8z5x6j+obJmCr6
bWahDoAWFcol1uxM+BOG6ld6dh72g4Bglm+dNFMgCv5ew5bco9KoTCBHTCTq/trp/dAZp7ulFX1U
gJEMf6WdR9KTt5+kQd3KbyKjqhe3Ivor0T2H3CSaGL60wZvzEqCpb70+UKvj+K7ivpPRMSo7RJLp
rNVdISbqjqn4aOXzFpGBEfi4aK713Ly/CXUNe/VzwG08eoeHY6egRxVFiq+JoPf2bPhsn4mTvWqv
xQbWLHDqyABTERzL7JEtURnGQbcw5FOQHqQ80DmZwfWEofKB46fC/XC5FDJ5KGM4TGGROFmPZJPZ
SnuiKH0lE+7PiQCp/BSg22zgkZ5+CwB1wDcSDsZ+bxLVRwMamqhpFaMS9PkHNWbel+W0dkv8rnaf
dFLLGYmA1Wj7R22i2aaOHIP/Udtw2OXRw4uTPTDIPgNfCZM8bdMyB5j/p9otUaOATidTkHdBlbzU
MuXTseyefHjrbBBp4QM01HWi6X/XJWcvcb87EfoAf9Vo/voDSGMVrZ05ZvQVYjUlK6aCQVuHgBRO
K94qNBTmeTLhzvuL75Q2fntqXEYCD3+Jma2GZReHOadJre3+LrxbhGN6GTzINahDaiB2XONXws5v
ankspu6QINZAB85wJ6rGD8E/rkWivXyB/DTVyokzpLPTCBb+7oA8VoBAYfAejCNh0zScGnx7kcLs
5OXOeWbw2FF8y3kj2nL8wX5myvQ7oT7JwZzLrOipu5iN/CPMhfOs7Uhh3kv4eqbGndM0oXN8txlg
dfn6czOq68JxMC5sbpbn8Ao7t3R2Hj3vuF+oPFgowvUsce3JAZDzM7qY7tpjna9XInpcUObrgFYu
thsIVGbOn0RbPdpsnNlsJpBxlE1pMIOmpu5Ek/6m2Jb0/xg5GwncvimlXXWtXGu1IiQK9Pzthxmk
sfcjyaRjZz509pDYEzcvjXj8F7XFGHNgTVm1otLUpNORj+xUSJYD42zFVpl1paqNWF/vqikJ3QHD
8Uvcp8sL9XaebETbdXhOgwhVhgyeuM8Vg71fkdyJg/PQzBSCiaQpQ/W7JB6Ea8r2AoGkscsxF8Vb
vq7J4hfe5hDuc6nAIU9qEZCTtqP3xbMNoZqaHRujTcqUYA8NmaVD4gKe7F9gTQT0pSLQW6Fb790/
tCR8lqxHHvbK1Mlrc+PvTvUAijuVZKVeoYyY6iJLCcY2lZICFaHQxt08TONmwZEXSazHMFzBfv5c
XkA+LFu3DV4AQ3cicV16aRziC66nXqbO+CprMsvZ9WlrLOMWemu+AXNryXRQ3x9KURlQGrPDwZh9
LfAqwO60Faua6Wdd+81f1fgQlXUDhYpfnariig9LR5yFC9K7ZAF/TbWgreaHRk21WWdmB0bT8vdx
+usA3jXibm1HDLtfXdX6ySLryq0cH/EL4u1pkMru6+ngF4eNynCOZ4MwprNRrbNorixqMawNxmng
JPCGYG8F8+4sM0LQUn8K2LDgXJVnCPcOlPzuih3Ipi5qNrMWjQf9wtiMwbXMJS17qakfcYqq/aCC
7y1qjHjKDEkx6F/LTknjJGJSVZaQqI3muF3kid2wvKGhyf/ZTcarV3iO6A5Ty4fNG1cml/3YLluH
IMJA0vldgK66O7vH9Eo0uZH013QT5X4svONWqAp1RJdXbyKdSRgrLNp1xWicqLry4xFpVzF2gDHj
4F32cvmC2KeSW7UYeofJWSU4uUmbkmbsr2CorAeslLcL2z0Ts7wUbHlr72WGHVBijuXG75gttt89
NF0iKcTnFdoR+mE453GVbD/LiuGbbUwgEVIgC+ylY4hcb53VoPzCx0IWFRvLWzUPPZHjF0Scldaq
iKRLqMM2xiq4o9K8/uRDdVh62JmLrr0pWiq3RL/pvZLyRSG656aJDVVoocK4YKbDogSPSOrMriCC
7aAVyfKvmc+pcAJexfw/i6WMkYLmXKkkaGXeSCVI4ywoL1oVcTph3/O5yxxkq2Tu3WNLMOsZBtr6
6hong8n+YFsKpxyjHtqPE28DFvNu5CRzqQr3G8ZyihKE/ejfuNIZslYYsNgSwsyrVC4sClTJVUKH
1JH4F8Fs4ZEe5JObwSCgbxaEA1P4xiZdeW9fBCoBcpvYerw+XPWmCLypjyZPycha6i0pthbG4UwF
K8SLriKEiBn5jw3/U3j6BhqFYXgZXsDxASM+z6CUBScRou/Btgr0lBb/bNRpG7d/P2CzMYFE7PSQ
WIoNEzIKhfEYjIKrdsjnMbWI0FE4FZo2NgtLNecgiGyJuL8E6yK/LsCvmLdwIpEyAXoi3B7F7130
vNI+3iUdbeic/D7gXGDh0H6JGMQU+6EYvSnYxg00hhY9ZmESsRxnYxrvRtzyFKy1gfQhzb2Ok6M1
/5J2PltslDJdHmC/DPG3N0JvSgHZoe1eo8FU0ioO/+ZT97TQkZ7dlU/L3j4ww2GoWbHKcEIrXzBu
jJ34jCDWT8j39Vr3Ru2xrsIwm43hl49xPwpHfp85rUycMGUR/zIIU1kgoSHkBZd6y0s525FkO9qH
ytnvGSpnpGNuJpYau24H5oYBM2ss5W6ebIBxfeiSgtZPdugk6B80+kN5ZUH8oYiVhzXK742D+7bL
biy14eZF9XzetCxI+7DGPtBN93BksTgLwMrTfbqon36FnJXOWVSjcLwXeqVYNAQJAM5g9JGXeKJo
v4YvE4nQ0XIgJDZc16zrABtSYM3gxZ0rI51qFW4gh/uW7ifi74UN1OdvbJD0JpFcNXPi/8ypnkBM
cWrauyWPqAEnBjx7Y/1mVcDRrpoeX2B7iw4gOZu0MKBJsEVfU03li9mnRWJQeD2vAHqbVFPMFh8J
YBRAbnLVb9OXykfJNb0lKqiI7J9oXSy6Dg7PrN2n6hcwxUHwNraP17hEtJjsT3WYkP1PIUgv4qyq
Vg4hnG1EneM9AhXH4I05DguGRvGDiMhB+jh6JQDUJEUh+jh2Xal6yPs51TMklmqiyBgmM1Uh1Bhv
2i3Uelnu8KjzZWkeFPGqWlL9UYGN+9sOfEYYzwagL9OUHkXVsoXZK7hFigy5NXQrkQlmHniFDzqu
w81iwaOw0Yc81Fp9CsfO8EAUygbonMS+hlAckYHnyqQCg4ufirBRx26DlF4Pi2pLXiD+5/F8bKIT
KP/zqiMsMKi6VRBkq1VwYwBripM2j+FxLF9f0T3SqHPQ/CQXn3KDpk5NOYYjlvpZ2f+oFJ6KyMfp
jphXt4sdtjh8TmRrSzoODdjQDOeULz7SwuMGA7WWOBHWFCv5OJ5hBYnRnkknnCrQuM++0IlVa9X5
RAOQ+oSP2HW6m284iVymgxadJ5k/+L/cudekCjm6fX+/1cISz2zpUNssxasxjy30be/Em3nTE1fx
e4tgksVg3hP1Qb5w9gU95/vuFS2h1VomuztUXIgZrf9RkN5JGhga0xiLNTzeIiLx6Il8X7C2STc2
q0TheAC8SlP501npWojSEe2YNobprvcQqFpKtZ0ONcRahxlfce6+QOgI6UsTWnCvy1jTMaHgg4cK
HvJaVKIJ96PHt/edApIamCiPalJdKu09fFISFW87YwyIj2i6wwG6LvZjMUabQbZjDb8HHWhDyiwv
9vsmnQYuQX+WFc7fvlyQnUDUmTmeypg7MRIKy50ftpZtRGYBZrWlkx0HYpl5K7zHVrAjpBdYtyHj
29OLiKGahK0nYwVkgKPUJwsk5A/IGTnoRJCktORwz59/+Mwb3K9+5nt05kwiA4l62XZpWEaqIoq4
BKedXhsHYOzELaIYsasTayQHuB+IfRrnU/0ukaWZ8YkbnKxMgYYU9NYxTWpa4pdcMSjQ75Z4JFb7
Z7XBl+DlaAZFpXwr0w5wnWfh8RGsobiQoCsjG0qewnCKNljwrTmw7dxhMtaLS4FddUcIkbogIimW
NYFz5XOXy7suxkomdnAbz8aExqYKIK+nMCR/Ddx2pySUjkRT9DBo05gutT0l+bzDL41ifBcVaJP6
AbD0zrBRqG3WcpS3OWCNM0n4SrFFtS6In8nX8s2s77Jg2wqZMGHku32+C06umiO+tLE6H6zkxxwi
a23X+7I/WSMhrXAEZvelmz8by78MmoRGLnsEoE6FCRsE57KnLijLwJfZAb7Ias+QOiIDLp/S0D4d
XiaxIGHfmszO4ltCoeooT4nhNJ9NagnrApNNyTd2KuUhmU5f/7TcxrtKbCiS0Ukk+yMEZ4LGDGa2
dbcF2eqYT/boGJo2jXEvA7SpsetaZSAO56kO3tY+gdhsDg2X+UxMctLLD5ATkwOcZauO/xUa/eXF
FAoHvuGAOoPZ92tZCcO5uj/t2UcMXfiDR6a9GkKKuFwwklYMh40nckAV/izNLbGu+B6xgV2MbMLp
u9KU3eaZIXq573mSDUmgjPhJhqCp/6Qg3GomVdOYi9T2R6rngkKdUB512JrRJuoaQ1QGJkQg4Q5+
rYqROGfTJaDsEmxzjzjkm5f+7l3BizTCuDDbrh4gtKzCv0mYBVbLaEFCkiuWFfGcFfvhlml01uPh
udT+ZkHkxELqRiSSqIrW4r0A7hxCgHfjxltzzXXtSMW54GgfzdyW/YC8ULUjqdQUbXtysyBjsIlP
eN3i0d/fOZpR0LUjU7OGqVNtkMIabc4JI66xkCshn88WAFxxC3MUY4/XETpNP2M+aacKeOf3S0DJ
UJlQv0x3Yt/v26uj8uWgM4v1fGbOiHd2kSIaMlw3pWD5ZOZFbcOVumEli4ipPsWlzJEei3qJ5YVU
TJPkjrtI1oPZMbQoDvZ4kxoqoCIxpcrY8umq+pHPQFllsRGDz2/xcLZgRFJPeXj9MBV3vZ3gthJG
70LroDLTVFYxpeU0NhbmCCZIzigBrGfGlkrwbbruvepjxzfgRNwSswWVQtt+0dd1eLGIw7JDNdQY
b/mRqi87WjWk/XUHAWBhrKUpV2UaPiBbpHLCHhVgi9+sEASJ03p+rzioO+YzLS+q/zQyqE1qQGKp
C+MSl/IRRZXYm1drC0w1ZLQxhRxbMShDTeSowIODxalgRj2ecvFSigRSzkfj2KcxNeZHbAefz5u/
HBJ2Yg81uIcCoOPgtHf30VlCKGEkaDTF482S4p9PQtQgCA1SqNL/FhCG3ScsA6YUoOp1HFS8S6h6
8nWBgfKG7G2DDv8AhFK+w+CuqW8h2kuO9mxig6Ryol20qDGuBf6ui236BULXlrzkkUu3wOtMkWQO
1eQFNgv/8qzynk7mO1oYYyQSoGKxgHvkkVFSR17QaEP2fH+cVFQ0eW/KPP2Xlc8AgAPBJJccfhW0
Io6dSm2FtN/UMiGYStdIIEFf6xf6USbKu/EXA2JOIkwygzrsU6us6nss8sPBu7H8zjezWvMJa8h1
3NAnGIRAb05YPiQ89p5nMIqx/Fe7EZiJtb1+6Ghug97Lj7cZ5feTaprleH8o722yFXZjP8hsd1CC
mUjoY0WqA3FZ3Q2fZcLk+hQy7GDeGyKHZNV4CCq6KpBvrHyFIeYN+f4RNAWHb8AgVmytqrNdVrYJ
ZrTIzhhJkiN09bOg/BtdJtY3dsR00OyW2T8rHT2bL/N9WSa69LsWMwWB5D9gTGa2bFskeeRbFp4N
5SQTMOEL2SV/yWYjOBTtHipNgXowGQrNH6ZxnDI+r6T+ckiQg0Ik0jVzjO72v3ih2w3N2l7Tw0Dj
XKdEt9mAHUQJu/3mgwiKMHyfQGkdF3s1OB7hQAnpkT9oS+4cnVcc8GQJvEuMvaa7gcbwV5ZsjGR5
3b/DCgB6zH+z7hTob6GLc5+QbRSm67Il/Cgd8u5Rq6MqLQ1LcxL78S2Z8e4WoFQLH82Tg5mjKmaV
aUVNgraGvS9XGkzzCF2Ovp7cb6WGBYZtsFNtlrVXufRfcYlYEX/upd8YQ0oqz6Vfp1d1DigDw4Cc
7sbkTMNdGAmqVi6UHiZ2jQPr+rdhXn3are41hhN45Uwy5qSXeYPnrk/DqGYApQ1Ol6biZ1zWtSRf
vG+N15XQcaf90oI5q4fZ66uoETPUYn22c5z33XS0aQjrQlZIUwCU7lmm8wE8aFBVClM7CARxqFZj
fqVrkHnvlZEWiqFGah8zdJIedqHSukC0tAiRrQyxNkOTpppAjcigsV/MkKiDKA+qzH/eA+nhl8d5
vPCjH3SASf+baHUvN+V35wVb0VB/OeizKYzKcHIYUJV5Uzf7sbSHw1C2h5jHbDsz6gqK9m5CRhPU
Y8tx0uOa1tNyK8mVrhrIuwFXwQIh+GxuHwogpXtoDDu9cZRGIU/FNnbhf3R50z4iVuNFD6HP6797
w05VIJU6OrOz0cw5jxX4lPJbKG1+BSlHi2BYiV2eZT8R38nFJ5Up+5Nj3vp17Lm7BEEte5ewsySb
4W8ulwAwGoPJNBTib3eGp5+QTMRDsJMC8hMQrtLq4SKZ5Y2QQ58uJtatWlpcXn/H3ad74kTKcvH1
4Z2FU0mlqkFP1Ij5lCUfcdhXoEQHX1oqjtObpVhiaRrvtUDYrrHWv1LSnrkz68hWKDyGObovUhsG
td+c/S1iHXDzeJRH0UxcgnFoqIv4UzzmqdHByKQozhvQwjHLeIa/MUTIS4dECpHiRaBEPQr+juwL
/CpdFRXOJAxLv9ZTbpEM6K+02cppU3AhCbprsT8a7QoVqFn/ve0XBJDTlnmXbEzxeHLrL3ROePjw
cMcyoj7C3tiVpnRVv+2x+OA/amvemNI8/1KYo4Uw5Dkeo0DLSOnYos7VjqWdZrRh5DI30ArlVB+b
2Bq3XBiXTJ3EzldiuKSYbRltbXyE8mDiByodtZ/xtT5XCE2tqO9inxZA+deSdgrgyrC8fG1XrZyM
lVh2WQMyIuddQQmNXG1UUH7C6DxTE64z8mV1LOgYNSTd+OGxB+sakQg7+yUDmyCYgKbKh8OzFcpT
ehpIum4NbUgjxrmiPblEStPuspbDFXwVI3fit4HvPtwbQYmwmx185jUdYeZUdee7pT70uwcP/2cd
tu0tuJFqR+yIHIB1toWoTzoOw0VS7EUP9S4dERRwGBkeauYfNo6mSkcE4fRjUiV5ts7nhnDtlP5S
NNWwOZ6UIeapohUBXHiS0cPqGdWuho24bxR7KDLAe5XWKhG+CXX8Q3/covwnhpUomqDHfOov4vRg
2cEgAgjAyxTRuIKCwzfnGz+hEKv/ld5P7s6wG447v4jq96DmqCw70NOUTvt6f3sSADRnyzfJshvl
hFtBGszTCr3yYIw/5UwL/p72iXnaFGjKz/Q2ChXko23UgWmMrxl7gOSqJHorV5PQTZjbU6jUKX+s
POiTt81GniVEGeCYK/AQnXz55vajHTKuIUodGBkkTtVCURA7v4ieEYLkHF2fXfDLLg/g7KQC/Fbb
ZFHxq3gv/Md5wuJSyyKDaqMZvG9ueTbKueBxjw/9w8hHdQEYp5aTbQLRT8JKk+ZN1RVKgrU+FupR
2H2Za+mH0Zty1EsFUmQAxVSb2KfQZk4oS+HyCXxUNxWv2qriBM6EyklK1tKM/k6I/3WgGnhwTd4T
7ghvIRXPu71OGX5410xywlQ/QpPLP3QLKBz27/oi1x1iMypoE39NWVCfV1Ol1vcPq+4fTEdLtnY/
xoQfvcNrRBlChBrpYuzZ7FYYkF1JRw70+qcGhUtzHYtAXGUlMzCANGrzxz6lz/D/7foIaqyEXRWW
I3jwcstXDM6Qk3dwEVWZxsM9zb6DmLdiKmEb59XN88QwuGkEpVMhNkEl6/pI95RwYnqt86cVAvD8
HyWWFB9W6+ksmGpNmspvgVKFpztjf1vL9svCFsL2oSLV4F80EbiakB3S0xbR3f/195FI1IpUVwYd
E2TGsxMYjZVNL7nm2DDAOdhp6oUNXFqCLxK5n+50v/fVYPQe6xqdOIkjvhyKmT6JKEgaSQ9nc/nF
qpz5HjYlnWdTwNMzhfjnyBAIR/eHLJrsW8W0TXUPZ8+ibbD+9cTFkI8PYBzIRb/wVzgZCitrafsf
E6E4JLckGlc+Ty+kKzVH1ACWITiGUx9plI0XjPCnfpknKDEFoeQi8gakqeDRwt+kOEruSVHwzx0N
ivulwG0HFez0NPZ08HCm0GyRu5K55pjOokmJYMhe/kfL1wW09ZyIsdTRMlJE7YLVS0rAl0EwpSLx
bNdXH1QZfGRLmY5qqVhQ/FfVlZmM8Q+NAKtmpslKFs0oAXmSOS0DUR56BjiEu1I1udQtSe0xjAKU
e6AKI/iTpFh8ENM2DLNGrramsTUBDFmR8XGjbZuQsppxJJkt38s+1YUtPf7i2tzA5PhPjSY/Hvra
JY9Mg+ke2n/7k1JGNFv2QKrashKCweNockf7OkQld40FAbgMmAKCS2I1t+anROGqpEkSa2/fASA4
IUUsEPdhp5IVf23p8ffE7/wC1nevMM4VfHsUMuff4ict4UzwyfsPVP5DDeAHEXhQvBV3z87Pw7b0
vHFMV/JhLQoWRJQ0dhCUkiSWwKmf/IG2b47/1OXMXnvR/CrPVQ6rGIq0XZ+sNzU2XZGGV1Et+6u3
65Ktr6SXdQMTUyORGZPufIrTflJROo+nsWjbXw3ve1GY7OCUAA9SCx5swHgfKRMU5EHjzH854IoZ
SPaELUSE/DT03hInXALr8xrKmV8bmKs/FIj2HrGGTkKr45Hl1Z7A+3t8CbMFw8IGY2Qx5EKPXCx/
yUHQeFQeoiG3TNQQJAA/g0gGdNWICyg3vDYBYkYPDlY1YvXGi5mHsoWPk1oDOgxPF3BWadt6ckcT
hXi8P9AQhjxOqKX+0P6ehyANdzBOT3e0rHlGvMsq9JD43uXPs+wQskYit4GSPZSpAgnd1Dg53URg
M/et3lI6n4D7LCpeTKg2Mm0AapBVPgcH7/9eb08zizKWM7g94aJoBoJesJdAWYVHNe3cAaWiO2Ua
DddilKbDkxr4iCICIE5xqwi6eSkbklQqaIPBEMz13m69/w2QEDu4Idc+12r5Ul1+YHj7xPluQSCq
6TAww0PTYXypFdA1GY43JDjQVvSuAm8AxXcbdH4GwW0hOaJMAQWnmfnLsCOt40c9A9L+GbJWt/lN
QbeFpancH7nbtqF70lWYuoSkhAq47m3Qr2FiCfF2EDHy70CncJAnvpNnd3BLURK78BDalGGw4/Ez
Gp7MnwM1di03zaOkGN9OGk8cKj3VQSFP+1hsIk5LZiXDKDazG4/X66ivgIaIGYBLibc8BeIe7EDr
Uen+IEc4Q5a5kBAdAggkiY4jpNU3ah27neMt/3EwmEH/hTAz9A9d4PYOzM0OsS0De5HIRN6pKnmG
1dU4E8pOeaXEGiVXd9cXD3BPV78t80SFJOI2ePMRpeGfB4GT/WlgRnfuEWfN3tCC8xL6zWG8TIqD
2zafxexO1kXhr//2kAA+li5XTaXvyhXEUmtdRUnQEJwlf5SJoDLW4ME6DCrsJp0mUMKTM+c4IPxh
TNfBElxYtqMu/TxSPhz3fE51f9gA6g1DfwuEAXOho6x6qBuxsDPRsa0baGIy00mFfUHzcmwlolVq
e7xJgQ5xnU0EdXSfdd+hX+2OiqEEhPjYeVu0cuAgdcPC4tGEEcY2rgkN3M7RV3ES7nKZJHNXXI9S
38fn0PynrRtYyL74hNZ7f1LGjRoqv0/+mchNvQ6WvR8uJNnL0DYfKAG6Q+KC8OFYuSBiB2SFk3P9
bd7vYgI0dyGVrsWiePA7mNkwroILyIWUTeiQ/caiISnzt2b+cXeIO1DWM7XIvexh1rKAiAIyJw4W
Yno2+Ll+VyzUlx2rTLaf5Fr5qPdm1h0RhSF9D22+XeEO8mqrocemoTpu+gYXnBotX9Qu0y71ktXH
BhisNJMv2LJzEa4+PIwce39ZCpSDzt4h1EDoDmM4M9mcfKhOVTFW5Ec5ByeZ15+gBcD8/k6OoZgE
D9Bozf4rslIrNyAkY7xcRL3ocFLfaR25Ph4oJlrRy+UtAYizRyNk/d+zFLxnRkHRNpmshmot6kxA
9PXSUZvQ9lRQQzf4cZ78S10PQPmrOeqdjtgQTfzEqAC+zpl079MoaX8CYJDXaE4B2ocoFNf21stP
ihmS1vdUNZA1SCedMcytyy9sDZnwHesdZbNxDWXrG4YJ0lbQwoLec0FF/YaTJp8l3/gtpNyE3Vg7
QaVQ+MlygMbLGCmFEIUACposLucZgbHZE8BmED/RfNoaivEeH0mpy9eXtJHtj/KlJ2lDXiIYwHq1
zKM6otdXjMCuTao7FiX5Dobyv+uMPbHVKCHD2aNYZMMLVqrZnYw1hGNvEItpuVy229eIjebigfNu
IJIDRhasp/U2fM0tZwfERw7k3w4NF9imUoxzzp9WiDT5tQiuYlhwEtTND5snSFRbrT00n4qowT3f
ToZ/02O2zdBWdAvgO2ICmk1eKsqwR4EWcBZJ3qaqOQgodp6KG+9SC+mRjIoodI8BFnx3ur7awWEJ
jTBiykLIgSs0lm1iZv+16lm5WDJP2/Q4PSWDQfXoidt7p5eyC/AFOXZK9oMUNAy2VhpY/Ged4eur
e7sWIvxBZAUu4KZ1VXVYzdqAki//fKn9DN7Oz6h1Dk9yMKeVnGaWeY0L8W/g676t7ov2/4zEnBt5
JkaMLwVOol1ev15Xenk87fGRGPov6tvW4t5qncuiXeJPQcrYxwO9KnGf1voYM2oOSqPhup40MDU3
F2ocTeRndmZTdJyGdPs7837ERhxIPA722nG4iL7Zd0gwj1aaR0YWbBactJCfZ7Bdah2cg8nHrqlv
KaqTY67ljNKSXIrAyKBuJycU4QH4cVM8dSWPcwRZjEpliD3GZF2e17+rpriAxbEV4ZjMcFmi4nTf
suxoOP9yY9zUxW7n0MZdvvFtu/V48NkI1Vw+cLFLhRi70xRUEZmyWayAh+NVUJHBnWFuYwOIJ9i5
7VAQvSKsSEpvR6spMm9oW0mfpyoRBDHWN6KzQcF2Jh2ifq+b4kJ4VgcQaaQl0DqHMMlP9R3EyvXF
muU2x9pKa3vifHx/CCU2F3y6qQxAYPWDG0arE9lryNAz86F5YBTN8JO2/XkBYCmpWCZiI4s1RCln
TbT3Ofeh4jUaBfwPzHlqNcIO8/m1rCVBrFNl7sxfdjPA+sX9SM4+lH0ENDCACNznr2YBGWP82a9B
HILq2yJZWzpaH3Jo52Phm8ktzb+hTK9QrWtkpyqbRz5632g0eI0SgrwC6ZSCblN6THOTPU/Fn2S+
l9BbJzSNTN+2dQq/chBDzajSMHfOyTG9B58pXKHXEsNV4jVEDciNtnwvx3Jiap56i37fTmpZmx33
Wa5m/RGYI0A7yuuuE2LzS5FzmOOJGlVsUepdxw8vrVUvZPzfmruuBzegxBfJLb+EvH+wb3oHVUck
vQbuXKYM+GR0Bm5fHq5HtSMeoMv6RTCeo9QcPS4DqvAQ6IZkOQoFL8StcftPkmpw3I0heNjp+v8q
VXZ0FApTfU0fa83S8v8R+zh1BYWj6dfimezfFY6TVS82gw93MVOYJFPt/sWVK91P4Lx6wiGPLVlt
9aYxy231zT8uW3wWfzv0NuSY8ZdIEjLPqh5TIvLXEfKX4h8LFMv5RQPNOHGOOwBWuxNvBes4pQ4d
TW4LTp3P6yGNn/ze5PzvBjdfBfPQu1Ia0bAG6+LV+m2PZIZuy/1PZy8vOND3Y6hbyfiWVDNz1Bu6
rBq6g3oMdxxyGxOxvfMtuCB8haV23jMFJWSJsDUEKW+3DjfbBNfg7fU7dcSxlp6eE4YddayydKEp
ysM4uClMisi6bTK0wi/w9cpMDhQX2UZ+Sge/hEc5APT5FJK33GnKUIB5UjPjKtQP8ykh5p9j9d3n
b/zXi8D0mPaASa3e+Y55+865wPDAQsXdlWzaD2Sl8ILsth+nTdOeRAbaBc+p35ADUxhxxG+TgUqn
2DG8hhoZ03BpPK7H3CC8PZUZ5y9VlgAR1Tgm6uSSD/9qbl/YK3Rh2CZSDP+ByU2lqxFAUFVn7qB7
UlZYpBJURH/B+a7+kjBy9mMkoyHsyK5PL537wJ2IiWNZOLWMHNAYj1j9k6D+LYhOwgTdUPxXnKpe
tZPdMj8PwGBG+SVj1T9xL4zHb4lPOP/Pcbh6I1Os1t2hY2mEAXi+z1eoGrb6A/AXBBwrXzDPNHKW
+jYTfcIQn2WdVvB9I0TLuGlPx97lBVzRlRmE/heZDtXLKXRK/DBbVPZW/xwWVWFrLh0OwSlUiw1b
jtbuZg6Yz5FsDP8XVyFeZuYnrUq9YuO1fKwcjYTuHy7jknwCeIegyCCGEFWEU+FWfJtSRI0W4kL+
7dVmZ9FX5EGgkr8vrKSswuucSFvo2iTTyCfTNATcbBwXV8G9NNcQ920mW6cfDLXxYkXyPN1HbP+B
DaWBZGxuSHzfSOe5JCbECrvJP5z06KpptYo7qtaI+Gn+PK/4wP3E9ZvOlcbRSkzLfQzRiRZMZYVS
gduWPJpylSbYBhSFj3ttXDBRBbw89MlfYsgmLQZa/HSRR46dNctzgcVH2zWkSBCH4t9fZ5FAfYHh
XFXsbV8XxMjmmiQx3Sz3yJ3pEFrrPlPinIWcJ9+81TIp4NfhlrqV2MnIdnhJSXp0+KXnVVKi0hnL
mP2AU2t0ErIjEeCNC7F1FpqIkwsCXVgRz7LoplIB4WT8PYkJqsWUAq9fET/2kUFMY0TkcXf7B5m8
wz+l2sHcXmKGsmpHwSAKGAZ7/g3TaQy97hCg1JVgoSm/4PoV8SlwZqEkLLZD2CKWlBnE9f+7iw5R
j9B9CTHTjcDgrq1P1owfR8jQB3B9mpPiwLQX+flxIMJMfwIr0tjOi99W6eiscbSbf90tPkQrLU+U
RYlMfT2M60lz8UyHPL/5ZeP1TB1MzSfxZ3VjNUYda0o1papNWHkC11PyeyoAkiCuJBBsQv5GcqSs
4DiEvCEBh2ad6PZHq25YpAUZUfVQUVxBky0DQWYRYdeEoNUyQyQ/60Cy+yvoVw4sj+6ohCX3ltCs
8cu6OiIYZRfJBsYpKZbqJwqiGa5h8s03BFaSOuVD4XWfFSrjJJuFsQm82c07r7td4n0QuRY9PBNQ
F7rCVeIaj1SILvP7oPknR7cXQDeyAnPsdDTxVal1y++K1R0zv+g9trT11FD5OFKhgF+WldBh6rBJ
NOmaRmfwsz2NVPxJmfTtty0napZB/BOd7Kuq08hF1poq5tXKXr4reg2a++Rpwu6nUBfqHT8/DVPb
fs8vUjx5tAUwL3x39kMwB+pr0OqcitL/l0af4DRNwNXNKONvqB7TnxzQGe8CgDalEpEVO9+WfR5U
okY9A9xNjkqq5Xdrt0LEYQwPuBSvXEKIvp2pgJ77qsdrCkuk994XANDp9G9XfaOoEuQWpT1AZYp7
X+6DLI+eaRSTb1Bnx9sjSHAVSKrFYiRqICsrlPpUjKTpbUP3NKxmLFH6PEmZOdeOPmi7ENOEMOZT
dmzjNsYrXH6rMM27yLbqY6+hildLmgXvamb/juIO3Ky+c85Rp9EocBYH+YFafV8BOlemUyHAMwbH
Yn+t9XkTtBK7CXEmusekTFdGANtF9SI91+f6zJd4cdq7bX0J5/5r3ijiuoqUwEDNTFE8Vkeiaohj
RpEbuFLd3V0gnPOYbZtVyasAd1tXHlQaff/tmeZlGCU3g77gQQkAzlqrlq2IyXfHc3TAisIqjmVl
ItvVZ0AMAmdkqnpy6I31bJi2hMxf85w0/eTpsNDr+PXY+mie6NuMffSkcuJ1+mJ6ghYB8uAj2YOf
+OXKQiZ+ppV8aaoxOB3SdTpzO1ieh1o3FqL5MhOopth6Tq5SgSg+DdzU6+44Nk2d1bN4Mh8xj0/v
cx0fgO/96Bi4kWyXTBRGSTlsh6bMJyQV0ddfQ7r4Aex1CCpEJ/VqeGZrO/izCi/YN3V6zy66WTD2
C0MQanjg+IXp4JRHt1fiTBlVlVDzDSSjLbgnyeEgrl4af6ahsZIcJNPXKCkBB6hP5c9PHc6D/Rs2
NT2fb2eM+UkafMNwVaCAfpyTLgEMeDZd9p6pDIa+m613tczEjq28Dx1PTLqS8SWgzItsHfi6tLaW
zNdIxr9DENKzpaBM30qxL4GOPqHybcawgHHK8j3q7Md2DEkYSTvY3o6fNT0oEJ29aPzPBWpcdr2e
Cu1ia3hpQL6+BcOa2c6xohqFJKlKm3X0umUtQGWGAp7SCs0oEBsJzYh577XLGVu98AFk1ndL5cI3
j6qXz/iBOXzx0chSaAmUMe4TWtoLF4b8EnvkOSiEYiX3yAJ6oJAOuyH5Hn2r+Dtipt4ZKpmsUrUl
2o6wZ948diMh+9zyv9XZcPStz24yYBfoJwgwiYqyXjSaC3+qn81jptsdusKceM+W9rsv232dKhau
Akb3JM2V0B53/WDb/1JK+xPXC90wMbUqScYeN+WJhG9zonmH5pkfuQg9B/cfZkMVCY6vS1SWKxH4
qaRnSh04gHylGqnrq4M4RZn8hgDU9bFjkpUl0/IVMMQgBrtWTSJ1/maMgSZBoMkfU93HZgSK/gjY
XB71ZIMoCBmuHzW6oXWMjTmVVha/Y7/K6qwTZHISqX2LTGIi4/mP8TTLshYKd99E7wp3S3W0eOVk
C8AcrdkkVzdP94YxhhgxiczOLsvHpj3wU56jFkqZk4IhXNls5aGJcNeE9VvRbPaiFAlV51q41dcn
nDcDrip8BwL0PwMkfJqii+pc2IIEM2kPLfC8rDCkquPmkfvmcs3zoffW2EZqsFmGndJxx8aXWfw0
oZjBViTRpYeGRRkDUG2/v8qRcPBQpVXCvnxJYkEaudGHtWVI186lh4C3kLtAqtTV161Zka62QbIF
oej+mhVfkPDXVH0aTMZwe+2xCdjqZJySC5t0ATrl7WiO04J3kzSa+mTcNVNFc8Yfh5cj8wlCIFGV
hIMCVfkAxmAThONNiUj7A+vp0W1hCveVwss5i1m7d90uJh7w0+f5brAgrax0PKvSwG6BzkjqPAj1
QPx5YFsow/k9cp4CRjSYmU2fdXU0I+YkhmuvtZcWlT6KP/uzOMOtjcV6xQa7jp3HJluKomR/3mlv
eh3dhZ4AvfbKEZIA2l8p+3CJW8lV2quf2IdUsByZVDIxbPB6c4ZS2yx6aQcG+gzDA8/6mPL0L/so
/wMtPs/1Ab7pXzArqkUDEciu20Dfwv9utbAlP7TXgtzoZiI29bkVRbckU2id6n5EC1yQPGpkR++1
L0F5IzTEeZFb9WwIELVqauLj7hH+1c6mU5LtP4pB5wgk22vPgJoBinhAJVFIaUghliLy/aqd61ct
pS+nOqzeD/qMlYnWLBIYggKMEWXlXpxwQ78Hr7rbFjlIRWV+UXtTr5+WsYGZ8dJzNrHUm+FxIttz
w+qHqmAENu6zOV4iENbF2qndDWZ7VUwP4ZYcLw4DYxqiIS2vG2OMirdABpKL8IgAaVzCCeavwDoz
dxFDpxV19xuzwWlS8TVmGGeemVrCXbVET/Xtzso2Hl2Jb7nkFGWpJN00K2x8pKGKaC9t55maD/9J
02panMbhWKA2c1jfBoBrM7/RarFKgYctmytX9B7/vcmbrFlgZHFMdomcXP3f5mA6E9Pl2sqG+2pe
M+KSMdfC9JTw0SDxyYVtd6S2B6wVKK35RC7fyARsrtJWQRFuxpslxU7dGexzURyav2ooG7y2Brsh
D8NOIREfyCxMB9SQ9rhi426MiaOv4TBe/LD1f9qXzibRBC+5Du61PJY0q7CeIpE8uHw/xr+9V3bM
Xckd1Qpptt9RnzExLJd7nmEElWp20p/xrHBRTLl+RUasgKmAnO+VxXu4oQxiP6B82wd4nIfJInoj
JTfvr1CMOAtJIKtLD9sv8SOypCKRU8fFA2Odyy0iXdzURkM2s/JNl+uPuuf/tm/tZM4JSjpt17Hd
UahMJ6MqzZwIExLYxjivgph+EsnnmRwtdNb4+uYK8/AFzk9kwslN1StRgU+qDoroZSqmdTkfOKcA
DQqWzZOhXFQdUXGVhqPrL9OnR70MVgI2/l5Cuuf2gTOBcOVRyDjrpQKN6c3V6UlWnJmntAW0qmmU
0GRpyOZbjiPeKVK13HP+KBPALTNCQ3u/f+SYn48pyea+shpzwy8qibikrvXI+GdGs8eY9EWd+msk
K4K1CQYY1MyjCDnYKwqYKJlHPAI5g8fIRyRGveQIPKPd5uQ73lypFUsICO99dsmMTZUDZbL7DQkp
yo7WYtAIHz7M8ET5kflI9qu+m5Sm/bNOA43SDZWzSqZOyMcVmhyLJjo12aCJNKciIIVEOJJ0qihC
sOly+LYrAkaSQe38INIFflL9jo4+tujbyPy9HkFzCMNZcmMj05T0vWfB7TRh/sA7v2hqjSsjyueX
08obzsf9LgPbpV0FLHcmhDKkePKuCCndjlVQQ/QeXODeumDBTr6Bti1vJC2XMulan84Z0tcsZS4/
iYtlfCSKL1SstiDk7xPWn4VYtBoEX++fA7hsNH/Zw+8Gw4GTyDAapSC552mSnsRtnEFMzArtdFR2
58cItj44y9Emxgry/3+5XTJU3GdfsHAE16Y5H+geeRH5y4JaONhu+9ZR3MX0jOXjBJiv5PwMwHmA
/MEP5OqPgMPjq04bDtIkZ2UCaFtz60oxyQ760sokL7hNgy5mUg1idpLazoxNX/6U7yiksxraCpUJ
sXM21fqyRjVANeeh5/jUwrd+ZVuR/eBIN8j3Glel9hbh5Xd0ZTAt787BgLQtS8/U1E2X7aNsquGS
cmyQEnBGlxgdoFTBd+s/y0UhIY3diFyK2aKNuPImW+nQfkUPEmqQSIjisA4Axvmzz8KujPhJ9Ftq
3AzGxsqpn+5qJhQnJaiTJARxINUgvnrzfCSrGywLza8hSvBBUzP9gP+tzl+RjQ6rTb1QuZMIWoOc
tw0TVXIPNBA0AAq6uK9+A41+6Ja3Iy91XogKi3iippi/ujMis+biBPV6pVcbO0524pSAGy3Yw3xH
/89F8+00/oGQW99BiojtE5BeMg0Coex1ob8+M45HA0FFXK2H9nJBcoR+Wd9sMg/fnKJXVZz0nuGJ
sEA7eir0Ib36y4TrBw091V9PXH42Bxc+9wmkXg5B8vxxdnGFgR5YVBuU4H2mFSsQqDoRW3ek8aKN
PvmghUf0RdyxuuUdcPKz/VYKGavSIFIJqWWWV80F+33e9GUykbqMyr5gkroXOrQf4qhfhF5HwhIg
ivmpxJGFUpPrjy8uvlOsgMymEdUkUswCnhU3h7jcj584D0NUwQsMa4ODa1YyjHO/ZopUC5RR1BZY
PbF3ECVAmbN1vrZer0uXXHJD/DavYGQuP3tGMh//cDsLN2xqvqfqShfVrr0OOyZsQATdV+bHeon4
hMTgTpP2PM9yO2KquGweqA32ouSK/vgXj6i9b/9pR2+SW/1+eEiKq81qkwd43cYoKd5xhNfMSckB
7jAd+6Nm5mNLwsuq22rQCNUvIK9nUzRJr0JOh78qdVZYCRpaRJT9nho+Q7+hNI/Dq7Gp3m3ZwFOM
JM5vL8Q8j26wJeq6hU1uQ9pkFyrwAp47pug0C8nuflDhF3F911mIXgMaevu5f8bDg7qAYsNczB7x
egns1uIQTJq/WwbweyHUbVU1iL0PXC+jc9TC0vY3vtbPIXt1qyX2zve7SfSZKZHoLw2pPrcdBJDb
wmNdmo73yGsbmcogWUzQveCTf0bVvoEpT9fLY3ZFHgFamEDQrpaew65k9oajRhw+oo8RfiDoJhEA
Wr7qxuwYw9C8CvCjVBaNKX4Y2aE8O9UO+Aw5uQMIQ2mclWBkCQvlovuV/iWed0PdEkt8cWM4lq8/
q4c+oOpiFkbox0yvTVF/Z0qGsF7v4cDJ7tyhXB0OrypZ8aiD7RRlLuw1V4ro73D/I/lmDf99qhSF
ZEyNnh8aXo6XpjKyndw1KIXIAQ7zlkOOJ0z54LZ0DJ3awCzNogAzMxIl4XBsdD8pucQ8kTxhfNOL
MgricmK6cwSt87+DcA2j85FbIb9x+69yI/yqVracSCBvTKCGxCPUIyBpXyTPvXtI7/Cgojjsf1D8
rp061NL3w6SOm1pyBB3EvWwgaA97hrPAlRzDRCADYo8D7aKEaAJusbTRtVCwFz2mCK1lA9OfmZgJ
hsvcgjdJt8llhVGbCf6a0RgRC7smFCNRvMDKc2vKEs03IOAi2CmMZL2wRg8LkSSEyyUB4iJdVH7j
NRH7XMbiqVDmwPrUuX/seuMhj/m1g8/vPseB7DYNODitP5AB6fwFN3funobToBhhHAZry+bnR0Wh
sS4bGepVVYbTakQ3eLx04A3nV1loWCEMHpJ3MxiT2lSJ8Pf6P7r7JSlbAQOYeWPKoEi2r5SrOGfE
xe8P+amBKlaGWuNCQCWK1olj4x6K6HjnQjnF54wcw283xplKJxXvvd6IVT1FXZJEeTiOYTOFM4ut
FbbDY9rE+kKsZUzZIdXkckY4y9pJvrB1+qH+n0Xgj+UQzvoctbxCRIjeaAz7ubRRko+dhwyZQlVB
eywwA/HuZ+ATmk3DFDt2OwZUW8ilEpMMxc/XZo94wI6cRaB1ZH6gZ6UW0UoZfTnsz0T/f4qCIctO
jbFkLqKrGzOdw5IlOTZcxhWMBhJEpbbQdzG1bqB5m4LpFM3O2J2n4N5W/rde1YcuYKEl+TiUFWKi
JNqZ595RmYB2+QFKB9vkSW3psQWZFLzfhzWVzEe1G2ag29ve9fA/1VtrGvtQ9rsWmSiXyHGKUxZG
pb6TF9kC62VYujqM+f7cK/DAI5dUfcNR1iD1BbA0fuBG0RNxgZjHAyvA1H2V6cpk0tjdpIS/DVkE
RGYd69o53RVgO5MQKAxeKOymJm6mXGSJ+o1OnsSt11L8xHfBx0p5H6tqtWC9xypiHcB8hwn9qZYG
4lYcL8CbkPXoCSYhZvB9hetCabylM+vBT8kkEQbziRtOK2fmtzy5bcb9pdml1gnfsCoT9HQ3s3yB
5QLVVwK9meyaN6RHVKF3ACp/StZpINR6jAWYMTD7X/9bsNa+zfMVuTN1DO2wOuos98/4SCy/D4DZ
N5tVOvV7hALxDOTw0NbgDIfNW9GfvrKzd11lXSAGGrAO6ZSPKLtIxmZlNLhhDV9O5/TRcqtvWCx2
b6C4wHCmeOTL+E7Hyhq9LSyhMNhAkZFSm0E3v9wXNvV5xYq8s5y/ZfvI/p3JDGDdlmPeaQB1VMpW
x59PoC5JqZvdlHQ35YeeMe30B3O7qXC7HsS9MuveS6NwvCYKit1eO3nC82qHEFhlFLmei8hb85l4
ibndLiBRrinOfTwUWSqrG9L9AVLjXGhYyeQ9AJo3P9EssElYnYBpnwZmPcj9+NSdkX2qHQ5gFN4Q
tuY8uBC7qnDIQyuU9LR7Ye1eXPJqIejjlVwNCgxWABiAkKZu33lO2k0pmLX3/G1aaHYGYyLIYHnp
4p/R9JbW+Yl1SRGio1KE5sJX+nMwQVQLNeHlKOFEeaFiZKi6Ii4tPpW03CALSrCOz9JeeAXwpHOs
hhUvRdLnTgFx30cY1O3yNZ6uC7n5Ie3413lQsBrqFgKgTyXQ9PUirmD7qdG7uQmM80nShpcr2s9Z
Oeu115RaKnV7V4H9vlurgI0qcyDZgu4CGQ65fggnSswA+I6tjXmZnZZ8PajK43hEoWMyEPWMr0cd
Bwxgb9UV1M1PtukgLGgUzwholRSDNNIV9pLQ0e1RiBSgcvQU6lsN+VnBr0IyYpXBYI0sT7iwXmP0
+VuyuzmO+LTjrKBqg8xwAx6ANKDSpJUfMhEp1zPFu8mEWixff2KNMbAY7/fcPZpHXz+M1UQRg+/Z
m/UpNzg+x/gvuajwa3dW3Aya3Ds4gKW2IVLLwp8Yi39FNm8bRsZG8+OiwL5yiFgPNBn0ofeuutB5
F73R1XfpbfnbILlYuK3ngiO6rOqWAaRMzvs3o24thH3JyhMtFTqFee8A2fy/TU683/Iwd6MR4Z1B
wLYr9latoIGWu1WRaMKfMRxfX/8IZOWq7FDHRlk0Gthq2uUq8OrsNmDTmiii/3QRt/RHE55Xwr62
yDw3SoU4PmYF13lyQezt0/bQcpsz3ATkVoFOXByZMl27OMchUHnghsZjZdcMFOf20f0/DMz0nj5h
Tg/Y3bK6Yo6ns5C+yLY8VbOHTrfBA9Dwy2pvxCIRXljWVnpZyL9qRBiMjJRX9TvIKvm4wtkw9JKL
0SF3Z8wfv2zF3FdKnpt4/YTpg6uhb7EyAEuTlS5zFNCReOAnlgMSkJqwSuT6Uf1x6Etk1Yf2KTsw
yGSvTNEvtAWEFYOlAF3Y9UpkFDPm3f5kaYRjNBfYLMcd2UOmtsQz9XSvsWXDH4KOG45mX5PsR6CS
hKu3kbx5gQKss/a1YdhsyLm3QUagOlaObS7fokw7KXjvNeIC/ubgwVFWlcfc155x+zly5faKTFyE
Rd396HYtAaz45qG9Ue0UobAbia4nbTnldYE+2OqBc9aZPdFxXJVc1E2mob0ltLMWFWDuwBbGX7uP
FnsfISWXLDgRTP1eZZfdHS9Ya5vOvs7+/+5NRwrvp8cf6BSEgLpZEjzYKjGXBTVerGNdsWA5dDlZ
KbdkTdlyiE266HJ37+j1qQl+6xP60h+oX7COL9yuAZXfS/w2/o+6Vj4hHS4ozrx59ME6eUMf/0he
yf6i/ttCrC8cyGIH/TmP9hiMahQb7GhkHXEf2IiqQkYdE3ycZEooDqooWhO4TlKqNTE/iJW+vNIc
C6B5MYb4DkYxQySVhsOkc1zPtLKTlmpG+BRR4ZGcfm5YSNVMFWz3kGtgo44EthC6DIngk4lQxSey
pe/yexygJQuPICQnwIwFtB+sYYAlA3ohlQz4c0RG+hDg/QmBtvaqtvjPxoFiQ9v6kSo6MjDH37R6
aVmUzUz3ZkV6SNHIXA37qdcS4cpLggB2bYcxG0Whwln8s6RdxHopYDZrU0UpuyIJlnLeCSNI7ouU
8YNeOFt75wFTkpMYC/GPOeDIzH1MnmwVlX0jRGAv4NTy6kpkwZUXJbMDmKdWCzNHhIXzilBg/6UH
6mWmQC5yje3ngH3FY8Dmd1TmkyIbuzXekPK1XsCjnoAxMsqaoYc+0U1J+81B1D2egToEH4N6aS+t
Tn6pynn3DTssFpeTNdpjxc6IqUGt+fyZ6v51bDWCBF3ey41gZ7rJ24oxEc3Zd4ie5PYEyq8d9ur6
1hexhNSZjhPHdyAIG7i6PAQw5lH7PFR38EkTw1JlrwiPgaf7fkRYOgZQ8LdbT3dlvNT/HvFuy4nQ
TkzX1qp2MSMJH20zmbMcTHgZXddDW59UVoAPhaUnY0w3sRito+rXw2zbyV07FyGJ7XEUYpP8/LGS
+NWHvOYIShh/etg0P35n3MKyPXbUX0vZT7blp6MIcGbqIF7dleTYLL6vBs7SVuTCncG5/uVSgWUZ
bz3zuKcRVDoBHZaC3EaHh9ULDUvMEbzaOC6h3elhstwGD1oBIpxsEHM2eEN0SdgqMeyzVvvTr/Mh
b49w6w20T/ODx6kM6lO0fnGfA5i4yB+jA4CV3O1tIQRGwPZXEafKuTY8kap+S/YnQosrm7mg0w64
/rwUlagRGwkdSX9aWZLkaUrituR1fZNv92bW/7dCSgc9cW/Sib8Aun0OrjeWm7I32PQODgqkPF9F
cxfFrJ/kqG9twwzXSmM4F1gQt6/rv+xXV418oUt4w+P/IGrC9ov7HCBBQ5Z4QbirVMGKPGcCT0Vo
XqQwfOS1SJSPZ9RSw4efTJ7bOZFaC6VoF8rUQvsFOR2WmdQkj5QITUe755sg4ReHl0LOtuVnIiU9
YczGDJRqux1HkigQ51VQ8Wy77TcQg9zacldCLwZ+VUCq/wXp3dEryD7/5h3zgC6PNFu82tYDeTqP
AcNHQsKfilLcq2iq7qxwiGZzmYq4eBGv8vsv1T/XdwJS3plJ6V/MTuhGXuhX210yaS5sYcFfXKGt
QILgCU5RaDRoBVsqQ4HsgPfCIOTgj2DHLIDZjwfSXhfgCn1nK9OVXsikoYAXbN6Vl+Bnw7q6yRMn
EuVVGHmISqfOB++fybcIsIpxgKDBnawOevg3ZiAmqugLBHMW7fTLWqi6RMS9gcXe44osw0kwWRO+
4rckPk14fppP16OZjeGhoxPhRpJDqIwfcUR3T1Z4x4PBi0S7prWUHTIY5CaL/ddF9OElCOQAbi7H
wTi3iJLm31Z2Ilg+FWwOv43u5PMBV7PtBd6GrMq9OB7dIx3xLQcq5Av6yjyu0UyPKO4jN2MQC81H
87YV8k7RZrXP+MSKmN1SofPkJA7TR6z7HK1tMtroS/SpyUpUI7DGTyyeva1Rn2fGeGFeoNcLfXst
hDvsp0b031VQ32PFRjwATq1EPlQ1VEP1icbFZyPVkVTI6q5AVKrHy9frsCjTY0YF6QETdExZk8qj
U16k2Cpt1+e9D24MgezRnYXi78odLRv4Ek+6n9NjfOzhdPfdKA8d3nhWcI5N1vMVeUugrXJRfHQX
Pevm8785zs4wnKSZeJ300VmBk5XUm1Jm9NaIZjQdfYAUKsSgYvkZxmOtEYJBIfA3jIhngQ5xkuon
paHijAglli6fOEU9RAVQEEJ+3IekOEi4vfRjOWZD/OnbfZMB5GfphktoFI2EwmPuT4qDXNwFVAqb
LIENKK0Pmsks9L6IC7b1ZllgoUJVBOxSnjW1HQob7oh/HDoWCAcoW51efluwaLUxVyihDntTFqpe
llbqLCE1WTZkKyENKRFYUJtlXNNDfpTSMiF4EotYw2xoYwl475ujnMVANS7dKO8UZ8e+NcgbiXcZ
WWWo474GHCxLsE6VfA5xRM7AWghPVFT5BxcKHf93hsjaPnGyUAn9weDmLq/2h0MMiJ9Qc9mKa7L7
6XsEEn2Dy17pF6pmip38cPmIL5jFC2BisyOzguaKPt7HXY5XJxFkQO+uaW4L9JiMFqtM995ikgqs
2VsS6wEOuhzMzRWfbG3ETB/aeSTduHEcIXlBwb5c9SaoLm9T4CK0yc8kXeOZ8Yx1l5lWTnKu38Z7
+Iis2i+OJn2VsPd/Gj7cfUtxlIW7d7l7QfH8ILKJhsqsVmWME/kNMDoUfu/p/HfAyt94nRJEGN/M
CoLtDHd/dRY8qoXNQQfLBFx+7YOhwtPwuBd0sVKs/ApBedcXfgVWm6VBe/wi4XgsBimggvP7eP/U
uN1OIdJHn2HmhlOePEJV0Eg/W35d41SrxgwtAYeIT1+DMuqMAEiCeeGlj6XMp4aR5U7IJ/+0xfWJ
dL7IUSpqs8WdddG3fLSDqfrNtn0LyThlwLlSp7TspUBpzYbcDJgZSY/iXplSpKJVUhn8V6++AVVT
zrdbrZbPJbjGHfdsG9+U0NSUDoYK8Cuf6tKoluq0seSVjPxqsTS/LhcBriG9BTFWMj78OyvWFXhA
lMyWv/YebRKDZs2X6tLnAcZuLD6yuXh9M0qgrGnmijZZpzYjiTxlpBFmmRloOzCAWqxwPUBfUcgZ
yCJDfOFuqqg77mYVB6QyX50EHmXEkFAhcCd/A6j5LKzX7sVztivai++hP/2wf42QLqvgX4ch6Kwq
1RLOTw9Hcy5qCtRFVrBsJM28KQu5NNxAnPBr1pEkfccK2l/dZyWC8erqFIhKsngLhyX30kGOkZQs
jbStLIVztWAc18dzew8+QGtwCPoI4AM2vhEhifCvplLTUhhMtXbYxqniAEhBUV5Y5myECj248xYc
TEVJqCAA3kOvPau164bSaFgLHutGptUyH5zSnkGOhqxcSU9qBU1a/aL8GosEDm91GucrEzHDcQ6q
+l4V1c3ePBqvHGWlDyE69Vo0WClgAyk0lqwundvFBL/8+pEh+2+GdF/ezaO1j2gaPiXfy1FI+z2h
fmMsgXAB3JeZDiW1aYX726/D3W8HFDLFQ1hnI0L8y82PmIOjb5Mw6MEzEdBHnlO67sB+g19rZ6Xa
5T7DzEW4s6xRLAIElJY4aIP+aC8kM3m8uip368AXFzME/2SLiC6C8DqpbqX866IhgDdzsRdtzypJ
9/6BOUh4fHBFDM0mGD5DDMP4DGHQ/jKTyR0mzQPIS452ph0zCDda973sDCGMcY3klbkvEP8py0VK
Qydi+q6kqN0KpS0abal6x+RbNa4xqCjecMJOYLaWqR1iefvmWKCexEGwGS/Be0foBu5o1wso6LjF
eeokhoXb/FY7ZvPzfJxvzCOv6XLZFL3GxUId9NGWpa512oK0Jth/My2x8ltFwNm81ACtRUgHDeWr
/YEr39a1SD+8r4BuKtkYa43Zbg2Wd8rFe1LgCm1QQ0IDQkcFbO9iLirnlAdWEpGmxggA/PM7uN51
w3G0W3Bsu32IZLJG3y+wX+9tz/rKU6C1YwBSmbj2tfBqUPlJfuM784WULUfWblrDYiXFVnpNSIPM
cSnEU7gCXkWWM68asAt7meHBHp1NSSgeTRgtLeovh+84kQpwjQvrJP2QOtLfrEx2fDfygoJ765jl
w4MIlR3WQpUJ3SbeMc9nEgeveckAwLQrHRvEBbRGyNsiDzauVhnv5iNRgNFWpfi7Ua2cLlq282an
8oCZVz6DLRuU1yfEomrxqewmZW5c/k4COhG5fgHRCKaDb61Zeut15yjBbjC2WsodYJ77wXaa0dqs
97fIXJtKf+Huoip7dhB8mzZZ4jHka8uwkiUEKytQ5zbszCp2wEcEcVSy+JECkJcpvxTW9Gjz1E9k
IYIIM2rJmxIpJ/xRF1EGRVxmgrrCqB+SbIdQh+Oid+9Fh9N8TphBTEI/yuB3gax8RnE6utnNWT46
UleDF+MUGS1hxFWjNIG+yyB7D7vgh1jy+L73sA6UoFOWexNkxIU38s5IbMVGaanU6ZVDC2VQD0PU
LZ7o3meiUEU5eDIUjLpSHonewmQkXqXdd/RZQQZ+xf2LMYpmjJDLEYMN5id06P2vUPkzr+qU+IsM
d02aYbyN7wREUABmOIyeYeQuFvwXcKQYjhKmGLw0tNH9xMP7ODElLV6XE00sEF/mWPIcRxOVncMU
N+sAeOBj1DOisxZu0z1phYrXQPv5kQctkypVcM25iZpEpMvxjeh7qy0hXTcpi/8a3zFK+pO8UAnu
E+qQSWhrcvOoTr74/BKUHrt9HZzcxwoWIBq3A/65mtUdthAzWYARS+osHI5tJRQ3L3E2mEoh7DIj
whs7QVcWMJ1uZvgTUV/ZkqecN+vqD/qdkWGZpkI3tTaTRQC+tedXy7IajL+AjA6Y0uF9QUMtvV6I
pETAuMqMDKRpmaTrAdS4IqBJoFVIXsUXxV6/K0VSIwuFS2eHosx2++kK7VkrvP7XveHDicQ3uUVe
bxGMncf2JH9Mbyx+X6wuK5+IvYskhirLxgb4fRnAHAuZdWvACfz7aj5CdhBlzokKveoQ0TaJMyLV
v4uCzJ2Ph2+MPvjw7zszpnXP9bG+OYN6NUPhR1aKTeGZoYHH+n+PqDjdVicwD73vgeqD+u+KGhIv
OR9JcuulsIUNOl93kbfhvqO4PKYusyKzh+p3s8BIHi5W3eMKeNRtYG1pGxFqN3IWUpUt97zilOvD
gKtpTPgD2s5mnuSu/T4oyxX56FBwSMcPPl5L4xftQVCvP3jlCe+xmZFXKwjyt4pxlAaagszQh9JY
1j7K1e9gnJtLEayu2CDyRtF6XC6xciuUoYjrkPPpkuPA4DSL/LVmU+pAHlNqe6gGTiuIfSxfmHLk
Hzj7wMKcaXeO55/WqecLbRGR85AqYrqs3cY+y+it9VsT4nxonPILwMbOuoz5TcKdCCcCEJwgSsg9
Z2407MBzTFH0whxcftSWHBA64qipoAzeTVUbg8ZAt6wbNPuGNi3dZsqxMiBgIYcV5g/DfMK8IrOc
FiyA+gAC47kLliK9wSCA/Hko5QT1qE41zR72k1CWWNbO4AKi8+3XUbliBWdaWMMB9RyolroDJwPb
ULeFipol3MCHVtia3dJJoM7wg7VE/rP72EP1RXpJmjJWDSQTEEoQ8pno22jW+oSt75R6kvceJ2ET
vpfe716O1yHOznE8p6fGnUri60CwVdjyyBJqk469IDB5vu/y4xw6bkscoO9z+RM0KCCx1Q5E7ibK
fidSQMcr7HuMPldxVBfLsG9J3truU2EmITz5pS5Z4bUyo0v61zxqmfP6quDbLzmPO7Xtmxu9YuCB
Lj1a0cUFupb3HhjuoQDkpreVfF0jVowZ/0GcrhQzTjxIUn6rJ0J2BfllLWSPEPYmOeK8V0aA4j9E
0VzRNht+IboE+B9YzP3gLEVkpVVN9Q7FdakfrokKDABFuUbMaRSYBHRCz4th1UjmViM7etmY8RPV
iOAuqeMvOGgiP97v9YwfdEHFz/BwZ6sMwDOvx+WyVc3zUgtUHb1FHxdgm2o64x3VdAzxWKAdfZ0U
USqyuaoPpB32vhIcdY01jnrS6vyd24joUyCsTcU8jXlTlxLg4V6gkAUi8xb+zEHZ0xksDaF1T4Vt
O+2US/RFvaU1mzbWWi8SIQyFxkh6hpj/1WlaMVd08GMApMGM/yl6s8V7xyTriXNRZKMfCgMivqy5
slLirkLXfNcJsmQWmoHoLpH3btJPdyg48XwY9enzR3toOhF2vot1Zs6UbDumkn9PGmSTVFtN9EbY
lAYf3liF+fFhdesi7EMiY68Pj8jbHtf3hYkj2Tagv6wdSNM9nQ9i6PxutOF7z/hfPQhahxYmQpUg
jPwLfaPjDxPy4S10MqRlGfH5feVGAQvnOUm4EOclXK67DnC6cfjL/RpTeFqBS+dpVm643Y9EFfsf
z11k9F6IAYpr/t5nY8rvKrBL5vCb3mWIDORFvVfu0qK2JRCjZBSGETvG/+iwW1jrfaTVepu7cvar
wv9OWK3LKodtpcqwXqzJ+Yvk1/eBvtOyEKIYdHgFGuPPXBIAmPRFrva8oQDQNU27qHY6aw6DFkgc
Ajy2jKlyrMTHUto/JChDIA3khhB/F66IdJal8G0ig8DXIZmhM8ZF6kv0ouEHPJaKEZdFlVSMv9eA
3XEV6vqlpZQ5zV3Ao3K4pY5kdOKTw1KuNxwt6CdPvUV7aqcNOcXhpeNzO3atqWWD2qVOWLA4Tc0K
3hWbxTQkcBy64PHP+nF5yqCpZd06dY9pybQqyod8z1/MLY22OBhyk1sPQBCEDbaGOL36rY97an3X
FYDAPoCdiUeT/fF8PaFguf/IgwAIlo/w+JNLMIbYUAOvBDmICA4IVWVcehOPMcTZXg4tyVgXXU8m
JtfNLT9gMEROOdjXV4GhrgjDfLK/P+QHS8G5FpVPuRLVmVLfMLNd2BGSuN22T1DVovlQOlptHuoN
W8MHJB4hYSYUlU16D2rAPPxt8TBvR2jwALHq5zWJ+Yt4JllEGfXkYgZCbiY1USo+ONWBfY5atpdt
ZkEzygmBinLKJqexrm0EiyDpQRnTeT520+aJkK88DShfoM9d68y0kV1BeIktgAfixGT1qjQYkxNa
tqHK7hFn9HGuEIKhcbyJM8dbvrd5CfFvT5CohMNRusHOwb4IZaJUUrEsc0yxGy78bHMdRn5lSFmO
VeVbvm9BgwvN8oesrHJSHAwDs9zeNQtb2jeHbwBMWR1oNPpG+cKnea54v7wTLrmWI1cc7QgbZmFi
DMDRdc/QrF+oF3g2Jl/pKVtrbFqrEJwt83dOJhXGK63BfUK6yY3efVTX3IGQgsEVzC1m1DEcAUov
zf7N84P3C2ofWh/A5Ioa18kXsolDAqTrTSpf5z2Ebdl/STA6fHFG7J3qbRY28Fawhud+P4dNKF/u
9AsncLdXBpvGLYojxhxEroxE0RKa4FHxbxyY8mywWZWisd2Lj5pgAnJJR+mebsAyj1R2m2e+boex
5fpomiBzzW1S0Cdm+b5R9qkZTOszKy/RivDKCzWFx/WAG/xrAGhKFxgWBMdzpinvcmWI2VO/7HRv
+0TWlAJJSUfMzBQnuZattmcGS5mVzUbg+eb5muPrxs/Q9+snQeHiCuQHStOQfvDeufYC+udWxP4g
a2zuZtzlq7RAMesWt2hzNkD3Dr7NeF+aujL4b5zYF+ecOdtosuPWhZP8NPC1fKG8D9vE9olvlqAG
7B+2vYPyE3NaodxMGv8HjUpXcM41iccOB21X8+lW6/u3mAfV5Wb6ivM8z8aibHYA3rWiavEl0ASD
w/V5r5EKS2Ipk13/wocze8voLkTrMspVeNMvuNz3i9L2DodrgHrzDJu7nrGWcFpgINmKSV7pjmY6
f7v7xHD8bkqBXmoF+FFTahCt61dpv/I6e+QmTL9L8Btb8MldXHFxVWXQWg4UMlGS0Oeb/H8LHYxj
6al23ofEMOYGJeltxVbzUQNdYrl6GKXa2JQE3ib0u70kGj3ZWWAClc+K4MINkP/oEpUZOKEEGyPd
IWyVfioyorD+L081A3bHXcfeazCIuhbgbzC7KbAe5V7Epi6naT2g6ANJz2ea6aQ77SeyyZThWRlK
kPr4SZfJEhjMFXnQ2t/86NBrG3TuEv1qlooJda/hRjhIObUrIOh6Km7diqpozCmnX+0XBoTGVxTq
WxPZu1SbxpIE706qxmILHHBbtW9vi17OUReZuOCfC48OUBYOmH51lKAr5ECuXUwsPUAXGcGsBHGo
RV9FqNAh6Y+xkixIIGD36k5n4xEpbqqnPLtOUt96ZX0TsAW8Vs/5w0wQFQzm45HSPtdpO7FE3meK
tlQUdYib6brpTU2Z63TQ88FZ1OqN2cTYyuztH0OLNkW4TFVPfIYQ19r9hBLL63FS/H0xcnWoo1n+
InVTEmz1JrXB8pAgTwnTZYm22jRonTUU6AdMts9urV+DwG0+5VBnq7+1d0bRffFmXtDikGV2CDoX
PYaN1pAaUDA9kVVLxnOWiNf+Kv0NaPLM2/VkKpfZc6vI/WPrLVc9ZNKBeF9Ite+MsAewHoiJM1ia
K7AvcJIUZ/3iqNqdVgbCxLvUcbu9puHtRx9I0UibWoHR3/rNAkIpd1MSRYlnRP8hzvtIQdVtX4Jm
+lhvSqtd+oWwVl8SUJvkpnmuHz7fK0zj21nQMblGW6ZziEnK8Xd5d2JnHuE6AgkOdg1v1KuYbGUg
MDwbjOlGmk7grBjlWcvB4Trg9eM6pBIr+S2r6x5XxDlS6J+AuUjJOsH13WHVO+EwXJHOjG2AVwuJ
wQ6rs96PMIf7irdOa3SXIYE1hNGeEa0t0fS603SbInDDdMJRuthT+9Y1jUBsH8V0tCI7IDB9ZDji
bmJlooBlZ6pRNM1Qgg+RPflg5r/JePAxeH3zE3AULkvCmVx5GFBoLR/vyLPbasBDLdRZ4LhGmj7D
jCd1WR6Il/0bVmYG/Ki9HDp7w4ahwG/QpMpeZwTNIgt1z7cDNX8Zhr2dRT8bwRok3WELBQ0YZty7
jcjxMcLTqblGDc2DXJd1GL2GAZRw8Rq89VTel7OEFPN8YyEJ0Aaaihy3ZTOVlm8NoV06qnchVBQ/
guEIjjRtPRqjXCAmq0aoRwpkxH+LEuflWOasevyLKnIPi/rUtklj6y2VRmx/l85XCZY6N2wYjsP5
DhuRV7U+H10HlWZOykGe08x6qKN75u1CYu/7+L87f3vKcsUk0RvGw2RPQIKUE0Aep7yN5S9rMyVY
GYgBxfEghGg6Hm6oz7Qw2UbWsBfPtRmhgNWbALC6k0dsLMkZTiauT8lyBipBC7PD5IDkpjiyJ7ho
1KhJ2v6dN9nQIiCM+HWrmyFUxL7doO0qH7Y6A0EnYGldzStX4vzU8K0arEAg9HD3X6y4ZYT2FCq9
DERYJ4/K5lVTCe2lWjGi7CEJWdipAfYq4aaf8Z7x6EUtfmUFs42dFE5zHrsbL7dJzNHvizXqqYcs
O0C4DpzgeJ1o2mGIS6uhDcdhyVoFaMNHv+B6138BTInFy+G5m9iD8AP1XpjkAvrq424Io8O9vOwC
3PBQlQzxzjf7pPUFsLNCOHA/03FOQuISWOXzCnUjpe+Z0KAlPytBCg3Ha6kKjr98U8DY0SANUkwD
wUN2aDZm0z44ACQyX4PQpPi0bq8OITEYKv4NrN8v8NqhlIFa4w5IW5sBYeEXm0cF18PxAzgF3k/6
V+vSNlSJX1o6DYUownlxmvaz/pxTFKJAoPxLCPw27ovpLq8jmipYyYk9CgcW6Gae70PLNWyWEtle
ddlIwCF6mBGjLy8DoNfmsMUfvcJglod294gav2krjrxU2fv3evThIkppjyrCsn/L+XwRExwxnVxR
3QiA7lwgwrhJfGiwnJiq5hSCxFlvl2DE3lKHpjLrc3FMWUO9GRc4MugKVlLWsmwejnUEXmixApUp
wagyDuqBdaw3IZ4hj6dxVgcFb9txcnStwzyvof3ISJ1H3aAP4qh/IsAscK9+KmE1puThkpWXgnCz
k9mFoqbPBGBLjozwJy6H5r0m3VX7SkL2CIWaAvp1110z+fdezG6Dtfu2PaSAA5QCpmzFdnuTkvps
XXkHNhzYBAEhrSk9CMdM+fSZt7I3Qq+qGGo5b5R7VpIDudQWWXU4W53zgBOjj+gEekl0DagszTqJ
e2rUB+H3+A3mB0nQpO9kZ000sPAS2TibYzAxb7KD0zZfj/JN4vj7wLx3ou1n2X5S8S3LO3pQL/1C
LvQiSXA92fzXTDdIEpPKo/MLb9SjV3aWqpuTfHZ7msyPNv8dalD/N5jqO0FcXA2at1+CcHrMfw+7
Lqs374AIWs6rnuudMi8H9JRG3kLr8JSzgqf/p/bfhY4aKsJeHrEvwH6gQ1dVC6vGhah6YcEyIQNH
+Tlv71nViGjQRs9kbpmzIwHAJZek+MVLTZlruCinAH8n/iLapRidTnG8CkPst/ANGnn1ncakD0so
Sq4RBycM2j/p/pGjqPhtJzhIhyzei5qtc+E5y0BPFk2NeeKv46n2S2CIFbhDISX9ujhrhclHe26f
2UtAx0TXrYlHATGphcDE6lTTfPP3Qkt3uYoC46Kwh1KJUphzSQeJAw+KiMc0258TE4grW6MQbnZE
V41Qwws4+mPRL6HnF8y7i/CSB1W5U3SLDHD/kVHR6wCJrLZCwuRXRQgsFVSrc+e+bPO2ZdJG6ZKu
4lCgs62szXdjFbsSvaCSPbBbPEdqYWh3+cmFvLf3zOczZ+vWgS9AqyRuR1dx6+Qf0duz3lSOzPQO
hiNGc8TuffNRX9b9tRS3+Cf+tyFzxoaaTsnPD0cMBU0dYpUXYD0yK9lBSishjwbo+ONdZ4HDVLov
6srq018wsD2ZEr8Dlg3lj7FLgM72FZRCc40mZuKvFU2hKdhDcwNsg4+Eqq9Q6++J4OcZzu1ILSZ5
iRq7xGSH7Pwt4K/WyomeuDLyxTrEgUdNjPtSRIXFUbrYMxCPRrMEwZG0QwXmdtYUW7ukCD9kNXgE
xAbFvf4porL+5Q2w2QgAY6tFjogPhrRgi5h8eiy1p5GIRXdsxhf13UELQ7tdDOWV2xLbERaPjgk9
jMNhazXFOHwxkC5uGBhmu4sVZXlUKMW0GKYiURMpyzTWLwY050UNXNUOPOiodHGZ3EENveEicdme
ocPkEqDU1OtrK8EYybYRZ6DwS3poNxaaaRpepxth9pUHZDLdTy8tsUiJy68OpvSd/pCanK3tbBS2
ctobgJB04b0hGBV1lpppOTj7zZNOwWP+8du/yGu1aoTY0NzS/RX9It2Q5q43ABxk0y5yT7AsbQr7
3oW+3y3e+AkwMgD94equ2VgyvrNhtLaIBKp8gST4+nCMf/JgFCBfe0UpoOPqS4rM7VJzfsWVEl1A
xpG30cs07SzwuAk0ckwY2ZGlPFfWkCYZk6w8Q7xI7b9pqs9PO727ev/diBAqScXtBz/3UYHMA+el
2e8yoKgRCqhJIL4Mnke7YlEdJsX4r0wywA3+/Xacw6Rsg9WR0Jff4pl1p+sxSnyjwKtyx8TrJocT
e83gYxw4FRt9WiwKELZim5qFcCMXGxQnd7v0eXIjBKlzl0KupufXeREEoKX+78DsMPu8x4lmmgoY
Gh968iOhYqNOSiPNMvXgAiXmTrQvQHWjvxCzI7chMoJhnb08SrMfHUPPT3zGf/g4JVGjTkqAoGJq
jDr3q1bJIip3/gTdofy7Xohbs9DmdeU2VsjpHZTdgb4ZiTFNQPmqP6e3aMwA7Q1U7VWNLGI+w4yn
5gZ+2thvP0rftFI7GlMRUXJP/41rYJcUD0WHS3ujv00uyyWxzJKvMnTUfWaUJo5Kg6rAIi4Nu1Bx
slRPpzrgLdjX30kYktNYbVJupbNMukGzN46Hr4QFIy3hVRi7EFqLQjDLyzA2FZNb1zGzCRQrFk7U
PZMu+/X1gcpQP8fwzn6Fmr1UzPWHMxAIDesveMKcz4lrAcWE89ROjRCTdhhq2441A7xz6CRHeM5v
e5ZqKTEqqNGg3E1yCS0koOIflJhoLAoznrFx4/LhK2XmQNX01ooC7TLwkHFyVKflVbe6KGchD9oR
h+9ha+sDnFS8unztMwGQAGaAdB9hFZNJiHEhnYv97P3spcRJK8jazqO0Z+aRsrGPbkUnTyVfoEEO
voa5tilRuH0fzKHNB0lWLVsVtVjxYg/ZIc6Wv4y2nC6Ss0NgPDQKZVfSz5q8i61TLin8GYvpknUq
wdTyp2PzBwOIQEncaEXl9c21Zv5s5GoMs0mz8wtJ8JtXZfitQz2uZWI9FXbR39SdIGuf/b7jaZ97
k9T8KQ/737ld7e+6s8g6O26GZFTzw6L/6QCx1+VGYxoe9jH1xt1qt6PMUp+nkNSFhwv59gvx9ofh
wDG5vMovRyfbxYgc453tU6fxo8UsiHxMuEbreylO+qAO+CM/qRjid5tSez8uaEqDXU7yE7JIBEG7
cr525wm/mY+u9Pk4vO1vBZjfa3yJ7KS4FiSnu14t3p29M7MvbCxIxfX4gNB+xjj06gT+T3s4NZsT
2DHWFy1gIyVQsKLNep9WDkpNWQmnt2B5iStqohx8lv7VksXQ85fNAvsQOcGpJucGPshIetc5AhKA
w5r9vXZtE9+P3WzBp8cYMTfsyEn8IAAYMFEA+gQW+BV7iwWIHei8JOij3RRNu046Dpho3YmKWLV+
XQuSza8an2bDCCbsIgx5ofbuNd6C/iCgw5nRXY0htZZV09VCT9PEscNeonBBS/OkkQjXtZ1hbh/d
B02ugAv713DcgFUfRva85KUne5d2u4qFMHjyQ2tQmKpJDFy0o2qP8k+M8LFRAMMuf+Ke/oj/fE5W
AEF42nlETpuZKxi5saC+a9XF5hzRpNO0on3vooH3IVLkDxK1edZjvkN3v8ZwOf7O4iHeJ//6Miv0
STVYrAbrhXH+ksJwavR9LfedZpmd4JWh0AMDgnZor3GWpcjpshRi6jCvkTpfH9osvu4pwGfBF4P/
/Mc9cirxeTT6O+W91JHtPBemBWSG37oOLmhpVzHDUrEzAgmFFgSbpz4mqlx0Jf2H7l4iENMKp/Al
0nwom6V9kdmjX6XPlEFnZOC/qyIJUrHOALT253hsS+tK2tu4nxySf6GWQENVcMs3/asXRzN1gKxd
Co3raxPYb3v61M6lCbhsQum4K3VRevehEdoZu/SYdqxOKzwKgDC/77bv3jGJ6PrtjldbHYmlubGs
e9B3up6Ir6xUwFX8PmNxaVO7lSt7LtUp3vomCLd2BF0Dh6BDhkCC3ivotGCr8IhofQ4gpLR3v9iK
LLtUbrrTmWEe06DT0p/FQPrkALnWjhItfzi4AslWBVugFEkxm23SpOk+un8XHAgSlCvW0u4JCDqg
/xOnJVxnsIw1eO7ffxu5NvWAZxT4xWlj3lb49kjN4t87X6y7/wk8JDPz4CpgQtlvrkPWkhkeA7xt
60tL2l6Tt2fbINxJLiL6iujuPh226xu6wdcX/qx2T778X8T/cjoFWI0R4TwRNR3QhUOvXGgT7dfW
cyKCxoF549ZvB+E0rJYfhESa8meq2Ve1WAZPdXTQjOGYyaeVNQpvJGd/uDmPNMvyiNpV+5PtTzxU
bISR6c9bTSu7fSWImeAyNOp5SIpVvcvGBR0LK3k+RSlpuFFO9IoiYvLx2LB0xxbXJypKsNFiHCgp
GZaqs03/0HbqiU5ss/f7H7w7O8/v1qSsmjUEqGPZsuO7KuEZRSxuIdgbC3wF6xtOFHrfcouw3L+N
dx4u1cUs9QIrx29jG+4VUdhBSDvIWsLRdksIz+zLg6oU8orfWdMViNZOkDuf5uhTcYepLOV5PwIi
JSvlTgNWqToTFsJCQ0PvEQW9Q7cO2RboQT6qLR3SiUiMBA3d+aPTOHo0Jjx33qEwXIdFwaC41vUY
o3IauIx2ypiu/cpb7ri8z06/pnjHTlXoO6ZxQD56kHQxCNCj2brfvN5zcVKNK8Kol2cENI5fsOB1
FXOoDy9i1rszCZekDYCCaw+7ockjvXQ+W4v5Jpvps1uiNOzE/OKxSKL3F2DBsNWuZUlut2AlVrgP
yEKq83j/HwPkMUEVqIam2YKkMHuOTpMZ2G4vqtsJpGJQ6wFs+0PAshBVN4bkMynP/9L/3SP1FQHv
IM47WWOVehOClKacJ16axpl+G0jsb4c6VZLZffMyA9pUQv7gy7a7VU0aqiD5Er515TMjhXBWcDgd
xMFNor6f8lWbGilq+ggOQTI9iKudJsr1Z45I+Sb9+HsM4C0KUp/YWFbVWj2KBMusKYXwizKRa0r0
7f0WefUjVRNlCpeydixhtkbSVEQxUCIqfpKJWvin8BQwNiFGOwXcHM36KsiRbzrFUEErS/EAwV5g
nkIgzCNxvXTqTsB3+bUKVH0rYlc2JOcRlO9uSv86uIN+gNDygEEc6T03Jp7vsUZ4HKmeIV1ChUhj
VNpV/M8cP9Xv0FdCq+QZR5wk4BHeXXqBOmc8JxmnhGldUjJHi+9pzTH2EPKt3DqbaPOu29xFGOpS
BHBaGDQM6bvIb1M83IugxPpgQCOmdU28ztt80xyErTaKYYNL0E3RqEPdnKz/Orh3qrIXYiUjqJbH
PmQmm2fu5F90G4Vlul3RjdiNnV4dNGxOAsHRNhOxioWMDBgAZTob+CfH052BrmlAZtBI7nsAMEHc
BE1aX9G0J8O9YfV9QOqkZwyr7wt8meN4O2QsqL0tc6NZgKu/LCKAaFPIQSXV9OU2eXXQ5WYVPmrB
WVDNdFeTB6QsOFUTrIYvNYpWEBJTAUxJbjNDmcIaobA7+ZEMTVtZnEn/0NCu8bcR2zW++7EVngwC
I/QZBAoffL6SAfVfByF9vnfCyFpMz2sq/Wo1hhrJ0MgHbhUJMzE7817RpjKdjlRUEgJ8foaucY+E
5dMQAnX7POmFxuAWo9TO/hnduQwOn4DNK7rZDk1wWm2CSy26ty5NgvfFBOm4I6C4uCGVaHrGeJmQ
1Llj8Y+YXzJ5qJJ2shh9XskxlUSy+WEc3WnTaqxNOqmIIXMH0/A240a4lX3M05U+CemG1X1sE57n
Gf93wA4+QzQVEcQM7TETEm2YYI0eLlvDgCbIUdggqBVXv5WWIc9OOCSn3wKrvfILOW+OqQPrvhAs
19xk9wEGLASugfjFDbL/4jXHBDIvwVcVtJuJaTHnGzvIFC4aofOIzXS44oFrCqNQEh4yf5jqks9i
K92D9eXIz2tbVthw9YaH50NGiP725LRCFliZRnNqJO1AyEsLQrTzHl5iC8vPIEy/vbOUsAPbmc2x
BwV9Rlnt5gBQLoFk5GQTFsvB0nPgi3WJy4p/MjBzptQoILewrlfknPQqg/FxR0MABQW0TUfBqvwV
kJxYSlCDymCnOeMgYd39/3qf1rBs9rcJoixt9fg/e4m42JP9nvZSrRggR3aL1eUehcCK5f+QT916
L6qeYz6p5ial9EAbDF30atsxf+hF6OkSEncanaK/7YfGLPqOXF2z6gG4MBLOAwbl4QYl+Pr1iLay
YV9um+KY1OR3mz3xjK/g7S4HiNwu6tkqjoN4mq2xvgLSG+XWJsthe7R+WtBby8dBd1oIxZTsYN0s
XaQ3j3Llx4zWnLEfHMCVrQMHq05nPw1DxMSr2wdR8YOyxTYTUsGOZp/om1VGGDwjgSyNHAFltiUr
nwKnoV/mZ5TGGn0AwJAmfDrB9HAA64NSjBeWVgbY9zloOLMUWQqIp5DDJkhiAwFglmwL+41rv4Lq
ZBza+wYiYLIW/1LOUry6EQyQVljrr+96VMJ2ZY3XsfxzI5YvuI4igCC4gd6bCMf8gkMQm4OCowZp
fpT1iQIsi9Rk0M+gCWc30neRf170N/D4psjfVenSeO4x5TEjJxHkibd6zUBl3qflxnQTW2I/1EjP
5uO62JVBM82gSpckNIiC/aDR6rHc+mb65dWQrXkdRN+Io+V2WiFSEK4edOa95ukzYSIuTquOlWKx
87DL8GSvNP4JjPhCs+RbkbfpyGVfPIXT6DRLPu/9ErbsMCLv8qnOcclRPIhEmU5L1PUZYEHx/tGD
xHBUqa++YvoSnlmweZKZRaIK8b8zBJUsOS2KPYYEuyEUV85NeUiMG5PkvuJrNX2BFVlLOE3LugBs
ewuy13+9ZjBGrH5ZRJVV2QEBGmm+B9FN4eIfr4S9BaRFs4j3mAEsk6nJZL+ZDYOseBKlHTqnkxli
pUAF8r77qHNnD3+44u4TgubR+oWfvSAQQLNyk7oYDiaNReRuWEky9Em8d3G/EL04lqME+S+5JXeu
3yZJXgvz0Z8d4ElliGRQ06zS0C1jaPVgSgs3c1an47Fq4jzQ2kLpd/Z+EaBpe5m4ZMXYWkSzbz3j
Su3ylPaZiPivPo/L45FuyGtzN6vf5tMh+W3o743CtKBdpK5b2lBmtYADQsNDuqi329jNOXRoNTJ7
+wjamz5EFcPRodlg+XKw7/fODB18GPMGGs6OrstWzu7NufIm1Wz0J/yt5RUqio89bT3IgkbfzjQR
8+e+hBPQFxDKzcHoHGjsfZbMxvNXFL8WkQyGk0Y9I4ph7oNG1q16jj1IqnHgQfpTFLmZ18Ctvm8Q
nQZjH90trfaRveu/tVvrtylMR6wKmQphqXxS0k5A6W7of2LwXiB8mxgmRh3olIbn0/Rd/l9N45je
GAFCxwy3kI6bXZ3i6rAApKZ9PqBVpHYNjF4QuGZyagw04R4tw6Sxn8aG+XC+grjzSIVGfLoyM50Z
K0aWzu5kYPomk8+V3ao+NDUdcNwvxmQ3zVREkifF8Z+DI65sZCVrNt+6RE50yvD19Xa1XNn/A356
hLpH/HsgEnzUyhNjmpePG6C0+f4yVFSrPbkUhq6dZL2OxweSqgBrlm1SR2qmdDIB/yAACUP042Ok
tKAwWJbDmIH8kqWNiLMMnNPhZv51dXwTwXyPotVejGkZQg0TMrsgReX2mcyaFXH5Dhh74Kz+cb96
e/f3XeflnV+JFvgtedFv/Jttis3c/0py695ALLIcYxWAfWiNL5D0VuxJ6fIg42GWpH833eXblSO3
xMnj2vk0lmMkDUPTZ1A3ok/eZoz1ddK5KSQ4fWp6peR4c16mjwzenPoxpyPj3ieCZ5H9M3wa5mVC
FN4xRdVJX4nJrr+yY3Lnd5xNqDYn0pyT/k76CfKtBijxrnh5/LiACF9nl+3zSPnAD9+hduOpH+Xo
p80Agrmqe7cbXPNyms+nobrgzKddt906QbjiqhMMvSZGuL2L5qP7i+IiROtMYoXS83H5jN+sZSih
L8DNuv7r10YQSjcu5Hf2ObW/3kvi8l5mWM7tIfAiocoGXAL0GK+5L7OEEva6KUYnLbDB2rNbH2WO
NwcT0IZK39dRlygirgonNxHIt8XYirIgCTfQI7DF1f3GM0UP33tyWKmr3vll01yUf+aTF0qbvl47
td/xUu3hpRmk1od6H27WpqW7jYNRfVzDKd+dM6nu9gUdMzlo/gCK3zkTuwRlfVl+j9ZOcSZoFtxp
R+PUn0bc8e2+yNZjILMAExG1z/mKHZ/gWB0QefjNng4TnVMvXZlYhtVZGLLiZmvNPKYScO1E1hSs
39gzpQrNZvepWWe/QYQy3/EuETc6JB4pVOnqBe6P6Jpz0agUgkGYisSRukgnVKgB4NhSGKs1Yrwm
vniNX4X2V8neVqpxt7c5jlbz+OF9D+cgLfJSaBa6lKd8nDKqWkL1aS9KGvg6ymKFOmdM2bBfTPQX
Xq0rO37iqyGYcObC4umftAT/7MylfU46cZcRrumG7tGL2u5hixOAjP7WJ8NG98uleDkBHiQxFE6E
q9jCvj0qmDMo3Ta9nxdv5yjSBKaEiJevaWYMPB5iy7cxULbWet44y3hlYw4RpyEmV1cQ+zsYSsvK
Jyq4QtvwjrudMEDJ/1nEIara39TGSpgTjAk10cG84HBnCLTSWbF5tQXolf5qKQfZQIhZAPEqyXmo
IbrMvx71jaczJ2e57zq/H0iSyugM4xnOqlrMGr3FhHucvC8n/pSTLFHd5A0exqCu3/vkE9fNtZgm
EAEaeqS49qcshocYdjcFEBvvoUYJZLjI7puYHMhD3Br+7tnYhKMDtGlOfQ93UPx2YAq8QUKINqUD
CvB5AyI4HU0mtZsXyTZCHhT+s/I3luubHZHpIF5GKVq+uOMONJoshb05FhI6HJbEYkARxfw8KNsl
VRHLP21Us8UeXlztN8x6fLYGS6WX4BW4IWJGzcA0VmvNFx31qspLna1bq2vstSdHXoBTCDwmUR2B
+meDJbKeQfyH744GUP1uGUdGuUwUPdEOuU+aFwlRL4fWVqYELt82/f/Fhgctz+wJk8q/29tFds5L
TbT7ZPNBmzpEgcPz9W/1b8hEe/H9NuPBz++a2LAV/7KS9L6tSDgKyGVz6XfpzDDt3eIAhEsmhZVA
PaimQfLCi2xxnVVGloyePJyURItuVApDweZvmFT5AZB8Txn7GPLAK565vQAKLCmAdgqZ4iEYx/i8
98rV7MkmBEe/9a272aBZdH8hMi3vzqE+M8FDL4zJw/dov31uhSsWUJCddbMc0D4sQtJvSdV+jvaV
wNC/eYkp242QH/OlOi/yF4lOo/O9Gj2q3aRDWc1/+5ZwkKT/DTSreeaiUBN8ylf4IaO14mZzIvlP
gpUUhS+GTRO+ttXYIfEtzPjMuGsVreCEAxo1lGxY4REVsZKOkcVcotRsIlTnnCFt77iwwK7u9Lgw
Y/ANymgBPtq8euUjyp2OYn6WON5Y8LCMGj7ICoE8qlWVRLXJkEEDQkh4hnP8LxPLSBXz4fCSciUx
D1BFqGxD0kimikD2KDdK1I8iDdISzAdirb3kdWB8DpbOX8/StIBPKBGdAYVJ8Fvp7KaFCBbp76ow
q2lvqC8Zk79Ya46BuVv8rVcSOrc5SlhEBc4Zc86Bc/7T1BpEHMTUq8VmS+uJ9FJrE3SQhbFrdLDC
UWm48PS41Sdce4Wfnar+gozUtCkJrjN8U2ZOHcsRanlnTtJTF7KIfefvxQGfdKZ+vHkj+0eC232e
jyhaLlkEsXUSJXqard4K6SY9uAs2T+bYpSH4qxsHy5k1rKJhd/CqClGSgIPYmDyRODTT7esva76O
diHuLE69AyvUrG3sJvPQ5nZX8IzKh78ytcumzm3g29jN0GwGD/wMcKjWttSedAHhDIfjahMrH9P/
sn5R0Utcwtct/9XT60qjE2EEM2YrEZowL/2O33FblnWV/zpRbNKEPgsQIEqhg9tyFnCOImYFtoTX
F6haJnBiFHjUaRE+uidzHemzm4JQaXDD2Tp9uNicbqylqCoSv+9uKL21+tJZION0RD05IH4vGNfI
sA05gm19x9EhJ95uw87XVw4oQuqgYBYEzdZ8HZoi7ofKwrAm9ugVKkqSvrqDf9Cbke6MNd3yGA01
NEPddDUfNU3vO238flAi6QGEH5A6W2zvl/VUYHBOOhVfpjhJ5JvT0crG1LYqqfTluXgjomv2oL4d
Hv8NhWI42eU5jupLLVY9s26gobL6m3SBaYD16EYDf8hev+xrplqUo1wz6gclayDW6CUrzwLFni46
HCyLhqW+VYV0zfujN/eOAc0A3zmpa0KRyUWbS0l56B5cQNbDFo97RIWXGD4o3TVgLphZeAcotbeV
RyzLwXmnqUaKn4iWUrkSo4iq6WFDu9Fh5erlEQNhP5qxILqgqWSPXRb/WjTs/8G9/A2lUjWqfdq7
yAPT40iyh9tGQ96bCPHpw9Mx0qo8Va8qIlM7dqxy8d5zqdtdoSIloO6HHZVUVCrnI8+a/uUmZM/w
AfiNyt0Au25ltZ82lfYAUk+jOvz00LH/PPzyFb1jvm9xJ5T0vt3uYDgHvOKu21EVgo1YQuIU6Czc
cUGov8BweSZrWtzRgsWrCUnkONZN6w3y7g9xiRD7zF8/DlB0tcrV+Qm7WdlS9cEivrru5+MDBOHD
OmzlhAX35D5dvGUXG8eGyZUg79PmHiCHuFyI1kjzHq61LSkqaxd3LUJZOAphuiok7YCWgk4YUmbl
3ak/qx2jFxScvKs3iNiOQ4UbXhq8nwLfh6eVLVZ+J32hOSVL0nqbnT76sjfPTi7KEeUllJWtYpC2
KXESQ5bdJhECS9yTDfH0dJl3sGlntDdSQaRHgHBnok6/brZTCryL8YNDlYBNivOLpU2Xu1eJ1bl3
+0HF6D/C8kHwSq9IeVNPxLsJTi/T5lNoxgpBJD4Tlhc8ZyjvhjmCN8M2jlo5YIZ5+Ncgdq640zPA
qkbs2aX4VDdkrhTi6BHjfKEfYtXiHJ5knBDkEyqCb8t2zPcPGIszusYFbf2FVxtxME6VeSuJpNIq
lfmAf7fL8WK4eKvnweBqhEiHmbVpfyathcNKL7Bo1z51C5wOwmgvZK9n+xBSfSJuFKsePMQSbmHR
7u+HwqrG+dU9659yPO62UC5RrCscYZXFqelnTANYaTyHvuSkC4ar5dssn4OqdmOPK+6CTVIWqy7Y
/KPq+Ko5aw/Jluf714GPS6SNqdLaK0X+FDksTUwa5z1Iwc/+zQpG6CO8F48UX3Fg8TtZNaBRYyUT
bgJRCRxHQcaqkl4D68Sf+joHeQzranxnXQ3QmytIDVonFzXI2Y81hXZj04nY7HSMO/NxvL6NOttX
cA1/TpGWlhcNnmcPUd6cYqNTJzUpzp7eFxJRflxZJbucRaj8r0LAQLYma5wtR3RqXPBPCdBom9v4
2xmHHC1txwZEcDsxa9OghjGeGb1UhNMUWp4pQU/x2BmLL8qwimqVrpJSSQMeSijJ5yUS2JFHwG+I
jFWgbQNd71tG+v8ALfkToLqgp3xWn2JPPJj7bigJAHmIS5fpr8sC7ncgUXaB0fYDoZu40OJqb06Y
ucaWw01SMKGargD6geVmm71ONDhWBT0/zKBNUaqEaaXD3wSatx5/7LbgpOABshtKIKsXAOrPBXXC
2cBQS4M8xk2aNMHA4Z4Ts1RMvVkpkViEnNYrhEnkjbZy9SV4S529fGvD1xKw0lSrtMDhYr1sd7wa
e2UDS5jEQgtYqwDH5hT+8h6h/MsWGhPUSMQoAiTk2b9lXXlBJa5n5jFzchY6bJHSQfyqgzlFyka5
GYDuYoW7NSW7v7Hni8swXQzIGeKhcaT26GTPYtdQ3LQp/deoBBb+vi11FBzUFqcdhY4n+5p6FNpQ
df7Mz20mcJ6zfun54/itCL7ZWlESCMe4LH0T4wp9CLnCoCSml8ny0NvAPIcBkvFZ5P+QKjESubL0
6cBcRLU7HJGcmUM2/KEU3HFeMpG7kfsdDGE5VoSeNqjbtA6i+ntHLUcXQTu9ZN415rAXNQigyXj/
2+BFvTBQi56Dkb07oopCach2DEACYAO6PM0rhcArgRps+QOKkDFNTFGpwkF40EbHEVdObB/ggfoY
uJKg1vEO8Ra34U5kmum1XPwkr5UGx+0gfVNN/NJG1Ua3nB1PJ1i03ElLDDQN4D6/lKkAXlICEdGm
IqmYwGpX4Ct1v/xV5tWH8wQIA2ml27gV/Kk/airzCzkhRUfL8NHt/o+Sj7zHsLSt683QR7Re3Q6L
ayKQirvgq77sxGmg57TJdqFR29CzBn3b4l4uIH2mHwUSpjzHCdPzJqLLFQyHl82tkyTw1zgM8Ouh
m5M6Ju1uSFabnQWrdEw4ERjK/UQFitliU22E8m0rMjsWwtOwW5tdbUjW9vpY51lWT8oiVCdajwkN
ID/ivFZaHaUuhxLU1YTdyceAHjGzGJc5ceY9ANzzoHcJ1TBZ6AauLZVlDFQjq4GhC0VuA2D0aZar
IFzetT1uQXyIrGfC7opyKlZj4YI77+4HFNaMmnTBVH2q8uTTAeJ8nPJGqCwEtQHMTjLGtH+MNc6f
dD412c/xVhJHhgJIYC9W3fN9qW4cZFyQeS10uyubg5TXEcGZ164am4cKTS6XOZPmWtZbHwxZy7FX
DjzH/W5ArjyCZd2xf/gNp6SJXeTdU/IL25U/g13XZ7vesjyZUnNtEH+mDDCwN/4YfSpQwGZh7ykA
cLP7DC789CbRLS/Cx491kKs8SzDxhOAF+Dgm/O2i29mogEhE5bnmwCv8WTEiA93M0ITGcl2UOgYi
+Mij65CdIhz5QUSAZclFzyWlbqVfY4HX4OCYxqk0yBRhU+a/sdVKFJf7Hrv6UHF77eHeLrAY051m
voTZ9UnU0FG14DUHDEA+OAy2XlY2JO1L4kbW7mSRqOtO9mn1uAQSYlNku8wKbhqyePanO12Rd+G9
LglsFfXk63RDkowz1P67yikDdSswgl9XvmSWCd0hzcmF9x6QtMZ1+BY4GrHfWSMUTQZcAX0wZu/n
ebdg9KFPW2ziyffuediW0fovs8reTMkMLFslp7R3IJVmktvIl7DnpYG7fJDjxAUx9KYSSmTvhyZq
FEIsiYNJ9RUJEjdpDHm8HON5GoG2shmPuj/Mp41MaQ3agmT7s4k0kpzmjQjww0cy7t8Dnrp/eG4K
BPJmULP/ziC138XGZPjy+uDJ7KQ/1vchGmLVlY8jYZAYxSr9rvB7gkWW2IfR3LiJ5mgZwBp0T+34
cUJuzyT5teWL2GIO0HPFzb25LZ52dqMVIcVdtsP4eTivFI5q4Smx1/SP/TGiGCU6p+aw1zt0Vbmh
GFVfdjokl39m+RQtjcpWsydlQBNF/cPoHwlyrA/M9TpNPagLx9t+pHykX7r/GHj/uy3bvLL6kF0Z
8spnXu51ht+XcuyUy5nwAV3jRtBMbZje5Q6anx+koI6E70bBPRpSj4ioi73JtYlQK82jZqen9nPt
FkkSOhHG5IthGYuLQ5AWO0PBZ/NO0onRfDS66vjfFvOTBTUo+plLZHVxcL+qVNe51I1xexDSlvqU
yVVgaVfLqtjM9BZYk6arTVwhT78prt/OAyZcieAmnEY0pj0+7C7Gb8gyY9JOLQE/1/h5bF/oR0Ak
cKrqycssu8McX1sSDjulCJeThQV7yBsDAJMfybJdetSqVS2mAV1992C4t5izp856goGDFXZkwLGc
R4HIaD58urqnl3f6IzjEnU6TsL6NxFqzA3/gWfKHOE63BowFxmzmfWU9R/gc7zrg6JNAyimX6d8N
3gdNMIWb7Oe08kp4WG55aY2weF/uFWm3x60G+C/qp1yZKg3W8UlhlMW/fxP8uBmIE14IZS6lS/CN
BnyHjwjf4VWfHr1WM+pHWAayBLJisrPFUuAfWEd/eG4ighcY6qYYSRVTYQKsS9hr825kJpxksyqr
j3p+OQFjfnsl6uPX5EU41P7KbjcSbBY/dsDl8PK7QbVD2ZhG/SqG2VmVAj/4CH9vJ+ngMDN6fkZ8
HjoAWs7OAUxboVy8D+O2CnIL43jhL3TyWTgsfjfbqACl0okyZscrdjDITm+47K4DeDaAcAUd+238
PNSYRCztADuI/gowqK5kGJ8ZaQp0UNKl5o0PfaLs5NZiCX5TZUAfSX/m4INSwIwiIeolpxoUE+4R
O4hLWRJHekBa6xKIErUpZH/hqWRKqUL7rdNcNo9GkjiYjMUqtSoQ2c878mm+g0q27okpfKkLsn8a
8zyOP1Fkrvfe/pZfP6QtGq2GuySqrTFdmodlJQi0fmcop66GS2usBp18knaP54gDREF2e4Id4i6x
XTknRAMFw/dpIzkyP2746xoIZeJB3zZehBrIQHmInr1wR/9qezhGbC2WaetM2wy0qVw8EFkTs+AP
G2bINns7WZmmtqR5Nppq8OKxai9j1WmKnAPWBfnv7Cqu9ZhzE9111dzcVyQscxr+/W57OMKsQs4m
SAS5OgYmHTBkEZCcBxg2vJng3ZKR63OyJQFjWFDYPc72ke/KzqB9MmsGQj6B83jjpNXM+8chcVaF
3quv/doq+BM+OhEMGSzRai7q3hMhadw36ixyz/NwJ47U4+bbGUgnACrbnaQjM0WLUN9A19OXjiMe
A6RimIKCo1gDVmGkJqGPHYR1P6s2KbVML68MXrRZBnw5crBSU+57TPiIJyciqsiGl5Iv94J2D4jt
cy5qfrn6zqvfezPz7q6P2uMggl0n2H5L9YiUVAelqkIRmF8Ic0IR48iP7UUjgLnXIjlfP9h644lf
Y+0Xjq9UVAzNk75YmSsAH7R/OZBRiemd+PVeMrx+dsFvcqu2BqV8RDn7T1lnb7to02VeQ3gODS/Y
jnZi3xeaguQqNA4LiMlpUKA2gL+0ibHPAcC79loTc7mrIEE8FWtmznPAnEbjAnL16dvz7REsOhf6
0ch3/tj/WEN2kDySDyUTVgG7ot0rueQPbZ43pPFDSbT6pWaM/O4zUS/SAA3E3FpAHqGUUyHwluGA
we3E/kIjioZEa0bkmIv3Id3piv96ytVa1jPsHoaZeBSqo47kx6oCcKCPdJSaNIzHQxhJTV2Yr/qM
qSl5MX8EBEZR+0pQiz/QcBScA004SrfIcr5rsbt3xcyj34bf4mRDWZc65S+UNo4SxnN7QazNqIbs
nGSOqnf8L9AZ+seGp2usxYtNOIAZITUl6gfzOh6H1aR4bPLflo/gieBoXbXPeWzAbd6LQiaLFweV
KOWMxnW1MzFvi8V1eNt9QR0esEH3SumanjdOnVCe6KtXbS2RctLWXizMGtH2EKPJKJ0PmU+ZKHsP
UgioKiTdIvvRU9WA9iQpFyQiS7xGUXjm8XXZiDUorIcwCii8kVMh77PCoCMUVWLAoMij5VPadLBT
LbA9BYQPdXMWyXYsSesR6G04ipBEryxqE2JCuPVegm75kLJBkXNqhl2rRrHgWObq2fMRK6/kWzQK
vg5aggTpCJvxj0OJdyVGcHYFNwoKHUlLCZ2bejvwypqTihL89p8jQyOwO3aB/Ll7Zr37/aDDLDBu
tyUm9Alk0iPUNoMvZ3GaEc3hIYJU/3JS72Fjmw7qfgjIzGVBuCdzRFm9XH4K0++Ki2bpYPkHVp7b
oWHQONCxtA6eBjaNKV/km6dOxcn8gve2GyDSXNmPsEdLTd/SpjFeU3WLU6JLEiZfC9RH7m0DQ+Ln
TT0Etq8vysD5ERs47f0mFkOKFFXWjIRhYD0jAziCMEbCuzOvTPv4nWYb9UmuFOioOzjiKYxJOsGv
NUHZzyO3CSV5yvgq0pBmIh3D6HUnRwV43bJbxXOLZ94SOcss+zA93MsgZcCUaIuzR0FAlTljfXWO
3OBz32gbjGuV5xX2ncPCjfQ0UYd3vltOOr/8SMyPp3tNOPHIbcSR9VymfiDjicynq3lQGd+jR8we
Y9+J57FEaq0no5wXpSAhVpxI/+tCHPwreJdkpgoo/Iqy6Ke28gEQbmPliDF/KNfxrxy4PBw03sIx
Oy/vkJ2HAZWDz3g7eH8FyRlwIqaNEfCDMWY90hZJBQC4nxK/+hvqRfQtrKdkxzOdeRpzles8NCdS
+wAakS6JdYFwrTP8vGSESVq/MM3NTzVxa2F1FB8ALAJ+Iksrv0kCWHWbP4FzcRChlRDoxKH2t5Gj
duAUtbCZy05q8xn7zLfobGfVOTki9zPDWOjFCBy3wtb90RrlPDTPWBGYAU3v6pS6eJdCkNj4TSZn
eIJyUCiiGBw/p63nH+WqTkFF7rbze1dn1wXInjoOyzVGfKxRhJiYEnU4jEluZGikhDT9/YMcNJCi
uN4ufgxvjlJdMqaZuc2z0T/opbkJ4JCRmuTuD5fUiG8AN/DtcHzCvjEqBLM9vocFS/+mUAizgxxY
XjM1RYNpfzA57a+YRN4wA/ZTS7ViK+KiPxsNid869nd923xiFSPUbIR6+nwZsIHcHjU43NgnXVOv
ihT3H/he315tw1Hn9MA36qpzRvnDDkVqCsxByjPP12KbKgLs9HVq2J2qlnuQ6LlR1QMEecNga7jb
CH4tS2l8LHPNxxvJalf4XACrYCNEYBOSE6UnEVp4Qwp4Xa7gTIxGS/Any1ukjtDF97uOlFZl+/wN
D+0gPi1Kh6qb+PPX++q3HhdXifUPm68wW32HqZugADOKbNr1W9vmhvqIXJWqH2Hg0Py7BXhlE/1D
p4ztaG6ebtGkDTX585vijefwfci5cQM8eRcAz4D9gbh0A49CyKCKNXlH1DE41BzesxrQVYAUxSfd
8rPMvnXUzraoEoj6tViFOuYaTYwO/ZnA23XGnDOOpNLI7wrq+H/eh9OT85aC8pmeFm9W7PAukPv+
X17NttuMSMsKk7fiYJMIgRP4rNHFXD08c9C0IpwpDur/VJUBJ3MewmDqJGLMiklOq73AwXwsCep+
7WODMW0b7glTIdNccLOfHUBXhHNB5I+iozk4RVyC9A6QP/0/ye6TH/4XGK62wT3o/cTUMAeLGTj/
ZJ9GAKMv41Yq0VW98X+4SlSMv77aLmcDIpjcHV1fiS8CyDriLALe5N/7aOPRhzd5TKA2WjmX9fTQ
IBLQSIYMYt+9rVim3lwpakBkJbOJU4XOVTBjpUsq/UnoGEgyaj6inPbQA3oQK19kN9CYjZ1lJGi9
ye78EJNX2/JqenWY2LUUeQTREB81rlxv4iuJxH0jUdnTbx/iFjctJbeoZ7SD1NgeTgQUQdMdS+TC
vR7YRP4TN/eMgibiYRcvVZ6hC7sgBmZN4qQI5aZIsUg/Pk19BgVxxX270HN3YDbQ1RZAbtg5TXDa
HHTriXhQPJEuiv5es9gTxO/OigfbqJyJMUmDNjfw95Ip9kM3G2EmVZ1ZFX1S7ad5m9ofSrw1TINL
B8nc50CV/VP7F7DzwpOB6ZHqlD7465ElzCN3EjNcu9hgeutw4BsZTTB/Ytb9CufJvklgNIbp7knC
NwTGQaq2DcI8PA61QgoSbjJT1r5YWbU8E3pTz6HUekcvT/9zVX08VoOm4N4VOeO9NmDMcHQXY6mb
uvUXKkJYp+dFG6uR7mwUi2g1uA3C5wwtjW9ZUhiKDwrJjvdVlA8sRfP3ISUdO6pZmsJVjgVj1oeD
UalTOuJdVLQ+Yk9gkwZglLWANujWtiVDL+ZP/CahhDeKjxlH8SAUicqwli4g1hF7kVF7wTWrFwsr
YBnoIWqUBpPNNMmK2az5W2vCurXG/VxRmQiyHe1wOL5095z0jfgeXQXnWCtt4Y1VEc67UcvOs6Cv
w8IWk8hdPjIdaj83uSrzneabc5Eu3P3ZVacBnLbO1dD7qXtbW1LMiz+KAPQ51xrwtC66lA+ix7nD
b3BNRhjQ4OAn6wepyZTrDe0pClaoPevqn++77RvZ27JCZ274v2jGo5DRebI//jR0G+K2qS5AMWiL
6ntW6c0hXewO1DzCMY91lCc/SvAMt2ERg13lVl8b0otNeAwVcyzjZNaYuvQmbpJL/jiG3+84D/Q9
2GZ1GexNCbN6Lg7n/Z0ro7zPcPGuDfFwov4xMZp0sFPynxbwIEiwV0fVYScK+vcwrxhZFV3qWI7F
VVoZm0Qr13eFOvuhOcyHuq4n1KVYQy0YiUpinGRDvOh+sCJlT1xtXVrf6XRBE0tJUClqBRIlr17R
TQl3Uqtgt6+463rp2cTWjgWiHRhf9QKBf2hUldlTQ5YPgsrgSbgqB93hDwE7065Ght1BxCuMXeSa
xhS4rFJLGvv2K+fujkQOjTmFWboIZTOQO0RCnacciuTa6VdQZvuenK9ICTRhrxabzPyLoVsx0I3J
MOr1L4eHLp0un1MgayhUo1c0HkB7wgJjdqgKP2W/QFJmp0PI9KFffiTVfZhWreGRgcqA7C51XVJS
B0+Pqz0xbzTDWvnZ1RvmhPHIk/WcScr1vpCpIiAFn0Nj++2L0dYTFD0Jsaj9jPgAPG6jlQ85yWXr
U6AYkzA2ZIL+NYfoqFrKD2yRueu2A+o3m1IdO4mt5FpMvj0s52qa4uB0wSfGFDe+CWph/aYAMp4P
NrA35lF8ne+j2ggV6iaMw/eG0qprdePOjzjlw4tnEofVSI7mrtf+gjgB4XuLMzGFy2ZnjAB7l9Hw
Mpmmxj4+vWMUXPvCNfc5S5R23pJwDWF5nGDan8irTr4zYJ3FkrI9IXdVV8miUr8xr4cyq5GuTvTQ
9MMK8hSuLYS2911BrP1Q01YMTVZaKZQBnjf5shQh5rF6JiuiYZ9H8sLGqAktziTnhcb9JEQlsr7f
uH0sLLqQbBTbAk5Iv2uu4dnRzcmiwJqCktC1qQhQkaLpLCjgA00/3bKG40BhfM+X1caQkKLjWEVa
ZHdsg2qJWSH+7aiJ7sUQZaTwTUToHrYPr3fTWP+2Cvz8rcCNCDE3H6BSuMGCYcjRte1j28jac+T/
m7UJFjusiHPxG+qzIbvM/Y0zXf6lL6UA2QnysI4ESn1r5pI0dgfA4ChwLoimjpUMMkdQQ/iD7+tz
aAj/IQC3+g0m+iiPqRx3vPmTUM2U2lkZFpQ4ZMD5/JSwTkoHZTQ8r4DUvFQhol8K2wiape+NqPAC
+Yx5hkaINQd5eI9t9GPwDIa/xWCCDz475D/2m13Bon1wrgHlABXrcVwt84vIniBRvF9pTL7rIadH
uvHQHYPoHRx+PoJRbJoJYGzSYVQZ16F58QmtJC7WSXRqcYWAucAlYrYwv3SCxCdJYSNCPNDihFB/
okPHREndpOAWdh888E0HoXaumdR2p1mUggesubkRw3z0+TgaUbYXakt2dKTKBNnsADYCZftEw0ry
HbB0M0qgqZ4nSljHvwpb5VwHlcy2+TNkp/J1mF3XNP/rMCA5gaC3zNL30I6Lz3HB/A/ZVg2TRPWi
RCorabhTBmzt2UHX6W8KHUtz8tl47fRGZ5BQEZTNQXaNrVNJzVjtE1V0Fhh/2+sLNpyiGzDkN34c
NvkrvmPzgvhDiq0xbEt6eLpLyRlQ9UG1tI54SpJwIBhTj48x3KU6CR4EUPB0EQ3fOwWcm6MLOXYl
QYV0eFWIpOLbl4Rct2WwxkqEqS+MuNT2GY8A60hNvjDmK7weGAsIiOhdlZOoxRACgknR1nu6eoWc
0YgSRsL5/9oxixTyNH/SCchYegB8cTYMJ3fBUPFzekgBONlMaxt1dJeX6+oF2oTvZy2CchzYlOLs
rbFT3EP0O7z9C1JODIVgNBVBm2KCQcggEDPU8qFYltMkUinpl8SeK4/jZZOzkzJTPM5V866lfEK7
dms6iw98An70gpOaFoChhV4Nj+DdlJOHvr0t/xaHcplYFrlBCwIwpnZ09NXEYImokOu+eK3kSMZd
0wL0ik+tAeu/zUTW2ewZsdKyksfkYy15mmK9/dvY+CZUhsT8Y23Sk9ftrQJPCn4qcObvoIB/U2BD
vYE6FSleT1WSou7MfkeFVdqrSllbEI/Dpqa4TjEQdvuO79wNyk2f2snWF0tnrFR2uQgVVOz97Xw3
zIa+fIiBgzU6DdRk8EAseGnyFhKNxPFparPjPV64LRRzpM+UTR31zFUS1clq7WUFrPFJ3FDyHP6X
BylAsBMsENiLpQKnkjeH49rQnZLiW/8zaHS8wyyYYmwa02+Ll5IsV53pBpNSFYM4l8RauU/n/kll
HawjpckpYKtEq7PbdMAlMm7JwFttINd2gGttmcXcfgG7phCeL5N3B9K8L0fwpnV3flITU6u+aHp0
MH9GbceCtXOltOH9jGmf3R0mwPFBRFY6EaM7oL+eK7MNf0x1wnGfhoVhAUZIdfOgw1dH4uFKZbLj
3oq4qyBVZLWmBxV9fI3OhHI8x/1Gn5ZRCMIfRpRZnV+10S8AgwWh2bni7tBKyuW00GQLZ8iDNGFp
TqF3yE8gyuNV5uPiJ2gtHNKB8SclQvqrfmyWN6X4IADVm0Za6k/QCka2+nv4FcWADENVyhVyrAsj
l5KxgykCbme6c9YRU3YnklcJS8Rir6KtQvm/3WoMqsJ8Fl85aIyVVlzFAu0olF3B7DQxP0njmOQw
7zNPCdvkAtw97xcz+27q/Q4f6Ssra2RnaZAQnSWxrTIm4XcwAl96gw8tKdpvIPLEhfFAUNasuEeT
EP4cgWk7xgqF2bOAj06ltrPVu1yP/+x6Sg1xiKJe3OM6cUr/UzP3zMGtAp2OlxlzSqUwkL2Tiohc
VLvhwwCrKPZ3lIsmu1JCs3YRAPhr6nS4YPoZvY05oNLra/W6PxTd8nKBW2mbGxUi5fpood/u5z//
O2q0SLwO0kdBAZHCnTbRKMvHZEA/k8v3AOMW0U+K3LXpUXJXoQyVAgZDMcvftLdFR0KJ2OPjxWzl
LLjyjnoQcYdChvuTQq4FOpblvDmaSGjvJHCg7RiztNtvQczdVGETQwBjN2ebVPg5k/fNDVwkuIDF
CCUEFXcX2oP0Nu5szM0fjc3F12E0IKSqqTN3yIMFYZxPbW/3eMo7VrbS64TpmJq+KIxmdmiOhzyR
WJhr+1dN7T73JszKdREMhFwPgPI14MPlL0AFF9xrS6EYw5lfunzh5gZdyeYMDZisPpmhj5hYQj7g
5X7ZgVQPi3wg67UvlD3MYV1apjWzusYVpLa28fmXFrdUM6CdXQ9mLgp9hKuDvzfLnWWCB2bOc7GX
fmkC/fSiEBYgchC2rNWUmyfLgrg18rBbhIV5Fif2rF8HxE6sjXBfNOjBQnJ4ljDVlVmLvVobzymt
XjsXLcXCczj2bc7MjWe2wW/dyIQrPvIZeVyW1V3N/UWH8FvxZXdy5/zfNJBS9Wg78bulGwQ6vdL+
E8TtJjjg0jwAL4L8STx+49u03Kind+D8t49SiI3M1EN6yQ6oYCk8ktHwkC15xVXJYef19VNkaLMp
RIwM0TsnEVwL/E2EuFqdZluHW4gpiLnRGvrdtneNsz4wuUAMSWmiS+DjiW2xi3qwTqxf4L1K8OaT
C5uTF3s5K0fq718UE1H/xfI7V+4Y27Ip6KDjW9KlinVK06wFc02ycNtZwy1I24ALa3jaYBEe2NyG
GNOroenp3hDV49989AgQ0LLKh5O3wGjivEKDRSCB7wdhZocpJIUuBkkicm0WlhvpuU76prt/M84J
VIHDhHMp6uZ/6mayG4SNGWF+egh+9BcSFwrDRu0E1Gh2zs1uVI2YVBK4vnD5UGuzqyo0uULFWn//
1tmXaBUI6LxqXG6n9K9DvCrmC8Og4p3ptufKPqHCDUO8Hqk5/Wf0hpUR6TXbUzZVcm1eJyn+iUyc
ivzX8jwRistudiSzH31Zx3dn+mlHGH5Yi5DqU84WJ+J8Bv+0npk+DVcYV/MhT6LSt4zvEojudejg
tmhsHSQSnq65rzsqKK+rVzGRoKZcrWLQrHOXDWLwEZwgZPhPFERpgK6NaH5mps9V3uuF321dB/U1
EiPME3mLEld6sp/N5hBTyw7HujY43M7mCV+TnfA9gtt+ukeRnUi8YiOwgxcZC9adqUkiJyn6eMYS
Up2v3cXmFrwn9NMfkeRPEgW7OR0fDogh+uK1ADmLtdCROmhfi/hO1oP6+bmYzT5L3Gy8ioLOz7lU
e3hzBRNrYgwJecIkEYGrdjrMiGiC2dAEsFzK+I0nCHN4lT1loejvOtmHd17ZluKdAD5D+qdMol5P
4PXEDp2MGvUX99Bfw9/yzvefYUflHOgl5fbcan96ucYnsT+vUp6mzX4sa35Tub3jMeMC7wtelAi3
hcUrpKsIyNmWIT/B9b8FPJXJof4podgvD1/xsBPIIcKG/VRB3+q90bjN6NVwZY5znZMraMHSD7Yr
QIWpbf622C0UkMQsyKiiRFQWKH8mB0MrJcmuW7iwbapwa74JZdzEtJ2u2v2SFKtFu8AtLlKJbrxd
L6HAben9PBavMwLfomi+NKSTN12N0Pt2dx3/uhUsJOwmB42zgLfRS5d2ltEXObpyoY+uAum1mw1C
uqTIe5BiXs2nbtaWtNSRR1PhIatVS9/uZXsapUOXiV1x2R992gQyZhyD3RceyZW7OvY+cnqjBkqs
CmWEu7fxXRJaX1uH+/tTU020W28Rk48TuHS/zzzzXcCBkrhKyuvc+TEdFr4H7dp92mb+skyAqtRG
vyovRJ21EPklKpbq7xcOvhRwE+NFn7+fA8/NNLCcATAW9/R+hfsK8L0vgp68vEWHI5TJ+Cc1axhk
dyl3oVm4XQf10uMiEeUWH0GbGauKBTEF+BZh5RzZmD+CJiO92UNi2LS8Xx90rsbv1+jsQYKK+ax5
YhV3HBRCTqxESFz3f4yobslF0h9GvEdPmz2kvDIi7prv3B2oopzJ2bFe3W+n9osmKz+5mm6ERC7g
AKLhSimkmS8Yo0FtFqJ1xQMXicAZ6Lcc/mt9FRyotS6Y8VzAZJ+jCiQJl3CpjTh8RXcPyMfE04R5
aeXAr3lui3hC8vA/IVjVb8sDhMLv8pZpiEHY2/Ou2uMogsiz/e8ERt6Yb1kAA/iw64UJsyX6iRo2
0m7phBRQPT81JuABtnyIIBUQoZKdxuLhZ6+G19ChXai6vhrVBkUR27k5DQMHx6ik83RgaPRzMnm4
uUICcZD9LdGyAeuZLb4tP/nzBS8HsNicBwCqPtbcKwTJ4dj3o5NvvtIxqvq74c39KjZfaihI2z0m
6U5NWo7hy87OIevdxOrZMsC7IQyGnm7azTodZ1ykZFpv+3DBnjh6fL10A7RFTFQmg7/G6SishOQx
sM/cez1vbKoxOFUb9WmGRTgn1MGYlUrMNWOqJU+O1DJi86RiVcfmXKm+0rFvfG8OhFSsSU1OunzO
MiPUeCWKOoDpoaLTPf+kKW67OGSXTnEg1UZY8q2HVS+Btopolnd0tzOAE/l0G1YAUdi8eoE8RP8k
u4r6Y+r+BdijbfRWforLlqt+GauP+3sRvzjvD85bHU2MsPIN0oYkGb7mvCnBiALLYhJQHSUuxpao
EcKIumbd1JpMAKl0syeaZMxwWuAgilDx5bp2RWd/hVim+ZLoWyoLUIxztCAI03A7SZX8ltTuDdyR
gEkoOzo2ZV//2kIB64n9HZ4Qb5thh4uD7eOoB8F+7XwLX3HI8aGkmyUycLYcUCqZviNegjZkAjhs
NUFOwPYi5ZWmcIAw0sqbXgL3l/6jZE/ml9Obwi1TutyCvg/Fk2D7SezkPH/3rh4khvqBus2z9THN
ayX2AkrrCyWIUqTv/tw7nBOqWDRgYcHSh6ON71cXD+BVywuDTW25wWWymp50W+qq3r2lBHiIq9aw
AAn1RFU9gcvzM0eOfbkujUcxbhJSMjbB52TGxHxKHXNI6sjqE/mvrAcYvNuyuhneYYq+5sTE9f+E
yfAw39/EsdWHzGdc5srXbTBT5xg0saL31w3Up/zR3MDHy9sw0u/NcZmZt3ImLu0Cg+rsi2J9Izp2
vPU04ww+qFz3UcBtcu5C/C04VzWwFUIGBkfMmLine7tzhKYTbqKzt1dc7KkAkufkKr4AlpBOFH+1
1Dz1tXY1vaxIyxEUhhXYNiJrPqIcsqmrc7xRLdRE+dX8O7NQOk6tsPyPSVT0EsoGi7jRL5oHBjqr
2KYTIMK3iqKxMgo5v4+bAqCiV8gDB4g/nYQuVv9SRI5UmULn7JbFh+w30rKeSJ3Y37mcvNUM22Kn
Pww9OPDogxyaN8hFEYoJyPrMN8Qmr9phWIk7NLNp/lkuBNVMNJxIISDSEwxL1fIpWYPFEnv0hYeB
68DS+9y2rCB7V4l3Ax3zfJHRHnm0DGe6Q30CppIbQVJGg5O3/O6smvpu2E+AlbLU9C4d/QYJH60p
wHhEfcU5f4CfxKw7LtrFnK9Prvmpmwpfbk2PxPkM2eEJUFcXK69XYksmoNhoIWTGprDSnFSX1ZVG
RxseDPTEQ3BzFUB2fIWc5A/sPPO6S5+2KM2OjtQwPYiaVRKwMZJ5TOZN3hEBYtSD0A/SVvqaALK6
jnlJtXm74ItDccYJUqr780MoVe1tPxUcOm51PAOt6PNUvFLr0Hlpagrb/zBur885cqcHUrreh82o
WBgpihDmQiX6KWj3ous7crqJdBoBfww5Hp7DexgXya5qUe/OLwudeJNaPkxoy7anM/VPsdbQ/bSf
kPlJGn/yGx9izj6Cs7XaMNSzY3664mK8seEiZUI+CyD6pkpLb+jrdoZJLWnfcV419iEhuH5yjqSC
Gr2tyxf6z9HcLpPmXT1pfTas6MhH5UpFEw3JBoHCBGuZYYf8sHFG/MwsP0SfQ5UmRG5lw6Qvdk2o
tSTxFn8P4EL4WpVJMWKChOMPQ3X52qsomqmjQtPpQoekefYGv9ig9CIOa3rZTw1NbacBXKMZ1IR/
H6iZYTeF35IjzRdfc/DN70CAB/4cn2tfHkkYjBXVA4Z1o7RCpglTM+/vlcgKW81cI0xeTaev7pJK
xt0uIaKMy9fTH6LHNy6ylU4dxWm/YChlpqXY6x8Eq7vrf2gxDOk0tnvYmNR0n4TI+dNF5K2dA3Ub
ikGqlNk6eszBmJPaEj07WtXtX9sm3kZnEcpPfMn6PMXWtA4sr49IKybkTN3TvUU41YrAO+ORRVL/
zm2Ag3T6sNaqLg+FSakePiwIqQpI6it0DqA9lWDQ8puFs/kE9OHqKu0g8gYno+ohzoN6R4j4WH99
PcGdVnp6QVruz/pQ478meZbxG4uwSUif2pULqe7cVvqEJRHrCcSs8CG+lfkCVaVQ2yBcSYplZ5MX
RhKdednsfxT2x/AiXDxHux42Rw/fNl+QwqN9s/NQFI/c6bMu3RpkRCzcdT+jCCmUPgq1Ry+Sah4i
OYMeBoS4JpDO3K7yhKpKqSC4v0w6M0lhrDr0HqJoAlK0y29ZFHXzIOHti1GrjbjlPtayMqgSyOEv
zlt+T9QbFLv7h7pgELJ4MBzraJ2CZfPpW5Z+ImoyM/0DV+eV4yrlG/d5A4Pt0iu8L9E+LBifyifA
T/3RX8NV0Qdx1noX7FZxa/jMdStOeVDLFUfyGbSzXc8OnIW/+sr3bfB++zlfaPB3ajWP9HRGCaMa
6+fevhqdR7iyPasIJeRze7IALS77rUmTEzwUO8jjOh182u7n7tgsIhJWrBrW7wAQISRUoYBB9SfK
9PQqB09UPcDgoz6mbyLNggl0KXSllSppPlOh65wyhFqbm6s/kZKolTxNywQMw2KPP5uBnNtoANJe
hDKez7yL1taGebYRSG7fI81mXJVh33lGGny/30n9rGHnUXBvL2nP3d/nQqimOtOPB3P3sGw88lyh
FPZ1NuuNwrND+6mfjGPFC2av/1LeSvHbLwCJbgrXqhqmnMUfzLG68pydy7hlu4nu3SHrHER9OE0f
9vri/eZ2lny4xIu9Dc1QHGkhZlZoNpXSESUNneSamyavl6Gt9RbQtGOFolcTAhfmiHRYiwn67jio
c7ASzvjGsXHKOOm3xOf0TLso7UNGSdAEKH7WrRznveAfS+PJCrjL6/Yl6pRtelzWVG9JH/Oiq8mN
0XXqRMDiqlddrPQdQq/Iy/CMfstrLfgAAs9NCQKvpnS2wJejcygo4Ehyu9zzFFm8VdFHB8kkGA92
5F00/e6Aed1HsO+6KL3oZeOffV7FnBMmeW8TzuamW7A0RNa2IKTH5JmOgVJ2cLR+5/u1sUf51pzs
rwKwo3fuy9KpRnTOeGXwZ1Psjo7dYXY5cgX+MIwytzMy8oCs2djh76bHi3J1pUvpaoJUn22i3Ba7
Ws1+0ODXJhTsrE6wZ+JEjkhiAXAQup0vZLNdr2xCPJvYi4tV/cYh5S008kjhL2N7zQBZO5okeAzd
JECBBHqQ0ARnxZF7IKq+nNRc1NuuGKEJGtUuBBJ7TTVHEV5D/LKckYjPiQ3egyyjXLGAWKrEvyOO
BsHtEEI9rgwAQk4u4hQrpCBFodHjfC6jL1KlRh7BJpHIdosTksmCRsDPDck3SZD2NnsR8JgcOG+o
QdZdxVhm8hGQiCNsN9LVSpZTIpMHVhc2GckrY7OyuHBKEH7+p8ZHoEisAkii/PZODzSklqERkVLI
JmrZ63B+qcvpD/EiKH5+tN0GObLscMsXHpIEQAKl3ycboPoNSmJ3bdBa965PB2QSWFH+218iBAnG
cQtKuMqCFxKPpzDisvSUbkdjK/ny9v3W/BYb3iSqI+sqmMbTdingafKFJSG8sIFS+qa3lNo2Hpw7
VkeQxjONBVIXkWgzQWw7JkDAwvi/2JCF0W7d0tKgh/6K+KxBZVK7MOyDD1M5RksbmPo4eRR5RrPS
nfUHT4iVR3fc/Bua99LzTMwN+TEYnVOYY9l+jDazLSVKi7A+k1leEq/F/LxmDBW0T9zFOYJLLSwS
ZM2vVXxew+kGKM0nbd9p5V5feRSO3J4rVU29bqIHiQfB22Yn+1Yi3cS5CJ9ISH2QqGlPw6HuvCZ4
wFiM9SV5AaVkluh833Q8jIZELWBBQpMiAHAVnFkhAf1msdQYK8SjBYyg+ZiHHRCuVC4NuhjfNolb
7ahz/k3SxM2X403CAiS94WIHD3AJVjIJBnxj29issWpCSPi80iPio3p44WdcCaiH04cSQNHD6Fs4
Tdd7S6OuQ8G+bKYr4RrJcaNKZI32vXZq7MoMr9EKXncroyAqyORdyVzhzGU9iyaXPnPvW+1830v9
JMIXud/ORVSAaBKf3XlHLTdQKRqeVRaXkI8eW3uFO0fI7Of8VcOjoFk0EkR28oT4SQ0ra6SNWMuF
TR5AieVRHXuVEd91tY2/LyjACjid/ketdtSVmbTUMcDqLb99wkvIEAxN8ZyKdlUTAj6HFAu1UnPr
tHRtb1WA9rd7SFGBuQYgBv6IilhSkZ2CwShOieQ41Jj6KC2puNHLsJFt0xuzBp/Qg9YHVFlyAnwR
9mn0ybYhHFV8n5O+vlnPey7rX/H3UFlowL9tgVKE46Ssj/VWhtB6Y4ZZzefUYTHxQxcCEjk1Gevy
KTgPZCZLizmt8IfppuobetMI5MZJKlDXvzOYLrb8K4q1xi4t3VRbcPJA1C4+EkN5BxU2d76LawZU
5a5FOyB9TV4QCQqb2DIS/ES2LIXiZkZT1TDQMQWnbjlfH9xLKKuChnSK5WpCEqAxAUkCBPzHB7ad
BEGik8fjG2Q32eb3DdB11oK20LeV+yQ1tnWJWoCaXXSVREDLWPs5ckqj9T9VTHdNPUyMXKSV0YIo
hoHBgfGsR3+6hU6DQDySBwRYy4BKaS0igSOOAjRh6LQTODejifLVEcg046rGaGL+Xu/TWhirjw1m
T4LoXz+S4xKQGDlzrmjoDVFfyELpfUBTRlNyHGNwGS/hSNmgHj9rujcG9h4h+lxX/Zttfzu7IZ51
J5TQk0lvk2eaotiSkfMnRlm9dXFww5NeLx5/NUjG6ZXx/9oNIpm+lEM0GUnTImqZ3MXzOowdwohk
SgkXiwWQJ5ASgG43xtJPf9lntJrIWRNkr65+HCYN62b3CAq/QHD12r43/gZp0xrO/sFp3s/DWciL
FeIVjN5mgNbIZCHVxg8zCHT2XdTdWt00Fwdeu9cP9UBj7lyljadbuehQoyQbnNd/W3mCO0t/XSkh
I5IJVtdz21ilcKhNpAKiM/3Ce0qKbOHOpkbHTSH0Kbxob8PCdZum5O5fVyYkvq0K93bTxdnxhJTC
TmVfFD7T/T5l+wmNlnGu7Olc2V0cEnrEFz4N8JE6MoCUsfoP/p9g1Os+pgc7kjwYWpqZvVHObFDU
cP1rlJ8AATEcSeZnWqX6Kzf8r9X9vqzVKskiKy/Vl/ZeQW9w6a62kFUD/OwqXGRLczisyu5IS5Eg
UDjdI1GcQCOZAb4u8LM60UqJPGFOo19XqGu1QC/TbaVu/r+PPBTP00zGZD8QOJVFkAaeZM+P378g
xwVKpcFebS9oJ3jAsM7HYEixOYzoEXqQXcHDO7eNbcRtZX5lL1Z5myerF1YswPiELn2UK3lwhxlW
M7l6kixkzRt3li3mV+kvmON3L6o69Gk0j627IVCdmk0OlLd3IrDTq942DCc7MLBpryc5oet8Ht6J
OzPFERushAXKZqOVSEejncosSpII6lKG9OvaSjTfbRbQ59R5Wi+Yvr1GaOfCGuPe67XLhZsSXJKj
8PplSEUxbAp7XvJvZhJNTsIApP1cB4pj1G477x6f6W3s9rPzkFevLcsi+PP+kAOjuCtHsgmzl6c9
5j411XgrTXcDhevfZAGXrn0klNoos+Qy9sB00HV93+lBgKcUdLPXlsdJnbDzSL4nYBgrSvAPv7bk
0rfA2FQjTtxpBUUi14Ba17Na2Q4bPRsbIMzTNbMm+I3lnj1XbG9vift810cxkC3pC/iPaAPKMpE/
kSdBqp45Lw3QLHfwssiq92/Q9Twz66oTopnQ37mMWVyiYmtUyHhkJr1u9BbCUIYk139mDZAYISrP
HPXMR2KtE35JQxSsAqqS2x/NFdE7SDHY5Ee4FZPSHTXkv3vQ7CWKgqY+wfCy67BGeBmj+OM2j2d+
mRoFx+lfsw4NA8Nxb7LF2fep5I3LNkrX7LLpL6uFbguwE58k+keIHra2kh/hym+C9pJc8cbty4OP
dKIerhfC/amzi4ehBtq5LLuKhS9ZXMauRgIMTgVnfU0aO5KNDqMRfyAHldm+PFL3rD2/hwfew2qc
zpi6LbqHmIUoE6+/p+lEZMbgrbonIHsMKCxNE66gMH0fSROFdPXoVQ11sEpENlaK3Jq/SkSqlcMn
cbbogReT7w6IFcG3rf8K8F+C2zugVDLBvg6wv8U7TtJ8xlzSI3rm5QSYWP109zQl5lRrfcW8yUXg
h9JL9nwVEXseQE0aZOcxgeoTWcEhz3xEep+xx/bqst1qBBc4AJhc+vnARMs6kPilzc8FPeaSdP8r
flduHV5iprzY///O1ZK617or6ZxgB4fboGyQyyFBGz6stC9QZrxrkRTB8lA+xbM1jgyDKbYvXnsQ
dpBxCJJjzhnU2rBoD3ksnOOXxaxYuNfPg0SujX5pL8NvdY0UPeS9R7s5kUHIQNQdXHoe6XNMcqt0
5cvNFeiTRm4/aknAuh2zvgvYsn8zheCwZl9mDDl6brGe+/FhEqEZTyNTQmAa0k2iXuAw2yM3s6t7
ce6zXB5dKQkDQzJhQcr/x8pR6/1eHQzwo0u1T9sVgL3xA+qqVsE1PCHG/qTdHkVqNBbhSc13+sNW
L4lrdVSnDItvUydLOv7bX7zSiDiSqWJHx19d2sMrFKVsCXs3lsFaHj6ySdLMh4RicKWjQszk8XS5
SDSiWzbPoqhTCtwMjSHQCv6/41ptounclpTCOXhzkNTg//JmiKsP2k3GDk/YnK1b847jdU1+alIp
saJRrKLnP5AW6YpIK7Ooi6jcBIq6M8aq2/zeEQ2WdxgZ+2QT9KxCKy55AFhXGd++DsZOFXAOKVOD
NlHQidQQgoSPuVnzpqQy1Xb12ltjZ8zBo9pm9+UbgYwFk5JnG7RebuLPRjWMy7gGf4hBP3nCWt5T
pRvMKnM6fIfrmFzuVQ07+i2NH3pgGZD3Pw741ynMHmrq97lBRIwIPMzqL6AL1JWjL+LorA6tMag8
CTUW6httyuAMv5ah2tIE2AVH/w5MkoCKDVKTzTVuSkZeNEWbAX1aEImZJm6gx5PFjeOCuD2i5H3D
pPm4rx4SP82yrSxdTcq3ntRAsg59wggLRqu56pRfhctyRKZGc5zWUXKDKzfP+T0QCUHYMGOIP1Qq
PLvdOhlvScgnMDO1HK5lOMrgtr0MZ+050NZ0fpgic6SArQTj/+8nC8KOpxmxk+2ZVdTqDE8DOEXm
hVXoEfMdFRzbbAlkNhYZ2fqzmM/oB7nTr9KliN8Y4WPp+g6YtEMePivoAXm6M1MTE6VuiPMixIRE
BFBTXFelKFRZIuK30zpEx12DMy+QBjjnUfFHu0JfqYy09Pxk2XfSiPMwNEhYk9jSDV0v9/ktP+EA
L/UZgYsgqYBwZo397c5neX0hVNxWz0AtW053+qP6dpQBJvpjkfwpgc6jZwxVM8kist54jn5e1YxQ
wlRGVWJN9RCI0D50yVr9WmfBcnxtNl3ElXou+21IE7/Da2SbgbYnh7wqIDS/U6EYO/YiqDW/Y3OC
zWtjsN+FOuSxBQ1Adpn6T1nAawTirwCr390FpC9PKN6Ohg2sXHGTZoHQys12lCDMx6onPUy1dP9i
g4tskz/XloIbIbRzgADxUsqXx7osXiUtqa1f7Q0rT7NUU92lcJPUVVX5nneWBpr99h4YNaGZubkB
pij8pBoJBdiHwPrS0QcYD0d90HMTltOyv/i1VrVcpK/EiqlEROmhzkTAyz1hT+bkzY6AMYo2Y67e
JvJbiqnfruX5b2CZgVJ5Ne+48lKmjMIh2aMUft/0viUtQ1drn3OJ8gIvMBd0UiGfsXFkut3R3+VS
5NGI7N+IH1fT4YgwtIdb82BPPHPLyLjlNI9FF1z0OAsUoBVNWmUBbF5arOdr6PpOvIftlmJkpyT4
QojG8P/MJgq93jPq5Wv1wgjzK0XP4+0diu+ulVJKuDYvTpUdKVsklqZ8locXtpWpSWExqeoKNTIe
FzV1bQMDfEoeQLWJx/vcOLS4kp8yjLfYjSw1jKk5XZ6lWpYQg7nE17rDy3tLmkoFxd+wchwOAxkO
5ocxlH0kWxXrlzId9jBfHM50dG8fXKRJdiSxdtwC9/f/oQU8YtK0HgEzuLU1D2NdmywNUfF65uYR
A4W1hNPXfJQH6LOeb6Xfyi94tuXkAzOvEQDGyyI01NKYefXfbsqTO6VjiHnO/Aw8G9nnizhDjEhW
bbuxkRLchYRKAt+oea8KBP05NgQepuiAE8V2xmD0jiYLQHUH4YpthkXxi4SaOjwgZDzQsyPgtJ9x
hkTC0zj7cvz3e0L7d+8Zo9sowvGPhd04kteEHuz8L5lfEgaA8Cm/LfJ9Xu+hKC5oadtmhGJ9tn7Z
PcM7rGs8kX0BNdz2+wt9LuHpS+mBdgsuffpETXvRBXwgj4W6PYWueVuv3GcNFjpOshjjTEdZcfPc
1VcSM2TQRRpVoAI1q0cYfbqWwvo+OPU4EnXi9JfbghciIU6pP//DtM4vh7CmyRXKCGD1ySDSTJE2
mUAWkl5BSli1BkPDLGqdKzg9L5se7PEBim2bhB4R2vWOyLXhSzqMCIVVbAacawcLM+1iaLNQBqQA
UoveDF2IjC1b9HcdBHQTkl2rToWqSy8EXzxosHlfCsnibPZ2H8R5DQN4fM54b23EfOz6/T1BmmPz
TpJ3VMm/Ie1Wy7coQOOtALg6cITmkIotbJahZmxU0x3ubxBc63IuGHtjjKWe8JZl0SOq+cetpoSq
R5xdPBbnjjaQRQnOu3mDRe/jmADGnqL3XB63EpOtXgG5yiJzIU+NjzPQLh6UlWpTt1AvkfgsD3d1
4H2UiUULW8u7uoWbZqLfrBzJx1htg93FMzb48WfZ+LDT2v3QE912hv69pL1k6nbvL0JbSftu4G8G
3Sqf4fcalLy8qyxErth9tYr7m4JRYfW5ThC3bBrLWR/o4qz6WK/U0w/fr6TJ7ru6LU2NTkKu0QmX
SkGs9a2w2Fc4VjfAEI27AKy9G590z5nofaDG/EESdmOu1fXZfVLe6FamOJimqnXkpxUA7YKkSr7f
qhbjpT2Aox5IuW5DktRixlDDSI4geUJ/Ezpozf5JCGyaO4ypm9EsXdwVvwFKJc9IyRljoWHKhcmv
niRTNiekJCMqFs0Krplo9C6yHPgt9xmoAsXbv74DUNSTICRlW6m6nNpYQt4lJ3SsweSua9ZW7yMq
r/M6J0EP8t7JH5f1pzJ9kwtAhCYn3K/MpdRyg/w0NX0DutZxfZhaGWLURL6TuvKf2xX0Wvvjt579
Z8/CQ6FGzWDUE9E1xgvFQJYD4cAc3tonE/GZzMvG6KJC4rls2qik9fi5BCt+qlOvFFdt1SpsU+ei
S5t5mEt4vf1nQN8yb/I+qdq5USCPpCHnZtvGxJTi6ohGjys5DX/mkPlX7h+ZknUQsABB1y8ee3nP
8f1SmKTEZaxWKFItYZQGi7GWZBjlD02H12CUvRWWIHb1cZEGqYtXHlwQebcqIj3OkNg1SOIv0Yyk
fOAsw98Z3b6Wn/m96wGD5i748kvpU6fd+5PgB/L92QKRRBN9RPfiY7YaBURIgiYt86syEnXWj+ip
9Zg4iIasG0elvVZWlfuv0Uck0j8S0HJMR/mLDgLgfMGXsNmeam/7sZ9n+CFWjkp/T6RgZgEVLI2S
uViwU4D8ZyqrmyZmRwn8ZjWmT4lNQZ3NsbviEpPSCqpznFy1kUrTtk6ee9B9Zr1PlFBH/iB7dh3I
5r5hpkWXmnzfcOK2akBQ8Qf1n4CvaYxtIQSZI6AsCKexfGqr/RoGvXe89dpO+0qS92bPDnz8eLfe
v6ky2RVuS0iDl5F1tm0mh3ZZGQqP34WzDKBcuvInqtDsZBaRSijGCxxu42rrK2HIe/h3eXz0ohu0
QI1T+TFquv/vyuxPA1kpeQvEO38AFP4KpmFz1UsKtx8IH5Ff8ws6Qj3cPWUmGPmALjHzwaTuCLTV
lx8i1Tp011jtHy71whXxQdar+pdYWi87IaAR+lfmPgaBJup8gVvGCVwnNzW9HkpXQcCbuVb4+A0z
pnIp2aHkPyHh0o80/XC5vmFW1hEsmnDmrot6T3w8B3f98CPoTfgO6saYlPWuswUD9mioHKUepLSz
+zLqhu/mvxaKDzQoOeYUIugVWb7WAhAhmOXwnpSVdoTG5enZtcWYzLmmbSQuM1U5LUqbVEQqUfhG
2WT+Cc5qvcYJBFg80dp1VlF+3fwFrgCzauAVgYmByYhdlairwm6rlIcxQ4ObWBPQKMg9SbHTUmhu
wqCdoB91DyGSi/OZEmBsAncFTmQP6otcsS/M8LTACHM3TJkJa1gRg9nXwYDd2mT8Alt5Zcd99GYU
uhTwWgPF8y8Vl4le1UnJEKY7eKcNkOUIRFBly3458qNY7xBABjeBKDs+03KDfXmD8e5V8dRSy02S
ZdpOiapnKRZpndI/+zRq7dfwdBnbv44e+Rop1l9KPKujqO4vouc0UTmgJrwm8uukyAbJcmduoaIn
5pxTUxO00RnoAZrLnojMjYdgg67WUfahg+4fl7aC1VBTeHolFjEhOicAfaPN7J1SqkSz1mWQtStA
8CVd0vNjzCOYgwDVAN9bVI9ZXV8yAptiG0CBYA/6IsJls+B/sTaL7l7X5LWx2bk25i4ZAeNyHYlq
P9yrYPBdysYK4EyBZap+nubzXi/LFeVJIXG/SxBJqgd5Dk/lC1JQbvJEIYrrfP8itHIaedvWMhQK
/w/zp/8SNptG/9z4EhBFsc3SD2ia98o2zqVVm7Z5XA0gmv+ZMZlyCmSz4jloUWjtuN68YtGjdRaU
4kPtNjTVjo/giBLgXU1IMlcW7thyZxuOLMTcozwU1arJTR+wibqMvkdD/uR+kyYq7so9i3lDDxaZ
69AuNBuRRKIuhlr5Bq4MgHpbXyH1RPZDv1X4077XluZuaCBWLEHl+Xdlxx8yCzDy3FxTTSRAEFOg
9o+EftfNrv5xnLqbwScdrvdJXlbtpC47978NgHUpApbSUvJSIxrMiFcfFnpY6keV9roGAnJ1xQoZ
USDSZSG2JxIcef8P/5w3GcVXdJW4wVQxPEZRX+ZJJpGZ/hiATS08aA/hCYOqqsWQ6Rsr0V6cV+3w
KJKssDVStFx0vQleRqDYmOSvpvIqHo9MOZ2NHP9eFItwQhovnFYF7pY9hLnjQgZ+NYCLMKDoj2n0
lE+KDVJ/be29IKWXCOez7mMewsk46TZB2/LeeHcUplXgmq4FldM6apid6Ggp7EP9d58RB2exikEp
WWbmNONxDZeRBX9VUek8zSx/SwptXj9P/iF42DzQJyEviT8426ubUGBPCnYB2AWTqd3PozTt9uQW
V+DKb0t+ns/KMdp4vMTkskjQf1115Fd+5gn3D2WFQxOAcYWu40vKYu+5FazCr2m8gRps+kzNz91W
Wkeu1Ip2xHQcF+Y8fDL33oPyS3mlawSgZdA58HGCtcSf/riygpkF7iUQBjwvidiTZDnoxT8GeOFZ
udLnbzNbCpYbGeupl2EcIaIvgv9NDAWUglwJQA5QFbqbjcS1Z69zO4ykopAjOKsY3h0MY8YdOLke
vK8JJVc3dWKB6hBHKHVsPquI4RAJ8MO1IkBJM89Bqck4W2q4+FwoQg6JBjs/k16vpf/06m9SVnln
MZoRh/hH9qGDAsKpCh6LeX8P1iF/E3J3aI3oiETMnLw1qRvnVYoBSVRr8rdhBghvQCkrY/4vxzaq
fyYqIsfuhRvFvJsdQmTEtJ/XEyzmyb9Iw0MUNsyp7T0WD03sTA9WpBLoMON8N4ISlYiELc0GlZ/i
2ukP04TapUDId7mcs/4XjgM4YUUP7rIM5gsYAkrb72eILF7pqAoGqlgkR/WKm7g3h6R9KH81DgxH
jhI9Pca58DRSSbVGoIfP6JEjtoXT4WNESDGUb4c+OqUWWzKU0xi7QshGTLnzlvm9f/1x2HYZQ9Xv
Z2CTu7WKIrhU6k3fyyUN3DHjFUx3fNwnYo3w5w+2ucmbWWF/Q3Vz8hE6PFlFAdBjXBkWooJDUVox
abXifCXlRql1bJB07jYYbLIVfYoGvE5Vb7rwIgCVe/i8+lOTCp+Mt1KYBtNVP2FnJzPRzbeVsz3h
TYunP0Ygj2149bz+AuqmJ+StsHvdqyrwlgZ9zwIRDyC3wxjaDKhxWt8Gz2VLrO0rAfREG7Q2aqX7
G0TXBk7lFDOmDF1JM05q8CBnVd/NnE+ORDWmCSitqnBB6In4qepFpEKmWcT5AeNY3eLBlr8zG2u+
aBBB/61yizbRisyrdd2463eH5ozA+4wYDmdNbe8CEXcYlKzX/WsLtUHzsvVD1/voLMVd7qsYQ7Mj
HQeJePPSv+sZyqi4uB/w9nQ1I2XWLrrbAqntEXQKzAOdRZ+K3Tjsleywql71Z+st2zOMCxRRsBYr
tcftZO8GDCsL+EyrcGsqk2TqVCKQszagXYOmgZQXJ+ERRpJbOAMQ72J+UBv6UM3t2lO11UIBL4xy
KdJda8AlwT4MgI3TdRw78LdQTND/G4y7/ut3WznFg8d6wztVupFNkF/mwwS2Nm8As/cBPHhuzIk+
Ih6lowOqVXg8P/vGvbAL5AFk3uNvTBuIaBIPVoUnyWSAbGb7SCS67NZErqVECq/R/ejkKxXyi8S3
mZA/1CfKjDtqP+u7d7mvQJA7X7k6j2fua/YL7KwdTbUPoPhO3Cz2ldxzdD55XzfYjdVmzAEqEN59
RkAJh3fc1Eevv5rOLJNxIVCZmC4S8+HSNvW5i7Y4kQ2RqRI0uA8kiAkIcJIAMA6fg7xO1cs/rn0v
E9NEibtZNilMvL3zfOyi6mcnoX3Lmig1X7UtMIJOUIIAfDk5Ee1fLwoFzRCo42Wrr4CGu0YwPWyd
8tmkCukpVn9rMd4bgON1TBDDEkrjwYt4LsUjaPIXKrIPpOqhlo1OcA7XZrsgxvOeCvYPXfQ+1g8p
/0XITE5h5FE7+urwk4dK9B7/QsO9Pd23Rhh3r5SANr6qgv1HXCakoapjZ7IGK7ax8cVF+08h69NH
e+WX3g8BA250wPoVMgf77ipoO5uVKROTMtlODAPDHt2E7n7Beboyf3UyBHZLrLAFmeqShUHDV+We
+cHL2MGJfxna0v0MuzqYe/JaXCGoQe/quVpqCv1tBYiAXhcaScRH/9Y74pTuCNyrZZFElQNWGiT+
r7xe3vxNJaj5jxX9YJYDGdfwYeLtRi95cwDmc+5Vlquv6Dk4uiSrFUvU25LqVL4OJ12e6b/2HplB
2f7Im+WhsmrdCBa4pIBRx7qTg6Zuqx+vSwz5JMxrbsAHHi5odgXcIUy8tcbScGETy++YG68/qADn
wdQI1PFzJVb9cahBCp6FCJ7bYLZLGaS7k8l809TZzQyk7MwbguUTC5daI8Hdj0qKlih53xTX0Zd0
CibS6WxipRWaNh384dmkBluDDQaRJxkpCWUx6OHQnxoL8/LNXJr8eJ+dpy38FhwQrKb72NV4q6w2
SLdjNwft1DfCiG6XFkR36872iCf9u8VBpPrDyEMGxfUDXbEvRri+M6njifa1jHR8tsCAELXKHbCP
iteKeG5rn36CUTaeDBm7PSEN92MtrleShyk2aO6iU7MIuZVGulyFzhH3D9xOE7bnijdOmNUWuB/+
hqprXZ7+LheP3rwx5HpquJjX/oZwdLOhmlmJ7P+U+Un+wbn98nCqWd6SaSDSKccGySVl/mXmGqaD
MM9sqSb2mEXGu1DiXdTpdIYn/4UVZGHdE0D1JPCldACFqf5vtJTvGYXetQG0vjAw0cZmSLiMoM8L
toEgyd3gERmLFRKnmH2/TCaRNnDFEHtdR0upCmEVkR3SVnEeZ2ggxRKVm9Q/LB2ReMpOehTgr43j
EvdNtPwoC6f2MG67+GxDrmWE2wIhPwk9sPHAHH3VM43PR+efnaD28nFApfSaPlfuzO1Vh7Jxg5e/
toEwuzzdF28dqITcZIE2eabivAECr0+otkoU//Fq3fCylENbSAByWrTY2DvbruoRjCduIDQo/svq
bNiwywRHf6vtTZDIJM3uoxuoPMTBn6Uqd1Ue5cmD+QPVkxuy4Ito/hQ15j/OxRnPunu+sxycu1yb
JsZ5ESgltbzChZ5z7/i0YEEv3DkaGN/X+qH+KyGv+ShR++ZHVHy/6gautpShUDC8FEOzleLh3G3E
vPR9kYMFGL3jAF+/m6QUJO6KT+Pl7dfTEQ2NL0bdtnc294p5i+KUrdqbsUhUvSEORyCxVbdJKyU7
b7S7+URdl5qdGZxUIRtmnvDXcbPTupKtGm7fWLWjfXcX+6eiDA4PXITvRytn/JRn1DgguagPBFZS
XjJizFDescPFQKr1MD2Gv7fgztBveYEDVgiL17tO9q9Ef5Mm06oiePVXbkTWmrmuW0tvihtAhSKv
Jpbcr2Y6VWb22exGRyHPPDXzILccxs94+0NYv0UgKtgbSzJuwES+2SC7dnSYwKXSLBeqdGusRxeX
0YY7rOuBwTp8NH1eDp6tvuocvPuGFbmWQsPgstvZ1WQv3+8cpkoEWdKTtZf71Vrh88KoJgdgsFPF
/2oz+ky+/heNwXUr7/Oue40zyrO5YmNtaxLUPOfMA2QiAmAvEiZyueuT/DaKYAwVXe6yBAlYx4YH
Lb4BXGnNihdQhqqVh+Bevg6pafoe3bnZH80YRAVtUKeZBAUhw8Xag2I8C4Werc2cfOKtMB5u3A3Q
VJp//fDKqru7xolZ3lecyeAS1hu3/eUxwPLIab642ldlI0hNWJ+jj7ZCifxw3R2Zmj6de1n4mKyd
zchKFWnLRRQX+aOkldhiBaDJhCKhJMSdYecotib52z5rC9TNDlgqHBQKjPpU6kzvBKUvsfTY+Pzn
rn8fRvHzAMdXywaDkB1w+7z0txNHIV7Nbjy1LcxZnCzzYcdkFVBHqcNO7Y1BpwZ9OVTzGrWIHNR5
97pbtyjwJju0N2BgpQ2jSr5X7R5MHaXIPFhK0yzFDJ6Ncpj+a0+dipYv4AHJbFJWFhN0yjYt7ZxP
xte8qbQeNaSVyaSD/WCNPfkTMRCC7MIuBw7WTsGGAKnNIx3yC1BURVWrUZdErjLwqN4d9aZfvOjb
m1FnenfHHwEeuRgMSoSnd8ANDrjx8n9sUbhKjh88Zzko0ERZAQkLS1GUtam08D3Vdn/EzlYQ9UPp
3Z2ScjeOatATyuw37fIqfWS2s+CwGWnZSneBLYbCpR5gXlkJnXSt2qNoX7Y/s/RwGkZOMHSvZDwf
25wzWx07Cd9h8vFoSREtuZ5YOkZIVGyUkRTM9/y9gWhSfej3WSl7j1oesZRpUnKcErkU+V48TxQY
RJXjPbuzsxEEHA28otE75219fdqFO5HkNxyY0y9gZJCqhMP77xvdM5kOzH8/Mlvhu9OiOvXivgJv
WMu2BvL+6PjzqgADyDtnkQIKPjypo/kM7gYXoX9yOohuYsEwTDXoWBAO3hN/m0vgx4cBzRqdqGvC
3WKtgmqPfI1meraNExAL51Zj/HWxFXF9x6P6uCg6kpgEBqCvMhKHyUGhIdlL2ZnpmQJyUY3YiO4S
QSPVrUqOOf7M+NTVa+RksJ4LF/aTMRUv8rGp9UdDLk61qM/KwMsph+f0m0fWDSOP82aa/QLzBQWJ
4pOPxv7DPqnXtBEzw5SHeu3cQo8hgTe+CUehrV19YGiDfFDvrs/eqRgGbs3gv/7hUWLOy49r7kOz
My1a5HBBK/4EKTzntAYV6NzodhaX3JtLyj3U8kfBgsa2H5eDfp52gEhrWSLky8flToOjkv7aJG3H
hHvwaYeL0Id8XT9r4ri4XYquf5pfafdzC6txmhAupgk6wJ2aS684dezNd0d6bt4GAdmf3fCrPkR7
KOMPLeRTdWdGHCPmuvC2wlIyW4JwTg9NR4Kig3LD514JkbZ1tU2waU9840fNBi6drTZcorUQhhsT
eNc9bN3haGNKzN3ieQDIlLZlw6B+vROMC61UdyeIJgFe3EYVwht9uokCpTBbSfiCSiyuf8WuVIBz
stL4ZcYsCr7hA3T0gTl8axV/es+k4GxnLRWa1FxcEh6CogGW+23r0fZl8xvdAFO12oTcX3umOLzl
oxYdfeYzKHpqa0ZFHizLLY7JyNvRvWlOMbvNUizlUgI+udd2WeHg/FigWuPs9FnEVJCtoE2hZ/Id
m5rPOKzKE6uOdSSZHBx6dh/EmXF/M6okgEjzocA+IaFYJggrmduSIhdizmrBBYSfRVTz8pMScurl
p+uU6fdYk7VCUu750/W83n0lmSk36lsueKHBWGyQ5mtLNp1hEFY3q5uBnWXrE6fu+0aBHRQ5WtXm
CXpwMwlc7xOT9SGsdPHKP+QOs3Molo98h7JaKMbJmGTTikbXpuZKcP/OfMU+lrfZQP9ma+pk8GOw
ClQzMNPDXT8EOwQGNngyh6a4ga4yDFNHyoQpsAudXKmtmh5VLkbCuR4y/ucOUMuSEJnIOLAJ1FNN
bV8O1yLgcX6fG3EYWt+bHJrV7mDKvcv7Qd0k4Vx+J+v8rQws2HfzMWWaIW9eGU5ThpnxWDaXpSVq
gAmfl02UnggFL1dsKpyHyhuiukKUg1SBAoPqUHm9EdKZ8ZYb3YGHYS1+jmyP9mnzhpdAp5fSnKWv
rU4N5bz0ExPj72bh7wL1+tSKpfsfFOLCNPfTd79AH661ng3j73SRL/mjb/lZtGn1qXeQVR4fGpD4
WsMJeUZbxhxY95po3NLymS2Hu0SVif7y2hA/HAVr9TL6jJfYW3W19p/MGxW2MkdWn07r+TnUyAyw
CanNB2lXP9ef+lrnsJzwfBoNzAcoE+hV6jvjGZ3hejo4BuME1+PsvXvjqltlEWqQW3uNaTnWebN1
Kv+ev6ogaIVbUfcPATUwFsHphPlu/9TDeT5NDcbS4/BJDUvD8V/ycezfiK2J4rpjfj0SzAMHf0TR
J1kFUP69xOTUnJ1iwadfbtES9BhuW/QhhBF8LEeaHkoMqX3D0TUwi/FT8woFzjDiBn0pPNKv3EVw
LM7kWbYZSKVWxJQ0HtWvTjuv+cM+u7I2tjc2emBmIOJkB61vxYdbsp0bWR3Ildamj0jgOgueSYqZ
TwYI4Jt68amqNmBBLVXqzclbOOBI3JiNFCeBlLfsSQbWyBgkgqMx1jpSUYPCtIJo/qm646hr+OqE
wzFWjPRU7YT27DjEC8OGQFrTOdldWsXRvyE3FQUx4CC5HjGTLP+AHpg2E4sPWmvPsEdZb/OVwhJc
dGBZ/Qie5LqLaf8htp4wk3qHJ6aQl2hiR/4meq3zlR1zrBy8yGfsiVcFrWr8mr4LskZ/qBWLXKaZ
ryR535lbLTdeLktcBhXdiLEO/OmJ3MB/8f7lvU0c2w6y7xbgIKHmvztM/CzwSA30REok+7HcCQQ2
4LSS5QY+FRzFAN/AMvn6xIj2e3IY69IdtHzgZyOes6cX/LgKUIbKxCONaSamAmoJqQaKl+TI+/US
7JAz1I8U0GkkPgKPUjJBB1LAQ0pn6aVbyb49oT/45ABViTqjEGOWvtceA5KjjNAlsr3QbElFtniC
bTq8YaaSixKp870cODhzbSwTUl3KJSzYfQL+uCZL1TWjpo1Lf2jVf06Dxh/nS7TVhIVGE7r+/fpt
n2qKsaV3JFlDNZB07diLmjkF1MEpK1x7L//HDHry8RoJbwXJCQxZJKch1HGWJIM8Sx4prLqBGPrr
CEg4gBc5u6n5aK8qJksSzgORYa8NU2FnJ0NAIfwkVXk2YbIxxoEP+mG8TZ7AQ09Myy7vpNa+g/RH
a7LXbd1j6IWYIcBE98nRFH8VLDJFR8yPRZgBB0S80HEH92rNj2HPqeES8Wkd+OL1SbwTHYDaC/qi
8meyzH0S6BjAEOfIHi0h87742IdYwzs1fh1mz9HpStxk65JfmTjrZORcH2TaJN9A50tRjB9ZgU1h
L0kdZdN++3J0E56MykRlai6s9C0Sqa1/sQnxbiFcE9GoZ7rNXkwgipbCv51PeqWRZMeB8aBNyN8H
aeAD53AOReNSMb5v0O5RBtppwr8k2JIfi4O0VIfsdocqFaToauSGTBvrdJ/KYAFMenZrUdpukTY/
IMDrp2tlzZq7bz2nLFHK5v79iGqsX+PI9e9xiqjQXr6BNvYVucYUkuM0fNHwg0I/FJhWPXNTV8Sn
w8fXohxHZvBbhqs27KtY6W6Ugk8Ki2epBlh+cWmaQdyXiMp1T+alerLScyjpfw6NzKWcfOZOoRTp
BSVN7LBCMLwviuc34sa8oLo41qI6rWYi9IM0xDTG9sUdeW7bH9ZIDc2eBZnIqjD6Uek5OYjdXi8r
keME8+4uyyBfpJIkNW5b+ozMkzWvD6lMUeJaCFQe2mGdTy/Q++kZXJb/Yr6HpMrFkZMFe6I3feq+
e7O+iFEgK5Zat3IeIW6NQ5JrOkrZWfiNwjDJXHTUDT5MVzg0VrzVioio298EkzLhEnK3xnUW1jt6
tTp/SxwQ5BjaFNSvDrYrVBU/dZyISfOWxqpr/xAsZ/4wYhislBv9xCPDEH6zQmPAa0ynE0dBAFr5
M74SpuU1Xb1QXJHU7/DEMjWHoXK9r/xjKjb7Ai3/SHNpCzaDdTY5nBa14XFfftUDXMvHDZ8uIsuJ
pawdrAMB4JBuBwWkzmeOkLx4i9LXaod7/WhzH0ZhqBE6+6ptacs2MPDvYvnRL2LdmuZX965Ithmz
GBc46yivbdrV7m3PMXAuKykKzJtErWzCKGOD0DF5BoKuwJaiGOGQmrnMBVC5dzPRlrpLhFAAm21t
KFjqAjgakYADn+Lu6ioZ6YKAHjIVTQcq/C8sICJMVHXEOhLpjH0kOvJPl04u9gzSD/DwSQ9l/Y8Y
aUZDPrAvczCAuajvOnH5yXiR236Gds1A3ek/csM/FQ8dSQeWaQDOXrls5wLAcMstySt34262OCQH
yCc6k5yjWv+eJlyUoovuP6GvJPWG8fJG9Jpk0maiBr/cMZiJcBUJEahKRN0Oot8vt5/3UTahzeKx
2Me8AMM0m/Nqf2ZxOe76ODcoosPj3pgpFf/Gi9SHi5LBjZfJ32WlwOl7EiH5MQm6yY7wT1/7FVIF
1K57/CoO071/uMLVF8i9939pSXFX1TmkoBr4XZ4kGremZceYfHKoPMkoHpL2KtwoAXslgnuOT7mb
J/FdWZ2mra+gbOwsIS9T++B2N+QhZQSNEwufw4R1YMvAcVQylC5gfyG9VJBqfbfpIgSsC+++o+QY
oGXJN5U5GXunUwacR+L4xAjtBCaApoOHISXZTaDgNar2FGglJgv0RHi/YgY9aHAJpzXq/SGZ74yf
joX7c2n4UevIcD/FwAz1UiyNy1YFx9vjm+Jtyk5dmafpRr1al1D48UCn3Qsf+J/wSL0FiLA/Ovof
/9wdjexN18vi+Icy6K6+CnPnbOhgSqVVoB2B8ndt3wno+LAG0n2+uq6G/2t9VYM8F0xlr7mZZfwy
Z6+6VGbp/ujSbzd34Rfsg/8QtBdV9jn2MjfB87/JeKy+IWSttGax3WaOYg4o36oopUY/cQOhS40F
UwiEiKRqyYvV5FlCwXCQI0QUC1NJMNIWt8DNqpBwCGKyU8+Roy5/tUNmQWznTNga7aKMn7pE1OO2
V3q3CWAD3DQPHrY2FmnGFVfGWGsklel4HuWDMIdq67jbj3FUFlyncxVejg823RvfZpVRU0IeUfJG
NyxZfFWXhnAX5WCP8drNB2/lg4pcCEnB42d2e+PcI+hNV9xRWZESXYT5ENE2M6pWXJ1ZAlBUjsIX
/RqPxrEzSr/DqwEOwenCDX0X6haNqDHGDGWAtZxBNXHkjoYQXu5fJxZ+Vj6ZFIoVDZvS4p8S4iOR
lMclfJ6Tuf09pmh82zwBbqlQLckb/S495qHXplbhbtietZ/YgMwXTfgreLwvltvczK5XxILiGjLe
jUj6IfkGHGpQkXpkzzn5uaOw3a3hQGm67WLPk6ydvyy2d9qx6hr7jzSga1EFm/BrDxGNhIVoDIJ+
vqaEeGW6JeeKg2iJI+upGWsrRmyafPycvIbzlUWdormo2q2qKHaGxarr9SOgWwaP1dsdsHFl+AGi
iokhuIf1xyTjnLsNGGXa57DVJt/R4nTcmT1Bq1H27oer/svc/gzWDpoNEzzh5mQbciibWG3XLGM8
Xrz8zhWa0bgg46sfkWfn0UWJjVMr/B4mZsP2B/QCa3+wykFPUwIq1Hx7ZFcRjunZ+7JGgawSOTd2
ZM57tgIOQWGe/+i7WJGsG46qJyOYDmSWswcmbEI82yaoQVYf7GfKfpt3ZwMoOetjJOBxc8+xW2+T
efqpUpRC5Sb0C5oQNeKSpaVMxxiDwObqVUcKzzBHJpK2BjgQsKVYZN04gxETRq+a64QAfjW97Bj2
mpQkGHiyYYwCMF0T5y6igjGeGMZBZSgl98i6BYvPxx4jTi/Vl06qLbl0960atLdBlJGI37Dq5WJZ
l3Ld+LlStn410GIla99NpwWwi9Z60SDlVZ/c/NYaelCXYwECHt1FvqQpf0hauwbFMfvyu8s5YP3E
O8Bk9eFUJNuPLONpdF9PV8L7Jpda2XDWVvauWjWlgnA2yLJzpXU1v/135/mbQ51XUkQ6EAXH86XO
ECYLfuf2OuwGljIfBOfGIuMKYxjWQvYn3rlWd4ZBCBi4I6SAQXFd6zBM3xFUCrXM+oYPFXqhvuy+
f+bvuoBS2Anucm7XqwRm/KV8gGTDa72USGg7w1mChi3eiAZQlTlVo8LOeyWmWDDCKNcnYLuYozfo
odjyM24z8S5mfIh6k/0UY1dAgTc9L55xbrvE+6sOSgIDbJWCodlJIKxV3IhkJexE4O+8YN+8q389
cwDjfFAeeH8dBGixv2tAl4eto8OtQabh86JgzQ1l+AxddeOPRc77BLZ5JFGKowAVO3teWgTXPXhS
alLWQgal+QkFMwMD0EZwVcuTGCbBAv2/gRQcp7ddk0j59neKyUFgeIQ9FsYlTKKsHOftDTMXmULT
7Keaft5BTKdIH00dG0sGD+Vbp7MjfBL7105TqLdqzaXpG12FEbMxHEqCbnN7kTWe/DZN0JmWecWV
AJb7520FYkUuBxm/K9TPwpuVK7fk4hL6k67us/XKycTkRKTRzM6I74AchUU3I7uxwywdnIa63WXF
e03Gb02x7FrGd+I7kABK7lOvrDMVVCAlKUKmdFozWPqKdyyd75418QxLmFO7qOiX5uYvev9S5mTx
etVf2cN1/RroTbw4jelccjkP4xolpheGDiMsSIY8WxBY1M1jqsZ6wQg28NehZnicqKW09Lh7jXT2
n74yyX8O0RWMk3xYCtFJ5LJRLgICRVW+LQPmy7A7v0nt3STR9gvh3lO9Bgj1ANegMobqOlEJ/74b
/40lXaxK0GfnnrXrPU2sWwLiN+A7DOm3PzuObOj8BhfHyCABKMMqICZtZgKyT6ESbs7wMteExx4x
ORCKEuhFAVIoYuZ9cEoQtQmezDZD3x57cAqYGjhJtGS7Ygv5kosyVrF4PuIEZVDzN1D7rajR1qQ/
hnFIgq0xLpqbktDWdS9vjrE0+MqIO0KdVaUogQMm+wg0DESyaAqurQ+1hj16dE7K2B4E+YPGcins
Plh4A6Niv/dT0VKn5fc0gI3BzMHhIGIr0tRKNmUNBHEgOEnoOE55TPeYO8wWF1cBjLdMF5C4ljiC
IDwMfIzGVvG5DXi/EslEKi64ozyqnqQJ0IQMjkrmdyZKD8ksAboAb4kKGrLH2ymYO3gcFa0ZSwyv
gLnsUI+gkAELB2NqXHzmq/BeYkY8a8CNFVazrYL7tJkGzhW5ZqAy6Dh9Oldl57GfJSnFrO+98rIG
TMooEhHDiuwEt1dwJmGSb7a1wnSIEBNiEabvBTzzDG5MIh7cPHrA5Fv1wHLGVT2J1KG454PrEJSi
p3cfrRiQDI4Rzq0tv75CXKLNQ1AoQoH7If+MDndDQiAE5hv4kUI24pZQGxhIQP/rSM5LMlUvk7jf
8alj8CorIN9GkJhHZob4sg7F1Bt+WFpv1B7BuQ6SlKj5jqJvMnnz/mRwpqpbt6dNG1xpHVkH5kYx
2QzYwZnHvvFab68pyHkxU6s1I/h8xAAQQqXjjXcuB9EIb4rre83W/PNXu/nOEwwohf33NktNoyRK
ArwrRRdOmuQTM+4bEX79iRrbGqOK2nxdPe3rxcCnqyliwhDGO3Ca9IOuRPxxjcm/q/NgkzFXvHtp
1MlWzc8VeWDKxtQUb85SeiIDxlyFSIHyFAUPx22QtzCt5as7KoNiz5l3o58/P5qe5h4+pjgMEKFS
FiHbmlCBhU8QYNoYfO8Zm9G8QK8EX9RlbbHnHJurkxuUFNLk8CdEpeABwA1LHwt8P7luNp5eIkEE
R1SXjSoZJBz/id6AgXtJmNJGX3J1mYgYWO6cBmM2A0aaEeFBCf4nY8paDwPZ4VU/YR4tE4B2SeAG
ynmXRpeaeHJNUuJDZHnzyaLL5sF3fQkdg/LUVpvmOr1PR6v0kBVHqDk4KJ1waFKCPK0uA9IgFoDY
LYIDCmQ5kUGVWybN6soGMMvaVHDYN2ctY6aUsc//n7jEmsYlMfSJ4Hc/GkO4Qu6ByOcf+BcxKoUB
59Z1bcEj6gVNttWOk4OJ5XpEKMDUCtDvlY5xd8fHap0ExL1L5bd5yzNFYsDivApPiqE2Y0NZmJZQ
n1grjkfO3qpv9mw71Uikkd7QdjU+XT/5Smhn2PsLRME7SMO8YLLuz/He4ZUTFrysctY7DjdGU3MU
H13bvwlyqt7Guc8xg/i+0Q8w1gkoSU57UIcHMaumSukFu5Kjm1qYljU/3yIseLBGcpksfGDFcnxn
oi++cl/E/Lrswg2O6b/WXY9SjlQqE+Baj/JO3avWik4JdfmzZV6mS8MdzoH11EjhJvKm0iABc9gb
oRcplps1MDVRNnvgXpkQ+o2oZdzcFcVjKeT7DYUQr+sDJ6/S8LFjZizQZI9s2zCKbJ56a83lwpcb
Pu3XSNbJrZdQsu0teluS/vrAOW91EiDAHID3DOoTmxWiMCVlwrLulEiRa2d4b1+IYsj7/5WDHXoX
GrStk99rhiw7JXFqk7cDl24tygj4Zcme8FFzrLOa0C+jMyrigIxUeG/E3iZjDh/zk/+cj7/C8d+D
dotLFvhHDXk4f/vTmeX97ySa4D2osC+w5iEWaEArL+qSMksKfHand4p0PyKV9nL00f+6jq1tZP9T
44zsX699NFEy/t3Mt2K2wwbYvBLjmi95ZfKIWYuRo/yI2MEgTmJn2yeFJ6tfdQ8ntbtikIvjxWL2
sqdt+YWX6QsG84ZsBvMgVemQDre4RUozbtzcCIi8GVr1AllEevavXZrPPPmg7mM7IxYNi+q7cPTJ
jA3rD9bA3h6aDbq8uI1T8nu8sypqmZ/oW/9gEQP4M0jQAKpGliR+93laUQ+VBp0wTVWrzsh38ji8
5zFY6k3TR51+2YxuzH97nAeTWZQj8bWkapPT8I3e1Bkaj0gTA7DeKFzqvJplhnxaptdzj8PxOb0c
2vBrUzTI4oRwZ/T6BM4/2nIC/wj+sPw2hjMn1rUTyBuurgTVRidrwFI57xREixBjrEht+eApHGBc
5B3qANMWeCvgi1fdZwtpfizLJ80sSzM1ZIAaZqAv4dFupK1zmkI/hFWU4+njfOtkyxKs5jFn/MQc
C0iwHpUBQgPf4rtl3Hihr9ce+WxmM2zzi6UxFsJFyvJ4pEX5mwt0nHvcUZmiC1dXlmBX3hYpBnVj
CwFkP8yzQ7FlNby/J4VDElLVSxgtbotWABW3g+edz4v0/K8fWbjDH2qC7y55/AbaC02GixlTpY6A
PrqVD/uQkDvgInsD7K056rSm41KXVoM17jenzE2aTxAJLzjIp9oZnoDx7f7ocNipQfcaXbqetH5M
2CL8LMTQ7qx4RT2Q52m8kwWB6t877lbyjFIMS3RPVqtvrx6oEuMx7O9N7k9kBjNo+tTlCTsY+eDx
vezeV9TTpGfCLeRvOYeHmHzJ0LM9d6FYXneEPa8IEiSYt8/gf+6U0g31erQqC+cezLKp/uryJ+6k
aogy1RY0gqsMYNWu7kdYOYttHOm0Bmin8ch3oRfqok3vA8HQGGSPP2bXtj1GawlQAemMkoMAakpC
6rf9px9dgWg/EC1JUSAPuya6PFiZPMpexNhBvDzgQ7Y6h7rcRYT1rD71uMFZgNu8IzMICU2jXqqp
uH0gLN3V83FETK8PZ4FkY2q8viZl2xwwMEPC9xwWkghtbYOHuwIl29miNRz3rNhlq3kaIexG+Unk
deyrNt5ffMZ6NNV9f5/hmvzoqzcL/NKSFcnvrhZa42rQJubccoeOtiFLC+gD0tukvK65cjFZ4hGA
egl0DP6nvgZRaKozGJCi9gACGfN/Awuf7rDHXa4CdPIh1s09IkWCVgUkC8hPvMexour+VSbQSguB
iiERYmOuJRJii7DBO98C9Te5N1KORfCRQUAqvi/UTzV0uAYtvVQ64b8dRAaK6EmmUX6dt1fbqxnM
lJffZ6WaqGabs6+xUJ5dyXNVRTVmUh6n+XjpBbBXbuZSZXN+ak94iNE53fJs/XibyuJAwWeYWAAR
ZeC/y+aZvuEgmlhjU0D7vUO1XtnmQBJS9brpT5obYciIU9JH7Hnik/Fyg9N8RQiVKRPCFPyoQm2J
WKnPnEl4F8DwiCxwwSTLALPsAoMN80hzx7WDEKwz+fCnj1+P4AO5mf7nWbd2Ad6XcNCLxduV/MNw
dta4jtRl7WoaR8uPUQvCAts+T+wuAiv7QF2cxzlL59KMYXy2I0QZNE6/Vn9x5FjvWegi5mt2YBzq
W1m1MsAdvvY1uu2cD9zFY5C1+Ytd8cN9KHkpp8EILVu4ebMHge9hMmCtSdBgCBcNITfkn52MFyCo
HtmLE+eA8cAYu9a6PAK1iNiORA1tUF2U7DN1G20qFBxXGJ+5RWWoWU7qogqsRLPCrvgGGWQIX4J5
/HcYsPA8lAbbFXOC8bwG93Vld77ql+n8ji5BW70d2Q+AzYSMKuJK+gsATd8KnBgsprQ3ieZIh1ev
+YmJ8ik5qN8dhg8vDRVEFOC3ecck9Su2U2Q1BWjyzSmKPL5tGO4KGSm5i10rJkOX/MHv1DDRF9X4
qaC7JOk9lkAbUKesO1xEbOxG7/kYfW+QM6HTbIP7mWTzt1RXWfRGbeU+sCjQhzOSFNnrybqTtJbc
aOF0VnaHPy7ZCEwJ9rnJvPqkVLFPEo+dobV/ZNVfiQnOE6IlIUu2MjfOcqPabfVom76Qxc9u/OX+
HySwAwyWPyofx/xNUBE3nnvpG+VLCd3dlEhVIz+fwvO05pNNo2RP0ZKgjFP3gAqdDYbi+nIgv7z8
NEOS0Uz7gzR717NgNRrgz1Hh7Xzx8rodMtkWbvVxl73Bmm6I9wawDTg+1zSzHVZQbYzItmcX341X
6pj6UH/TEG0uXR3AndhGV/5lttxQBNDVWVDTwXRESdTXvvFzcFiCuvxYUIGPeV8v2iqSNRxFP31X
X3lBPfcndsmbtDdvOjQqOT6oEdrx1+43RipKxVgf6H9O1cxOYUfTv2M2yIk5QgC8kKdtYUrHqCEV
R4WwXmIKUbx/p0cAXtttuQz0yXmJuki0lrtbiCd6J7RvSe1ctzR2zYGzvj2BqzbdMr570VaNfTOz
zQvz1zU0Ncp++TV5PqEMtIbBNrdDgMHqrXiD6DEv6DS+7y4bGYtQCTq4iL3TbVHgvbqMXtnETYDz
+RW8TYdqxEIhWKSRRPp7Na8W5WjWelnHbB7zawbGv8YQJwrgyVefkDCDynoeNP+llwQClc4mdL+T
DlmRwb6yhEYufmC2sX76UZ6UFohvHC+99UjnUd3jdTEqBuNFAaSYr+835CAMS0OMzGU7F2tDwrIR
g8dRL0k690o+D9ngYPmtM96QCtGOtdUZ2CmEnUKnepK0VpheFrF5y3n/uC9oGx5/qJs6Q+E6zztU
FeSFdV2LkWJ+BF8CFLoWAn3OQVttR7OhcOe2JhlSKXJp5SMvDHEVU9JYkaJnNMfrFJZm4kZl+X9P
KtfJluBaSuF6IIEjH5G78rWRIVHVjnRTrJNrL22ACDcbldGrcx6+43OMr9kMZ78PnQTUiYAobxOq
v10T5rlBLYec2e1J9jCIUX8IgIoIGgndpZHkuFuabgH1IdDiicN7/YqmX9EaZIXH/vJbnKOehxMx
8Ov7z0K9HV8NO19iNmxotGpL4/ZaHmP/+jzfz6Qxiksf9Vjsc8X6ZG8s0CmvOql3BBAC2oJbb+V9
gzoytnJ+i49CT2as5vxXBIsg3vfPVPS4Cub817awTUzy9PHfjcFh9G0OPUKtOKEqnFIpo6fQwzU6
zDqhzpEQf4mq2PzGxTas0m8P/+e/Ygpjn7uNn+sfbVIfZx3P/GU0jxdc1CSGM6S42ZX4XLBp0pgv
LXXMBI8Rr3N1z9f/ZFySYIuD2h8ifP0uqKAxxmP6TQe8DhlJa7IBVATqNSWUGyVpc5lZGSBauarr
iv5fI9G7zxQvLI85kgPxklgUKDWDfSoGQPMpq3HhZINK7W77RTM4KiwHjgBKz9rrUQayGbOBP6vc
st3+lehhh4zxVpm8jnBykBbn9xHv1upLTbh9b0EUDGt45GxPCztDDC59Z9hSvrHqRfAOzGW6nikL
+8n+xrPziE7wFbnpoJA+MMiBjkS8J83dhpp5fnzv2f8WuypdEEsKNd+BGviVWt3QOEfPjIY9TVKM
L5qaqdP0CRuQso456054ooC0yrPgpsxdj4fqi/rjO7/HE2Pj4+9FH9vCMeKXtZWcbyld2hhQTykw
AsdSGBxbGY/EFxpiWzai5IbCzwep4hZ2jJDFIxbezhQKyGQTctNzXIewlcnPYDXOma05OfWl41VH
w/gdFQXnKYCd+u7JoJkC2mN6srdeF9daqKFm2M4kjPiKer4IPF4/0JDxRFpnF/TFrJd4KjrfatkS
eKR2A2j+xvAXIH865+cd2aoU08IKYzZW/nMihG9IAe5bkvq18YTZ+2idM3WcspsKi9GtNqEJut+r
EniI8Pw6tANuk5NAAHoJ2/VnAji1jVONldmL3VFNn2eP4un3o56v8JVQCWANrnXRkrCRLCoNpL/H
AenLQuBv0G0I1bW8d31ody8vyhPbHeCyEbcdLnIQKBN075AuMCYMb4DdI1rOQLOBtE+W0hrRNVv9
kjUG2D4EvyWO46si2Cq+qaExGOhEAn0+dTK0Bq6t+TZ9ME0kcCPSMBy2wKF+mBcsznfqg57rnyGH
SexHUed/OA2kXKAcbNsxCX4iVIeSgPNqZ5bA6vWFIyTeYmc2Ex5Hdd08NQTK/ReZlcP1C2eGk2Vx
Qcqydj17N2HaYCVAcwtu2wf31mOVDss/vSt/DCNZ76hrXXss/Wz2Jb7yOt5jxEHIFiQy44vmVKu3
YXQrvGIasX5nR+qpZXz/tDP+BLA/fMLyJ8UImpVBUO1M3rxQpGVaPmhmnjuecTjA41+DGvR/yya9
ktJfk2NYzkg1PnPyiFqMFlBofAGBS6jMIfkb6NBnNygfHl1mlfzLTnKro9/4ZcNRHToy7yFcJ8hd
h3+ApX+Z4ys7siZXiqT9xLlqm3dytNoL4Anb8c4lMknVwrPEgqnXUT8TOokp8FxknztE25C4A9m3
qIPrr+xaNAebrwLhHCXDRgUNeufrqneP/pjldOr+QqTWoptNfeirWq5874fYMiMcqmGv/bd0icLq
MPV/+l9FuppMCr7hz9PvIlp/SmBlS/+96gP9KQbblcVZoCq3tT7lDGbmvz4DkSvJBqy12zxl9bmw
CM9ekVZuQeg+mF5UHygh3Ipa5EHF/8cWDrwJjwamGLxJCShJrvs4MAr6Nb7OYJIT0PCYd15uRMq0
ErdIuKQxWBE95m6xVJpVzqfM1aZLI/ugbbwT0D4DkNDzXB0EaRCW1JGsNVVlQnaUamlkwWc5XWib
aYhW8hCSSc9or8MzAlS9l6hCE5PK+82xBVIi+teYknzBUpUPpDRRSwOI0rnoiPOJ0OVAZgWNZtNJ
AawL8J9ndV55PhjckYUPa7eb5hD7QWFFRjr8U14ezaY3Ikaue4HKhksND6FKMJryHyKZ1dWkFuKx
TPNwhNNtXidgkQg59Ik00NiWM4uEha5EAGLTS/g043BDxbpiuWVRE435o9GWF6t4Z4n7RW9Bs09k
yTnFtHW8Fnbndf0Hdcs9ZGqNDOfdzxSSfYnXMIR1RkOnoEAzRdc15sdf9xIIKSe5LnUFtl0s1OS6
WxLJzk7p9QHDNtlxSdLmEd/53JHw9ZJmccutd7LtqO/CmXnT2/erbPEuCI+W8YafbhmT18XTi6xx
KJSl0RpeqM1f5azpk2mCjjjYchMruBPZp6rMSlAqVG8h3KvEXEtRcSsp8V+tpqF1MRRGIoprdoqZ
hZ8zmlJi+1XinZpmYEkaeNDXCecHWsJStcuCy+BxrPFwZkod63HQUtwQgYaoBR8wVLLVOEQd0dWD
QgDJ9LZ3b/xC7/gfAiFEH7799/OUWjzZv3BqJhBRHgiZgXTKAI1jsJLZe5ls4u7kpZCJLZYuAMFL
Sjz1EO06NqPet/YPJ1AMfdhcMU82Q4ijiQmxx/2hy01lcvicsGWdlLe12mR+qE+COHrG0uNcOoSz
NpSK48+varOzRw/rnmFF4bhkFybJyeoiRou7ttKMTe1h4pdb75BZtRbsqpywvfQnHSU6OJM/OVJi
04dO5ilCoeXI96mrSq+5ClgEd5nH7EDyGpAD8drn2Dj6lNZHgQm4MvJ048lIbZ0XnRictnk2WXbP
sBkW3n+nAZqIqZWrTrd4DEbPtLH8TZkV3urbRfrxr3Ym4auuov8wuC2DRmTbCkO3d/VqDNDM97Di
8qs/AlI0RdAx2f3zqPeg58hi9mRlBZ5E0FLQHMjL36VKXUq00PxpJYU05EtpQ6ipi9qtQW91qyoW
3m7yRWJMSfmi9ti6XhW2c95/Asi/PqngbxyfCKwNyIbSy7aGvzZK7kySipbViJkDTXf+7hupcr9P
MysE4ieR4SFpEbBcq+RaEiFAC+auGjzbM559DQ0M8CzXgTGv1A3J/zTbzFVuPB+QCU5xQ7yDgnU9
QZ4rnz/PgNF/WOuU2I4qi3/xct1N/6fUv15bqvmhFQhtSKDx/7aowFLNNmLfy3LgySQpJ+kCBL0a
IvoCpVNUdIAC4wM0yl9Eli62GCOM18+Bnz3Pil6i5evd8zisdNynr8KvKNBKvgTZO6Il9L4XphzZ
V1SyduovQ6pypuD9WcOUPoQFVpnJQ2U9dKk2l+PfwR3HvHxKl+MNu/8JDFjpQJ1LjeszR01HsMTx
Z0vEEQor2PCpRQYF0qGS24zSLeQcPWnDcuoGs2YStAEN24GQRNijVW+2CiXaYylLThbsAZgSYC/y
dFU5w2zqG+k/aPNrJi5rL/+qNno/tcC+O7S7aSi5xHj/beRicCT3IPwadQJ8vy4uDOPxCNzqDoF7
XGedMs6GwrRmwRf76BMILaYnoXXPUO9FmILk8mSv+hfC+I0PgzMK3S+LQ3gjLLqHmTKu+ObYb15F
+C2Avax8F4HrmEy6n64RWEMnroqwqWlzz4etpnntFc2F66oA859b+kmQxBh/kj2T4pcOtbu/BVLY
5e8zqf2Rc3ao57MUpe866l45tJNXmgUIhZ9J67B6LVtN8ST6salq2iUPqyvMxAxNlwXT2kXRStoy
cTyvp8naTGSBX7lBsxszXb4wVijhY8kAG1nCdMCFcShC+x+mLiygmtXUigbhxG3o58tbgmHlHTLa
JelNFZrTTn+vVclhqfbCr9FBwUFTX5iDcANahvri8KvtO83IC3iv0/L6oPWkUS5T21RWIa5H0IQN
mnTMUl55YKkDuMOyiBgaEmtSPX01P5ZcLNi5Q30QSQ1hrtez81mIi5MFwDogLetvrxo0ubd9vAfT
EvDC3KMp5x/hhIp0yOHC3zrSjLDpp7e9uVKwplpHmkTYNNw0raOL4UHa2u44yJgN7Gd5ZNhlYPQ5
GKYXv3GetGrBxkUGKWDfkMsb14EWyyC5NO7a+59gJ327jQhP6mFik0LfdnjyOIA9ImN+wSC3oq9M
DpLFaIM3/KloLszhh/JAXo/ydDF8C+Y2ZFEGQQ2l3Eeq7Wk36WRFI4HH0KDdSQMRv5//FgWbQqMS
DcYLl1ysgGo+JAV+ix4bRbhXpWPcTs2NdY9XYHJQdPPMy2y+GuM4k1mi1kY7A9QpQO+H7b2k7tMR
ZABnQEujqYvVfaJ+BP0C+/7fOaLqJ9Qi58nyoNlpJpaTUK5UGY4A9YnnLIHkoPrBAtdr5Myi0CJe
XCIN8bx5xL0okl61cLkm67ob+G0zals7+kulaA97UNHpDBM8UyO6AAaxNZQrqXYvfQkOVtsym80d
ZLFXiv9EVXhhh4Hx0zjz6lY7jdt4dZW38184Dz0W3CKTKO+wk/Ubs1BI++0o3lH8MrUKlb8W5sY5
tz2Xheca6PPu7w9p6gpaNVrF/+zQvc6hG1muTWFNy6n091UIRyxiX25R7hfKHBTt9m7ltqGb0QbQ
pe8HHUI5cT0sZfqnIH5i+uDIfKssxYnlwzFrRe+Pk5pqMJGgvAF8/I028NUpQTuzxszK9WR3wBuD
joyXGuzH2bq07WZrqaZUhRMuWuNZxRuWuyxkJvNv8+PlHJhyQ33FIYH+kM7Syak1CcmYz/Wv6d7O
xRQlu2n1OK1HY5nbDa5Dqfer6awFU7OMUQ14JSxH9OQ9247DAjNReROEUA0Zch8BBHZ2EGM+MgPw
nnlovrb5trrRGcA1pFXIdyEunImCjThoWJuzy74935XHuEvIIyE47+l8TNk/WKAwPAiadQBKsr90
hKsSVL+NCXHsaT27y6T0YlSA0PhlU3KuJg++X4fwhYY/yyOpkmwGRc6F2EHAJAaXxccjw/LNQvsu
+kqBscfN6WgB25mMMvnLP2rXf/peZjJ6xnNCGEK7nBVEVkrJ5/hFOvQ2V1QqbUOVH3UIuitsQ3Nq
FJSSWY8R/EbhetFvO0hFrGH4nIcRahErhQoeeRHoi5jBAI8Lpjsi3Y/hvIn4FKQ9aiXZBJYAjOHh
zbSajeC/taTei7W/wA7KchxM2V+E7xhY8AWh44EjWxpalXyhgJ3LbujHUGF6JnWXiZFZN6P+uGF/
e/v1vKZ7s/23h8t+D6CsDBDDPUUgZBsTbBY5nE0d4B3rLQVWRnbrMReaolOPLJUXMvk3k4jRRDL8
Z1m62qKNwgLh1EGH0XE/jMiV/tyXM30N5vt89eO/9gn1Bv8oqDkGxy5BiIkh1W9Ld0P3pMNL8tnJ
WI6BOPiJ6wpwHKrBI/ysBnLgwbnoN1gCCnaSZaC0k6maoEM0cQX5o0+y4QyKUG2ytmXUk37Wlq3n
V1yBIIrQBwf3oS+U/z15qCT6R/mpEb7IwsfBe9faTRXRq9CJXqTDAA4yAb9LcVLB/Pu5paN/lkVP
i6g+9fpcSBl2SsjKnKXxbCmzUJRfdUXLw1IEhFHr9ree+mOhFaDXI4ja5J/GrA9/JaLJxqZG6xMs
1DHZlGg1BjReJ2wFt5Vcs3HeqvHMwr47Y7JFNYgv8Xmw37JUWbRQkHEWzpHG8Bsu4w/JJi9Ip36a
vvSfpqwYzT0X/Z7G4tMo0gCTubn6LCUEV1oA4/bUku1+P9ZOO96aOlDapTHwpWrKTXsKVXZIilKC
e2BgcPEt4wGk6p9thgCJf2usG7dTv+hxb7JJ7CXjd7GOD7MCIm7HiUvYtLxxvp9pXHRm+HISj3zm
3HOvI9YyPRuJE0d6Gpr9iy5lt3t8DkPRztrUGf4H/7UMAUSIfwx9iuj1DmJsb9VBfhuQ6vQBiMOd
Tp8f/gMZXu1bkvOsjvs7y6kM6ogZshxgYOtPvjvIie9ZGT5ttAdpiY/8BlLDcrchycyayq9pq9Ba
SFOZlg8UtcPgI34fyeDPHcDtN/ZASc/338nmqSsawpKcBKsALTtQY2Yp9xBut7BaHrh64MgO6eRO
Yu0LZo4gw5wk/ju5zHkgrX6081YdMgMrdudiaHdYJkQssl7l5Rc4/nony6t7q31aOmpa6k7Y/LEO
SUqL5cKzLEHidgXPPWND21HVG94QU7ejWk3eNJyQVU2fk5GB4BrsZbeo08KGgRo/eu0m/u4cXFm5
CH3fgIsIzTZAHbcUG5T5802vD1jEJhQPgGI5nyqP7AcytU+Y4BsxpW9lGjylr0s/iAHPfyLXnAXY
gO78EaxZyVTpVjDfSvybHS+I7xgxypK9SlsWW2W+QPfX4LAIk3Vc5e8yuKGfsrmZED+9KP9Lzko8
65Dy+HT+6cXi+9CDDFVmpKE5caLPg9SoF8Tt+8TFl3oI5ZFGfJr15Bgib6YO6sr6t+WX7Wcogbmo
Pa2JjbYjGKDJTYGsz/2z25xA6CJJ6pclAH+sIzYw/U1rlEOILbinKOhiZfa+pi5UPdJfUFlcpVqB
oCxvcyHBGCuE3xWclawg23VTPpK+G/ojCIrEvRC3c2tU/ru+Bk5KWG8asSCDNBNk9+zJcZVoz7t8
Fezt2SuI7sfoEToLlsQje4eir2zy47nGZ7J/Vyn2aBMU3qtAmcVbRMEsAUjXdYjGpQEdJfOKSecD
8OHvR8ayImHBAAD6WadTnpvUUxaRh6EMpELrNrXg/Rpw5OutfuVpqmYm2XxBr4xg59sFl6/sWe9R
EskBtB5b6//UXujrjXcXoN3Bv5SHw3wy6WaGVH2et2DLnO4+auoU39sv4n1UucaQlVc0DPgC8ITT
/xtKAX7fBNQo50PlxA4u9fZLEjX8OWzfnI6CvCFLyhP4CQMcHylRO2zmti3HDaaZEkSsniEqHdjO
NIWwj03qZDX5yZAibXN/ZP3gufi+InGQm61VqWE8LzKS5hDJyO+kFo4BSo3LfIIdm0+UBdoHc7/T
cTwXMhryeNZ13GXx0E6RJVq9ywWtlvZrvAo/iW92IEfbHdY+gZB4vJJpjRQ6Nrv0ThJBcw+BaCiz
VcMuD3HZ88/idGvHz7fTQcFT7mfW7mzebAuA7EsWAyPoSU2FDF1oX4BXkADdl/licz1aMTA5lAMW
vJ4gDS9NLrFWwAmk1Kvx84LutvuNlxNwHtexPjHGfFOE6KFGAhygtlDcZGGo/D5mUrRH/8Z9iJ5r
aZqxCRavIOQRq3j0w7P0Mw2URg3MOwLyc8Sq1e3NzPZmUwzA0uOo7bPXY4wLyZ419KgBM2vInp28
gEA4fj4nBXvXGtnwd/Zj26sXUaYigeZhfT2vGJbUQMdJS1Lu/BUvSrbIIBESPQVmKCn2mfKA6Bdp
Z/MpavTxlKXGARzmia5bS4oF+bipoI6xGkCbDFWGnGDRgkg683kug20O0+oMc/5MRc7q4DJzQIB9
r7UVipdv8jY5mHUf5c+7Dw9YMQeFo8HODIOP3OswL5xQBXyliyTnQL6iGaliXOhykxGSJIegSsOG
fagWgyBCcoiT5KFfrwtgyHKvmps7K7qjSEC5S+22jJgChfaOQN3V6tkccTYfEXImgCbcZa/e8xIz
uYZb09hz4cYbRZQ0onVJg3niHXmHRdk4aAiJBw9zqE3qJA40W4IJfeWZD9YbxXckg/qYDNFWJjnj
yxfEHURZP2pCQD2U7sHDMDVG9jcOEocsjYpkE/LUJjpnGdBqrvGHpWGOSMI+Da7bhMkfWGGirUgC
PtvhapeK3wgDuY/JU3R1aZKcIn401NLp0gU9rYsd5o5yM7+G0rfXMmyfsweUTY6mcb9X0dXUvsuP
ymw65aOqKGelwuPiyTl15jvIF0Q2a/d5G2VXMQDdBQbBBTSJUoFLrZvK15u6ZAdm36/VpH905tOt
LQx5HSeObqV8wjbJvMfV4DQcW6R6LGGeIguyc5QsxdAH4jXEHFD10E0v1/VblEr5JGKTpRK/XK9e
QN6FE1UTumsa9UW+jsiwYOVEBljSFzYDft74wzORLBINXYIYMpMghdrFmUhBCyz+3+EfWbWN1Gkm
MDnJJXUIaiToVNOEWIzPp20Hv2n/VIwWT55ajHLMTajXuu4P1/IzBrtODrc5EwzdUGOI5adxrmsu
Ytdf4HzTviZzI1JflqYLzPaxJcxb6yzZ63n/6jBN70u7SIuWT/ZXUU10SSUU6AqclS91x2mgY8JN
1EiRtBhEFcdvT6pGjLI90yMnboEk7t6//VWo1qiyFFmIepzai73rQMOycIf+qIMYMhbqxoRROV/f
plPPHOI8svtrFFEu4v/RK+4Vbjxsl6CIMtM/dAeU8E+SQa8yg7cJ4VMzik/F5EahgJLoVWB/eelI
GD53A9xtADH3NLOJe6gxeD7828ggqtuQ4IQNopdEVE6luWJfwgAjodu0wklgRg0UbjMxpL0Ex1+b
4MBplL8fYSZYwg9TnAR9CBuIl1mAX1quM8i6a6VNA9SCGEFjaIhIUPC7m7mnlChFoQaPHr7Psqrg
tKe7ykOLFXkwubvbrL7gDkegUHYABWiObFrdhh/5LZrQKN8eCppSa4wTL7pn+QUq8FnbH11yGqcq
oZY5unRsORpvRV7rwVie8/dJthJ4Rm/moOQUbpNrT9Bzaoz23hsy2jzAenFjkWkcqehv5AyhMQ6h
2zJmmVnPy7mQi/++qGX2hiz2ddAWw41jY6BF8vkQKdcCdvV8zhskSiL9GbGGyOEYtxyKmfA1e6Jf
t7o8bPr7DAVe8KTkjXrn6hc4AVYdlZbMHpeOmrk2NZ7rVLm7tfbCiMT4mfH9Y5uPWs2vEq29CWyN
QijfrWQHR1sVKVz1sJzVVz21O6s12xGidOgPiMBdPh6JhlpIEHKeSrDjRkqOWydT1Rki9uDyCk5c
FMuh2xKcj196Lw189dI9d1hV6AECHLFMSTREO1hKliFqPA4dTL1QQLjSRkJ7ziSFuZCmAgwh78bw
Hxe8XEAIwCIwccH8S9pPhTM15fgK8CP/wp3Ur9U+rQjPyQAQFVkZcZJgZKt2CxDO7JzlRWWwcXUb
aQnVedCUOPIUjzBh5jj85ZNnt61aI/wCpW/LLbWqa0X1jsqgfO+IfEWK/2yvWxFQTcP8yK20VKiP
1/cwdREkYtaBWwWsMbbxdPmtxhmJ+7f3U1MwU90PJ4nZIP3tMZj9oJ486aHnkSk+sQk2+gxVVURJ
o+Hza1kUQrzIYllTg8ZEefBJp3huxqmKmdTVTrkoOnAHrvflmyzHU7rUI9h0po7TlH9qcfxsTYGk
fZ9JOXcGs2LhjX+qzccnEcyaTjm4qaVR4ZRmRTnxrqAg4HkQwA4nTVgjcXjb86tlIHy9a6Et5o2T
knWBakYREwESp4mjJ0L8kZdhSUc0zgrKX7Aw9m+xKsVYB6LqynZbP9jf6pnxs1WyTNb2V0FetmIF
UaWTeyfIK62juEBb2LatuWDa2v5IBqA3RkVm2XzkqL8A3B5JX4TVXrnyJTcazvkI+zdVZNsxbs73
FowFcEF6KEH9nqV5djg9EW8fgJRflcFd5kLDwIz74VdIjcH9lJIf+DcmNlJQBEPwuwZuM8EV+o7o
36VbFgg59aq1YIqj+NjCQdjNxo/caCmZCSOf9sMdYFsIGAyyaQ+YpHaQ0zOmaxdaTWGVyE9KmYwB
JFZaJXUztj55CIEiPK5t4ZPza9clfTUqxfWW05QjhlnLOGmSBNMrzBE8nscUqFwZCYh+/YwpPf5J
AHFjDAXTkgAn3VrDfnF/DYhs46gq2Iyeb1Etjg4ZXpja2QlLklC1/Uw+upUCEkjtsEE6UbWNrTWj
wSQi06T0FewOKW+/L0Hq6R9zBAz7WNKtrUVZasf1lJKqfgSY/EwTVgqV604oNO8dLeUhlxI88yBM
T/YxSfI2huWHhBIajJfqM8vji7ke1kBENiLs2nBgHXXMIO0Q6+uOdaqpLQYX5EnuD20X3Wk5EzH/
NCzsOrnEHF/S0XNvmwsvP/szMcR93+EF+cR2NP2SaGB0wne7BRy8imD3eivFlagihwAqTAoMuO+0
a1LXZW8Adj4x/Ep7FmBE8xcN3k8c2/dfF3HmJB4hcbhLTFdEAaoNO+Z2hSnYK9BVCK9YAFCuC1zT
QZeiJK5v2aS9JVZCU+dOnBHbREPHLr3RURdbfQ4t/Pq5cwEOj+ElxhNA9OHWHE1i8Zp7v4Pmeugo
rJ4DW6x7vF8IsX68B/kHxcbvSooVInXbLgJ4D7BXRyYhBHrjSLFhPww+1c2sATntmuhXBCjAQAE+
2FE/bluFy96KYX0cW3cF4xZfssVEQKoXeFJ+OqVfG+uhEo+pRcxn3n0Ns6RKOYFyQRDWu623KB+2
DXbkKF/uMyqTrPZt1MXWIUk4yPkbXd1GCAFsXc0b6pjYGB8NEl7OARM/qmIUN5s/98TQXwRG+Ko5
NljqaXR28IohRI63YigdNnjqsdXH8i9fFFGe/4byTbqMijUXtrkMAh2C6prCufBSJPIkCFwARWg2
iwEiDJXr+KmgSRJAXG12Xl4iA7gswlAjS46dGC8ChzPMkeMAqcGUmwLhXfLloQsupvFrE0yunStM
3d264ET2Ih06Vc4aakclsewj55zBNQPRKH7V5vsRKoHQNYuaj4U3ClB7iP4mySP7kGf9VnTTcDtI
eLyd54W80/P8BPUKQITrvPKvjgmAAaTt0xUKrCqtPlIhfgvGafBTC3rBDRcI//f3ABobTvq2MFEu
OfuXEwHXDR3VrCPDZKirPX4M0sdM7UvOCrZkv6iuRZIa8BOPTZmPPV1jnqBwSKinxbD2UPE9SPfe
LlHcc2JcACUn/nW1uHaZJ7O74PeGz7M91DkFsMfche9a6kMLTg/2GFj2AB32aU3FQwL1RkfgzHEQ
5Ef/uebaAMTQPjM3TlCkWzpdpwYM85GDz24534+sIu6cTQ1qJ7KebSAbaSWfv7bx8m0H1ijgCYSw
Uf5I6PfFYXET3A4EdfE2de/yDPuOsifmfOeOb1zGyjGwhiDZ3yQtamk44RijIyzApXORn5FiWfrB
BRqlI+BYizMUz/2l+TgV+TLcC82x+Z8BiLL1QysbDUjuUtQVHSVG/j6diHXnMuRfzfvdT9Vx+Eb8
cJ//DCOnszn5XFzaPJtWFYdhlCZMwMDlyhszziyTld0DoVewimaocmz4UZrYIqoZEBK6FddMRgwC
RDKjf5+kZ/HSRY1b5fLcoyPfdMfx7s6GQi/w4EPurYmXhSOxVqQRx3eqVoBdppQZOR9ljgbukORN
F+ZW7dJg+edFtlyszfnWd3vGUEOWlxGFVoZB34uUJ5deYkvwlJdOyoAJG38hzFaZT4RtUWxo7ZY+
4dYkvyZgJLYAv2aBfpvMcTqIMMlEJAgctV5cGm+Pgpb48wOEfyGZJVElnCDxbIvQkdB6xy7vSC2z
5FD/id8gwtFKKxvvwhq0EQ1Dbr05yPKK6AIK+ybJrNTv5f3zbev/T7u26ojFt9bUC8Hqgvcu7r9i
fw3nFFpVjINy78my4bT18Lk33sEnm/rLbumcmzpQwcz6uN0352Vd3i4Mwq3/2voF3h89v3W2bcVo
eo72WiltmT04j+5o1F8m3Azk7ev42eMkywYV2gOYOUvWGoXIQwUmXUQdsWhOLfmxynOUXwZ2JQiC
pvSIc9wgj2cJs0Y8+ETK/4ppQ3kSP7Eo0n48aiumNr1kvZFVKh1V8X1JrrveSQ4neDOm/M6IBMsi
uYjLG9Co/h/r0xLOmd8FNxQHLNBYRuj+ILud05VTCPiD+xV/mT1XUqdHBzFUvD3oYv5rHKMe+6zA
oilwNe54URtjemOgy1lmGQezgH6+tMzmpm5nrwSpSkKq3nZDNt0JIXIEhX3+q9CZONaDyyFrJ3ku
GHWFuVWFLQQUiM8G7pSPJEEN/tSSTKUnZ4CXduFVVvLfOf01sbNBxaDSDnecbJby48s2gpX+mTqx
3NPe2TwO7FCLPup16LIeS7DaA/h2cFLAkYmtNH03G+73/wcMmnw5/sZv62SiBywFwZ/wC5O2+Uw/
Ma/xTAMNPC3pnv8JQtWGhSsinSlRwT5jj92I3THpDbn5xO06UQKlwdKZ7o9tjFUhcOWvrcj6wl+W
NtsXpUAiLMGqH3BxZLoGCH/K2ANV2A8bpiQTBe9WYszwH6x/dm4NqJEH5VLH/R2RS/sxU++B1EqL
5g27/tCDFHn03Wt4fwttrso9+/X8YJGo/Zb5yUrSuPfnnYWUVhzzSQXgiXjUeVrvQ/hapxOySjpv
YBgRjhBiaumg1tbux7zMTbiHLZqokXOFFlq1BwCsVgcsdpOyYkcKtTask926Ua4q9D5+58mgiHq4
W19VHGsYhrWeUM6tXkRdO+ryLwfenroZKY8xKPfIYrvAenetOV8TaK4qxQ8WFNgrnRYiwh3OaR3G
t4H1pQF2Beoao3iDdyRdor8bwgXKo1e4ntW1mfVQJo5ah63itAi01rB2V92QZlMR/GHwCYpg+DL+
j8oIU1ThiAsS6/1Q4LGFU80aey2dYpt3aem9nwPqTPOHF10gdxC+z4Idy9zA2an10apQV33WEzNk
FqBi9YAzF3iDYilMx3Uxrc9Cx8Su5m9/Y3Vt4f+UT6OM3GluVGz6C4eRbp2hYKEAgIzGjRwZOJ9g
IBKSkb620J8rT/dE+8voq9ZnlH5ghJubKCmDWxBWTL1xat3HWFJUEJPLM1mj1tk4E07XhR1uF1wm
WUS6wj2uJlEscAZhU4vr1yRLGz7KrYim0vrsEfJdfqQlMkXEus5RLuItI6mpEmkwpEML01WSiR2i
zO76w/kSNaYvwIk615HfDryju82z7p+pvoV8W/7WCtASGSIeyLGf559aD8b20IbrkNQk+2mNc5h0
E3nUa01ZlEgA/uSl9A2Xdd1156fSRsVoK5ewlEd8kal5yKX92VKnXl2/uBX2Uh5T/+fSr6ZcahMN
gFCnEJWLCiIrH3LJpB8+Hd96zaH1zqEU9gPctFSb9blftWGZdeuu/yFSdsdga/383CVfxRw/P09d
nOXQHTqzv4/jcj9nYuLOLvLwxGad93IlXKF06y2NOt1TlhdfNOer2uM043kbFAPIKoetBkglFMf3
BNi4WvqVin1QSKQRNoSUstaBtvZn+nCTFN0TuvnzK5YkuFGBPjF8Q/O51tcFUzzfvjC2rxlzk4PU
A38cLMqcYorkHPmk02HZFifTDBJdWQY0STKDog1iFebOqyOYxYvMhqG/BTI/kBM/HkK/zvl2f01h
IBF0hDEav69gBr8NYQjxSETG7u/HKYdKuadUcf3wAnpAmcHIOkR2Uz0IWvGu61A/u8d8CcabQVla
NXyClWpMpx2WnbFhicdV/jg4IkKk39CVs+y0Uk/GYPA/YQBNx3uS3lEA14txdsEHv+CBqGugLKN9
BhdEMI6/azSHOqLjR003P1+Bolj2PiS68Vbh7ABQIv8ONYkMoMLv8EcrDJgSDBUU4kyWZ0nKSfU7
/F6hE9Ihr4rmb8UyhXXrI7+Y3J2YOw4i831m9ICXoNhILsWBjXDzvOi30JbHn3D95JdatPm/Ek5F
DyWooq4n+32U2znzaolCgwg1UBIqZUsCyisa1WlgdIxpsPtLZLmqNwgwkJ7afNlC1KBI7o8G0dy/
Q4St510/KyAhNP5TPDXLmGCxGhFd8AhOMfqeVdUSihRDrAZRs5xV+yJoWOzSdsAiP/zN0cjRsgew
AvkiHNA0kfRe6x2U7iZzo9kqn9SGyTqv1omXqaOoJEi7JVZ+6Vpr9nkU7/KyXBtYfKxOulqPV2x7
kTb5yBMhEdFHxAsAc7zcnNbXY6BiOgcks9xYtt4Cco3zTlxzVpmOvkoyMtHncC5aR29G9H9K3jIJ
wJj9JZQKmmRtu2zVXMWzz99PurVRLWS/v7otYLH4IvjpEgp5YTXzu3jX5xIH4P3O2SjcoUEngJhU
rep3OC285sr54WPQStXaF+QPj3lmwvC2Bk20HUy6r9lukc7vjbDismUphLPCKBQ37CEYhaX+imC0
NgG5+vxidjAJDcSsvR3p9YtLr4fvy73RdX0iRYnEcARRSfxiOff5pc8AN3y6drRrUxz0+r72yV9F
FDFcoS6bO7zDC+hI/pJmNxyCTru77lZ3ho5c5MvIz52Sx7nW9fgs+/CzgEk03KFkTSR1S8IWLfhV
GE6DUqUVdz815zCW5nCoFS5FkoFKHdilfQ6q/QDw7Go7KdBgPElGbaYwEEZCgXYGfJxU08z8pkzb
3pdGUs4Xj6GYBGEPjdefJ4NVbxYV7grNjWUzf2f5yZV42JUwfaN3tiKfUnoI4/RS7IB4q5Psq5gw
jkdvwUbmy2hqcDkX9CCVs8JHQdiR4FykD4fUu/uUygAMEcqlbrCAkDZdc3p3xQ7/iSn/OUjEEmmP
zyEvSdELgjVYqjky0Wacuy2tRPBnjA9jtzF1aEpheGI1XJHIVUHq2HsqjweQNuok2pfsJ7l4T8yR
WNC+RpP+lQygJJ5nz1ofuipZWODyXReYslUk+l/T4zXXmb8KgHPUorzdBa9HqZDS49koIuXZjoFc
Wo0jA1XdVvH1+Hnrkggydz4N+uWUllzFdd+TIFbpaXNki1IJR93Pj0xITVnzRhUEIZ/5BBfCK5Ng
CgNI3UOCKz65S0NVJlXns2yV72e50f68eyWPzmW78Ea9WTqnYn1EoE86LW7qWobqDcVi8bfCgTcj
lRj+GS6Wb+sROnD9WiX2mXQAX2pShUAZoOcMJqwi6vRlTQyDPn9tR037wooA4M1NJYYHRwdIEPRN
t6xcT91AC4Yp50Z+VQRmJN5Z6I+EjSwv6Xm8cu/GfBrF01jsxOYn4tQgGMis7aZFmgFNBtL/wSCp
DCP4WxEatuY4B6kjtohA4Qfj4bSWtPUKG1GNuvj5YeVwvcPFin7cnCJzShtPbskwOqxDz+b5+OAC
LXfWiFrX8EWRO1E1f5KuTpj6Cqs09a6G1ZPeKAG3fdHxzGTEmLwNpTL73O9CA3E81U/4fuXP4Cyi
AGZQZGcyWyVADgbBVcy5LYLNur6KFI9+NU2Rp9kvdFq+DEL9KRuz4uURMgINb3InzyNjzRXG60mx
KdggORDLsrRwFNURnxg0TxXPPpGiabPZRF8PPUnvWYQiMtUeZZjBjvRr1HDdT5HbV+mQu4f10L5g
LRjA2opsJaSh2VgnhT7NUysPHFsXBeRouh0s0tkPGqa/y4j3DSLLNAp2TyZ5jJYFlE8YsknZl+vI
o1BHIqI9B2V/IuQnl/+4Qzk5wV/zyLh4zat68qkhPFeG/xcrkpR2tBZ6EBUgUjl6zHvv1outDg0Y
Nr77MwwTEDXwgwF5FvnZgeNYjgWPd/OM1CHWEoRYYobhh//DIe1bxwvOwABa+1mz9waDh7N85tXW
tjYbvjaIUWev8pl+UUN13hdsawM8K23JFD4styCgMO7Ku3n+PLPLJhaXZFMU6diZkD6M9E0xEKwh
6HqXK3haAcq7sGW4ZwsTnwsTk+Tmv7RucDRmDKWzNQGnSMQnFfxPJ02AI/+nQ25OeO+YLx0gxX2C
YlMRiTJABdrH0vWkFKlTnvpaDOE2E/GiK57i/qrfdlzFst0HwzP0CQa/yRpWE3h/xiUDIA3DP/iB
7k6yT1qr+ZIUSPvFhqukWCP34MGo13048XAhJtCEJ9sW+/QIpgzNiqHSeV7EfeAw5G8JVK3oCEEa
16GzpamOW/8b5Ci4ONBxthjT2JXOY4lE2A6k0LZF5Ls/44Zc+VTvbI9NcMX23khLNDCEfk2J+4+h
HAb5XIRA34W+XwFyWBWt9AVjyW6NyFpNvKY8+oLpYWGAKVqgT2nx6e9BdVmyFXa5isv9DoGXgKY1
LDw8ctPaqdGmGITKipFgk6iYGqKUQp5KCnM46HpP4M7MxKqHhEv2gfItMN3NVQ4JrcWFn8mcvI+6
mIY9f7sRa0w+yOirE0gIbAM3RuN11FDaJ7UTFwgFhrJeKAdd7JrY48P/WR3jWSh0H0RswvrjR54B
2PUJFCTO2TJV6tnX4ey5xOtQgjfT7GeDKOk5UugyHsn9nq6dnAzWh6vAw/GS7yqe5hTuCu3f8JJH
jX/ErcLcMFs2T/h86w+1a173s8OS27ApIU/3HWeSmU3aB5wHuW0ybS/Ke7LepUCtefeyNVD6RmCH
a7wlYE5lo9p8H52tC3XjYr3N/I9PE+JUSnPY0vq1iQAYzYI6/YOHmfGAQNbIW9B3rh8YsjWBQLqa
dGE2Bl3n1i8yaly3i3sOaJxGh9Y1OzV3wJ9a2TFG+JdPjJe8+rtkei0eirRUPEc8DySpTsijpLjn
lWV5OMpUArfrKQAQcPzk3eqemO/BUpo8yaN36Fj30Xdd6Dms2oQtCrBsXWXxW13vQd/Kd0C+1biZ
eKaIyXHWvjch5gCe66ktlL57IJv7pMxe4HjwB6sHJ4JVnl+9KAFfRkaqOeGWScJKR4XHGcTQ5Yr3
CtS0i6s+i2ovQ66RvaKxaGKBRS6f4dMTywZ9sE1fyw2/+PAHTXGzto/L37nNb8If53QO7PLb0ULD
guce+Tj2yf+GCtOTq1SReomU8ue68lTkjQAL/fAzQ7kXLyJsmK7OCXu5apjCITeC2CBxY026rf0Y
jotmIUXZIRHtx44i2IRhMfsfgo0nLXeXjVrooxDj3IkhnzLnRr79vUbxgwpNHy2HJo0ovtdU/wJ4
XNUiZDTTel1rCTTzvEsypZKnPYFnEZYrzpzyfcRzqVcz/PEydnplSHNJ6BiIEHMLQwjTZCTM3E6z
3zDLwxZ5uxU+kdGFwt390eyXmEeaBmUE/ArzYd6n3fw/R9y1/tQ12jAkWA+ugusZwrBm1/8A8SPD
zEhy5zdz4p3spQdn+xMPa5zW431w6/Z4jYnVSDUp1xQ2CIRaTg6BBk8Ci58AdNnUt7r8SixuYvA4
q8avBb/KUAk1Jvxuy4kBzB02y6ndG5FuoJL1B9ZtYoU3dRV8tluklatcnArZjfDMfzvpAGGzTYCZ
Uh7Y/JwV8InLFy61TVdpSFbG1A56T2JcUuJw8N++sqH3VnEiuJ5phAF8s4m0iSIM5Md8A/Fa2ncX
V3oeMmIm/ODYTSbX2IJlPeGzc3YmRRZjBr9AfHPnL6yaKD35rpvsKOVCwWBjLFlU+9ADk1c4WrRD
PV2tlqWhAPDE7Mn9tZ0wvpWjkxssY0+gmf7s0ZrETxXVTQ6fr6OErmPum+e40gWeIkAu4UvvWhbg
KnQ6AOtW4NO7rBcVfGnBv67CGXUJAc9encpLVtKDM3yNCTRprl/A2nzeHRh+OuEjWc/WFITQivhu
0VFILGsJlEZQZh8AdY4OBhOzq9k7B4MyINh8T7FQebmfW9xRiWijBl8DCWj8hr7toaWEN2HpARCV
GCsu7H7Qz2cu+T8GB4TrcXz253hPrxBY4Ff33muVo9ZOWby0UTMZotfSwJfYu+EYcl0blSzq8MYy
SDfA/XUuZI9JbRD8CSYjUzsqvY6jzQtgbgkjH2wacnjqRN2mpgtgv1/7TuhW4FNt9FWz0LEiInEE
CT87d3sUciB7zfYP5vFXaa343RjXyHKanN12G4puwVKAtv+TnxilRgq9UoNmKuRqrdn45aDG/d0y
LO8xOUubEW9Ft5PF+PimpcHNpysAUzcyRKrP0tYbD72teJGc7Js7YExZacUXJg20SeWJq3aRqz9v
LYOhhIgAhx4YgMlPWYVI0Zs1tSfe/7LKVq5PYugho36Ux7Kjd6eRxHMFAe73jmLT3TVkgPQDzC5h
TwwfgTocPE6oY8PdzFsQs4jEkQWbfmWWL6UgRWOfPuseFx/ZU9mLlFrlv/gDgK+nQXR4OcsTUNL4
Hp7DhCQFZJVEOXHKQObk1U3DU0DBjO0osj3OzGDGVDXMPOteZNzBYBooTP8mSwYafljErMPGA6b3
0qZmir+0YuGusQQW0uHGurJaUdBQavQaxMWZ73kDArZvah9MkKMi0eGAsBk+KzIcZkGXN5EjU/DE
faeKjwEbugKO0slD04W6XNLYoEcvHwBgbRNEHF63abcWVC+Rzhkrj7rcJMJuQG8eGuI7nRa47zzk
gkUT7dRQgTsu3VVAnnShzbxWeuTlNrhxeSpXfdCfc4CNaweMNMr8S0ODVjG9vb7ZWp0Hep0y5ntf
eZSAgn2TetRpRmeUo7WUCJGhQJZBAtEY9B5M8UMR63QGTsFtDQ5QP3KXj+A5jpmwzQXl2if8FoHi
4EZ21kA2PinaY5NYwg56W5aVxLh15xxXyvYgRR+QYnMKy38qioKodU5N2MqvtJUfEzdcUJRxvP8i
Sa+awfBveQeoprwZpQTJ98A+1q1sIGav0nKY5cibpzFOi82PfzrP+eNdmZ5KYbFVBE+HSbPKoSsW
mU+pnQX5530B7BeXhhEMTyc87Y9LaCCjeCQftHl1JCOheGGVzkSdPVrKdn1nGxnIS2Xe5VuhgNU6
DI9pLHhvIRGHTNhumt9+xCap9fu+x/w+/wtVLCinWFAprhl//BQL9qZFUfnKbSNNjuZlE/178Mhp
7QqH38MarITc6n1Ie0Rx/kV1hujRj8PuIMe2Yv56a4kpJtW9IuQewASupXyLwdqFqyjmU2zvmOoV
LWj2PffpReSHO1R4Tlh7XeNzN2RH9J8f6JUPD7uBf1WvoV98G6z+HpkpCrhLRiiL4f0U91FDD8pW
I9s6WkfSgx468qSbCL+fgSgzL0Q5aleRWI4aIEfyusUFcJfWcTUZGy1LGW62ewJLyZl1iKSGlUze
GNnMNf4Jqk55aTuz4mjOn1ZWA5PlIX/gEaY0RCad1gS44yKGgejom914JKXdaJ4IIkLj/VJ03kRH
WDMDvwWL1PwYE9H7DtAxrdXELFxyR7k+6974Bs4yeXxVa7+LpYLEDudVHTbgHh8hxJ88091ZawmF
NiEMLtdciwsCMchTBwC+ABonVDw0MfXOKF8qfzp9AdxAcxD2WC2sIUHuCpEndpTE6VhFE27nkPLP
QVovFRSl+m5Erg1YcuNhErjTKuBsSDquxofyd3XeG+kYM2xxHA5LcEep4z1elAeMSd0AwCYfI0EK
qlznJR8thHS/EsCJ9NC9tkFJVCjgcWVEtl1ugaMBJudrYRdI2vnsohteJVajvVIDXmJ+zq6PwZsF
p2Tt/lCSJMwzN2sv20N9cYkDtu085C/n88ZXdh8ytxhSq+4Ie4KLUfCB7nYi8R7A27NJcDdtP0+U
1MLT7l51bkIB9XfpthoThaCDuYXBGaupA+q7x8cfcyLAF2QIR7P34nLCZT9PPJDxRMHuQNhUr6nY
a2oy3zUsvJg5Sbp4yyddZn80xgxfycHkc9urCBA0A7DaIHc44BZmD9qtp2I7hbOPlWx+9jhPwBKo
Ygz1gdPDuFlBa8IMjErO1ptjm7oey4sjSiiIcYQXl68c/ehF2p29fS8vXa4wGyNK8b/9p3lgeJuO
tXxD3Ff1IdRTngytGjBhjlAu0LeGi45TKEGipDmQfqWFvy3iBPmdZEkBtl4wZ5x7BdHptrdg537P
iw0tGq6ugXjHapfEFkkAx5rQaCv6NlWseX07uzIjR/09thiR9TMyLqOYegt4z+BmvJeVbAmS9pkT
/XwukWIDImLWN85qrIbGS6MUrqVjyK6694WrnqxQ7Zcj6SH67tUW/0XVVLJM2OqULI04cEqEocwa
zjVzEJIA4F3fEFESQS6K4sAidP5ht4Wp7DIexqfTQeV9ftmoOarA4b16wdjoJqI+cXgNgu19bD1U
RKoOJcvCJtmJXzP7SZUU3BzIkTCeJ5q0sIA9E1A3SGwr/7Xw44B7i262JMaNn+joVe+SKQJWXGg+
9ySbPtL6B+gAeqb3FxD7fsIPrRTGq+t8A54L2G+7n3YqqDl6lFMISnnpauemFE6H56JkI3Sw96hg
hIDWMWOHkJ4IP8K0Leswc1AyG6xykK24P6ZZlQ6+9/93AffJ6OBOH9f9R+hySRk9EyD83VLPy8J3
/cYc4jBR4nHMDrUQK3KTwLN7vU1/k4Ki2XbkBHDy3JGhJgdpsEjxla37BhglXvew6boQsbbb94z5
/pSJp+rl83LcS+yqwJufL74k7bNRR42rCSxZk3fWsaCCm+xnTPpewGPwIni5oojQQVJZZsfdt1+O
TVJOg/e5xMAc/cQIXFQYh+KzWLcH8i37k3QeyGIM+3hWiYNYtOSem3jmv3Rq7CJZBo+f6fvu8ZJ3
Gy6mWxTaOEpq5QK36V+j/25QcxbFWLgsY5BASUKau5d7uepklV34Mg68Wo8dbXvximzn9+TTmTiO
BkNzJJ7jelpt/F5kt3PCT2+BLRpUXM3xcft6YoCq9Y5ZK4g9/JRsJQBiJmdUtx0+a/+NYgx7h71k
bBm+zBloPhm01yZ8MvFsmXBejBozdZ9e4NVFpB0ze9UAGpblKVRzFZRhohKpWQj2cZvu8I0I02ek
IeMwJKKIOgNhWS5P88kFFfMC/xDfaiZ/1ShEVSIQCbG6QjTivVTElk/XEdo2oWfKFQxRZlioKUW+
KIiXfo9o0LwRQyAu9L29u6p9wiQEpfYVyibCsOae3DJoINDLagxfn3rKcWRCaCoJgPE6udTCaCmX
wjALkhGB81fn15cama4RpjJ3T0+c1VTkA8+ehrb+up1yTx5yp1WshpAlbK8ZckOfbhkBf1idnhT7
fcPxRraWZ1DKczotIFZHhpmfbSD5yV3bcF4h7rlEZvhvRYanRX1yuLoavmJTM6jQpb6u5myLQG3w
0USXFu59oU0vdH+07IVW2UkQXqljWydtLwNiM29k3xM3E8FoHun30KeyOBqSnUVX55LiGjhyjr31
ABzDtzihfdD8Zv8DLCn5tzxus2z+uh5Mtj0a4pHj3WQGj0vrqGLwlj9cf2biWectIHA+Qa7X2xSc
JbFY8UJZDl70rz7ARZfQjH01GA5DqgebEvekG5cyTGrxlnCsAJxydml52ePH8e1hJmTC9fH3p+g6
N0J9REfVzIIe9zEDN7EA+4tVJREQzGL9wzatzRso9l8CKmnyKfW1lazvZ0nROL169dgKblAnGeC6
l87uG4av2SfO/8/ZOcdoHITIihwAe2HuHQA6UvNomBNKb+2sZ3zXMY+UMapUxztdrMRCRqBAXhBw
wQYXdpDnqoys6COcfHsvMU4aqBjEOu6AUM8FoJcNlmAgBzkIHVOXIaD4GerX6xMYSKYkGWVVpO2p
8nw6C+yKj6LxsPSTrjunFTpfzBzzEX5X7XtWwNGYtGmvGTbd2UBQrLjbLHZBnK8XH5ZD3t2Sevmj
rDNcrZFjqx92JOHt8/m4mIlr0Dpk/GdCbmMHZ3l85BeDLDjCE+6wUgF1nr9ySBmPDfhBHUwn+r9n
KeO7arQp76zxmczeLjAsn825GYyQliH0pBnWi+pPtwx5r5c8xMvRIymh04K94JRIhn/FHbjBBJSK
kqTjFxFQQZL3wpQ2FYZRf3VwLvXbsBQpTuiPJXX9RXpxylv1zfMBtJQRUaRBkfdNBvbNySd0Xhxg
aMIqbp9FSsdVDI0ScJy6hJr7rv3H1eI+2Iz8Nl9kLxdJAZmsfOjxiNwhutmuK65LneXnAGg5Ue6x
f3jEjnjPA3kXBI6oJoV51HhNRGUDrGayQ4pULXL0qZtVir7rRfkPvH7lKPPcq30wJl6tCH9eRwDz
elfuVVSbtrhPQzmFFuQxL8C/DcOoSyEni4i3SPt7+p9i6FhGQUoC4mjyUHWTGe48AnNc9tQElkgs
2QCPHCC2eSa6Mj2xAPh8yMZreh4nV8uzNIaCwBUXj9MUaRMysNgtIcEttFbn0hRi6s8bvf770EAQ
T8SvQ72VsYvJWhfpcTYqTisL85HO+rSPTpDO5VsQkvctfW6MhT8thzCQ0aUxOkec2WGZbZ1l2a2C
yK/TeFaI8Rk6aQE0B8v10XV0MGhmSmp/gUTkxe5fsZNAs5WNoyyw3tIZiIQ7b4sFFCrAn/vOuIeY
CAexK0g9ch6+8hsFjOW9k4ch35wgxKOgpe6rVa7AJbANIjLvHdka0BpwAp2lwJDUaczn0G33bhJS
b++FOca6Cb51tchALh60713F9Hz1Ws510C3AhcSlON5H/T0s36aN8tHAsLKbEDrLVft3jN3Eovz6
M15MzVkVN7ZKOO6qMnB5AQ4ekuhwIFqr6plQRn2hUwVcAPHpLLRaAaS4NtHXkNKAn7NaJ13E5TO6
oPBNpr+PBHC2t1LNZ7sPJb/9OaH92aMpmSJ5Iqb1l0SJdZUxkUtnTP/h396MzpLAphkUame9v3Js
2rGoGQAncfivvkRHRTdXpSLypPnjJ/fPKTXq0K11/4NcmfPeDO11aWEmDJCtnnR/HHKfCXxpoEtM
WwCeA+mY2/XJLBoFr31QPopP/yp9S7bxPX0DPb8Bol7VJXlSuFHEkIMFX7Z27jRB1LmK+nnLFNI+
yA9vRYUwx3Ncqq70fAUyjWbfWFpvTq490s3wrP3nO6JF/DwB14gwLJUUaZMJQxZ3RH8w3o7p7vKj
xIsHchSuADjYUbT+rFlNLD2uc6bQrW7n2qCx3inz3m4zyW1oSv+tJeCajIJ4jppw7dL22VGjX2Yu
+RH+0tXTQI37eslRsW1bG/Y0D837HIsGSfNz40EnTvK6s58Kw+BrTcwazWNG5T4rJEANlHuzRZL3
rZ6vDX/e9qeQvAL/rkRPjhxP9UpeWUKLcd2/Ze53ITPIsgDBw0LE91QkLWfG9Jp+LbXKWcEP6WDY
fcx03PN29/Y+X/1TGSw4wYA0pm6LOv/rCrYKhzBE91cKp7FLgy0ZnqO6vRIFBs6k/lor3wFdLVWb
Vcg2Y9wAFZ9JxzGAR+AKPNAaBXhvsBjSLPeL1LS9vqYbGHnrdpWTRu2L7X2GtTsuJSSAJ1pXgLP6
yataGlAkFRyx5lLyRNo4Zd1bQgKLLrAAdYPMt+5mQt44jL5PQ9xTLzyGz7/L4A7kjeLCrNjf2PVv
DiMm3/qgX4Yn5edWFdSqMIJs6+LidgD5hdWvB+j+T+QIZzD1/7h72x2HTVbA9x+14GV/ONZUUiuu
8gXYVeVD8Deyz3XqWOzdu5LttV1e36S3e3qUDJhfhu20IB+KiClTOENKCB06pN2dHY7wbYoOpHbz
3xiJ9TfHcrFFF6KnXlLRUM9NggveWN5prjeSDx2nDFDb4SoozAIREBRJ2zN9jWrOKrHnZUoPTf++
r8ArkZfO3f1rINrVWOpqMDTLYCzpRYt2v4oU/YziPgXNdKDtiLd2HZ8/y/iQZghNRHmflvBueJkn
3Z+uC8+TVPcmGTBXWPVypY+gqLYmLFTThGMg1EHYDvc/mXHHQ8SL0MzSGtNgdDXCein0GuYDEP6U
AoZr6OAeWub1FanV4aPRUw9hrk27gPV3FDssivPij21EyyRBwXkoewcFaRUFQ7WqyfmVBh/QdHkM
qBYWwaD8fsczOUib7kekviVhU7Iu+jFbbRuh6bp/CmMidAQxbOQpm0CISWJfaUOPVhshZLKLasA7
LycvleMZ3Pij8m7nxOz4gl7mV60LIXw4KPYxqx3086VksDZOwDMHhQTe/exInG6O3Do5U2yh6GWA
SGQSxNJpL2sQOKmzM71iMRp6DyzW6m5xarKZ2tppsQ5ztObRGqN44FXsH3ZYuRFejnnnIrhBS74J
sdq3iUI/v8W/VKY3VwtfmWgSikDuz5ABO/SHSicpC+vUmzb933Yh9bEMrbITiTLf96gKzqU93TQq
ByLAoYueVxxqXvKpbj5b4I4wXKUM2tLteZL9/wHGbQJCxeTbnLSqX68ZLpkV75E/j2J4/wPz3ZKj
+DonJpsK5KE56Ojba3Bh9LxNKbiCuY370HuSzkNyeJnKuKA29USXafYGHNBBnDlN5rR1QDtHImW1
d2/d+q/Z5lJHJ4lJ15bIzrzyNFaLygjtVJgKajzOmtS6ZCYPz0vuDa6fN5Tb12M5ydlGhYwz43sy
1/0A85XH9KoXs0JdgGAlhg8cHetA0aHKDSt7bsie2r8pBbCh6ewW8LX8VwtXeIx6/D7N+V2QncZm
expn1C2B3q0DGwA56hv+aJfniFiYtlMnEg/SbojMAT2miGJ+5kQE9Wh1TF911F72L0NZuiWONppB
VOAacbsXUvCl9uURVXC7TJVEPBh6fZ1Fz0kCDbNBy+ANl7ryquo133KW4pshApvr0vF+K4TN6/zd
QAbIPMaqiW5yHZTG7QfE97ByRtgfyqZZGlQ6bO6efF8A88ZpcrLbSiiH4EmY0mOZZo1itAUqFIwS
JgCMtEPNCUf5IKC7kLeaj0Wyj9Cv6l4wWJEwZQASd0v0sByBh3qnYPA8QcCxYiqSqlACUmmF1EoF
LVgNkEHmpdCdZmAPmGbXmerGX7gBiSdvJxoUjntayc5LOlBtSYZ80Cxw8/YG/Yg8XkoEEP8XmUkQ
fbS93YIDY0xsUoRjTEXYxWQ2ubricQzKzy3sIT7vetNGA2POQJcQBTmz6x3XYH8v+b3bAnnjGN8m
0lOqQnH5GSleYJyjBPzgeHAL1DZf7eQbi4zohqr2K906E2dVmxcAHhiIS8fzOLyplqCqgB3NlKHc
+sdnF9YPGO5bGoDh8JKZFt4hbecevIfL7sgKN6Y/KQLdLkzEIHTMVKQ/5vPY97KyN9ujOpun0v3M
5qFkHn1LONcvdUdNxXD2BBqvA6nFlJKjcV8pWusbsmhzufw5kdy3XJey10n5BMneJMDZjgTQV9Lu
2yKuaPmtSUygoRxXBV+0vJZRrd0jaxNVwmCvCoBoMMLPhMwNdsLyN8lmnRYXUVC4rZR/mQDIgFhp
eTUvdIxGrqYZWTXZYUgfaXrbImEqnRVY3eAdEj9e9bFbwBNuy9k2l1pOMTVaFQwUZwdaTYdVQ2Ig
cpFl+h5D1LvMRG65UNS5xwScZ7odVVE5M0lo26JBIv4Zu0JTKYChy5dRbw44kteb+FWdTfLmHd5v
l2WP2t7EkdOJ2aSfA5n/+GXXULWfOGCuxlQJMQbr83aGnibliydLM6qFb9dkHJ76l3ZU3OzV15bw
aHmCNqzNTankIN+5T0f+5GHCcZCE5H/uvHz4R2hlAmXQUqWv3fAWC9qFiOtYkUdm7x5nTFfXGXJw
jJ1cZ9SatrfaKbNeRXYyXpCFpiMXmYs6TK9SKb5oiFZd/7IUCqXwB4NDpvt0YWL+99cUyVBIVT4H
MFKS0kSA7XsHnf4D7x+rKCNBHbahFwH7hyVytPNMMQjknblrMoxaD/Xcwx0BT823ci4pXm1andq5
nnakwazCbSxA7THxqw4O91e+hyOd13ltz8qGjakQYE/4n6RMz+t+C3W58MP6VbfGrjg1B+j6pbTc
keeRBWQxPnWi1CnR+qfvxU7a1hPDKPfymaq/kaxkRRvvOu1idnn79b0BKFwt57U7HExlij/9FRVp
oekWCwNYbvtdgqwP0zQPFt7ky0LVnQREkEFi5ALboqbWIJFN/HwuAhdrO+2d4qg8aBZYMkkTgUWI
QV0erjh6zPfqjzFcd5F94elV7VZ5DYtXqLxSkcfQL6z2Tyj+MFKcCjfvXFkXq0lg6JSF/5Xbl1uj
HsBdiE9d67SLUVLSwvIFZU08zilo/Nn2ZW+5oZWcc9VfR2OUq5LbdFFSLySV+71Nm6so91L2GvSx
tCcfsByOt/rOzm6Z1Zp5Z7dLOzUb4EDRy+kp/EnjEl/Ju8a2RbLYZSA4Qn4o6Qhq/KJHGhklhiok
p8nLlGhhF8+UCQnK1KbAi06H7DqfS57Zvj1ODczPTp0SRqXNip/xtIRgYD7bzLwkReePPaOyLxYB
DfcVs2v7WQbmmMO6IUhR++WYC4ZmO7LW0yNtrZuRi81rBdhyBC/ZNARd8De+knTa59WH467h6v17
d+g5F+4R4qr5AqEfBnk02olla6KY14CC9y+1/KFQun/yxp27Ib08So0ZtwDpZK1IonZzLZagdQXf
ZP/7hizHcGRHWOQ0lN+RXGERfEKReLpeYQmi+tPdDaPE8MD8DMOmrUQXb3w0B49u8Y0wYzsfN94z
st+NDf0ORQa58Jwgy8ZmvG3T5TuVFeF/btcg0atGHnQ8RiftQia6GTfttfUAXkKvV8J9LBZLO+4g
3jo2y4SKQvtbl/ZMQk6tWhVG7/QSVuGouecL6EHgkwR3PZmeMYCPB/gGKq8iRBREDnlEmwyMUz8A
nlzD/VBuUQI6eMg7QggHnXSORAvqtka700nu9+AwhnXGKIeiOOTP5CVOWN4v2XIhdeYsvbAR88n4
OU5/rm+CVASUhoA5ctJTiFwEoeYD1wVM4SGYZTqvsLeaciwinWPp0AEptQnV8mw1BRoku2rHgq4B
1Xc5IFer3XnxLpgBXKS70RG2/WcDmMDRRDdCfTX3yntj/JCq4Ji0i8UbQL0gG5CPe5NoBoLVtKLl
YbrEfm7ai4I2HCa8Jml4ljIkMijB3iCXhNSFZIu9qHqnG8MPlqL6LoXZz8lbU5sjaE4oJKQp/Oen
+9p04ffhl2N6yd31T94ySfpmkcqSH4QsNHxkpQiKVjPAMY3+NiXHdOT2XD18bUt+t7pOZKPK+3uZ
/DNzMkrwnuanyefZvTGsi0kxYf0aFWzQBsp8G1SvE3tRa/0uAuMpiKMZGRz5yyG3N8GvqRofhgVX
MV1jFhUPJaqarEQbJJ+Nlfr2+eIw10ma24a21piQP5isYt1VI7ys21sPOu3b3ePZApfL4Ljq2V0R
U69Y7BFsOri/iZfU06oOETqy7gYi0zKHgFMCUOQFDQN5Fr+VFiD+/aIZwNOcXziapoGNwxFS7OV2
gp2G/OxhFnx3+TUkh0GKXpYdx6W8kzVuSWMkFw+i74LcZMZipVFbWCNlsW5sXlBaltuK21cKnHbE
IXZhxYZVPTETbujbAOsb69VHPJOW8XG22CgecjiaLLJuJvD/baGvohipJi72WL012Am4PQNJtjbd
qqzyFqGGzqSbDlVEyCVJ++vv2iGJ7dCZ96yx2zP832TJsGcvLJ05faKVvzE63S09fazO/SqAzZAC
U+MI4cHdMs8PKOPvYDKK3GXZ53GaX4ZQP+R2MEgBeV9NaMw8CYijAAN+VI62SWoYunyhftFr/li1
iGgigVxv2t0+PUFZOFdlwQK7kz7JCUJijiqSY9Qjb5STwxHXyrOYkdEXFjx7dRjxhDgRxK/c4/w+
gHWfmusfMN4He9T6C2hPuUo2BH3Y2EulxTy7xqd8vrzshn1D1mLoh05cYDEcTalLVWP8Bd1wrMPK
Fr5Xqkt6LPAmhO86nsM8+onVeFVJ2QlAMg3rte3WEzVL+Mugy0k5zoYrDkLyhziresCxm1s3y+wQ
xhmIYt1mKq5iF0z3Bj/1F43RsdwY4C4qwQjcValpbBm09qQLU7IfuEJ64dAKPMENcwYzJ9B0Z4FY
5YpsM7RP0JwiFFu0sX3pkbLrGWEdwMxgxDJyeDjoAl7xh0+BNItwXFS9ZtNrlC2qqcwsTpnQYNFQ
GhUJv5WZ2Ie0Zq34UjBXRS9UiJwwN+tvOz1pAsX2XbXU18nVaJhLHMXwV8f0SnFkBCsvACc5wotb
7XrEtfFNwGjfwmh5LnboILSl0oyi99eZyxYOYrxXKS/xnSXEXiY1lX09IgfDUvZiHrXM4d20cknz
+4EoFebsC4cQsXVNqa4KeZme21iLZBtk43fFApdcYTB69jMfAF7SdR4VeMbrPxlMIstYMfzwDEF0
ReVgTT/IvR4epJh7pj+3NioheKvAEPajOcmLJS+0SpWem06GempzJ3LRT6KAWUEea2NKhfbPtXpF
+9RFuI3CvbffFqnkU0Sr1Bmxhn8qnyhwluj5uwWg4E3wEze9ZXxOmNGi+emtvO3g0fgqq0RBef4u
WzcoXAlTwG0i7eYHESraUGW7SitzCIpgtqdCNzCayg68a93mEJdZaod2pLIL5ebQFCSKw5DAOSs7
W3UrzTZ8isuX0/YWc9u5c8M7sZaymQbkUvtHyoer4CMSVcvWts5H37bJJSXLg+nJ9Z4bvMDq83Lk
W1+WH5xUWwhvjRV14MGHiQ2Xci5Vvr9N3dZmP8dRSybKWYcqNysqgqQXl1Y0G2wS+9+hH1UP2O42
+YNFFPd5mce3nk6ZUR8WHSPMavznGdO2k1k5adWSUuj0ek9MhWgX/YNwEUEIfQiNJa2T8SfUCEHe
PbY3iksyoE6/Xkarcl5QUoCqZKHPVwmEjY3CIvDQ0qZhALcbBTA5RnLi9It22wGb3/LuOoJODQNg
q18UgHfWY3K9gWU/++pR+EoCzAtwiw2ukDAQRfOoV6vRxx373V++XqV8y7CKA5yF2MwFgIZZIrUf
4rqwRZa79mg7FQFEoFJaZxYotZgq41p8ixQGA9gfgyXV5aHXICTzRPeELsYGVyi9++ra2vktBxaT
w3GIw1E719XRHe4IC2WX2X584E98rm7e7gGMkfMxujqjK0mIDJj3jQG5DTMhGjSd2GdhkyLBpI6A
oYwDA6DfTs+EV7eJeT/NufdERTAVa5ayzzrcLQYEXpSecCNRqbCBh3Le/IqjlzXHXirjaskEwJqF
6+QskFL3AvoeXA8Z27Pfsn59G2tmt6jjoUvjIef4lUHc+zU1LCez3WBQsQ7ykewsLYZ0ARGLuz19
Ecfl8MYUqKuWN4BqKZXpq3ZhbzolaT/d8s3SnEQ74O+IGgWNGdugizTb+KAxq/X7EnDj3+/+OZYc
qi1TVo9125q4NL5XuUwva2kSCqOLxPBYevGH9tH6YDiMHzh+3WfVQfic7lZlbOwLxImM5asCm+R1
nWW3ANGMOScq3CitIR3Y+5BsxkdggN9/lB3wXru3IiFl5PLqZeBx6tj3gTvIQXwkrTdoxQEAIUCy
SE3uGfHvnIqmRDNPHpmOq6UkjQiURYohqbxdVya0WB+0GLagalwNcXlt06jpnbRZAXr29sOpIdMr
mSZp8djSAMsawCo29AxXN38//DVv67JIMaiM8YrngdARGf6C4cjI0cYwCP/QVfmBdlVnuRCCy/MI
WJwYBDx3bs7Ms6DUpZYxZXSOw1Rg0Wn4bKLemQDrZEdQwiHgQBPVa0/9dXDSY6srjylkWcx4ko3T
G4gUgeL6bapOSDeK1XWo747eZsi6SG/mA+tCViirvNkTCRPIL5QZxlrGF/VqC4HSgaGCTWOQco2W
DUNiZcnLFQmwlig2ykiMQVuK1Fawzd5t/IkcYy5o1A3aIqu0kNVlONf0lagYqKMEo8TY2tEGRldD
tsHGXpYTIkcTPRw/GjFNvAq4uWYGOVu4SfwZDC3/RLARjOq2m08Zks3vOT/NlAv5MlhPOhUQkHIZ
V8uv6Pg8pLl/EoqOPku9o8YzgV5qn7I3AV4mk29GA0+a3gtOgX0YQaUNgJxajzDocVut55R67r7o
CFaUzLDzvHSoPOebcSfVRqj2HtpMcai8S4fhrPFza8AbHWwpXw0dhPwGJAmpsmQbTqDX0/DjrWtf
D3RRm9IWKfDuponTiGhnjIuZfRgT4qpliW9mcirGmacMhYQajr0dLZQNnU/q8h1r6JoCcAeFzC8u
FXeAb5/OKQJAzNGS9rf17P/OeBP2pSVv5BEV+gKMA6wcZS5u4TGxJ8ThciIznxHRsc8Q6RCk0v1e
uMlTdP1AXfbNjMn9v5wGFXd51LAsLL2XrA283dpEqxqmMd/prTzrsrnkahqkLwO/QUchZ3vuFw3f
JpeULXDu9VYKr7VqFXOMyBQXKTOmVTDFfFuTumqiiCId/uDi/P+dxoyGmgE9/VdAHT6iIZiTeMtp
jR/gQttGzPdpeloMX7MDU73Rbt54kgGMTlLR5T3blcv+AXuRfRdGPMpjL2WrroN8J9wouOVSuwiP
0fWDnBbbceET7rwyVHebsKy5WMjXwY3xadDxjq2EoJYt6n2dMrSnAm5AF84XFD0PqN3/ZFyO07zv
VR2mff99Jv+jtSK6YovM8Zw3vyb6W03cSNWPmEscLSSP6TriwuovO1Riyu4uXMu47I7q5sUZ1m1x
dES9YBWnuLcrsQ3jGDqMmomwXDIKjD+bVy1xMIXQ/8kEY4YBFft/P6ZL5a36Ra+zS2wdm2Z3wV6O
LctRLNc8SZ+yiUxYj0Ml+YLJoAEU2LsybpPMnM5r7g6aWs+V9TxB3HaPMtkgPN4nd+Gj5bgrnloK
tbuaD3h+jjCZDIz3ezgTxYkRoIInUnBsqJzrpcwtG7xwl2PXOrIHOrdwgVzU6uoNdBS3dg6tk+xa
rTExMdEcaMLl5dEdCIwGXPfQv7hieuoRmh6yceP/xLiend4L4xTU1YoNNgfA6zZYQ0oZRz9svzDB
AF6fDjzNiJhLWSeRcsG4iz2kBDm9N4+06gvp2+wP8++4T++4RPgpKGdlaHKP8XOYQjqFPZpW/PVB
iXg4zk/auxmM9bogkLt5xwYQql6+/d6UFeDIPm0Fc8T2sXG735nUOkOBtOj+SdCQVRrG27hiloBe
Gk78dC/4dKwP1JYL99EwEPKZanYc3jtL6IdzdGHjZzM5Es6TbfoEs/zh94HIZNRs1wb6E3lo257C
1GyHpabz6poPIBkjwQtJ3wkEt6XSTSPhpYb7ta1drud57VBJkBJnkVZPS0gqgo9pqbvXwE+oVjGg
cBrdEmabgT2Im20SjDh668eqDXt/uNARCn5ui5vSM6zLLps1F3jWeMFa+iRDn2ZyHZlYC+RsC4yo
Q9Ti4wsUj6+rc8nBrs9JfhDAG6vw09O2sSj6HARC7xf/fX/F3NMT1Fo2Du67bDoUG5jxeFTJcm0F
/5S+KanTXMRvjrpk0lu/DMWYqR7iTp4ieOeBC1cwQTg4jiuhlCtOgWrF5k9yejRdHwcviBghhxyy
h7BqGHkP8h0+/lL2ws1G32KZvTAzsvR+NIsBbWZrKKoTldPUZzwYIFFDX6QB/9STY5Zo1SZjZnX5
BBkv7wTi23s1YY4T4E5k3yxl7IcKtbAFMj8buEY13Fz6aR70Ppw5JnvZZGgM8wRjQwwbuYWc6iGH
JrF6b7bLZuYwUSDtgqBEu/VIiY+w1K4Sh8hpfFt3LUmA3fBpgvmVJg/hK3Dav9Jlu/aR8SdHjA/W
6YN/RU+P25Ng0aRWKxAbcYT/A8s81Mq3PYLQJgc96bWTfxE9Nw1ZDjTf6DdcFLculd2y1EpoZfPy
1r0fnvWGgFVIzBBS5aR88efiAFJfRCrQNwPQoLyhh84IBTPUVmesXQzNFRRNynnVHLkeTnQhvOlN
6ZR8Zwh4EIvNpYfImrNq5pJnCHZOet3wfHsw16v5+5qMRp9TLXDom+wX5dn6ksX/eUXqzsxEi64A
2Ao3iD3u7PJ9zfINOuW74ZIdViSCa6sM+3AQZ5whUCQ1S12duQA36tNhyXMBsA2hMagR6qW3WuAR
79of5V0PIO4ZTMYAW7dzkQO8SMdGJBsljjrqEC6jM/rd38oPTACosjWNA3slWbU0AwosvFSb6bW9
XeVQvuGogWA4MoGj4zmXVrL98jHwU+eCH352uwyxYeLlOynu4Pij3mfFAZUXP+X3Ah9HMGcfzoTe
G9+fboe2DNoieQiXLAicsmppLxe/0B66y3bNPp+JW5aYWRnZBzYRJXpgkey19dNO8J9x6LlFYuhI
+4YOtIb3pTVcUS1Pq9VYxVI/l/ErPN+fzcn5oywqgqMytypOOJhNvV3s37lnmoRm6usspHPim0s2
jOfE6Uzqz0lBG/43Ok+CXx0yGc3EV+hrrGrAAavTxO+CeAHgLIpXXGx5x1IhueqvnT7omKVF+m5l
UBnGUGaQV2aNLQHm5A0iDKFOb8h9Bi4tDQ7ozZS1vG0cfu2SQpsND0YKFfLO26X8rjWXQZ1jyN5g
teJAq4Z6+YwcfdD378olU1TlEo56LeRo7WC8TIFk8WtPPoAjPYnEqVIhI1xAWFdHLoROXiAb8sJF
IHrmkFEwup6+mwxLRjnK27h62SnflT6Cary4OLz7BT8W5RsM9mFT+oD00ZyO12PRmFeTEBN43RkZ
SPCIqnYavo39Qa/SwnUPvnvHKSDfFeE+6E6fiN30yz6MbyDSqeb4y4kCaDARg9IMsUuinfWOi0vm
wz986rPqTNMPW/suaN+lI49DEAEpqNnrPTfeaSnMJ0cS9vIf4R4TiXxWi+gjHtdt/rKkD45Ginep
uTqvHkyS1A5Z6kXpF9nt4sV/XvYGaUnL3J/UVTjqFn6luGpDKSvy1Lfx7nSTyu0L03WZs3n2pHsc
+WHtRGf5wsvv6wSQ+coOoihDBLw8WL0wZgqDgcq0ehABOAjZaSOWvSXe7z3vajFZI/AYR6TbYki2
u0IxciNAHM/j4JDJ7iA1CRmg8OSW7SxVknVJTuzJRs8gkxH16eD0b4yeYEAT+V+n+clOCr1pKXKO
pcSoYU5ySYyoNGaNSPQJ5nEVoJufGQZOihbS/F0GolKVMAbzBKtCidG3CGbOqzZM45ABnjr5OZKc
HaQsF6UclLps7oOxtD6ld6sifv41sYnyYBzgwuaK+Qv1a8dhi7FUqkSbhYpa0XAnbfDLJICNmzyK
+a4Yic6GoXFJ3W8AYD64OhL8UntA9CP7MBWMTGP1cymP2BFGOtPTwjcpwlDUwjcJlFCMTqN7DqCH
rITVW2zrlvR2iCIWWCGICuwBeZ9EY5vimgILycVVr1bEe5fVJwy+h9IwTWr2Sc0jjCIMLwgZeNEG
FvuL72SpB3j6PTlqovMh+meU9UHsf/HkySDknIhhvfshr9jk4AkYH209skXEYyCi7lDYeJEjsYJ9
e6MfPDj6AIIE7XiBVLIYD1VC3V+H3ZQQBQkfCxP+UfbxIguVNGZNEvipEQwCinS7X2o3e/+spac8
gihJcan2t+pxiaSRtXCIE4/Mxkv4dRfREmRMpVXZ+BxQnqCxgwQYX5Q0fLR1WufElITPPGOaKkdC
8bAKd+sNqBQXtyxSZxxh+0ADx6IbvK/o0ebf+tY7UnqHDQ7EDSFrcjN8MyMfCOrhYBQ7hbah7R37
Exg3q8RZxL39EMdURxdk+NV/hTBGwiMIfAf4VFUP97bv375TpKx76NG9uRe7bag7yeZCrCi2h+QM
vGAoN85o/WzeYld7dPsKcvWVQssSRjYheT7jElFU37e9FgQCjYwuwb54CzmMwR1AUJZaAzlDm9g9
BRvLpobuOhqkNu6mNMxWA/bk+knVYGjm2qOWtu/YOqhq7MhSoO9nXYJgjj2q1LhTJ0lPYpawiGpX
gvoi8fjJElhumgY2NPjgBL98oM3a5nxxMCSjz65lDwMWDKr+N0FFZs2qOa1fqIUwWHdS4+Gq+k6R
zY0E/jpwWom0LsLabTbdPVp2G/n4DJ+3jvl43D8G/ipPE8xGoGqywrp12PWo7j/xUn0pIVY4tsLw
yxXGvSpcOWUSt91KJ2bhoxp+YYoO/gE5NliSYb/lRiDi8ChIdy/cd4dDLRiZ/+QHiuQjS1zrhsoT
mSwCmTEJZdR3V2O9uduxXPAEiFMPReLDcy5n/hK4bHT7w4laO97yFxgaAfPSLN1GjerhqBt3fJcs
RLZM1d5hwvJZgeoo1CFEQN4Jsfsdr0BP2tYUatSLc6HRXAKS0G9RsGNBolRY5yAB6LeV+E7JiNUy
d+tb1CecMtNoaOjVFp+hW2Dt74QMYr21yuI/ogusU7epZuMUqbOFAiMJT/78L3nfWhSleSOkd6bw
LGjZpGJQMIOtlOsdnLBr4re3MJRtah5oeKiUeV2BdKvfSca2yfiqHYFFyBY8z6Dsl3/1dCOrqgMK
7IpY5zcdFAdhDZhZbukoFW3FKIN4eoBJaNxDvNN5HuQ5FZG6x17ArEgZhjwj2jW/icRBbnm0Q/Wt
m+KK5ZOzhUtYL6UK7ZVKdsxPLTwBjujx6CXPaQvb4dk6QK1tmYXxxsgB7usTtukf5gXXQq17xMbW
CTVxDvGb22jOeTRhE5Mwak46iqED0fnYGTxfps3ndNFS2+txZePK+K/XVr+O4Ay8ywFHdDgfLzd1
bMX4Vdoz97KPzWB2pVRumeMJCYbPU6kxHZMxwatW4ADkUNxffMjj9h9Dviowd9jEUn2eb4cw6Gsw
nCS/s8iJRFior0eC7nLA+XjEvZFWMVBUlhrAIdr2TR/bdZ+WKiBRGz3qS3uNta+6HgG/idK0dxZ3
o2njQkbd8m0bSN8yzqvFmJZQdyZyYAzEJWaf3rUv1PWjIwOP5f2t3mSyeBdy7yRTDzTKC8j/gpfq
r2H1NQCDnKXDx1FCZ6iU7F76lcu1dJQDy9IQa85WRvQ2xqvkKDdpsjDVzcd2JYxmL7MIXtj9r5e3
6JlufsmzvSvJI/PRUE460ML8uIiAv3f76w7amA6SSkZ4Xc1VIdE/1SQx8f5rbOHUZDW5UaHF6jLs
GMqmNTvgndpXn//m8wu2JGxtUIdhtNYlzBKriio6pX9W8pb2c1pSGdUrZJyHq/iTVdEHG2AkTNE9
xB/lko0mtbbkMHobZceo04suASIpj6I2qumxpV5pTC4IzqIkPS3BiTpCFHn4fmtB1NKNAV/62xqx
Hyd5HzxXctq3gdDoPo2gk2Qc//+gbaB9QedE11SCdJDg0G4TlfHiFcD2y1hdYbiu6AGXXGz3nFXC
oEvPNTqJ5oyB2yuD2kkxqV8sv4qHe6rWgztSVmbKk45uJg6PA0QoHVm3GgzwsIHC06hti6YXC7T+
e052mtTssFVIvJQ0pe+PG0Sqy3VjYfjT401xBT7JZjnTKXKNFMPwnRKrKvtfTyFD4t7r5IhaYlSF
P9DpM7vBSoaYgwZnfC/Nu/c+Y+j08XAgONRxyvtaOvmy/kkHwlF98VO+SC3LRIpBa9xv28u3nrQT
oIXRYtwx5/QuGKNWO45AvNe5lp0rdp+AuEb0RgPvf+t3SdYGcn1Y0TvRrhAt+WsX5AYyewchFInp
xbBzinVX5bhzEeCo744LGzqV77YXOSl/WA5RbMly92jJUySzIXLpf6WVSlYTHvVKV+Tx12cnQ9sp
9aaON+h+XqwuqBKf8LvjhdHMI31hH/BAbS6RiLy6Gc2C2uj/Ctt96U+304a8MtwojwKYDDnJQdBr
w6gEx2JU/WKDcSb201s0hxr+0fUtDmXyQqVfTHOQ+Ed7xsu/fg29kMtDAq44DtxEBrwlh9iNbJo9
eEoAwjUFbhjh6MilU53xryzLjzaTIBCjpvYmqZnpBc9+yuCaamFN8EpK9ch845RWfOgazVzV4/8B
LglNvye7b/vL8ybY6Jl9v6l3BID6swPvvcgiFQci/k4NixG8K+zJbdjU8nkoNrsT5AcVYy1SNsaG
qhNusCDgvsGuOVeAQZ68BuaV1ECfkjBqzsSQzfcF8DJ3Fs0NZLp6wi4UAAHIAXbdqwmSUPgZPJR/
ukB/9oNtE7PwfPnw+Fu5nyOlfUypIwdv2On97vvetMeA1V2hJIsj9s1A8skYtYJPm69h/ufB17VC
j8EWoR8kAfNUeDXNwmJUL9y847SlmgqEqj68QCKBlKx+I8L6CdHYiF465UrDkJlCzMD2esVOYlRh
BNfk5Q9r17f/MjvksodwbylwmJDF/pcn4a1VAQ1Soo9vGSKq2yD+TwLDbD5Nd5GqtbReAL3M7XVa
dQSUoyU1W33qSVWKv9KLAyfxk0OCPNrQ96iZXe7xaSC2gHUPcRjwYR6IdgCOimyaZs3BvYzSlMaT
S7+caWD+nLk+EtcjeHMBotiBEbeU88ypHHklIPQpD026inS2bkxY+YL/UV0lSGj2cNwh+WBDE9Q2
dU9+vlLK3e2G6/dBXJzav4/+VrZf/hVZ392T2zztut0eTRF7za+ncYg1y0VKT53k8Bw7+YpFik6j
1+k0zO6PZozK3DPn88raa+Rcluw9PmDUrc754iU9TMVYI+kKO5iEqIaGlNd2mul52gcilp+uVexk
Gw0AI3VTWv2CpDxLWiXHhSFVphYKbC5pbXwH7b7tq1XRcTdvFxdSSf0K0Qe9eIu5fme+VO6nj4Lh
zOhBTmB25cbvltkT401kjZFXYbsu1X65WG9AEQwQ4qVJSAROzzbtu1i+ep8jjVgkWGdGq/J89Whu
3hC1ADAsSfeCOVgoQtyfC9Be/6+HMAg60V4RpxazmaEN70Yc820lXOjDrxx5mz1cmsC2M9HrXdWj
pKyiiWpQ7dQ4x9kQvtHdbBzn7rS0zYI0fGueDV13zE0DsluWAOO1COEkhvNVQ3tFsWdLQ4ds7xV6
EIXJ5haaV8EXEVH1lvSdJm55aSrBoBfhZ5OkDSdiOIKmwcxOeG6YsPAUY7JDGeBb+3jqvQg1fizA
+bdfiq3wECmbaTKmpL7jukzJFkx6pfagSkdgEzpj6zCUFnJbnWm/wElAnzx7m1XTGVzeWcKTqN3F
SeDwhW4/EdOc0lc7rizbfmRBQITFAhAB2evNe4f7v2iIPDsNkTi+idJWYK3e2U5guq2MYhX+gQR9
mXRoHptpO+0tJKcL8XOWnR5nI+uIsE/uipuI7bb3ra9WZ41Yoloiz/ikIP7rSbjDUhcdquYUrxTY
eUXVVG8dFSRcO57uNGktgHODA2ODHf2yJJb3kZnb8e/tBPDtA/REgYmYbnXvqq3/4W7G2W3U9UeH
85COwXfW41l/bDIWf7U4tsysxO0diFDI9loHnaLDJFVGxumUXGdw6qA8fEC8zUrXBots0r2rLCRd
bhLlGPj2/xtZumwjAynbY+BX6YZIJ3JO4Lny4E7OAz5g68i1sJSPhTiLdjQxrGwbzwvY2G/jh0BO
nmf2DYIhxGO3oQYwCn1K4QpPwXvyY73i/Yk+Cjx173rO2Zt2zF7+asAtlta0Hc9V3cG/G8pSSKlY
IqLrtMim02/RytumLZtSMK2O04Q30FD69Awe1D+62qipEnb00mbpOnD/D4fLZ4ad7BxFaQo3H8ih
dcPR9V3av/BNU1wYoySckXt5uaw45FFBiankfItV0SJc6/edSDDSk2n/RhdD6FFO26YTX7vzGVMi
0VMH/PMjSiDZXVO6rVECxQZ3Lv9oRpG9DE5CCt+jdIJ+E1yRaC9qm4/D0bcGRu7bquq6r1ez0h3b
DAlcIiWRR0luys+nNC4bpov2a6rLJgXKgRF+vHj5IajMocMF/Mrbp6WnqoJcLoXrz5tqrg2I8ONO
5elv9PIrrb5xr3s05bSEJHb+K0s/pgfJ1h+wGt5KcN3RoIJlTqk++Xfchtm0cL9VSTUs1WZ8lOSv
qVnq5FRwmwto+f4sB94yo8v0ygRtkKb5EFXmOmxPgRlwe4734YQLYSjxMgRaBRYvUBiEHHAuBuA/
9UtH6whM/QVmT0V1vP9TQfmqo97HiqVKIxkDI2dGFbct4pUGMxB78+wZGZgGX55lLMoN9A1vVxVl
Vfu/SP+OL3ufdy9cNJF+b+XDz4rOldU/cvyCMMH5lONXr6Vk/0CaC9U0kMclit/EbaXjmMDvgd18
aNQbqwyzb1q1UqtcMalEFPo8f4IxVO/P5Aq/5hgkXgqRpryDXqY8T9YSO/ePDNSR+FD0FwRlCKdA
w+2mY/zA5EnymTX8iUpf5CI9rsgcz3zLqq4xsW8Ci6+/lDv8iaQ7Tf+D+0UdC/irPKb6J+YJVWDC
cOumDMBmAMc/o8UCwxlrSnCgvQPAgaa117wqG0ZXS6SE7gF9bb35L+c8XJ9RNg0+8Rse9JjurBXK
j0VKJpCQQqW9J3KJq69C0rANs/b/z3XckOJkVxTafosCAD4n1J8CP6ZAoxBTXl3G5DAJlNqp2fYs
Utf6/C2PezTwLywkIzJfbNnWDnuftVlzlmyVkbSvrTN3+i0kjs0ZOFETP7snvHq0aefAAQ+E4Vcr
lA4+3RDNWlXvPU2uY2+1JSGTi2snjU7mwWgFYcI0gYo4tkIUmJZzyy+fBgGeAxcCaOSyeOxPH/f0
JOGY2NWX+F5RLUwh4Vl8WXFn+qR+cwhNLhi4KE3IlVxFcqHlIFk+78vgrDw1JYsEquG/U6hnBk0b
kRcQscfF8a1s1s51KfZjtprcZ78sX8SB/grNBhyHt+rXYtM992FqFK6Hm7mLM7co0VS2bc4g12tV
24vcvKTqCo1kCZGZ571dBLBniOQ/hTYfpdqCDjxInMJSlMDcCHm/aN76Qi0NhPJHsjgBQY7Abnv8
wMmZMgggakFPYlGWK/dKJb7n/fd9UXWCyWrVsUSPsfEYnk5+iVOgf5sCxsVp4CsK15JakT0Jpgwl
yreuO1OThbyGOXNytnTlr3w0yo1It5SUN9f1RqhrN8O1IerX7PgHTZEp4EK1tKn8STiQoXJyzSOF
qSZWJfTDAsfN8Q2hotMxt6GK2MHX8xMANAelDOA7alNM6sU4jOETDzcbzPxwW2aBAs4ywRd8wjSs
aPQ3px6003dytfX3Hi3H3rDIa9AyIWgA7FOqSsB1cNTs9VVPFI5ZwNJl3mBrw8VHSYR1uZmOp2X/
704o69f+sFgkmpu1fw/ixUYhjEHN5RX7Sgk1Q6LEe4xpD6tZiNdgGTWvednQpKzPCogz1jbmm1P/
UXr2h9NVMmq14UEUK8JvG9ED0x5ervzCFE6e6pQ4wMpvPHsSNO/Zeg3jkFxAo24TYzpTpRmw2x6K
aZxY0UYK+0PtYjuAB7fbRCbH/zlYozWzdM6r3ntLqPcQAlfaKyJf0NGh79A13Bg/OVtidinqWH4c
uJD4a+c/XR5lOC3/wEsXdvIDgXH289fC9E6rqcv8mF0fZyNa9qvjgNxiulAKUPUSsFWt/4y96Z+9
Il8rH2H9jr6iiS65q8pzvkELjv2tL5V0sxvwscfeeflFM7Cwr8HSeUAUviyG/efd7DPr0owvC4qv
RS8KN7XHYWViZN2bwY/L2RZn+RPCoWnK2WbE4VoW23B0EGNHBsSBGLHpvtWwZ4XR83hROZrSMn/b
tGOesjtWK58xVv3IM66L8mba0zBnAeAr5BqbYtEniYeZZoEZYsaMob49gQnE0FF8t3+c/UqWLCi2
UHrsclouS2Is6Pe86KIxpmZZMQPp5qmEyaYLB+qosPFR8OtK3M5VbQ0ulkK/T/DO84dBpRJDIDdx
1CdRQE9hMp0NXGrNgHum4QlJFESOesv5tY3QN7uZxgpVSLgIJXAPmQIX1jg3en3cAOX+8F2Z6NE+
fPg0sT4lqolBxozNZF6YHxV7FXa2KgGbOoXUcyyKYnDIGJqhhnJ+5SSU2qz0P1+5MAvx4Xsdc8jD
sxeT94sCyhgFu7KkRb1Anl7S+irupu38LK02VLN9xt+FcD1bc8NNCx6bxi/1YPUnXHnx+MQfGGXK
uudWgL7xNsfRjpvQ9oVaTN1W5Mw28JY/NGBd8MM3Rgk5bAMLp2BBUMmuUiGzctKZecxCDJpHEGE3
RixXdHiJvTYspp3edgQgKBm8ps8ID0OmHeODzPaTJwnxDao+Hge+KAJtgg2VbeBu1FvfenYNVoMe
fCy/EKjVaHBGv799l7ShcOR2KOW5ymZNhQIuGEg8H85P4w7n88vF/BvU+dN9OMbdsXkqQijSk0UM
LkaV4r02J1JJeJyj82QvF/QkrCNuOqXQ2DdMUe828l6HSH7NfTvd6UcXU57yjf19hLSdApnL589v
E5Vxk1+4DTdY5/++ANbJcbbpjYifGgE5pPO+djCWaLFw+7WAzFWB9NQrmHZtNoJ55t373ZVm8wNr
Au4UZdhO1TNRSSX8ZUZTgruKnmrx/8mwq748CkSJOPF8ioLb25u8qJtmoRVvRo6mh8ejkkI4JQ54
d9SlGqMVmqqqmfuBK82QT3IOreyYfRB28XIoEsL/m7V2yhVL4ygowYs7uFe/i0ua30VJlFnK/Fzi
+tHQFTtcIoD7RZyxF39UrxU7VF3M4Bdfz27FXuq0t+A9fEuJsqTVrfIYF0ehZwN2InTl4yasxEno
1P+cY4kvZXhqr6BY0v8dhTPMSsnDzwbvMlsWFZxhzVqqEtAozBZ/rWCTm1ZBLYj+qazJGJL3cg+r
QeBFakxGXzlCjtRoCOlHrt1t/VRjkAxm4Ycd0drgnawAZjtUqcTBP7ol9ggERIcYSLH4uCnl67rp
yUGqekoHm/MiSEG3P9Dc8Q/tyDjYRDegS+3mgzEkr9YVb9aCAKQI26sil9zlWdnqSnIyf69lKcbU
WrMtWmml3dlO+QUG1sTLNSBiU95BGuovW0SBgkI6me4H4H2FWCPjJ4A8Rwe+DbydKk6w1oghPkMR
VoGfZwPKzbezSrV/G2DVgHX/9zmNA/rf7v/GS+Tgz8NLF4j2gWCGG84CbEyaeRRklFe0/3mOyfo0
XIU9xtsL7nkLks6wvRUpQQlAiZi4O0Rco+LxzHcDrGJuQqT0enKCcbaozRL5+ZS/XyQVhgUsMzCk
IGKw/EUhEVjn5v+6DaewbBcUs3OEpy9lB1EHV8RRojQ55pLJPQ0WQ25hCgKrG9uxP+zam+OrkSQ8
viqcMkMM6zxoTJCrKeKyWd4662kd53jOHWu4ZwlleAoOEduhnYNnL/bagY2zgIPSarzK83VFQScz
D4A6s6R1NF5QK7g/skVT4OKqKd8wYkfXH5RcU4SaPvpnBVwCAs3huTcZJnKuTJCRY9CeMAHCTamY
B58LpqHdrP4q7paXmWC+GMrNmzFUWyc0QZqkEOVRxJG8BHshQ8SmfOTQV5e20amy2Y6aVdEO1PaR
GG1L7Y1kIC3A91+NfPhO9vaQqXHi7yu3nUvCQe6dGFqSjoL8cRUq47+haKYQ/iQnwzePUbROqJn5
nYdg0flYziDjJb+hDIt9HjCDwytS+Sq5yx0AU9ue+8o821xbLF18/0lElgdLf3par0/rLgyaG3X5
D1K1N7p0C3VDDzP1bZ6dhYBrYBDc9L8tfbrfNicx7FAWtsmGYzRvIVVymYyzeit3wvTN3STiApgc
2Js7Q5RezpTxsyxs77+mBeSYQnd4vY1Ymnz5FnHDYS3EqCtaLmq84fCx4HsyedW9WpeX2matDmgz
JY+jdSAK5mqhxd3wVM1l+hscsd7LBDDmIz2yYvl/JIuBtT93usCqFAgP46h1rPfOvXURz1KE/7nc
Jt3dfbwiJ8zLjxquawyx2lNY+GGUF7nutigrpfaExU2Pj0Hcjn1JZOeoGwWGQnnKbCgAiD+dHSho
EJlEPt3IxCIWOe1JsikAYuFFsrQBWwwLAWB4blrdbH7lPdWlvQG3V1Cg1s+Uiw7ckdHoU7l3ZWUu
rPhQV1aRnM5nPUDDOqoT7BWm/zHCm/p7Fm9XjPsDHu16HRz9hM4U7C0Co8J7xt1cV5FbgC3rvq29
UfT6VN3EJ1CkZMoj65B164jTnTxi+Trdh5wDGwCe58QGP5b73ck7iVTyk3/9xS/DyJrvkqNivqZ5
nT2oKb1W/NoK+bIIWRj1KKbt5rSStTMgtGC9UKyF054S5BAIl6avBah4Fx9T5ZgrIv6XDKtatgFi
0jvYmsVCq4z3OslVFBmIgaewdLRXkAHifjWlKbEt1tPtoFcpiuqIr0Qdis8Jc6hJT9wfRStQwUJg
Cw2BOtx6sqSSbXgsCpm/Id+6NURQUTsnPNOg0WOMMryjRrUlA3cxHUe7pWMmVhljJFA0HMWf9+zd
9xjTb8il2gC2Cbno4mIvjZQZCaGkcMQS9hu/lWDFyrr0aq/2D/p2rgXmDtluRBBfoJdEOSFNEDG4
6eOw0RKevm1QmGSNr/6xSFSP+KLSjS7R6M6Di/mFvwuF50NeIniG/9sonjPrCb8DRYLk3vyGu7Z1
S1xNf2l3uOgluH6Alh+BQY7Sq+m2Isb47cxmWTVLADeRRgpNDWOHkaFIgMLFpxNLhReoq+o+5URZ
5vzIamCeucnxCNj7mY0Vr7hnyBpTKou8BnWAcOtV+fgkFjT1igM9Mp/H0TCH2ujVtuRVJZf8dEOK
QQ3CgMmzboDEi2T2gHNYmfzNc7nzIMXUxpEdu8klHVXD3XtQHvdUaCFpBTv8Yma8R9A7wrkFhqyT
R4EgZDG0krk3DWOluKcq6ZFB2xKe3af9emdKz7FSBpExBUY0MpbJMNLxkVrVmLfJ3Yn0JJrDgNJr
BUgxS35wJTV4ShUBQRKxKcV9Z64ekK0ebobwG3UOlvgTUJxLvP8mJiNT6RRvGh3IxNRlTTICm4uW
fCS/yd9gNKWw9Ir2PRzVq44RtxuXS1nFNMTz4i4L/FYk3FedCXMaQu7ht0gWI7EgPqg3rAjmvXpw
aXlfCgo/KVaZHhq4DVDaKuhODcdrJm2qYfAHPmLLIeaOjvNtG2sTvnA4a6JW3IapcZL33hbfpNzn
6LwFMwoMpBIOUaXJhXroPOpDU9sP8g9zrD7YFBrS9U6q/fQ2RNxe2FYAZcoJn0Al3G2p7AetPnpX
TZlvewB6ENV6zT2S1DfcdYypDcw3ne5cJE2DeLLgbWScPiE4fI9DdNxEkzMk2CMd8b5z1n9cIT12
whryYSAG//zKvQeLxknJUD4EyySNSt4nnP595xH/kIUWltxr1BgN2pwzSKF4hzxwsS17aUHfWWQe
zsJgDXBq1HRm5/ZGDaf6tggWSX+MqwbGKQ0q8soJQ1WhzsNThAPCVBcw5VI0r3sUVq4PFqqy3Nzc
7UDHFRNMvooI/uGt04kmCBcUptFgBQnpLn8HirfuKF3jHtkBo6FTug6NI8bIhHTxIyCI6KvEikR6
iuOXgiOmVJHMEG4sgOohfULsMQzOdvMkvd0YKawoClDWvLR9ncY9MLpmL0tx2gQu8O/ZeKqCwZfV
fmY9qpvFTGwtpDTm3VuuWZu3S09av3lOOfq8y5hMoDr322Zb1B2Hmg2XE8YOApRN5CSjZ9UDRBJg
YV2li4pSv6eq0b6hoTWTKfRirKamuoZcFlS63LNFJSNYmFl2O1jYfBBMY2HxhGjlmeJgVbg/vwbJ
eul4VbDyP0Ub3mynim/SrsKwIARSIskWRrAc+lQzm95yyC116CPLlli2y3lzmn8gIVzHTnBBAcnz
vpxur76zJohinClMUqNcT3keN9Ui0ImsRMashPD26+wu95v1raSvtVIXnWaUH3BpbAiLU3wQ4IBO
WCusmmKOC5JKkHZidrs7cLXlyjM1DFlRKDDCyQNDSeIqOElYimyLW+4BzU7wDoIJc9KjhukzhywU
KodWKlBGJf2RqiinvWeUNhi9fnBUcq8AB4i/ENeWmIM9Pfj+79LqxM3ureyjDOQA5AG3uRM6xRF0
qgy9Ttsd7mB6Yzc5wNrDa4LRJZcDMeXHy1MK0wnExSC9Few9B5RjlHzzaRiAqptvMQ8tKWasEmCB
kq2verJ+cFQiTq2B8sVDzbZ1RISlgWkF6z7t8Fij01ukBRfLFIVXJe9QIHtFp2mXhfMPhBJTOXU9
/C38cH5auMct6N21b0H64RwOMBEF2vk82VD67qL01iRcbC0hzoBFGzBsAPtLOlOgOtKeQytooNGc
hsbIyC3+SuJKQyHvgnHuQtZNOoj1n1OwpNdjadWdSV9tqAGfNDkoFMotp9etHYs2j2FskmfBXPqh
D1fn1XR64gKMex8mBbgPaahslQAPJsMglW662aQckHiDK6hShYLNVPPtnICgf7DR4jN+veNgsXEo
ICHTuavPNA+8XGCtTaXibnqXYQdKNaJc+DrroNPg380bJywwhdFzIBTZMaTl5w16wlom0+jsh95Q
v+wOPvJuCn4LwutXRb/hUR+kXzN/ORzT6WPfTMG2+vTa+V6ey34SbjqLvKwtAftzmtZpVAf3l3dz
mci8jeWQQELN4FY0QtVBWd9TH3UTi2RKOUjjUv9eBaMbM+hg5TFR7ivfADN8PfYSF+Nn9lelnPf8
WAJIqYOxG9hhtzrFO2yrg1pfXHfpK5SYNG2kpCK5tTV6NGkgMK12PWQQl3dQdi8tZ57YqJPOfeXv
M4FdIFU6akDqRveUGmkvlcmp2rgnk1Da21wMJL0PuUgcrEO4ReaFOsdhqUvX27VsRKU4mx2oYSp6
OfMVCAXbuGbgRaSQ9JcYyRAkS90ZtfEYVWrkkQIiFzZJU8B+44oJ8U0M39O2nVyaEOPvy+kZP4Zj
wFXtCvced7Y1j435uyAqHGKOUBe/UJY94SYyoSaTBHWdGZLIwHl7sAKrhf01mROrUVDn2cfY1YP4
1WP+NvzIeSfGXLj0hqhCtHkduIlkeiiI6TwOnb5x+lpVqch3zrOo+o37fwh+BFzZzsOajrcrZu3I
a7KoXpw4XtpLDUpGlSSZy3o7qhy+I03ksj95bQtxTUblicGoImIjAysAHW0n+dC2P9+n7zH9RUeZ
J+O3gTxTXRTSGS4E5yTV7HfEJ3/TyGKuFiSSykCDKl0ehOqSHTQmQAe92KYUSrDDTLuffzQ2jGYh
uNRDw/t8yl2Dtg5IgDg46mdvSbVpA78XZv0dhDouAgNs7KqmxrBqj9Hbdie1H5qEsruoG8gbbu57
XvBuTiKU2W8+nu2yGEOrhya9+6E41R8xIoKQ5CzzJAY9Xj0ti8xL5x3PA0WUyc19PKBnUoEkJ3KT
zKPjrIVYAqf75tYaYhPp+w8/Ecvg2aw2iFYkSz5QdDX2QTlsotp9cwz3+rgqhZ4+X4TrCTEdATFK
pV/ta6MMll87mqnV8hjl/6vmqLgwLme0NazJvAZhlRrsO8yn5nnHenw/uASZ9+tPIg1kTn9pbtx4
f9Yy1VTpEdSaFz38F/DSqR9h8cCS5kDX4jPkYnT/Dz2wur7NEhlQ+aReSMENXdBjVAZUnKY8pTJw
jx8vC1XxxLOpni3HTdI8xe6i8YHIuKZllSAtiA5wDD0qGei9sFoGPQyyZH4NfQOMhuXO4Pny2K0G
IOWrmOFZ/7JKxIPtFmR7UFpMsvyrBioJaVHwhrAnq98dRiBJ1Kqp+7vSeI1O+Lc5udcMapmA/uIx
8sZ3FJlJFRsljnRR9ACw20UWK9psG+otRMa5jN9z2Fe3REksLgUhRoWO23Pplx3NtcdxfHcEIURy
kU8SR2M00JuCsXzIo1wXqFwLraf49q6I/CI6nDqpDcvZywr7+KJ2ER15vR7baIKZYXHy7bOSUlf9
zfjJ2LvurHpbYVqkf1gc5ImsZBRR25a2sshvja2XzgrM5VGYQ/vAsHbQFxoDNPUCEQR2hV4E2LJw
9bM7hm+jWq3NdH0o7DmYAga7h9s4SQ8cZsVDAaVM5Z5EotXGCH436gU3Sg3U/haNaLi8RXkGVlSj
4aI9Kk+Lclm03z+puSzAs55jWzB/GC5Fbpqk++yE08KSBgcEdWrF4qSZMOfg43vT/Nh6vXM4x71K
JOO2FAhFU8IuYfsDHK5buvPyOAgY5efxSCWMo6SBLoFqksnOFSro7gwT783c30xarJh4OmxecQVJ
NYqB6uEK245j+S2e4HrjiWmkiIDx5/BwLkmEHeWcnzQcfsKwioBbG+nTbvEYyv5ZbLLZlDsTVwUq
Ry2e3Q3u63EyAFJbm+E3VuByrpJnu06Yw7EFFEdwKTGdG3mXskYEl1TpH1qQRcycOBMp7IZZEIJM
6sl4T2k5R0i8mZG4DBBNdM9Fo1OJ2TT+gj91NV1F6E7qsPz7cz9oeUqXf1mzGw85iGJ0i13rY5bG
6rb+2QWzbxfV1wI//pPOUaswxXKJSE5ARhBzIgTOJTlbrd4+WqLYTE2pYNguOXSYXeoyitrFoWQl
hTmTwzo40SU5BE77TacS2M5Mj9kW/JhbaEj/wd7JgD8GHx5Fy8cHkqXQCnCE0YNiRjsJ7bgXa1fa
asmjZxbOqUStHZqz/USEeMI+u7F9XIgJ/9drV1FiR6AyqOCEFyZNAbjEUlKmrYIljFr+k98kHsX9
P/LXPLw5ik1YYqRw1bFQ7VEveopv/OfAGBZ66vyhZLcX8jibdlG98++WQN6b0XcgdzO2NlBRKTVZ
/qB7/VWplMPFMxIqekTA5nLY8cFlEfU6x0CH8+LCkylsK8fXUh7qbQy1ypragaBUzhI1g0754cCV
HDEVBTMDjwoHIKWmZBRWkB2ym7BSInJ5xxLFK6bTwGJ/Aub6o6r6KaoZzSSNvqqqQ+7gV4Icgh2J
gHtS1EHUoG3kchXlfq7smd+3NkpOuhm/W1/opUREj3/uE1FD3EbMIJe7vrjnibFylIRxT7YGlGjD
V2hLs4mLkVky4LOaUQE/FqUJMniYApYHXDV2dEKvR3J4bzHBrRKLG65h6RTgYq8Lt98BIMSFQb33
a9si5DxlDC4fb9wMtyHO1SqB0OOyLI/28khnBf/VsA2hI5g1VHVbR/oTDOD0XYVnPJh/b7gMUQ3e
5eZIuQl5D/f+zEifKQuAJ1phiBg+mAMQ6wO8lAIHgnWNfnG7OAZwu1QJrFrR5S80Zixzj6GMF9Rl
/qpb9/JrZ4cyJ/kAOYP/v/3qLtrXEg6BX4RCG8sh3eq6gnOtmRJsSK22RdSG2bB9x4gq0Gzkj302
GNDcFY/VKihcj/KEE5OVXV3ZWnDXkgLHXQuVm/beP8JHJxfY1nVDMQpJuOZQMWAZZBxQfDf1fqj+
jHRE07lpWl8E5jV8sOma7paUYM6UBV3EeczwHrohEDlAISccuIheBquF+OF302QtI5i/QJLN+6kG
oRjPKzQz6QcfjAYxT8E2LTrqOf7HPDrVvVhc7Krg+oZ1IUG23luLQCxoG036hVXFJ+wFHu1qbALJ
VbSocvdkMcHMoi9oSWZFLgTA8+Q1gBfbiIK4wXCWs7cqi0Eu5Xar1eq1Lqx+Y0ehsUFkHPkcDOjb
xgz+tgvr7OlZIUQ1NAQlkDaMY74uUuIcvf0eBMA84GOTn/NJBl7a0tSHN38zT+PDt38AaHG09A9c
Eqnkrnz74b35wUAatmwMTQWPvzFWjxmbRYhIHWclW81zDm3Zp9XAEpFip9Wzee5PkOqaU2KHZnr3
mSLs30/KTrPZSjmqXBcgIRvRJFsfTmcsvUFsAhXv7yLv3MNdHJVRvaTakKOEGq/yYS68liY834WT
9FK/liYIpWgeXItFHo6dSMEXFNCXrGAZg7/xq7OpsqPvWL/f8M5g+qk1ArrNiuusac6hunGQDveC
wf04vM2plke4FpLAL9Z+qJxwz9p2I/LUOUwv5l+CqlEtKfEMAPSKrG52q1KNZMTbsxe2ZYtDCTFX
bkRplEjqEyor8mRyBg6zcuruj2gxGdHqnphM2AqC6YuzvhQqgCap0mukT+Tfdfv9GMjmzaT9RV8a
WKFb39lle4jy5m5fuILSwxEDeKjs/fYjVXvpODDxMeRzQErBkuuzAb6BE2YS5MM7PGIktBbh2TjH
aP27JxmqJTBpcbZZXAU8K3jyvRKrttCf5LxVKqp/1EMYtPx2xIlY7UH9ue9o69ZofFqGEzIbMNDC
3wyq1upiFbJ3NxJCWco3vcxZ/mZfM2vXzsJm5shFj5ffXxYWGAE3Usuy7gh4xCTEWVkJjyjWmN35
INi2tFtwT0AilMGciN1IuuzopYuyDvEnsONFG7gdvMJ1LVEYt3wAINrFkMxC1CSwEXJSap0zEB34
jEg3eUAezcV3hgmJNfs4AWYEKEsSnzagTMt/brJor431Z+kUCqFFZDb84JQ2vP5gY99WEhPBj9l4
6QcAJdTmDbQ33F6X5cRKfe/u8HP+bvzMmlEdhvsLMRtJhepT92VtlQ/aOb+r7mEeUnfxmb0UhLj7
GKr41c67qXcF4z7N7225RH7KThX2OqoUCzsFREiOgTYTapL9YtRIMVIARFeQSyfNFCaZB1yIWaUF
+bHNIwkpRsIT15pdY+zoaEsahb2AWyZJRomdZPQC584vEY6+SI7xa+otfHPFwg17Iugvg3Q+c1Ry
NJ2nYR8f/B2pgwwouT+Dt0ri8cF0HuB5XvdvYQ+VgWHJR9yi08d1XtfkDhxy9z+AcXZ8iJtAVI84
zc9F24GA7M65jFSTs1GJ+4SGR2euQSA8g0GZ8hwsHKQ5PdavnJFzLtT1Va/ziMW6PdWPJKJa6nS0
Ht3q9s5q2m9abf1+33zLR5yr7M76DblpMb6kMN6Xay//AjYCP2zb1bB1KY5ZrC/XuXUAavqiUTA6
Lva01fgarfrxmHgg60ygLYpHR+ewvqhjFHihsXWXFLwNB7+Ttm4JdlAvR59cac1HbeKcCZi1cw++
2YavWIbxkkgFe4J+a18xSAN7SfPRSFYebGjFnFDRJNsGZVw5kghyVaf4hPID871vIM5efmT+8Dk2
i0c+sIx7oqkPn9FygcEqST4ViHaNgrfb9BCCOoal07M09njQVmjIcvSFEoWi+BHYCmYR3JcrckvW
2JmGlgFtesKfLOvVvfkyRjENLWTNKTAhBjX7oiuWuVMlX1DUICFHXdHJE7sw1lmCM6XmEdGaa/2p
3W40lM6jP0WFZUl9oRztEEpbTDqFP0FqMm0ORsP8hKDGjOTaUoU011hP61VFnStN2HsBcv1HCrg7
SIrHAOdw/1EnJP72TzkhifRLId9i/OcQD7k8mElLknQQvsbqBiwU1gGOfuvnIOCfLtIHcLZApAIo
UJ4JeCT2l7t9M9Nu2Ay6IK4MQliBavPYSgE2pBJ30Ueuma3N2X+3Tsz8K4+fE9F90ZNYg9dqWRMl
vLPQzLl8rwkfb3mSuuse9gfevMbxYzwMRougGv03kT2BpmGSCLMSJRE1jQM68hmD7oRJr3fZ9gTJ
XJ5VCMxaphvCAmy1xUIQp00np1WJWs8SSjBLousz1g0AOUIF34tujp4xXHmBXl2lvXmw9jZgLdYI
K4rtb5dWdmUrh6FMxR6AZZmKqFGsqhKtIl2sYgrrFDPINw8KEktVu7Sjwa2VAmHAkAWbB7C0Tu1a
GO5S+00hAUvjuynr8F/WkKNrh4tK8prDByVi4a6d3E3sXZ0yf63XyI0l3pKHAD2Y0DMUFDfrb79l
9ShRmZRwLbbZBEttFQuQgbsnsuq18rOM1Fa0wtn9g7nRgWHR3pZZEdCw7lwK4Q0ACnNO7Gs0gipu
QPFbh7bhC55bCA4RBMIyarVoe21qyCEjihA+j0b2kjjKQTfl4/9GnDQAsau7ZfPtcjdapAWT4XLP
PTGzsXP4MYg/8w4lIPa8e3/zUtq54pBudnG5HxQiUpVZBQEEMBFIcZrXlD6raYP4pFZfad7wSUV5
gvaxifoOeXGIokDRD5+6yDw+ck3/nYVuCfrLV4hSf9+yBI355PgLfmgBuYxfH2spPNeveS2LMi7m
vRKQ7KfgE8BnykLrbp6Du7f/Xjs5wueMfIpdVY7Oafc2wStrTeIdcFfd9CpGxepp7UaazNTBqW1m
9oGzOfo77myA7LIdYxNx3AQY1IWCRxaZK/nWeQ6cdW2grnFYi8dpQ6gWs96ywyTaVMxrgcQWyAmN
IlzHJQxCosnt8BYnwe8Yl3PTr/VcuMkfZFyHfgSH+Amk0MpBv95hvEGMJug0Nn/7dca6rg9aM4Mn
raNiri4DsuXlIeotHer2Mnu37ggswftMLA1XxJrrqfR09xwsJ1Sb4DMiDvfvmbnlRgiBNE+PWpIu
fUzMEIerrcxGwgBHnKE7bSNyGTcPW9p+Bfe0UQ6tdGrqrfou+cZ3+hWUvtFxfTHxeXPgXPoB+VG2
oQ6dWxlAUVVm2rXCAVpcg39fYoBpokbH/TFckhS9aZvfYm2fYR5lyl9tMIXegcO8ekuXLBN0ORxR
CROtc8QyXaywPh2OBDogOTmNHW9zYYynt1nhoDWW/n2dR8XFJPLz/odmdvOGX11bUZAFqAHScBII
MEBaKDeOADOxuAJo0wT9k1ePlUbSqq89UWBDZfHjbbmb31vDInQYIo4/lC+7FGZ7p6fAzvcjd+a8
gaYZwRqXhc6dQqccgO6njFYPvmUJhjjxnKZReC4KaLdc9r21SzZ6m+Mhtzm7zQyBJIdGnkIYPSSG
ChYXffaZQkIyHK727UR2098XT0JXB8q27PLmHSQRbM/8mceO+GvqMzFR3oPHmglOTboWdm89GteP
pemWvd9CImW2g8Lzi8d52zWX/mRSwzFeUT0cg9Cd7tRFMm+saw219zDpc1JxlmBXiy/xlu2Uy0Ub
CiqyaWnKHa0NN6lfLjZIHuXpf9A/Ao6pDcv8V0DACGea3FqdPtl1cH93cminGCC9V9tWl2qOWtdW
oNmUu7+jtPgPtXQQqcf7OEbKo0uGFhYcTsMdEAhWOrNEsanHwp6ZU5BtrDs7oAUU75EmwKzFMV1Z
tW/KDP+4J0PpxIjrCkIqKOawu7xXfhhKkowKCmhNpCsNoJafSddZz4PGmORU/y1Aihj82t89Lq9e
DYzD9LREqzCmG8IfhYYC2IqStIaVgzXd1TyXHOpWXKzdQei+3zACAL7m0t6E4tzNrmMEuHi8X/aS
UDpsumnLXszwXhHCVTri/QA75hWVFR8WtGejxqUJypjbfa1rUu9N4Uc5/df7+jxYUvlQiau4ge1m
VWDHDAwrDEj6VlOUrP5nP4WXXuy2iDo+NCM3TygRT8xwTYAqbikaHvS6/70ut/z1KIpdsdcpT1u7
SNPa0Ng/DjI3eT1nd5eXAJt9LgfMI3PTOL1pSEOWNUA5+wkSU4lH1/1PZ0+VoSfgYDwxuZ+PfMrG
lPHm+dckcg37Vumy2JTGzr/yY4se3EGZt287UxyD8OdAPXlLSU1XfLYdXkQ9vj93Y9d6jPt9QjCJ
76oxueeV356eaf9ysCOR5wAoZhWwLzuj8JCD1nmXjQsiPVSxKR4l3nTPUaissL1CW2ULlbR698wi
YgWvwVAsfWlKEges+fViE2PPayqjlY6iY8CpPXiqscVeultzlF6azqDkBx5GsOM7+iCKwmu8rEq3
VZzDhNKeVToi2k+DpZosO5znZviyFd89e4DKUAOyLZ1p4gl1aJ4xI9xPOQZZ9Dn3PRRBgzuSASEY
2/kVzVKnQrrUywNSBZAK25InFoIpjVuwcc+hydCOzZ43psCAJEjhIOp18qmSCEo8lDTyFc6EXjrz
kTbZ8tuVKU/3hz6Z3yFVAJLsj0LVh16/BQE7vHbbcpoURqrHeMNsPm2pFxbUB+EwqjH/Vpg5O+L3
qeLw24VIgU8BbqmZdIv8kfp1WO8dDgMBYbAxMz6kCOhygPN9AJ4hXJncuoKvMdRltMWpNtFBI07Y
lhx9lwlUpUK9CzvyzSqXdGJPJg0k/ua9qZAOSgvYOb8xfFfO/yP0sGVI3Tp53wJaRbjoPmlMmKnc
m+vUjaP3NzsCHSKxRwqCiT+iqoWWLPqlS0OzBzivz9KC1loHmlGRUaEh3uUNITNGPNkJgGSmOZQR
FVPosMwZh3QSedvsyQCF9Zcq5RhuyXGc0Z6WWfp/PJIYk5hLyux3L8HZYYiH2ap0ETsJ9hYR7exs
XPfnyVvyz3eEJ6iQC6WZwJaUDSlgHRD5o7+FbE+yuJsGlfuOPJWCiFru0CB0qrKX7k/eJNuRmewG
ix+VDBuP1jGrJ+/TU0f31c85m7NqDI42kGdAAUgzzvAsrAe2M/0P/k2urN+dlFwSbqQLmSD2IAyv
iQKpmXgQC+FBwxPb92LFA3Gdxj74NxTVjlxGLpP8eOplUsSQeaEapTuXRaUeAA6XQKGnWLFstNEc
asIvzIEgHBggV8YvCVi0kiw/H2mZI5IPFMBGNShZT+igguTSVu1rSlYJ0f0nccvW/dlVJz9E2FW9
YUMEuaWoztSwuf5aSSMtuqzEalCqBHOoZaA+gDcwVxUj2Wvcrs1sUcEyFaRew61cJr6sWl8KH8h3
MnMD6JM3OSIBUU42P/z8UsReq3L6LbR57lZ0WXuPFiWFPtGHJ34jPWPYZVpKdQNzLx2b6ku/VV4j
I0rQ6zU18w7t6cZSrvZA7+Vehgk++tZzDzMr6YmMh61kY3F0sSPmPdyGg4JXJ1yW1MTpzg7U2tCU
PzJAaPeHNDAHmqQaFgbPYUhaG/cTY5HfCucrC0aUi9ybehQtg1xGK0hQI+xi3YS6bl6xxGfaRVkg
I3mj+DjhV5VmhQyzj/iOzIFZFAm9qj50VjSJ7IcXDORnDK9lcNa91/O6BQDnu7RSyzdgc3jU22kp
gTX3aMNNAXZOY92ShKfrDembmcBzbAtBnfUhT8nLnevJuYSU3eg/YWywWvrh56ET9ycYYSgbr8Ue
Dk1hVQVPJMBmKXcP9JM8wQttiJSIKiYwTkRWJgT4MeHXVfqmkrj04s7YH5hoGfz88NeaHfQpIRnP
35Ri7b5ZmAyVRXQFeSVsySDVfpuZmgOYKktXHox3MsepPu7cWgqk8VF5mhguMGH96hEPdKEq39yt
1LBZ/PrQwWhrxMsD41OnqdUPC2hgzImFWo5j8KyF0F9ufJ3bFZwx7xr7Oz1zyc8srq0s5OqIaC3D
P4JJGw6btU9xOxU1iQvPj+Ei/cSOlqyFIO02enUhs2vjOXqdgKFMeVcktGVZweOJ9yA6JNUOGVni
3Ev4CxAJDExH2IitIp1XqGCkAIpePFYyFMZC0cbKzrPnnQIQRW1DnmByfkaXt0xHVquaB8MsPjbw
MI41LumdCgN3yh7Mcr1UFKVUHQEINtKrjamIwLB5YpPssXicy/8edhkOQSUSh2x6dBQ6Ci2fAV6L
bQNMsAG2Ah9+OfCkb2tP3/VNpMLPtc8yZLChAIOspug4d3wjLgfEQeOXwHYI1bVFj8CiIu3f2Rzm
Xog1k2kFb1pQA/wlDOGG2dRvfCJhE6D5vfFIDDaR9/XPfyeH7PKEXQsa3yVV9TBhYLQb12ZuSndx
fQnb3Vcdak/0XZaPbOdP21kLaM4FGVTn8Q1EBsq0lvLNLvZ9pcUCS1o0K9ShjCeAmH6XxspDxuCm
n7xGOGoQN4J4f6IQfqfG+PZHaNaE/EhKI7PmsuZD9dFEueHHZz4YCpn2cg8Ux7HfJkdQM77MGbND
cevW93EgCxXVvUxIE0iJXlq+7/tusbZafblT1RJRYGvX6mLE+PesZ6AwRs493HkX25YQI0GCLpmv
TWVwhWNBgpiomHlx+4mlowIO5wkaIL3Ov8Qv2OQygDu9RnA/0uulArdl4emOA6xF0RB2Tvr7492q
E0uUgtqCfJ4EBO4tAZJQWc6N1O3BKAiNmyjYqPmVZJ1ATeRaLPh52WkljhHlFUfqpD/fGz/LU+xG
7tgHH2B70dGGdtK3Kbh/wn1dpPahcZyXtkmm4+20jQKnNgiE2aSLSHND1Paak3ttOEbcot61bM6l
RMRIae/Q/DTN0d1A4+l9Q5y4OIXVBFBFxXRUMmmmop4/LjZHzFmS1xvE2FQC9cBo9YX8FmOd6UZa
RlSISgSabcM243e9jD3WKvqHCDdhiO45uSEtgHV21PhdBrecGjmCCB6p14hJW1lYvf3/bVrkjiLQ
swzmwp6s+eiZynHKbA2bufCbm0UFonG+FjBiHxwl3KCNLRG3j/kXR6gw9r37l9sm7u+WA59SBehS
Hf463yxLIIdF+5K12jrbPZNZdLS76kAReisqqYCYwDRh4cqTMZOoQwK4uZYksEqWglg7zH/Tz5Sw
AzTLhlH17840yccXXHBDHoNvd1qoxSd90P71gWTlAXprVGJrL+9SabgByn4yINQ55NOLqkjpgb+E
5y58r7/Qdz8CKfSXQqMzCrikpPI5jsCNZ+U83TrwG0PYTN9K75BlX1qHGDrVjUOPznmjXeCersVI
rJIHQqwMdAQBf89VZTovj08t3O86qe/e3fL/2RN864CL2ldnGLd9r6U7V7ovbnGTySKn8Fvz0sI5
Z0PWQnwJvCxDDe7S8Kwg2UajKgjjVjm7EKejzzn1T+RtaC4hiqONlzNyTMp4S8sRtriNzyELQWem
xdIGf4xghBuHcsq5P/tuwFZ7BOgfA5YofBu278nSvliSaVfg0ObxE3fF578wS1iWLrL41fm4XKLn
xSfjwNXYu49VOIBDN0Zu4z6Dvc+6j46WgXxpMXeKL682TLhDh6ZRzBM3RwTt4JDCWhYC52owWZxp
I/eGPRriy3L2rzj4ACqk4FDDRVT4ywCJ/8Lw1/NLDBlif/KwrGeOGlhXccydZ/wygd8tHEqOewze
E3R8CopED8bs2W/Scu+7lL5HPzpRKZqT6p+Zaj11ZDFdEWyHs8fuL46brwcVxtTMFdYKFnpEEIUK
hlAlbYIOA45rg9XPxOmaV+x17lbbYvGXdPqEV6sl+WnF9Ya/PBAaWzN94eX6rSH5ASGyYXQwwQ+C
2YI58ATPPAKuzV5lOmpiTV10Z2xWtYOAsYLJrWIONqnvFMCWWd9vDG7i7dHcKHf5Tf02RvNLkFTK
yckUJG6QOUJr51Ap2Dq6lVfDj0tbAXueU9WLnVVTTUxr/qKYFONBLlwAu4LeUT/bofKxIfwviQMK
jfF0NYTraC8ZN1vO7gKIqq0tMtMxGro8Kv5X6noFgV0Jj3Yxqx61TDear0CnSk4m4YRMkotF+DpM
67z4nIkz0GJr+0UYJHLGV1Gzm54qrghjW1RmXlidDeZvopVTnvm+BmnfKkubEBfY4XWCl3qUXYYA
O4di0xH8k/Koh+tHhVHhCIWzKiltH1E471suErYRM1lgD9RAp2tDtWsjJZXNBYlKAQK7jpHqDCmI
utCmJT9arJ5yKQbjAYSaXKzL3u13ufF0mYqvYPzw/HcWP/E1boQd6dH02DTm/enixdemMDC2DINv
zaOZOhY+Dv1xdJqfA3az6kqA5pkse0F8n/YmpZ3U1sl+96/EkdL2jpmDywp2u4VZFH9Vd7Uxr++t
nLIL8ig514HBRpqj56axBplhle//ujGdbQMZtpq1oYyZKlwJmxT0CZFDy8M83wELcJDB4qX8Oism
fnrPjjKNJP0OqAx+VKnt9PjnvGFT+52I1jwKK6rX9RI7fAePb/fzjS+Tlq2XEmsExbaZ7V5yz6mb
xaoWZiteHWgu064h/BdQMJZg5o25Edg7QbawmxX4IUKbjlHgQFvDcrxtZyJ8UAzHFAIn8KV4SMfI
ASWCdmfocC2drf2LxbB/yHEPjkbzblPAAn/BkADdU8aztbMJgccuIflGYoeWuzkEnEGPjkPtBRfp
E+f0qPPb7IQ+Yh9QsVKSO/4gKzM1WPBDKG7k3Hq7omFpy8Y4xq1v+xUAMZPEbJ2ChVPIjE/mb/ep
+pD/awyW9YQGJfmBURRIsPTCjMX2bjqiDVcZgq2Zb2fuWEoH1QZDNILF5zODsONwbBhOLfjvL8NY
GKnuLapPb2fFpaoPupb7ffABv3mNAGT+aecvsbM2vcpDCPwZ7zPV9hZ1g5G/Uh4/oBMXvFdyPBXi
wbf7Io4+iACVvWsP401FWGGJa4TcigdXOnQpOYDrPaU+HJTDVs8070tX9zFtklqn/nEoI4zJHG6y
bVtURn4LIyNEBW29t0Y4jnwP3rDafv7D+aCMyua+WfCdZSUdvbW/+nE/Pvy5Yr0UF6xyrnGv0uWJ
1YFekn+eMOy5XKjxz8xdtdZt8MYMpAXPoiPLs8p09THbpluECREfkchZJWyjlmaXrFsY59zEmtTz
MN9JoFy1m8txUiEIYyqyhAYt3RTq0gbDmths1feg17e/tpRk3j69K4cw8xn4qwFMv4Qk9DuRQDUE
RVOwQvCcQKgtyd9Rto89W+yxhfaIYW0wHYt6NRoqJu0NwCIiHcUCxKVYzQTVnaJYH5Cn2p6Y5lRt
cuFD7mcPVv3DFfndg5shx9TiID3AO961NW8kbP4MmCGvMvpwXP94wv8lb8joLCadyyvnzr0WxCMR
eyN3GM9WizFAg4HYApXh2APYVlnFc3RN5Ts1v/fOgRTNAmcoLOi9Ma/ertWH6GqprpbWp8p4JjBD
1PjxDWzh4zUZhL3jmk7ClYIN1tFAeECHfLMfkU8hs3tiwDcwOFattNR0XuMOnb4TVmt5g4dW/llB
LiNplSBnt3LtGyKWpc/jaHdb6oHMU9fQcZKfFUMYJ3f3GJVU437cSs8DzqAUm8rgnfxu2b5mnh19
nXtsUeGHYl1KQJX/diHD9B1P3EW8bQG6AxcmOCgpnERowZ9emU5OpGcC48ukRVf3myCHPfGrgoGM
ljtyWxMTMVbTL8Kfvq41Dtc9U/0CEb/dxdqFM+Oy2o+gHWjum551knBUHjzOAqm5TpivDhl+fCVz
08JTtBKOhwt6N45tjz/2PshWJaiw7URHui7TjYvLDcf/IcVnBVgcsG4fwA7j4FiRVmqaVNbieyvJ
wvG2K3KYcsYT291vVPSt0I9pAFyunENbHa/ZNx7AdB84mlLGdbbwt1FPmr5D/FtlVh2Tm63CTsxN
3tdnxMPx4jw6owTKwKXBwW8pVOyx34O5uDpEUUwmz7H+SwDj/EIrJ7F9JHPXmofFr7QCHDR33zfN
wJ/+wRrQpZs6QQ9mjc40XWGJp2ImhOpvf4RlTeqtDQdT5MjqKMfXJWOstpnM8Zd+LB8y79JPeEK5
J/d0phbfL5gv8IoY3rZ2tL9YT83F3vxuYwBA/7rbBukJl+1tI3EsEEuiqMyQR6acsHvm67iuJNZz
K/vmGaCkWT1HZxTGuFxSwlTvV41f4n774a4Gjw20xO8eTJRKHHMZODuKuBg0FQ/vXLcWc9V/OsUo
zclMTQIyqInBCfpj1fx+oRUqODkPpPIOuyhTtlqQGA0vb8NkMUUWFHG3n6B7pSSnUWqsn5w74Q55
6Pf/hJQM3hl8gY+KyCPzDbNakbB/dsMIPkwycu+dZpWSDLVOrN2zETJEKmRoG1OQy/y05a8csWpN
9ctgrs4jZXDQL2e22Xc2OZMuSe1MjBoltAhwSXKhptwrc7a+X68qWJx7xct7ZUSicwt5DgaPfw/N
2cTsK160cK59XCbar8jLpPCuKpeW2krJa2F2WbWKSCbMvWiyQrHsHdNVcUKagn3Jb8LIx+pgnMAJ
59ewVgUTX0ft8vkrKsogabl7h5IQ1RIj85DnqeUOZ+rLb5gDoAk2Wers3pX+1+XYhPz5AGUDR+9/
LK1TCXS3wcDeLR3H7g3ikCO/SYQLU7fbKLPMMOq5YXTwEZxhO4x/MXj4617kc1kaClPoo+OC9L7L
d9Qte2pHWudRpOQUoiYF9d5i/46JXHroKyKf893tHmUf0S02if27QjVhDC4rNKdhc825VS4WBd44
Oq1s8djerqaKc4G34Aa3omW2A7MZieHuZ9UnrM8JLkNNR3HaivNoddYWGaOIkamD5EnPQe+7iosk
KV643mCsQIWh9JfMn3k9MGC+REO5nfcihgeehVSO+lg4HmUAgPPKTQbkIM/uu07VnVXoga+BHUcr
KodJhCKxMh2IfVP4LXpIuxcYdX6SikZmgzRG1SolXAYRI/Ik+AH4OyU8SpWYrx2L7H+uRS2sXFmK
zMoMJK8ty4KE01D1iVKR6nQpIQn4ZIn3gPn5phusZ0bjJXPkRu6SUj4GDRdAezK3M2CQ9JxLWJST
wITHjFskCA6RUe/PVDtJ/Gcur0VDwDOZnLtHWaX/bOn4XroKAEPvn4fed+8rxq52aMYbJESxo4lI
yuzNKBNwLLeontEHH43kBJsMlUFPmXk+CvUQYTodjBXNzPHRkVO6LXR6bL6CBRjVxpfjG11CVC0T
QJ4/Lo5GR7vELqR56BO92CAsJiG8JT8QBnEPN6VRTwDP0RkExbLY1qeHbMomzGTj416jsASglLFK
/zWFv3zA+Xi/RZUSkoZUlE7E84VcqV5nJGu7+LlAvKo4bfVI4rDYaReJh7E6t7N0VOnIXF6f4bzw
dqGwnTLFTXDgHNApmFTPqkgOQ4aqYB1uaCdYBda3CJnYjYxduLZGk5oRBTW1r1hbt1LPr2F347c/
hDs9mPhlNVISbRmNg2Z6Xut8KX4u4mOoxK8cN0JRvgH8Z65JoLCfeQbq8PpoSBblXf4CIuGPnnF0
JBuFaiAPqKPb3I0Jbmb0MYLofQ1pVG7Z13u7xE9+nZOuAKh2VZw9qqPx4ES4NpVcgE8m8HOg4Bjh
1K4cDaSj/49ZpW7Lo5qXCf+Y1DfheRI8Z0kCj6/cMnaV16JJTM6CFsqiSrAZfsN+7OfsD0Fra/gK
xTGRb5S4gvqikdkdj4CaZlDkCO/0ofgwn8iIwO2+AGO4YOFCjn/ZEnPsRh5pbP2961gfE49T/95Q
CuCeGljvchN47AYhe+RNVWcK2rBn650by01Ew+P4eCDjBKs2O6+U+ZgCN14FI0vSttWcIBhZ7J9l
P16TjHsKtRiZuD0rWBCRNKDydZXatxLvlMuNVj/4CkJOQh/8mxxp8zr5dKi+6434gXJh5qZdqhp2
Fg0DK2dk9eFJKXcCSL3x1XYtzVEdLpSt7a5TjbtSxwMF47YmHK01b8cVmh/SgnnUiWwFejVXmCpN
5ABL6wzWU1rBXRxdC6LSXWo4AomqPSvmdIJzcWyfzM/vd9HTOhHyWsowao0laKcok4kP/LN8uLNr
XWeXd3xl2yoIJB4af2Ggau0G4GgonZBz+rQNaLzlWSzs1Hjl/5iIFAGHWrO8LvZnRqDImlNdkY5B
LckKGhy2HB4UXchY/8xQx4cYzpNljd0LT7qUT5Tu0Mdl8o+KffOxINLNRS9LiP+E+pFRd5Yc+Ucv
RMZjw1jIs6Glqeaw8BzW5H4sIPCk4HAnbTseaWTQPwBg3SfqpIVzkDnaUHPzy2NINTTmEa65CRAS
sn48kFy1hY82IDCNCchoiQBhXIeBRIYFfqYDpOPReEZCAPhruzSWuqRYEQ77rnXQ0vFUqWJBv0xH
17m4mbo5FhXWlypffsl4PyM17lq3JoHXxk1Is4d1+Xs38+gPnXGeG2itYpIhFzwDfcg1htq2R/yR
U7dhDjTZzQbKQtom4XaMCB9SPd9J16KkVqAQzSvL2WMJ47OHpKiBR5e18tizF3q6FWzUry1+N6sO
hdC46bKCeH3TEcVNhLnpBF3RqWPropIz35oAaM4VWKPlkWa/S3/LVwieANjO8jcA0yX1NwfX6kYk
pQydSyXWPMn+5hhvvnwp2C63986Jii3cviY4DPGlUUpeshDrNjrNbpbefyZ3CZRELTpklLniYsP3
TisoJnbFbl1R1S/0YyHbhKrXFFyK8UzZ9/xeCuYk3Ov4oVVZImZ5Tm9Ch7v1DzH3KXm0pmGkCXKT
8UUq+D6Wt24GfXr4j62R6UJiGbDlhYmpBSuqc4gVS1G5VoKYb2ZlUZA+nraqVbU6PQo6DhrJBdNV
jQDAKCXsZAGRth7PFj+e5oR1/kU1ulPLJuJpedCeiKLWmfdtbeHgAtci/wvXEneTtwLngpmzR/rE
fX82Atn/YjDIDkajiUOqn5UOI2R/Gkf/Z/tUCSQnjRgKBu+kVxDJ7suC/FqVj6j4ewbzHnnVwBUe
kJLvbt9fwHvV/yJ2Fo8zQjv8mTOizu61KcvJZgD6jF2jirxFB0GPEZ0G0y7aK1o04RwRQl9kq4Rf
5FwOPujV2qhTB+Bitd8OOBwH0+xF7x8JFdT395ps97nC3pnWoEgZGkXHfKrFyJdmSo9RYtQf/TiA
ZZ/hVJcaGJ34MUqz3e+sYJYP+JWFUKpgMqEgIwTRf6pbDszkHTzPqTbOY9E+GiR/mRpm8wWOjK/d
Zw2iDi0vr5HmkT0r3juUZ7sSPa2sWh60HN67hL5iJx2SFQGI9e8rbvfpywjfFDlbxf+02NkqeU/f
NAgNgTpit2aqLlmOl1d/5HvCA5tryKKo9JlMohphA7pWjzqN9fYu7Bx7Oa+o7+f2CxxBzCKI3yiL
PUN6V2KU48BFZlDFxkpoZ1B+URe/zOKgw+DZNrOxu1DCsiMfQJR78L+/BcHUbIaG6pjvDQCeN9DF
+rz+ohz/Mnc9tr2qmD7GQ/3ZwwAKB4LKJjdLAT1M/XQkOaYwE9SFBsz9+qPe4LAgwv+fS40keFxN
7u2H5DLCn1AFLMc/qWgOj9iOLE0Ry7e0A3UhIH2a0mBcJ2NOM/t+ReVKQ+SSdg8N1AWrfUazs1mX
Da3VewYxmgvs6TvgsK7j1ycqVDhnKrAdsNtrdsIwOrxDgGCrXZAPCiX86fyRrOGkt5kQK+uc5jWy
V8WmWFW7abd6r9PJu5819tg+EVXYzhXLgENqnMpCpbXijSx118zkjcWinkndrYDqxR8LU3o3n/Vn
8WhELTPP0qYWZu0p99jGjvuULPzCFNaK+phbI5knbkxRPNC5MAMYUz17fDHt1OmlzDUrfR9LS0K0
3lULvc3ipj4+mQkIEjnV3hcm6TbKi3a9rTw+Am+UqwVovUHrRZb3OL7f74GcMn2sSLuKPz+h/J6B
hp2IbAz/Yzf7PqsR9a1hrlxhr5vRtNaHJoq+Y4ku8PJQrbxnI4HbEE/NJ4UU34vKcXlxU/Tx1ZoP
nyHu5Sbs1cwNBcDIU0WJ0xBvsoLF0u+hk91ksaLdAuxErrw8FboWp3VAv8d0IEV3hTz162DVLCu+
/C07GvuTMPsyRf74gqw3lvSXNXkWZVkP02KSA/+VsMae3bn0hLiblT3omMil/8Y3ZjXj++4SDGNV
MnDUEW9A7zZBRx5wnw0i4ehMQ7aNHG15/FTE6WCZwYtqt63Nz1vAitL5KREh/87PyDtUXTfmKuEI
ImEeLSFf//1ywK+GW1s/FeXwkq+Mh7Skz78dniCLrDY8UFPf+P2B2zBF4edsqJg916aWSFfzB/Lz
UeeRz9UnhH1c1s1z+vXi+u7NfquK5T2Bm8OUSxf3RF0MIam/L3cO+23Bg3QVbDTEHa1kY6agnESF
ffPqnex+r/tE5/zwWYm4ADJEnToGHfW3oIU+DP86GrsxjpwtQCSWnYfsltYzTuGuZv6K/gGfUxmO
zurU9Hw2vhQG4YJ0oCpfKBzMr8lWHSQSWELNXQ+KYQhbxzCEXB2Y1njaKUAMySOAz5yFvdgTdSWE
cUIw2wg3qwIVBJ1h5RckNuh2HjOJyyTN7KXqmP/lkD37k/TBGwOiPEIsL2HGOhBwq+LMBWI0JWJM
u8SXdrmBm5u0Fd3i0nH3Pp51T1QV10NEOwxz7HWjsYc8rKvSv6pz0R58aSl0p3m0vIrvUHarK23r
KP6nSxUjBXEJ9qQUcbr+IQZ6RQ9NPrTBxGw2JgkmTGrfOnrioNihJV8/x7RshUB1t0upZZWsvusQ
MZngQq1GPESDiYeACW4i6aZfHNrZO9YweJ7wBtWSKL7FRbD+NnSLGWOE64H2Wc3ldTX+DCwCzpej
ybsDLyTJOUoYLzSMSVri9ud8O1vkMR61wh4oT/67I5sIC1HvhnQeUIJgyiV+16L1she8PF9oKBsw
J5KWexV/7FewYkFq3CxikOlNPy5nO5NlJySjEKOYtLjuC1wwUVIDJHp69Thr5MA3HLw2jRqO/kLH
LJo3bugSAYbc7Ud+kwsJ8c0UqnXJbaLrSfwvhX6OrsiRGFhBVT0eriU+dTTmHXwzsPzYmFgndvJi
hjAwn4isZAaCfad843hROw6XziQFjwasGUqbIw14rQM78odiVKneTN/HExP0m/J6Q+U9eDFCPBIb
sqtkNyBReBkpeOiJtdtplhmeRz0p5sXFT7KjI/i+L4g3mS7ryiVM+KVKqt5Z7gC/IVazYCDvaqX3
Y1jD/7n3kiq7i0jd4n3EmJ8C5xFsSSEVDgJxcfkzXixcwjvDlkKk5piDikYDUmqBdlKz6jUEq7MD
9EslpaVB0vi4rvtZy/Kn8D/ymjvHrptzv7rjZ2k/xt+IkzGaiOtP7An0WAQOTGqDhPV0rqclGmkh
bRKpg4I1bcS/IZPwQBYbMjt3Yik+7sYVFFMUflVzj+oSvi/t7H6N95tjW2QPkboFOsP6Qcchlilo
/Xv5zV4Xv9VUzGfp4851GCAGXOhu3GyniCI6KuI5W3giR5B/2gg88mdEhRrtTrBPYJ62W7DgD0BT
Uf+Q7WXR12rXtqh+HvopCN5x4qB5g/eJrBLOUm/e0PYKth8KXgktkctg6LWnSyYoVtBwXc7EMw4U
ngdlwOYc5qCkDWD4GNxpFtJUyMp+vEAg3HkLa/9cSWbzm440gSIKgCF9ORvsi+xfYAuzSB8vAMNy
TRBPWWUFk/+PBzFsAO2Deu9DlTHkK9sA/y25vxRkW3a/I1tN4iFHMkMugtfm8Qlj/4d+2x6KM/UF
vJRWY2NsdD2/CuIJ0ZF4NCci11Q992kw5CbrYD7yHNk1PDt8hUA6bRd0p/CDulXZtMKDuWScJYAA
3wKYrG8KQzZ2X2maNH9qY88PYy+Pi2PNy6E1ELAhQ4PiqcqiVuRRWuMwxoftCQeR0fjIB+VPQ5bW
TWMI0pYO8RprMGfcIxfF9R8P0rcuDGL4dXUQPJPTszjNlaY90+9BCNVn+g9eNB/lShNBdqhZMuEF
UYtcZhNCWmFEBnQ6/P+u14f9+yMRNJc2LFsOHBoPp+1E38HsHcd1rz8zK4/8JisPR2GeWbowHQ20
udNdmDfzRcrC3akDUt4W0BEMe5QOpYmuM9v+fKJqch6GwVKJ4iEHQ1HmMTPxzTKI6/Mip2BdRPoS
sEtWxknbHnEakWaaHPA7As2HsoU6xLfSmxxKDLzqLYkivFOX78kw6IBl5cFj1XThLWm27UUtmWyQ
RqELidQo60juDWFnbThtShZEpON//cRQi9EQoO7fFA0d4j+7uR9qp63n6yMrHvi7PpY/I56c/Fez
CK/2T7wQMUmgQSymKvG0U0gaED5KhoQ1emph32VcF5S1HVizf74YJYxj766ks4inTICOTZghNslj
MKJ8tdB7KrWnqZYSNDh+60Xqr0ja+eA8GcarPyfu36rCn2C2vrbYyufzYUbvdDMVjTYyDRTa7zoZ
8zTz/kx8iqzKcLGI9kEh8RHvn+v0Vhf6N2iQqRzg3CiAIb+cnj+hGP8LeJhmWc6dIAyywJht3Nea
OLi2sHMMKVnbdNL2AlRavc263nbS2WUsLSZimffNALQStB9rSS3fadALyvGbXrNjBlwp0CKJQVB9
ecbBV/i8pnjuTii4CCERvv0u+lAVVonysaYq9MSed5cxMARH656CfxXGc9JXwvyPEi76G7/OjDTd
DTto6H05NwFKUdsFbSE/cJB2pvM30ZfXbiozjwTAjDpvxgQE4v36pDZiOPeq7ynL8RfO0bc1aY0d
nGXjILMu00adJzNjl7p6eaxwGiawUZXQUrlWPmUKUmc8zuedfUcomDDHCGdTFJybLLv0vdc6Ibjz
KBmnB1f/qQmB0mb7Rve+AsgUWtKE2VuYrn86LGc9WnJqK7G6lwFDeRMw19XZQRFBov0TwcMcILeZ
u1DWszU67BTWFyTiAloTV9qUE7K2qLY12kjgiOJM79tzvU9+dfE/G5q18AHyvY6XlrrHnFmtFYFj
C4RtTaytv6BBhXagI48B41/+yrFobnu+252aqKqMqi3kxQVpuzo+grXcbprMc4oEYsBGtzs/tuiF
CrKguVFa3v7vdL0W436PgqEz74AucX3sAF2D7AxZqj2a8SfEXdQphfPhCFZvRHo7DKwxO4OHSGQz
bnNBG83GfMXl2q50lQcXpZNeTLpU+G+H0XMmCmmb4NkDpD2jvcJ5J19xhh0rO7j9KNJAPCnY8nsz
g7I1v96KbP+FIRP7W3BgmGnsViZw18ejJgcZJdj4aF0frrZkfP3aSV/Hs3kQ7N0Vyzr/aP96Muxn
bOobhXzmj7hQp71DUiotdKZO6aYsDOi6zSr3HBhFFAJ5nNJOgpbN7pQ/maJnVvjdw+jTzSc6NjU8
tzRmoRDcsCLJxVxEKlnqqHAc8tCjl8IQX769IiKU9FQCz1joW6UOV98rt3WEJdvg/Y8EMSe7QbF1
6LN19GBsojvofueOcl/oQb5WceDx6uYWY3isLeB1zw/wfwmvRhsB2oMYBgXbFpjq6b2zZdlp5I0s
COu0NE2jna7Qz/2SCAMeVS7/ckyiaQRYr/ZUZdIHKREysuQpymwy+bG1oG/Uc5HYth0v7J1yxBYy
3Lz5xXnaYVfKYSVOEp4wLfOA+Bzq9/yhkgGBuCRHSKXR4lPXtk49MZ1lPLd1sVVM9qvneO1jXBte
yF9LhE6S+uGPmS3/83ealC/P22Kqiv1fyAhCZzJEqxADJncRxVNxPbOBqgww/E6SG+PmI3KO9Jbf
ySEmwz+ibqRdrNAy14lGROIytkRrJHcoo9zg4jwGaZAfbm8+0nBoTtp8Lc0w0y5dnpB7HDhwdOww
8pfSd9b9PdVw0uJDVA5xjMh5o7w7UjwhNBPc32HXHUYjOVrpQFcCbdyEjwlVIKcu6PAPc0agP0kl
KCVQNeHh+lsLpWLUipI45DxUu3u8DxqyAj2P92iGRtcHhtq88QzqUB4IhrusPtN4FgbobYoRlXSQ
VLMaz33uEdarFaxdGPg/GJT7PCVdGmgRxJO35kRJIVADuP0cMnnwknUbfWd0WrAJt0CvhdFkmlZE
YCz/imOpl6i6aN0aW+T4ANGDaeiLwRbSlqPr+xpDl5kMdR0tRzVR6yj2+mu4DS6VQsr7IHiad56u
nfReUNnRlUaNsJdH1wsBDTCtslo+RaQz1Anwm2PQHisElWyATEoTnIPWXJdwbfu4ky0xkUTeX0+Y
X+fAdfawhzSYfzt2+FLTs+EnWRDVjY30NoCABfr8Q3B1rKDTSIMPs5VcJB7I2rHMkrrNak8XumPV
lnY+t3kUTQi4t2weZ3v78oc+gQEH57pt0GgbTYcEfzFECdYRZNej6dL/m+3B36PCiBw1Zo4KCiXD
LI5q8pv3sYHdCKGLmXP0hJK7RfPoandEcmAfNcliakXLHhMsNxtwGoyDwPObjFV5at0SgdBNRGX1
1DTi2gpehy4ESnjuKkU9PJ8q2WuJBfShca34s0QbTiG2dF/1UxJRlnjycbsAB/vpboeR0AwUegyX
6nHfEDnHd46KBatcM4KSAngwBgcxw06gSr9fz8NdcnkGlg6tBZWIHiXbkSpCIgLZYGf00aS0fu8j
jnpUCt01WAe1t21QMgyCJ8ARxn1AP5vThZ9YmmEywVReu8ucgyiQlwKxZQDjXJeIGIUp6A8D9ZMK
kdXVAZPT9berYnYaylKpQF0NXVLM8CEdVTCUV+7b8I4eEdPb5FrUY4fMjsaK6ej4gXguUuNgbVDG
HGBnDAIK44W0BQwoG3bNOa/FjnO5wK+CTO9ZlBf8QwYcyEM+JGZhWchy1ojvBSaGsI2OBKlPHReA
OqqLYedNmh54TwaaW+Y2sogmMjZyZ6WKXdMe3W3wLTZx/OE6S6aXLZvqLFt0+WEZ1b5/8Mi0ZdGA
7Z8WXXItGgKYI3Bs0xUWW7S5XSq9GLV9SVIHMvZogz1y7KBHZf0RmyLZjIrs8d7pxQnO2nONHT6y
pTE6aQXXJbeam9cQzVDQxJ6Kc16UsP229MdCEInxPLg3637aAvCoG8yZKxard4ni9YY9mwj/Gvro
7r0ihfN1wRfMcqj3FFX2MqqKwwhBQC4C/lQ9DxW89sEGkwAs82+VKHBP9x4nd2xHeWhcxU+JEPd5
hNSwBkQInqM6om9X6vpJ8s0Z8mzticleMghjAckN9UJBKTQqyDtY0xs4nDKu520tDXzF4kRR3dAu
gQn/HaCOeygv1qTP77/w2wXgMTqmrB430hG6qOHHR6suadTB7i4fdPKWBeoHpOC2NsSb/jH7vYbn
Wz/IzsvAS/l6K1KAFvhNUPtyDRizE7Sn1Defp53CHrrbP/uk+kARIJIHs7imFnfvkcKaInbQuRdE
8yX/z6vT6BV/gmr7pI2HctAR8ox5Dvcm4kGUxHWvqxIfaRbYIBvMZgFk/OL1xjzCsWkhyxF4Gx/O
nY8hd8D8BPzT07g85NzAytCu8hvotstr+CNjM2ZzqBL09m53n3hupGC88j2jZQ4l4TWdK5FzVjAz
X6UycoVOz7ZHYIoC2jFLXbZb/hDuoITvsYjnaq9ytk222jvkDeWxcNhR19ohGEHE02wEEIC4ds7V
L1k1MTSgZDItDLi3QJ1Wng2C9vxt/0m1o9qG4Q67+szrK62AdV6MckUAY/1Ap7n1xdBsTarA4e8W
0GdBE7clbhd7zRxyldl7GMiLuY3uI1sl8bK6gWwYF1N0JONP71OaNcQnqzBxpkT2wL84BWUNGLhP
V5P45XXHVbT6mEH0r8r+cq4GtmXiGneuqE75ov4pcuMgymbkKe06rIXcEPUiaNp7tYUvKj2ujKDL
4rpXki+SsAfxNvf2Ihrn/1HcXw25czFzHg42A6dvH6L0ZOebgG8OmFy9zlTo66t1ZNh6ml7R08xI
blfoHhr8I32J+sXcIQUfsRSaFpzzS8d7gW+kotv5h5iSkX2S1GqW6mU9HzILtraC8DuESsJU6juq
kfRVxhGM2QInjntcxt53flS4EXLOAM3JPq92+1I8qmQ4qPgdOXRF4rzwPATYflyDmCnG011bbG80
pTpUYY3rJDu+/JSNXxcAwa0NV2K4q4MwSZgx810RhVT0VcM7IHlU99+uEBIOZcu7jXIY1d44f3+p
71br5c29rtf0lCwp2EZR3KqODxMIZ9gEWvFyj6sxQoWeSHMKD1POL52XNYdy7876Supit4ArYHyt
MgbFGxqDUIv/qa02JNPalejaqHF++CqK0DOyReP5aeYZRRptq2MlMCCDAi74/TFJs6iE0XaghrJz
5sDip3ID6FLwnzS4FbNYo5eZdFOANxdqQyDnjLvaAPJ6OwpmWLRlo/1leC8a/ChSwDt50aigxfjO
IxxMM3hsVVDEhGGbTgl/ehYOPf5QPL/+O/Wn46vReKkUCxUqAJOoKWQPgv1ltrhtMSy3fYy3QDyi
sLn4JskAdqL1knkRj8kw/eWMphVC4NxPGWDR2TnY+fAcdZxPPF8mBRtXYGDtUTs3ADynW/qhnkKA
AQ21K8A/BhEpVpIRTxW+w25wZZ0Y6bGjzdrAk4ok8DYf0fKt1rNWLKHx4oQI44UpKH0yrwd7kCWK
4Rja+ODT6zgOxa6+FUs3R0+fNGzs5/OlDmtm2t1YH3/iHKHA9k2FeaJ3DZYiXxgU/lOREA+ktQt4
rKDl14fVYbCXXlDN8ufdMKH5plKeA34OAVoCTVLpmZpzwAjFPUqvgx/676QFtfIDyLCkCFgYI5+g
OHo1B2Ex5ITA25R/fQZjlfzDFeB3qDX9ckcOFEdjq0v0JWtMfK2EeW9vmkKMzqBff4ZYoP5f+vll
YEgsNSfHWkHXWRdqvMQ5vI50nRwH/T+utexEJFEirc0cExX01jfHRoUQfCCf3cdxVtEgSHqkrqEa
zhK3mL41f5B8u3eg0KLego2HF5bVfOJScnY4qMy1rC8WHSNJh/niVkw7dEBWVJnf8SL/CkHK5AvJ
05XVoGy95kQkOlNg0Fs1XZPaexlWBmaxwbw+CmcAf5XcvApx8Mfs4fF+RpUBcmwYETailOCOy8Z4
1F+adzwu3N7KovY8LDpI+a6Ao9wjrMpgzQeX3GryP7ob4Vc1lnnrkvc57jx5zGiKf41V8CvJpVXW
vlNO+lNce/r3VXxC8Acqa9WgBF8BBI81Oe3lI7xQJVNok2vB2onULH0UrKEMcxW+D6P2Hgzv+OV2
himVkO6HcogJhTQIHe/VXDZoAtsy6fkXY0eyudGOe+aXSgAF4Y4EgwLrKm8mqHLuBs1AIWjjbHXS
955iDB9TfCVKWgWdP3BOuxgnUBaz45WGpTGZIpgS5aDjDxTL0AfJWnOx/CA9bfJ9m6HmTfoaP57h
AQ50BC0/3keItff1gZBGe8hVT2KJyBeLU/dRzj9RXD6xsx/fP/AbQ2iy4PhfvzQtb8L9tcYTZrKw
HQFCUStfnRbgNscgN+SGNPZnxlg0uH07xvRuaCA1uCJCGl9ejPRR0PBUk4dDLw40F1zPjLA2hB0f
l3NOD8vqMlmaoKCk1dPeCTMzyQNtqxSgc/M6fLVxfEtCEXtix9cwSi1hVqXJ+WJdcvrBVIUYlWqg
SRsoekuM+OMapI4mJICrEeDdynw/ySWwnXvT1Q/QpIpyJ/Y+yqCqcRXH9pg2n7nzifceTOnh5a9d
gzvhpZJG2Y2n8A8ARiLN4tLLaLszVHZim8Bsm8ChPBuqRrVCss+hU0U62csF9eP45x/p+/Vci3Cp
z6hbavN6SLyZzt8NedHlgQuDnEHR7M0Z1y0U9MKIPBLPdsgFg1Bv9+Azt2TYw4jHRPc6u3tEs3MR
BsAHDY7lqYVdnt7IEQnO8wf8p3kkcVN3cqswb9U6e0OUIEIgwr7qqMQ5HcmFGN43hW8cs48uKfbu
vEHbXzE3LCTn4USTsQazkpw3Dfg5NKNIOsB6M2+IbMETxzDc4+Q99p2lr6tldo2Ubbkhb5Xvztwl
4e6Ya4/BUy3W5MCLDfj9T0M7uidi2zBo8aT9zHSicK6jxM60tqdWJoTsij3vaSw50UwPaYBoHmMf
M5T73sT96oPwMx1MEmeQSSrc/oO64VszApDnqWpr10IDGO51eVxN4O/DkC9baEcfEFV0FuENAEpY
xcZbujloFG3OSEBDS5/j/o1T57GGpLkO152zoH4sDDvnRWMSZvV4Iik4JxNbLchW2BqL7kbjmQ74
G18eAzd5azUjkbeiZTTgKptVKsV7cnx373rstTBDf4QjWD/4UUFXNow20n/mEPnKPwtHrdx+XnBY
r6UTkF1GY6qDNGNi0w3iwLpcUMfgEzfXec/jM30Q51S3QoQj9/C0QhnNueu60xsGBgS6QvJhNVzD
Etujm82meYglPirQq6US4+oxk7Iv0b4cDYqnYDR0AvhQxmHFWPtf+Ed+NcDXtFt9SHuBjBIDtuHL
g7tmIheeudIlKDKpj6nxcU9Qd2cBOAPlBEuD4clCA5kCeYsq+FQ5cH0yrVzFPRxKzgo5jggKDtvE
LhnlI/nNajfHOrYFM2tCXJeo2nxs5IYTMYAWmJSh3lofFmCzrbCSMVHe0mcMfujFtDR7kWVmY9g+
38kRVa2kiNPYbdHPzyd4Q8pvkKpN+pSTHNESob58CDYrO3lv1X6kHPYQxeC+zr+U3t5yMq//e+G6
nbJq8TfOMWEmjaQWkYwZ6WcxoQf4JzhhtOf/scXEDgjl7Yfb3JdVzR9dS6aGFHeVKMEKw82jxgV4
lV6Y+VRl2y4Jgo9UVFhoVAU/9vafZC/HQ54FoOLBK35bKmBRMG+AzHqcj/XtDuepetm+4NAkiliJ
vcJhhD9OLV6LIvEUDgcavau2vcIU9x+SMm+a3SCdnX6SWdRbVa43qF0qmDIPQx7qa5fjusbbtBKD
Mj3K0asm1qqCsA0vBIwTQVsR0Q/5ulPwBPzp7fAx1SnTa5yr7HUUBxgyq1CThQO5hgI9dTyxm0g6
jkd/VlwlfxvDUBDyiusxlacx8XS1yDt2+fXI1TZQfWnZNphbjlmK/SPybmjNnd+js5B/yoCLkbpQ
4WckLlF5ZaQY6Inz1xy5f+6dYMmWqTn5bBBY3cYJzMHLFNOr63nrke2n1bPfpY/phzbRNLsh1etN
/ANvMt8wjv7QoqsWze3G5SImziN2p2LFS83eg7xzc5tePm/txXWQbR71yCTvZIuQ85tfN8/5ZPf/
achJeA42gmDVBbBSWn7Yzoai11uJUwZn6KLtAhVWvRDMIaFY0oW2nfQ/5IllwahmvGbw7i2VAHgu
80lf74xmkrs9Z33o5+9CTLpVGPgC7jvjcdWzxLKXwSlsLKJS/b66tDOEhFiCV8pml3MEEyWrhnMY
XWCfzKvoE+oqT8RZEygZ6SchBInVIXK+dZBog1xa7eWMfGkvCoGs6SJrga3rRmfDfK8WpYAfuyvw
Snli2rQAk18TJS2FG7n7/hbpgSXbKBkHyYD0tanzx+wOQ2K1Yfq17alaC3rW8W8v03kq7ygmuvpP
GXYQdZBZIeyoSDgghFzTDDtI9AxsEaRlt8WZ0sfgUfwWcwWz/OB9hmjnwVcrHHZqKc2JpHQ90fbu
d3jw63R/YUK6HW0uh/1GxgxLD6FtqZpy1We4PSPjSO1gzdFK8qC3BRiHyZYtQ9uuSKHCYpmdQspx
6jq9IvpO4dxlzZE4iOHLUpk3wz/6uUIMtfd+YWpe6nGw2Cu4VSYqXm8JvlN1Uqck/fTG30rDq6Au
85ho0rGmcT/E3MRgYrtr/idsXjkrcx/IUeUwBHrxN054lvsLwztRrnpqb/5FDJnWwSvZfOkVdPBu
G5GHVEN1NFoa4Ah4eyAwjVA0KfNBMZmXw5V8o+E9IzB9vuP3MAsip9Cyh9pepkj3ckjI3CjXTSg6
oo9k4xKv4PoKfFZAqSxr58/TVBOEdRTrsBW4SV4FjWWcaVqnjzZNnZUhSHupFgqexVv+fzYaRL5/
bayD3PTkqx/mDX9VR4CsbOCQhCMASJ2dOFDr7DWb7ba6b9Eh5CVfEPaH/quH0ifBT5L4w9S+LPIJ
QFc0EsvDRUT6FgTdc+PpOwmAcNTvbPEFs7UbDEjvx9JuQn72GMXgnUMPGoDnEl+zArnhdYOcbtDM
vL/RxybVBSJYj0GpEP/TCkqUReaOYTI1HxN/gfEruLJIchR7SX+r/TzQc/8MNWKl5UgA5CzvDvIe
nbc0EOuBwUdqcLbeXI3DTTexi2ugGwzlI3zFlgA0vvK81EwcV3F/YavEhp8EzmykJEbk4D6krw3X
/ADNxKufsRXNRP2qmWUAe09uW1GQZHF69cWF5gcIanBd+HrcXSBowMRLuV2VKjn3xfRVsLLXh3mi
6TFJvoXYcatHQSSFdzoji1iogHfaFqCxHtdwHEaE5pMCCTNx5n6y9VbWCdUpMcW5iNAVkb6NpwGe
tti6zaLl/14tUryTBXFnacYJZ7DeYit6mDY+5gJkq2++lzyeca6atZ0cOFHvpeJze04JifwXSRQz
If8Pv2c1H4sygGDSKRojxsq4hPnigSLNOpwvpkmui9Vd0STGjPjdX8AEK/eL8YiB8F/T9+iJ+rga
8sG992VzW09nPt3Eeg1ZGlaA4cXp8r5KEpYcuGKePoy1fR1FKXIEjl446OBnUvo0latPVFDuN3R2
QuDvZSLzHdLGvOBul41n+4I59+bXRiYzi+IR9oK2eOkJmvd4s2V4433MZ0DOU01svVEalPK+yFEd
j+AveZIpSiPewdB4igPI0Sw+Xz6VEXC8cq96uep2HSW2Z9E3Y164i++Qc+Gzv654qVyCI31ZV04R
ADVFmzkwREE9lxmeW0+uMNm1uHmHeISzzX9tSnREKUxqJ20WYaWJRp4MIASjrDlIdJfhU+fSRbJC
GM9SpbzCiQHae2LV0IvA5DgmRNfo/OoWrpZS8UfMrFXIWYmkJmkhMGxlnbtwvBNdYR3Ew3cAW/H4
relakm+yIzujln6oCHpor9ngOACyW0cZl4zpURiCqLgSzFD4qxLle/kUAduRwSg3j79B143lxG75
qoMMD+cT6SmPJX4wL+vG0vAZULm82KuLNxE7cB0zYPhCnAv4Hs38SR3oA/xwT0QkOjHsocEgLYMF
XjE0BP3ufhGx+Fes2Zu0n+S75jEn05JCMV53hrxGY2fEQwx0vJglqAxXa8xzOxr83ecqnzdPWeW7
VTAd8cYWsU30Wv62oo1HXJvYUYuhTDkCMqhRKl3yAIyohykY4Z03XDp7q029Ys2sGjAmCADopsYl
mp5SBLYe1hJ1Hh6lXqHGPntKW1s0dmXvSObtoCbh37Zb7oG3zQtTPCQ44XKSlU6ZpoXGl4E8tCyd
2SapxAVH6YWcfsFEQT9RGcaj2SDBhFRqPp7eD4Z0oOXVbuY3rwxjMYc2dgZHxX//3CKTO7eHs4+d
gpk5ZwqtSH8rfMFOwopZuFo3cpEqJVKoyJ90YVr4tezypDfX0MzwefeOiujEwzH/2+haatWlxZY+
/FwgZux6wUhVvBsDMcKrrnRZnrjb2if+c2knWCxwMsrUJBp2077TI8cdMLAVgyfEt6IJbyoWEj9a
7sX9ijkwrDKTADxclfjKT6GDYld/Lr68jnd6URkn09dFKpIjWmd3285PS45OGo/TU/uYlpHiVTJI
khgWNDFNoK/CYtyHxCCKG6Wxoz2QPtnWJQO+bDLVlEglze0+hnVrUaJEBMc7iBAiRjAJode1mFcF
uT/Q6DC+7QFgG4IBxpZgpd7fWBho5K5gX6EAcVrvFIVMhE3W9UJqBOpzLLscUXWJ67W/AXhNnKG2
w+Pk0w1saihTqE+6mjV3ASctSop8ITAbfsAbssYt1u4Km5iW+tPQJI6XJjrgXptM6rXKpvdeCOTN
LGz9Ii+etRC/xZmArk852wbc8Uv1PwSAy1fDj8OqbEgKOC1OFLwwtyT8izfVhryqkOzWZWVK4sNx
ttnux32dWDIi9mZELuwW5BcPf7/GGKVZzlIuUFZs0r1V9SOezICRXx4+nyORL0FkvOXZviDaiUoz
PhLzda7Du41CN5CDUJDjMr/7ZXaromnTEbDhgnnOZJxjxpISkghST5FUn01mcAXtetzv6imlEn+A
4RmzgCOLQTrXnC8Sf+eotK5V0Jy0+iC/T0PsuLtPV8q5hhoEErREduEKF52veNdyUkVD/qoTfsK+
xO/PdLyCOx7UF0gNVNRPcB9U+E+tmvjmiIQnlzxKaFdqQTc6Xic6Uiy2MRmBSniD3xtLfWSvb+oC
IS1e/WN3TneJRQMG2HTonLCFMU1j+CEsyawfn7Mkp1L/0xWpSWZ5DVX5iO9esA0V2jye30fNrqqG
ICXFc4+nOvSN7IHNHNZwOpGDs+opXW0tsf3T3Zg5XlVnnbBkj/CA1jU6WcuaBB8xnR45Qa/0YhTA
VEB8IX/vKjXQrH8zOEr7zPvoC8WjpZ1Six9e6KHoz+CgGV1CiCx7cLo14biVCXX3W0Ju5uj0ZlBY
lARu2g8jht2gGui7DDoFhyTMgKnUqi+O0L18W1Leqw7i0LDj5d2GmpTijJCcK/lC8niOWM72hCrT
vzsibtqQAgYAzJQmyL7jyET57Xkv3UNjC88x++UflZrOMCVJ5rTzcRMhdX1MjrVuKtyzFMMAlGi8
KP4dAZZQngSHQrT08YtbT96shL/ZEHLAq8ZHl0S1BeMqK/YOuD/0I/bXCyJ1C/fVJzhBAyATLung
pFnHcHCdgie2D0Zj7iDXRlv3AbnDit/g0qIfJ/HCmEvL2/LfagPspZU8hLg2XOoGGkoilAmFYFzu
0YZ1KupAH82PaZJ2Yni3wxDZFb3MbzjoFrRa9LfBVd9edregyfjbQKwzeuvJ+LC4pIITPNMR1b7y
bTZv71umH3juJbgCXRgQcmx5q6hq52fcKAvdi2tQ8ojkaVNQZQvtnYrAy0XIKm1luF1gMbtDv47V
vJBBIe6mgYi81ucWvUjWhpXWwyWNCOzoxDKo3kMSZQn4E6/sPZZogNuSveGxZNoSe3r41NeoyNH8
xL8dW+OGixxn3zO6GpL9KiMUulhBeeoT/MX+eJGjVsMLd0GAWYU8uH/yksGo16grt1wWZx1+ZH+Y
EBqBP+KqkyWFWCY+fgwLEHY7vIOKg/QRd6275qWcAT98xO2tskSAVH3mRAVxcRiDNXxpFkCzqJlb
uUQwjPiRSavDJgk8EDLowU9YKZdltw/WcdPHfANxoqUsVW4sBgUya7dJJb+mprHnv483lq3lT5NB
xSHlNtIM1zqrpFmim6AOv4AvJZFF/EYY+6oGlI11onUIebjwjv65F6/EgYNo843o38S+WuDXe+ZD
EEkI95332sZvHpeZKarsx/CVRY6aMWJ+00j4IJMKp83VbgYnmhV3eroMpt+RkDsmy11TrGi4Q29u
sKTC9ft8IBOFOnJuZWQseEndz2b4uzFr9np12mnmstVeDn5uCIB+NY2JtwPSirU9ZrGdUXDenNVI
pfx/ZJhbEDt/8rvAp5Ft4vaBhdODbYBVGcTXWNlhsRP0oLYzb5uwbxx/tCPSpBaQHIe7yoLxoGQd
NANzIL2WbxAHWDVfj68XkA4OeYAHC/uqjPjzfU0N4vkrKVTgWTGGi4vYPzDJNovabpIxpmR0ZTKe
VAKJUGVIKzOMkXVwsB1nGHRu+7y2LvGCBgg4PuD62Ez/j9XrEgpnZEnTALhDdRuiMy8tvZobFMVc
fwcqg+enXOyMSf6Cjka2GeNRbRUNTo4v4Kj3vahFMf2AXxbDqkvXdyMbGp3ZLET6oG478zoQ9Fxh
ZBXh5bXWwqLVUVJr2j85gDT6pouuZhZmw+0Rl5PcGgRjPUSqSqGfuJ6b0BUGDGW6RwxDXb0w/pie
0ofH/ESBMGqKBIqZkoQD/34nm7R9QUceskO9vhiNYktz4Z14k9+ui3Oxut5dbcXe+9s7IFFj27X9
9Lcsyxz8ih4xDA4r6IQiKZEpQfAtLnrqd9STsmdMKTTthz01+Df/OxIVjBjkQSIkzdSkTf4t4x+J
znFnWhkfJ7+TIDgXEig6qshAfLlRZxiBs/yVBH2evb9pAuxBtRELOJ60R4g9lpwhuYaZCNP9vaE7
Z23URrZuaomy6GttdqRd5jy8jMtZEnDPKNO0Qz5lFjgzZSm9p+OGUza+vkVeieRQXje/tmWJubfg
m/d521XIqtNmWdXHlrgwKKyyWb8CnRcHusKTHoFMw7rTff4VtQSzLEtbXxlbgtHHhmVE/kQRARBZ
GD3pNKUztjmV26sUqSHz5WCMbF8xblTAOsAjxbspRHtrizyBTsiWPNei0/Z0MEpjh36PwlwrH0Yy
seUrSR5o8POZWO2ogRX7Ts9IyIeFrb/MvtxzEahZKqo32Bow5E4Pc/7JblJuHyl7+qIEfnmLeKCD
UXpjjnAf4mwT2QJjsNY9ik7pkoxg3f0xv7GAzAw5GNbXahSZoyPkWg4i2ar20/vhG4sBtCBhsGcF
UxwVfBIdqaflEA+G4c8GwMni0u+Cu40LE3Z1i4kS0CS0y7JG0SWFsF+jXUYvr/JfmZOE9CoXDn/O
KtpKGEm2GxcxgSA0uqV9shqhPX3TfiiUiAv+93p25qKxAcKScr/I9pywF4+aT5mVbvi3uzIRaPRd
g8/RjT+cx83o4eXHtHbl7RvkalcG8ZSxPyrLTG+Hbu5hUg7vyD47zuBnUF9vGgJaHsuOW01ZhG7M
J6Fz+fnQi0OSNP8aMqtGxbaqzUvbQo0sdxX1wek/LweHYDK0gxHRpfA/CpHKXcNdXL16hHAevoJf
swqg1jKlcd7HQAan3YyVU+Cbw5HgfU0x8rpalCKrlm6v/sUxSiOK8mcOiYmgJD7Fd2kCAAM4Zwxe
q4savYKoipibp6bg3vlhQmJZbNuseBtInmglC/gZkjvsOkk7XDBCtJc1bF4xndv5MuZyvq9f+Q/J
+GvBIfmvurJLakir+Ll0RytMoyOdxbP1/PWPOuOiKPkKyQDcabL05wa1KYNyuGtS47TWEkfYvnDi
ZnjRi72vXpxHa1q4kfUrzNSDQ8imVAE4AmBqNTe4p44Nr66qMmMSPRGOXCa9a5ScEGsM3yGVFcmw
5a3iYrKIBpb4abbEW3isjY4Ju5/jj+A+EgJw8XNC/WIDrylvbk6bRmYUOuLqnlDErRIGykBcwu4P
5wlWarH7Yn52RplK7wPFcJMxakelQfIlFLEp/cY4yBv9UAA+C7j8+1DawmE3/WN0zuuRKCFy40hP
NmAyYpZfrwVTgrRb9fuckUsRjGF+blFecSRe7DBu8+hRP/61orww74AqUKR/B/XMkV8YA6Avn+5W
vjdZSxto4N8VRUsmlxc9U6Ct11e+H4tLi7WH6Yi6lSLzpPcmGxHXD5POdNlPfvPdg9qm0A/mkgSv
qXKACVW/ho04QSbKNlaT0lC05ZP+7SIGpkB2lDUfQ+9oHTPUKKQnNOXVMxRk0d2RbW1Fu2ON7grY
hJ1ysrUvCDV4AJT3E0yZLq7O/nx9g+OG5eQAjicSPIHNgFXWG4taMwMF/J/++eCOv0RvXYntACNg
9Wq6CbCHMKQBAQNpoWqHPi+A0osmw5pOABXlTsJ/YSjyYLKvs61d2fB6lWn5ijufm733G/PO1m8l
eXTmNKvPltKDYVoLeR6fdi0fSroRLDhZGOdJcmHiHUFz8R+I+9Zy53qgl4eK00ctt/Et23TLN37Z
EctyG0jadp47sLdluazV7p2RZrwVZRUwsHlVgMLaeThxN/K75wiO3nrKbrR1DZf/P/jtCWzdyMCj
aEbTx21ofCmO8mnH35ioGIklTe3pXXOg/TEg54GhMACBD2jqComm3wSKyGdHmwx6dHEl8d99mcnC
5BcqPQw99NJH1sjYAXwxopCaOULnTFFxEm+ljmOhLE9T5HNqTbjAROUJIfWZ6dj32rES1ZYKJmSm
5IrUA/OQB/vCgRG2dNjwozZdAICcBgS3TGgv3jKpKCJwukk5OYKD7jZbTdo1SsrrvlNGTh0cMdSo
23WoXVjL764+SbPpqA71KGBhnOGydTOAz6qv+YbhxM3N+D35/HwjnTrCu9p5H6x+UfO7JfvdTZoH
9/yJrFlxySa2aOUQID7TJkNUYlwsAN/DC2DoXemPfFa1wZH8hePGmw5lvWSJENp6+YW/oRCDgvfH
YyYA2RbEDJvcBM0peYBztDzI8F6YIbxylEiNCWI8kA4diOaYzTO2T/cPW+P97QATqYbpxqj1d/nu
deMThdtVfWH8MUCJ2VACjTfZqC837R0aOTAuWvT3ptIj1/XOO3Hf9wBRJx7ZKC6pXz/VebodZ2By
FOw2wZSoEUfSmaF41kTQh7RmELhGmw71qxP9B5incn/PMNsiiM98rAzLYnub88o+owePV0oL+xjf
f34VU7cWJsRlPRD0dJGkgoKdnPSWpxKiprDkx7Piu7iFyCNclAXbE5CGqmJyIxfKpneMLcrT/Wiu
UJZ8Ks2iR0szI3EsTsZPiZpRjj7lIEtD3VvkQeCZ4CoeYTp5vsu6Nc+6/wxqa2acWIomiSJjKzZQ
CPHVhopzEgeMG3ivu6jf4MoQI6Y3jHqXg5+horsnxnZgga/pJQaNzHQh6KFcRgjDWnImIoJJlyll
YIY7QxdHgG4qHQ4o8FmZy/s4ioO6gXZB1FogMU5Uswu9bTdtlt/VkosqhQzT0t+CZ8Sk/zFuyifE
m2mxtJ7g7H4oSdiucN2EFu8AD4ux9m+BRAwNZK6KL4M3zrRpoUwCI7bokvvomxWNSzYUq6MHpqk7
g3VwGCA1n0dNkfyY4LS+Fj9htVA1kEJjlQqQ2uU0pR3lVp1Wn//biUnvsj4uS2iMXEnmVw0wor3u
j5OQAXNRDXwr2Y493IXY+lxd7rNH0dc/x5ennCu38ZWDOWC4J9jaNWcCcAVmC3q0dZeI8CacPGAX
8/iWDUfHwCHs3ZCAcrGB+gMsXqyPGPJvy7wtX7ujQTuiB9BScwN9fcBvKu6fYhhIFw2dbNNroTCI
Zn/JStL13n1SlsQMeVAkTkMIaVzrOzvNkENYsLObRqlHsGEl1QdCg8l/ZBiJzmQez25F9XLRB/mC
QtnhPB+NXOn4ZJISsEfx+4yJrTUFWarkjRPxsZ2SUJr/pu4S9kirVdzDAj8+gsiJNawjvCS0a2+4
23C/rZxHvnx0L9VLfNuohuMI12QCIIICou4S0psNhff26Ug1lvAwfD6CNYf3UWrDzVnvTsOdSSxr
CBFrDzupBDOvQiTszoUBAxJ0WtNdzA5JPCTwO+DOilhPnjACtC5BaO94MpfxwfF4xQlC01aZIy/z
w/SYYFEGkT7KbccfSGgWN8+oAit/vtoPaVWKLyIw2aQlvUuI+dkO4cCjMoSoAVWOJKnc8dSmpkyE
9dR5pT6nLINYeCzi27Q0XXH8P2uKxYfHRQONg+cpHYlER3D58XTdXzWvw3z91Z/GsajGN0XLteyr
p0X6CVYMddWCnEixIQCDGZlN2W3PNYhqpuYpUTpUhldMke0baUzJC4kxY3Pqg3MY0RWHGsZ75Got
8+EiaEOZJH+oNuoEzbpdM9/2kxvIeP+QqIx/O9BlnHCD+jU1iG/1d5Bs6nOxyJXSnEm4bIf+Y2+X
eyvxkwbmyWEHa+dY2EQhi+rOvcIdUdJxepNwa+Q3DB0YAGAn0ZUN04y1nXyYrUIyck3KZ/CfCj0X
ML6ooeP8WHFE1Z+pC+O9Krm1ByXruW/SPLYidAs9xl/AGlBvE+r7/dvb4TfSlvNXwK2J6su7Zp78
HBwfjuIdS6cK1WnWAe1ZwsBoXKDHvhLqJw0XWY0LTbrlTBQnjD6I6Q55H5dHYGoGPl7dXQ4gNnwT
Ey16y7A6Pk+BmPJ7ZRt8IRqDObEvGF23PBmExWQeAMVWCBcWpSa1w4e+6rIFRKKWCjds4jpG7Pfr
/xsF3wMA4fYxffI1rSIPlF23iJKg2rtRPrqQxpTvUgXAtmdxTt+IIRiL40WMLyHCdUUbbOc3ZXRC
jPK+fnmxDicW/LRmUVc/npAx+ABCS2dKiCcCD09aP5+NSIa4UAVNNGogDqhtd9vj7KDj6O0OVu5Q
cieXBNgoOcg2XYpRk+HBEFA1NshxqYcSX0k5oriYFMNROgdo6gttBBEEf0mollk3wa0wpnXqWO5d
aryrIxC0TU1Sc+dWsrJB5QH1m7Ku7tVO4A0Tvofr8AgRux7QW+TzdBXEtFmNLaSgSJNdQ+KurAsR
U0XmvrCs9vJxFhWv/N2HBsHKbURSfdHBQI0ryc8jGZCWxENWk8htOaKsRrDrMxvM82NJmG7edkRR
L/oBP6AS4FTKgyDoD59LvYAJiTz2pNjxf5RLoIj+tAxC1GWw3yX9TNZmSXLx8lm0//FZrCUVHAsK
okSI5/xzmjuKpLsYFS2xmStz/8CtJNLh86b/j22xEe6H6hpWh1qzSKYYIHxspyPos7+WafXFURZF
+veXFplYRjgYewVBdjTUMbUEKnhWwZpc5K4Q49rXs4NEOOqQGfNBXBFOgVG3T5ag20DQKCmMXDqL
RyA/CII18g4EYlvtkdFOwGNAQ3UeujcDgeNOHsNZRVUHwUa/mdIOcCfnXyPgCvj2Ogu2h4Ca2Oh8
B1VvYs4cB25uMq+gThet2tMFeVmtRzNt+FmH6OGEI7JvraNPVPxCyEcYgEyazFy9sW8GOU9FazbX
OefcMd2tiCDxg90KPT0PvhvHrL28MQ7iNpZwaod96/mPPe7POKHEqUTeyfzlu5+8Om3GbPnvx1wn
IPBWG2n0Bh/PLFR0F8lgRBLc23438fvAeHpbaVYofitUzG69mWL+TBKaGjncPQziy9OXsusGkt2r
B0SW9tDODJClKw8R7O1iPByIqzV522U0c2fk/wL8HVUVKvQD8WuIS6Jv1uTbxA0tdSgSApdSOktI
6ElvsB9FK3HkL+omwbyChhyJOGLxmYFoepOLN0L6T3xzdIc3J/UEaXZkg3gUu0YK+oBT1+TnWhaf
7/vz2eHZbj6aYIHWvMD9SH0IA7lzH4wZjvSi4r4UXbMQQhrssKMlU22qWAKghCs0/pf5j7kvcH5J
1SiDrSodTqALY7yGN/HGz8C2FrwkXfQ8u8dPqaVEr1BE7XHS0agMkrghcKPSVJEzkOZCVrmiscny
aeakCVhJefzSr2kB5+f4B9BpCMJ6y0gb83pUYZ6Fywt6tjJbur0ZJUY8hjAS4Yk4bGY8Qru9JwY1
y9pS6WOc30Se/TUkWJqEPJWvH7JJIC1OaWI5sGVrNnQn7e0+CG6IFulIDME54a2nwVYbAWgqaWIY
yT1S3kSmoVLHFaQ9JjhZ/QAPS5Lg8JTbwwRT/TO/IZaCblQLj0ZAghNHWATCM+Oc3ek1kDJ3FwO8
ImFnt534Nds7wCgyKNBcus3N5+KA2WztJG7usD2zHjp787+bC8lDZqeUMQYSqa1LVDatwXd9PEzK
MGzt1ROqpPBfpjJqZFb4I4B1oSOXfZjx+78lGIhqdtOCBLXyiYfSg/903S0k/1mFpvylDuqq4BgL
ezDeo9joU3PuzYt5IoJGcpK3onTFekfnmfPs2LjAcjEkHxcabJmhL+XJsYbqZX22APDlsJYuzZhf
2r4ezXyREGtHQ+KSN/XFRZdw040OnRxFFEJz6HEXM78i7ep6b/VXX1M3+nlWkeGwj2Zc04D83ALX
wWnj/EcZlTn5Lbo/bCTlmjtu3SzGZ9uNTzh9bOvB4cyr1R4ASeRIM7iZuIeloxooYcsizkiWc7jN
8E60oYZzfty9bTwhp5ui5qJ5agWwde08wIFHnm5h+nEGn44UIAlaGbCbPQgFOyFeAgNVHfiUIKgP
AnpMMRzAAD4J5GsO+jAmv53TWKbWzNhhzbm6tIRmD/SGJ3MAO1otp43/8vz3reRvquw6uNC8PMTw
YpqXBfWgNJ1gWq961bC0h3tImm1OM+Bou0osVtOSHsIECgh5UU90MWhQe9Jg40YPW6MmNg7Cm9ya
zhviKLMlRq7B0WjmsNiwXIvlv8BtscOtd+Nj+jIRcpK0SnKbVYeCh5CtxCryghE8Z5a7+wsRrrKE
HoyfJ7DHpLZS08FFdMUeF2i+1l2gxWwqwjjVVLq+SlnmirNy3F+jSrdjyrAGNEyYVwLLuY63Ds+H
J03X3jrPBf3693bHDb0KdRfv4NsrpZLOFDmeUrQpsiwaVoS4dZX71GfFcV9g6NbPvOyGjJ1wZ5BQ
Djdm8fUU/bOaIsGZqG/aNTQhA3w2heZS1SGXxFHEbPZ2iBpH8Y0BPK6TLL3w45RVjM7NgqKVk1Wo
IbiXsbSYd/uvIy70NnnBkEkwCrwEdn8/JPo15oPl2J0o/6nkdMOi9s6rH1uqlZCuOo57+az+mfWO
ZPDtwU4eZdONtyiNcAjxCqcAHD8bcx6eAix73+pDq/JoQt9G1F+TlB2KkLwko3qgNBkEw8dj/NIW
c59dukdocreJr1znLFTGVSZmP46lRx8qEk1eiiP3IUKh4wJqJBhP1aWx5nGVXTtvTJF6FMfWInmm
V3ezk6HlGG5FURhqRdcpUapt3sR4rJUOiUpuT2BobZEx09xRGPrKEh5VizAgMKhLiYYe8ebGpbyZ
bDRZ83HOFUCRJkOHXec4dhOtHIkQvv8BVTDrgUgwFO/L1ltNbyB1UJDGq1B30HNTGktIDeanVdWA
K60c7C0i7vQocwOkTi3ZGl3OsPIgp1rTU3BA6JZD0sMLF3yaCQD5Kxf95g8RkEtGXFROS7wTtAeH
G0b8K2X2RpgK4gAnA41itwTRoV4oGsW6LgWhmphU34nw2Q3yyiUe2aEnEG3MPxjaFXNj7fL5NipC
pGhJmRcJvZIzxcvEOescq9rRKFGoBEb4x4YtSv6Y34+ygEdUR//PpeKUNafHnYmvj8PhLtapglA2
MwfMrVTh8i/jCU3iZkhwsSOY30M0nsVUogZ+V5J0eX+wNQR6cT4blQPs3e3/d82in/safhYUhLT/
IjnPdq6M1q0bL6UzBniaREMiVwjo+SDgDguom6u2M7VpMIg0cq7QzzyqdN0P3nsfU5YMV+JFBkO3
QtPUdo1g9SbodExTEv6i3/e16RYboYvF9nFwjvmCMeYRSBpTWh1i+CcpKTXuxIouRhKXj9+ebJqQ
bQtCz2Ra6JxJTX3QVZNCAQmr03n2EiTwgnhB9GndjHMtXCL9hqkFAcbCOhGoRY5xltRJORnYqotO
k0oM8mfbLymejheq4TlYUQmYUjV8ZiKwDmH/kRhzbOeglU+DbByesDA5/AxZFXp8akSHmXxrDIQJ
5TBcgjYQsmzmOU20ZS6Uwwr2bd2xoFEa3B/RY0CpgBXgfyb354/cLwuqTUzJ75aMOSDykJ4Wv/Y8
ALGckw+Ra5sPsLreMghDpc23naJL9AUyD4qQq+qFgbsArvxwziOj+Nl1AIgnfqup66I4dzWsbIML
qWBIApNmVFWeNClMRgN34U9r2MYMStN/kBZ84S3V8IK8YrnXyunRi1eyGKlK1ox98fBS9II2sMVj
gWv34upl4TpajxXtDemUYon23LR3GNtOw3s0WuVbS8yuUmGB2RCKOk0BdzzWMaxokO0+QHylNRjp
1qSsoud9uaitAaAkdIJvV0YfxsooISFvIzmVDj41s8TdOZ1uue5HQl5yplD8vSxT3Sw9m8FdjzXL
229t+yfNi6/dAsXrbLK026jLoW8Nwjr7gX9ZChca/8fhtSLRoPmSUNPTuWOmia8e6wa2exhI6fGw
b7ba7zywL49XLO8BL53VH3j5hBhBZtY8TGiatCQKAq8FZP3BJ1PByTftsZB21m7A6x6z7d1+gADj
Nrh8UoiXizvtbLnMwfUw/qsR8Cz96dUU+5aHr6ioIaaXvNUAq12Vw06uI3u2trNfvCHdMZJslSj3
I2IpEZI+MR7jcQjh3/ie28eFJMDbtgAf6KFJbQ8n5zee+67tZyj53NP0LWhUaYTwQPmuuIW2Ku01
PPNBXrECR9DGAjNdf90NkYDXAIHXpNRtJ6UtPslwPVTx3bOhVQ180t4MyI946OCRe8AF8SBiwtB4
ryD6Vm7NNl0kHMIDUYQjLDRUkXrVf6iag69bz3mqq2kKRW26/0lT3VueUUQza1ywPOUPfda+pWid
dhBUAACKU3XKRmhF2IBBTPw72PooFxxwvyjT0nyAeTmwvzcCGZ6nN7hjR3kgdCPsx+U6YV2pidmP
wGpypj9xZpIto7PavoH29SU2V2ddQPrNl9qseuVzB8Yo3QWj0UTpluLAsk+9Yw06+eGje9ddtyCO
WRLq6cTeFtJ9Y4VaL5wHhfKgi8Gh1frdvfGaq6sRZYXr/NizoogLsD82Wr6s8K/Dcogl++T9NQIj
lq39Fw3t+4E5PGARTEn/Ytlhp42z65qQtO8M4wHXE8isB+DgH/TLcgn1j5lZmSjB1aqyg2daUcfo
OZCGyXpCJIqB2t1A2qGVv0zDjj0qgkYgr6oVHWklgQWgWcb0rftrDGj9PBTCRd0osrSnfoPNBhm0
rvQ+sS7ToDsDmDpQcu4znrWHdfzpjKD0Am2kxBf2+Zu4yvlSHJ4fybni6collHG70yErIW4SlYEw
C3kEVJxi4SFOa3dWnJBI5zRt3zkKl6ASHitwyuJ/ZPQVYYlUTycigtEA/soI/tyIW9y5ylblrZgx
EKOgYP0XvV0jHwbrYhEX2lJ1t0uKFRXe4b8seVlh7CYG0fXYNIifFHLTeBVx6YStgXOAmnQ/Q4Jb
QeMpJ6GqwUwca/Upc2TYdO3Jx8JCItbWlLnvmnptg70k94F898//0++QpQcNm1QqbleoNLXUB+G5
gVIaDJCXHELCFr+vSv+Temj4MYLQ52X1/UtnvDZy9og+DbyyE0wAuW/4ZywK2IATOTnm8tMwyZeo
pAfxNSrq4xaTZi0mbeNaMAl3aGLFBuv7v/NUG+gTFRWC4RayvS6HiLRLKEH3pHEthS1/FI5Ji7zj
QTwlwaePpT88ax9haWO0Ury6XiWpqsA6PRdfgK9WMFbq9Kp+xBYaYqa1paQ9ippREYjBaYjXWlP+
GXjvSA2NfWu41eZm63kVchn9byCWiifb14bgCSLvnxT10Nq8bmApB3Hl4Dc8wRYTo5n+FKbHvoOB
CIrJSuxld7BeDBS42aPvVzNTbW5JJQKq0UiJcI0BsXfxvYVxvufR2F9U2ha11HwfEvUMc1298mc1
Abrmu+mjIRzYfLIN32Pn0QFdU+NsiI8/KR0d3+xUMof+0kpvaL9pmE1/USEUUZravpgbIMUkNaIs
+vb+d2f/cY9PUALGtfbxpSaxV/YNW+9/DWRuXrQ2Ykpi8h8cD9w+AGM+POSBZ2aWUzGJlvTfSf8D
7F9lcoxURsDSEfvR4hccz/SjgMMiP9fcbqU9Iie5/VkJCnD0ZFIOsaIY9L/nhWZLgYycsbAgL6ii
G/JEiSco0Hi8vzGnYqRmotC56hz8XEfd63LXW1KxyAov24xDsOVcyoUZSZrl6sLBsA4gat+f48dN
nfEiEPBZ1NiYomKTo5C9bzE2MvzBYxuYLQ64WNXETP0S4Rguv1uqYVVVDY4CkMrZHXmNs46DzYBv
gFNirBISmexEfRXDMH6J60/U+8JROYuXR0gQ9vdj8d6pwH2qsnqjA9Xe1QxS4/YxjofD+j5cBGCG
pYpFK8gtRfFzReoCVDpGp+vJNq13GLZIqeCwGSOGIINnN47X8rF/5qbIC3LUxoI8rzy4mX9adw56
K1oSZmEmk3MS1lUPRzjEBjQOWiP/Ke/Cic3V/yRYEMx33SzzBBNfm41R0ZP10ig6Kpri8PNvBqIH
MvWTImcngxNBlF+T3rsx2Fnyo5liKc4Ob/rfE+qODt70WSAcOPuuHfdVa92rFFgxrBDhe68nDFcF
zY2ys+MueKFeuAnK78STifSGA3d67Gg7Mvho3c1ivAmHw5s+0xGhCt7WlXUBf/w2c1nj5UIKfuTQ
0Pv6T2bwqYnrwMABQL77PFl1eUdj7UFsaKDiPlNhxwcLdeqqZlMN/eSSeN3HHVssAvBdYk4sSnoE
PeDsBgCWsiI2yk7KLBbO0BQz9vnxQ9duit8gb6UiEzmaqNLN5YMb51M6lmcyrf1vzyPLTdLTz8x3
t1uRxKESeTDKq1PfXCkG+xYrQzMfYp5kYCDt2IAlKeaAEGFcjdk+dNbCD0v9BvWyX4Ie7C0kEkL9
+9iRb0XVtUJxCyVvWkHpqBtDJtGjoBku3Ujw3veZ87EBzqHwnGU7m0/vvFlrdrcYg64JLUVdq0VY
VB3yMjokedH+yttWnAVsR7Pbn5Rp0zByXRAgxBAk/2BQ883ibb3xa+fFO5TlbDk+BdJZ2hCABUwN
vG0V3BbVq/46p9HRzWaUBA8vLpyFvBLtGgcONk5keM9d02N7gRToRJ8nyiAltnmANd2dwZI9eVOx
tvJnO9i8iebjt8atesuJthC5RmS8cpYxhCDITi9yDU78EcIAonUxOFcqUfdVus7zG3NL4H8LmDTT
2bYf5ZhctJguS7MlX0GsOUJCCGqWWNxiiCswQjagU+LwFXQ5EDN8gJ56b+9MWpsOV4cnmIt6Ui/o
uFBdaZGH+HycprIpgkd+JqLZJhIeW9XgcU268cFp7bY4LlhTB48s2yGZzdMrYD/uGMgjOvoED3rS
N1jUuuJ7eNs4ek/QgqWFCMZAqCEwxQ4Oa0hW2AIHXb8j87vU++NwLomIQ7iZyuyq+RoB+KbftyzP
gPYQcObrPjeTFsmLEwtPAM3mZEB1UQ2R3Jv6KjjxW7jK0rfUWgBatqn3LlvwO/KeWyQXFmAqjxnh
RGEHNLbr03lFcrBpqcCxokuKCJFspjmzIKJDLrfEzNt7Hnaj9NDG5jpj5wsFSgTS9QNu+Ws7WfxD
OKEhX7jB/9ba5Zdat8qEVcfUCX59l7iRgUYu6+g6f8KzSxjPefeTtlIoATPjgJIr4Ylc287Zf2Ml
sa4HLWIt4gHnv1aXyLjMRbGBFiztwBqibl9BBA/k2N1yp6LPBvDgZKP4AGnjgKrf6mm5CF8sSi9Y
7xkcjsJQdyr+4KUriYEa1BpTCzum2kGMXOV+LARLMkyGzt3etugR57xg73LzwJu0vxbk5bSd7cIL
alckc4ykrESFsdVktMLwrLZcS2p8i22V+o3mApYra03VHm0XDdNPxtcSDCQdEhLWYvsZeIE7SvRq
lCyEisn7/rAslCHdiw10gUJ29jDP1cEezTqG10ApWWCt6g3klQA+P7vpl9JKRvm5KjsNcIx+CqYX
C9ccZcXV4G+Nw18XpCgXLJPZWOphajLfqYL6IQUDBS1R+yAYpygiQv4zAk0iEFF1XNmdbdI8O8t5
yLDH+dkXN/CJCTdIeACjOpdWAeI7I9w41x2qPoThkcDU6ldKe8pHObhirv6MHR1/P2MMQDSLdJ7O
OBQFoJ6YGfdO8pIecvW+Anu5iBgjoZSFyDQiqTo1G+51Uju6IhLILYRFd7QBrZZiyWVvoLZu9XbH
O041jH68CkxdtAhhSDH8v4AM2jHc0Ch4hMqkQIs8od4PvnflTScKd30/0z6w2wGl0Iw0+5W6nmW7
SPMxNdZHPTRLb74y7r39I92SSiMFMT4JVIVjbG6w2et2bkRwGjVg84+CABofjhRSBxOI3l3kxuL8
taX6h3uyivOB8AEw2yzLySC9wX+wIZEbtKfsefQ3SCo3HEJmBqvD4dT3bb4vYhXE1KS5yNhYXhnl
BNu+8mH1eYT47QL5ryhG/miWVBOwGLrznPfiWlmDYBBoQN4HDg7krISoHGA7bmlJ4Eq6gpttjXRP
0+YSDQ+HHiwJZ7P33sLpSSiI6uaqf/88vbzynZ6xHkvDpLg302JQ0RZFP9IoKExB6MPj7eUM0ilU
8yQyXKWc/RHWYK/2WmZcr6lAemf9FqHhtn46r2As49K8iGtlmj0JW4HNAy9nukCKSuTLd5oLJY0d
AoB9jvMXYa7OVmAnfVBgTzrI4QUIvWBhsprR0DacCraYB7hyeyq7eKW1kwP9Yp1c9VUP5oSpwF0V
bLk/gaBhuEHMysBdpbm3kV0DB+1+Tk7hcNB6poxddJnU2IPzqGeQnFxVu2yPeLC/TJ43Z4SJ4QtN
fvKwgkbhX9uayZwKrCK2AWmW2vYCIlXD8iaJqM56RL2EtV7YM9ddpzcyDogyUrSc5xfKW4FZLGFv
i63Xm8o2mGnQWNH+1kO1UlV/EGVsQl4SCKVEAcxPoX2iSGat06VswnXnSuZobf2jwBXEsVm0PVzx
1P5lqsO0cHJlESFV2VwcFJ67yQfjDjTmDbft4ccHo+QDg+I8FZIZFzRIG6YZosL/DsWiS6FX/k2A
mTxJ3HD8zsdg0swBipwixRYvM4dS16RlwmBLYFZYfBLPK6arPjN8K/ViAndmQBkMlSxNqoocEIp+
99lKVyGhf4RC4NArav4MxK9oaSigHwBQg5yePmPzDw3RpfNXFJQDDCy03eU9G+2GjihgBOy84Wfm
/eGHw8NW3oc7kRi59Sj3qM1dv2MMz1IUfWRN0btIrfApbNVHVM9H80hrylzyaR6JMtXXbQE4LIPG
4cO0zspax7Bk8d4XmbBiHhcGfiE1i9uI8E1fEl7WLdH+3O6VdHhQTPQIHeBDtyYWCph9ewjZVPOv
LDERo1kM4F4CAzP5d6P2YoZMBDIrYrCsDZt+L72TMnUBJabMTPF7nXIfeWIAO9YWD+SiIbE6kpa7
QrRkEV1ooqhpqYvFdQk5NRL1UoNUAEa5yHjUB1d6eUybLSXURG9wlzNXQ3J30hzw8FW71QQaNXex
PSeMH7p32nF+yNuoK9itOwjJW3Gg0EyqzE6+e9pCtlIuDNzQ3HbYVNYN5j5beIUEGy5+tVe9dkH3
oLA/FvbhUrg05TUL9EU7KTOEtmjIbcvyZCXN2spA5/rLvECnj6oN++hM9786i6Dzm0EaZt0VNrGf
mHKfiQ2GIwOj+XEcwCElcm6Ei+uoJDivcMiTJZzzumTvKROvAwzBuc19ETCS7Zs3CconeEtYA9Dr
ak7LDRaZ//DgcwzOC9fNxFmncg492Qk8TuIqVjnkF7l9RHtJg32fg51jBcrpcKctaYayZZ9SDo8g
Q1rPnwnDu80k08c3OiUei+MPIthdsdLE6I2bugdJfSAvxa546Xeu0HonEa9tpZAieHmD/WVz3D7b
IQ7aJETTEuQBNRFvQzjiXH82Jib9Ew5YhKFFyQJ8EFszwnN0rqittHxNnVwjwCXqrwihdZsq7KKO
2r4opLE8y4DcnBx5T1vUnp+bvDRnQ3BqL2snCE2D9uO7oE72E6bLrkfEIindN+AMK9CtSt/2y0sN
Uk7qfI/sPIktvBkEKfntwfD+jI2q7POP1rl+fL5n8wRxQ2VPhVnNTaP5xLVUn3KcFXJpy1F0noZ/
NVqndh7HLeqBTXnQb9RMEkHnmWlfMNEFd19my16WPtMKzFUAqv7SH9cs0DVYr6MydQuYCPPc5NNa
TPUaozMJikZAmFsOpQf6khwxC7ZmR2YppPc2XnFn8M3hRAhRM6ar3aLw/gcpKdR9Aww9pQuC89oL
9fj4CPN1HO0jLMBN4ACaHpA15rxL4eHHo4slLoFLyRv/+smYu3AZrkvNN1ss1PQYOrIKo7UYm5xk
t3/4XzUHIHQXM/WGPOoHBocz6FQVXsiNP9ai6ga0c6u9u0bYNteyzuBRIBUUFViYWvgxB2Gx4y86
Amt/hI3VfIR+Bpg3M8O4FX2SnPBebybicDh2Ndmw1w/6+O1JYyliFoe4LUTkY+jDKp5Hw8tdH0OP
nOyJbbI++eBXIPXuAf7gT3ScHKZIAm8DN010fmLGbco0SvCfWHVGEvvQo6JL7vAkZnNdJWzRc/TX
Z4kiHq96+bRs2z9k6NI++SZmaAlTF7ONweOnXe0sT2D8Duur2fYdKjbdsJQK6xnNfAC4caNih/4m
/4setbHRiw6ZhEbaylK9J54w6ma5xM3k/GipJHOn7Pw3UmlE/werb7UpAB/Mc1SI5vJXD00ypDAf
kLLaB0UK2XLpX1LzsSvY2Lbu63FqXHmPDgcWi640wBxeKykcv/GQwWzkqyd0oXLTRmTpwCZxSAtr
Hp9GIVfTzRYlFPc63hwbVqVkBsNo3de1IG3kISwieTqxLmN1JcEYlqJB2G7fceZD7sNZb9NuO55J
SaNsISTRGazfyP/l2Fs+Yf7pdgklvQhdIIIRvOVho1vI1LJPBY8KJ1vXgnLz74fy3vk7PxPbWaEd
YtcS26JZqCH4cRFc20dBB5Ls0HUYsaYKNmY/G7if1mKrtQmhdqfxbPAvIjTkcaBevNljDpYZvynv
TzlNaI0DN8Z8nAW0CdCeOoPhw6sqRWLnYrO8CJvZSCD8osb4kQvvuNhNZAGX7IZhcr+TUi4rbLfk
TekelFEjMoiorDcTuaL3J5bHSXiwTKcHZMJvTJsbmviUGA0BZhHL0fxx4bw5zE/N31ggYRf8wbiz
QZGGvzRmjLya+mu4Ygzn6uRQx+ozkA7vC59UJillfjsfGuHsl2AvWYql+2PWc9NiLlNsNYJOpWJ/
8U6VEhgxTTHcfBV6sFKjSKnwV1iMvIQ9J+oF8dQ/QH3sJbtqr3OSxLVw4tgN03gSwMqFUa4UySiU
7jrU3e4cxJ89Ra+ArTD0T2Y+gFoCHG+HGe4L5ySxALcSzmZrYFc+iEbYB3avSCoGaAPUE+5h1Kr/
483n15YTPe/UX1M8GSLTN4+w3pqW+L0HIUwQcrqWdd0ClQ30aAiKFgNiXSPB84hK48f2YAmuaNct
5VGTBgpqRc8ClsDllSR4I7pS3BiLQsdWXlEQOWPpzKX8xkSdVw2Xk3KrjXUE87wR1L9xrQ04JRfY
oHUvy4PeIfBDtIqjhs3QD6u6zKyDJEG3NwGFeBOeHrBNwClENNKwugugDn/Q15RYXnBer4ka9S/C
0w5VJLjvsbZJK39Q2CwaF0bXIhHtrdRkUuF7HkPx1PWwlGyyjKrc3m83f8nIFwhsin/maY+YAtxI
Mz2tMHM+4OhX+3HuGC6tWL06RAkbCdTL77JJxsOe1WtTV5JObjLOzvXelzD2TODuqdq+bCfQfPS1
CQVg3N+U677rAFMijE3Ac/EqYlE0B12j9ficUigqm5GHTzdUfDXcZyfUss2TnVmqB9Cv8E2cYA4i
GeuQHVuqqep7d80nFHITFDa5KXXzuOJ3opVyIgM29NUpsg2Idu0m6YV3ntbktaw/fod/Ck/PTnJo
ILpQ73kcGscPjydbMGCefig7CrP7nxvHDBOMXiQ349+sMOTdcrkfRfjFM+j7IOfBgZKgqs5PQtzW
F0zgzmu2cGvXzA1FwWTg+gvLlZ1Ecj7Ko0TVUvrQEl5RD40VQWX9J/Z3WX9se63pJ5ZrmX6Mj4xL
NsDPcTHry6lb93RDUUXD2vU8yAchnNnXuFbW0WO8BzmZBllbYy2t1LLuFmeCBlJ94KrfCL8TpvvT
0PW4FmIypZ4cvyUj+2X+GGUHAaJm0U9tG+2fXk/lUejQu91naR0PtiKtxN4qpUgRLyRDSNTGIx8J
B29GHhSGa9lzyVnjaaxyxOwCakzgXSQDnqgOMENgj1NNnv4Ylno0juSUZRIQgoYjOSSQ1M2AZAgJ
ANoDw7IosPjK+KFN+h+htF1PByx9n29HZFw2e84WxgiYGUZZx7pjZYtygHUeB9bb47OGoPnccq+J
CcokDFEYwYpc+SG4g5Xw42B2OwmYqKu2Aes3W4iYhLJBifClOH7rR8XKuErmQQ7zmKtlKn9//JRo
wl5+z7mU6VG30scPOFMtDPjEJV27cJSPgS2mOG1jl/GT5D/XDETr3rrXg01SMIUrbKey/+uqAopQ
qceuQ6k5a92KtqgnnyqPW8KyWMwni0uBh2sSbMPbFA1/wMjNib2lPGVwp5Tf9dKj5le93kcAnEWN
POHS+ZiOPYKC8ojQgdAAI7wXt4xoI/KDE3EKET3O7RXP4eBLEYnLMfjBKwX+pTvPASdkol2YbWrh
6VeiAdt1au+W1SDaad56BslMs9LcQ9odKdJuZcD0lQVEeemJjNiJV4BggJg2IVxqUshkYvQAuHRz
RGrUG0FbmQtaQliaLQVuJzoyisgS7ICORpBgHZt/p+SOHDq5+RBNYux789u0LzT/nK4hpPwXPTzY
ZlBTUqlRKjzTeUNHBphZ7rTpIJz4nry0aiR0fH3ui2rdjzVMTcGDaZ9YjXNQtCUfmiQr7RyXfmnh
wEBhNNPxeeY5wFwzOn5tnRfaBUAzDwrJ9ETBZ4vUdou1Dtd5y0/gCfUASDja8rholp/9ub1mT5aT
b5d6ct61lCTyP+BspPem+4dwkN+Lw+7DbHjcdLRq4OtZAbkzcS2svojG/v0kJFN4nCmezwbVzc6I
3A/mWF68D5JK1tHcM3DWEvx7eOEDWX/lcfGBB7PTML26+n2IFPfvwnZXNEnmnQSWJHN3OUclxTk1
4a2Jcm905Bp6dUzMv+Q2GGk/lzOrhVyTf+ql5mSEJ2IvEqiKMyrYdP60pIrQfuOJyMzwH3I0CyPe
E7VC7dYmw2aAYbg+WbL/AWEBvR361s0lsBt+ntJEprx9jKfsaNX6F4f4KA1/QB593yMZaydEnZEi
d7q51dwVjErsiVzWHJ9QhPqzRwi1UncGfuPp0quiekqSF5Qnao7sTMIaHMrUU/zU92scvN+0UK0g
X0u47jvxdo3LmSxYCkW9/KbrltBqpnBa5mMhS/oum0imZEa32CE6VPreQt461EfoYDwC52ZbkKgn
JmxN0/EPrZHiz2kl9+2CjZZ0l7tF7LucVHi3mu/g2ZGWUu9kREoAbUF9JhWneQI+/91G4N2ABktJ
4M+fLgQzTjQl+DJmAIcL5fKqkdvF24re2hkoGQkTbxJQOZ2ymezI9JncWCk0ZW47RNLbNLYB4CGJ
VEBx+erAtMZxhEOzMDK1KlRUkFcaFHilHqDbppUYtjKORAWDjm66lwgzkMxFcQWmtDU/R1xTAeMK
qIXUQnrFXDvkmhtQZkgEaK7n+a5hp1p2Ap/c01qC6LyMIjKPjojx6zXQoWhHQxowftlNBBJEYOuF
SSVMZ0OMl49ID0q3bdwpr3NnPT/pB8E2E96Mz1taah0yjv52QEv4otI8o+JIG1rXbveYLDJ/Y/6j
7MYjiiRTeIwQPFba6QPNdaV4fAlcj1FZV+Y95rsO5KUDoosI4z/pXXwH9ZlpkxQ/iy2FSqdpnJuc
jwv1Oov6PiSJr7lymfxpjNtqTCrFi7r98TYsVpLsTytBA0JnP0jh0MBRIGV/SKlhOWGwUHHcxT30
ZpRnEkZBro1zSOwtUAklzpqwSaZ2FANsbWiIXPaVLVfoGXdkCW49vNTlzPhjRgCO2Oxyc2eYP7xf
5NLLcRUyTZmicZmK9Xu/s2pXLlEC7LZ2Qz1as7bYsjKXB3PHwJp38WHi+Y6BRJ+E8vvUGmk7VK5D
foFDGGoxeGfZBT1Z6JG9GCAgjkvTBWk/UMQlvKi4bkPNiypztVo+PnmY+1lESy7H1rG86Wy4wU2r
wLNwEhfBE3a74L1mHf177meKQA2fZkwdBv+T+x76gguLBLkm5M8ujWTSVQEymy3Qgol3yNpYAhUc
bFu+o+6xJlsHNoR9bmld6VvWXmIrQB5ka5mWEL4gxEr77uO81opukB0jbR/U2X7oc3qM4YbXqWD4
PkdSRBKLTIddRBMEeiNIj/i88z2zyfDZ8xt64ocR5o557YTIfCPTYK5KgTthc5HmXWOLGng4g7sy
oQTt+XoWnoSDM+A6o1VRca13MEZOteUYqsDc0WE/APRfnhb5CDULlEw0EqbUYEiXyj00D66zJxGR
YSKFpE+2Z4t9zUQScmYOHYTkOiMnOFt2rTsRnA2lv4+/ZcAeSaPzqBQ7fFcrlz6M1vHm/TUZe40f
r7u/segk4cbtBpDTj14n7GSFx/jZh7RIazbpbd5CK5Y/wzibzRZlgNb1TaHZld/o95J0AXZIROjB
fYE8/NiOC6yGDKif45dANh21UTUovnXvpNfy0yvBW3OAx6Rg+n6WBdMxcsnPznsKXD3AH1U4CeUZ
U1rgGE3LJjkyPsKT4vqSla8M7saf8NZZEs9w3uZy/Cj/nHjLf0BWLNYNXdJwqs4Ltb+3Dgsq6E1M
iKWBLn0hx0tQ58zeTbC1KgyYGLoWkuyYNeEf28Y+Mq3WJsF7n9p/NjjBMInkF0fKzN7rz3/8z4p/
QBQUh4Zz4ZDenINSDBB394qdzO3CcAAQWFohDyl2lpUED0Lh393r8ySPJEOYtLY3ulEdldswOvdy
dnUfYQ1w0LQnujy1DecoKqo6V6ZONtUfdFOBkJ1dJ8Szt0tojSKD60RdxL59gc3ISyETtmJ6JaaJ
T+MMOwPER2mzpffEP+RE8NDOmIQcz1mNctJApqASb8fWlb44prMk5IVdzchAgpXO8WsJxbX1TatR
fRGpnMuweHreEvpmUdaPiovTWfwwoE/3JiDhbYESV6vwKuxdwKiGGOUyUBEFf441lzf2SNoR5vuW
B+/fT6BKrC7TDAGgNdTNvaowsiRPMF3S0KDSU2f/44FXzfJuXpXjMAblvTNzEizhXlFWvXolUY5F
EH9Q88qBwjaPc3dxcTrqN/MWcns8WaHqwsAPQ1eZzgmeyZfQIi2go+A3/yC18O/ugi3IVp6QNRIj
7b/TQKZyuNtva4HaRHr6Q22nIz3ascVsht1UYDyUSAmQFZaFMwdstbqmh3U7131cKd1g9XGarURi
zLwUeghouUeRk4M4voST88LSsTiCU24s/iRrjpjNUxr+WzQNlbc/bJvy7KydTxdmqlgULnklDFFy
IPVPcKeMSkAb4D0yaWlOqYH46xXj12pWZbid8igoKc4p+SVhdugVHmt5yxu4PAb26pPx65m4YT3j
sThsk+9Vtwztn1SKV8IET5/o1j5l94QcmiDU9Z5SjLBA/L/e6j3bPYZJLdoxEfkrElqrp+0hMxkt
toz7pFLPRAFeuhqFW7OLjgmPXkqYGGfwfsg+M/f0+xM1MRFUXdCAOhZSyaPR/Ic92Nok0aHyQdfM
s6llUYCLQ122yoetHqPLBgSXnk9EheLK5xy4enCqfIu5AdoaYAuqQ6kB50RMpq0GfZ3Ee99dZeLt
7eFvptdP5tTtqrQ7PWlzGPaA2eFvckNQQK21jF9YhHAyEDXjkUHH2vcvBdaJItfxRagzjPF8dVyU
HRoNnwm/+Gfq+PcyYWw4Gw7LDNVo8AEwre2muvwTmUH7AcJ/eUAICtXdsBmmZOeYiD4ttDO0uL5c
Y3fyR3QiBxFObkIF/cJMEpztfmECi16dHbLA+CPPGkMMLttyAAlguqPc2loI+CWC3ttFpolV5tws
6xXVcCDnxnwI7P7rZCXPJQNNEaCx3LSbfs5YIok1HmY9jomfKp9davjniDlXbQN4cu6p6boxY1oK
K9u+vJJP9qphVaVBmt5U14NWbSmfreaWsy0Zjs7YIRWILEgFTZ/V7GtCgid2Zh1FRW81PywOypei
M1XO9ASjbHOWBTq9cD6f8OGRXTMj2WD8LOXbrHwagZqlL+8pinHT/PjdH82L0jeGT6ds3hzcCcuA
D3H/ORjoitBvLsEXcLVv0gn3UihMSHOJWgJtomKg3ifKtCKv6iaJc0Q0L7dgq0WBN20hcfv3DHW3
KJG+EITzARFIa6XAoH63+yPaJkchdZcJ4DSLDz5JxjXlt8s+sZNg33iuX4+qc0rQ+4w27GS2DPgC
18AV9t6EW6Bmcd8cn4bvwhOq+nHFmgXWHlGsuVWKHDh1rnN89dgEYe/4rMZSNS2L3VieLOhXPhsH
bQ5AiEIPw3pz313++tKDIhhGDmYJWpxRruY7Q2I/qvj2BEyPcAqIw/57QtGqhkmZjcGXwVuhbocK
bZntqhN7+8sFi8+ZBYzR56t64NAZGOvtmfkg7D9PYEU+a34osYdjCDyA9uUMHIEs2Z21OHzyH+X6
Pgwkhbes9cbhupR8axvi+oLEWaYPITa6rJYPXqfOmJ2UlR7+BkKCwVQVr6sBByp+m5jq3+vfeStM
YpWe4ogXH8/e/xsNxSI2U4ykHvdygCCTsTnh+LfSp5141eLPakm9yxAGIHIrD6Kc7RJcuRCkGqTV
cYkMoEG+d+hKVUFljIybxCRw+j/SkSc40MrkhNHD4tyQANTHABq1hoCKLk/zdFU8Y4nVx2P0tA9i
ucUYa8XQtMFctxYkclc/lee8lVyTbz3k/zK31ilGn6ePPIANHgXBCMksOduMM0yR37IdnocRUFoQ
O0VIzkK7LKJaweT61lmpZZoXaNHWh7e44Rdd7dKP+AgSvE42cUvA5lFiF+ZRw7/I4nNH3nZYfDlt
4EhhARmd1crvLgRc8yosW4Dj5WwzrURPeJ45JyQEHSZ8UON0RYe0oqRqKeSAZGvfd7bx9UGqMlHD
jFIQ6lgS7mJQcTSQ5BFsN2UFDc9GRmVcPfQr86AzrRFc2Jv3yH/T+snYmKtt/xHvnkHkyAZ/hkcB
ZOMcZtL6Gb/YPB7CMyxHN+IyvXhcWo5ajzO4h8okg59VmU/62kLoMBY/QRzvRJbtd0goz/RPZ1fe
2neam2KpqbJfouefawcoMs0Q+K3OHXTf9OIZnA/n3vvzXETADAdODWz0kiVqbmqXY3R1fgzwVaJ/
107e83RTeDLMPsh/uY6CV7rzjlJPm6MypX+N2016ZWOQtsFE7z1ezyTZf7h9Gp/GVhrfyE9b02eb
rRS0eVKcOxBhqPTV0HBBU/g5bplnuBgiFvlKx2N6eIcFos+/D5gZtHSM1HeMaQEeLUJVjtJQfs+x
8b5C7QHfL0xEOuxuP6JRwd4dQv/58IZw/DoLqsAb77gjNSxL5q2PQzN2W5i06HSEg79erdReLJY2
VzQ1/3jsoK18a5JtXqqtcvnDuXEfx6s+d8vdOh8TgRUhzA7+IIEsqxYVKLe5e+YgUJnMjSh/1waz
kEtbnvsBvNe1jJy55ZL6gu7GI61hpHX/2CyzHMj9vBd06lyqWK9EEPbS12EvtWbI1s6MlVocQdwx
q9J9GE5ju9eBXXxXZ+mWyXmh8iZBWKnzmnOH7Ev5WiqLmYGhIlOXnO8KQyTDRYLKenSVicMXu5G1
O8vEu1iO6zSSBXXaffZYup9Nfhs5UhNo9sJUpQtNYr4cSr3Jg58B17hCB3LLavUBRNbKBmig8qOn
5RET6nYbBxkYNDEbAp/O82sfpTshyWXbY6oMsWZi3IfNieLhTo85wzWGSm1oofuy0BNjNRmN1233
WpJeA4uSjHthBtzrFs1iafwcBwYWaK+VIgDalg+2i+T7aJ891P+zgPFGgCXHRMmrXwV48BNworTD
+rPf/vmshhR6ggHBnC/HzZn93ORKS97R/pzwgnWE2TmXisoSvJY7hDUFddJtyOfrV1+HvfwvPdZi
cQcNaawFP4WPWNcm8ixrlh0BNlHwrrbnYvvUjcmBdxzO5CzUBrV2mwrNjrsqKITy1/3+tQNo7nrK
tC05yWRIrzMTcbxMALA0yIzK62oS/kprpTZEXuQRrmNYRqyY0aK9rtFMtugRLc3SexA1uDPJ8V61
Gj67S4d2tdJMeyeHuTjxXGfN8UZnwoyg78fdffebWzkt5Jr4BnWekRCzci0X+wbzUa8/pWdXSnda
AtgCpqfMy/jJpkw1q3w9iS0KkOm8PJu1QwO75M3wz5Odk6vX0+aCLw+8Xh/OPps08LkCdvuheMUA
sDuAgMFVNfNtvnwgV6asoVfPhuE2FRpNtvWsVtfzSH0VbEirRPLnE1t9YZyv1LvC8HkDP5CVplqY
AItjK9xGnwISc8v+L15Vx9+v0GySPCHJbOgWXI7I4R0SPOmS3FMQILBFsGoAHGH9TXn2t9vFbxWG
c5cEAiIyP3Q83iO74ypm3WICG6DJokEd1ZtLWUgDA8BlzIA6IW1fn3zhwWI+tRhQeNrCuSvA02Nz
zn7aHvM82flJn4Asj/U1raLIdeTi62EeUJdaxkT8Izag47jl6WqFzn3+Fve4XWM5rElZVPjgCZQA
gBFXNWKhVvnQl+aRR+z5TBxzoOiDSPhL9EEwCGS1EOAEtNBBKdYIw/eHiI++xgIpQOJ8NVycL5fG
ijKWAmyOnrxd1wiKzSjj6A9OBPr6LBqJF6WziuA2fji8ohMjshOhCqQVDqognvqXVtrRGGiO+HHF
mNMGeWQaZCXO32+hNlvNKrN10YQqpkSxVbFtcMQLAW1M4lYAbqbHpBPdHWxHf+IPf7cfTWlRGJ0K
4tlK0Mp2LQAWKqA11WAV3AMx0X3bKVXhEZfjg7yD3+HQM+cceNvvPh/KIja9+nfDUKxqFTRc7UId
76v9VxsV+G1uyH3Z7Bbo/RrXg0J8xAoexRZueu20xam8gLAb5r3qIkduJqQscKmT7k7AMsAz6Y5d
jke0slSKhcWwnkp8PYvj0gAgfOwPH0Jj0IphRQ3WLEXz+4CQhLQoaD3gZoV+IzZvKt6aT0LX3irC
jQsT/N6JNdvgXfaxjK9vkNxoQk8td5HnruBuPh58q3havqkUGofGinZZEspFYtSfxTnOhUV7tzcT
WcOXtHQPjtxh/C/d2fvu/dKWBdpIsMfg3zqXytFGQkl9zVqM38VTB3eaFAjqVddbHmaRIB+H/Zwq
PrgoRqvNhhn+nfJ+pRQmKPfneW9fUy/0snhR2gJ+b8IFKHahSZtjwTGESe+C79BlKVwRTgG+jpCf
aFaKbQxglz5hRUEL9vmssjWApbd4guZ/3MCgJNPEgcLSF6DDBO2uNa/HoO8lGVQDX2VoMjw7ADPH
hvgFW65tq9XW1QfR+grA9Vkf9eI+3UaKofytng/Ws1jeE3lcTM2O1894FpWzWccMJ8KrxZjBgt0O
UNT11+LcPYQKX8J/N/v0Q0fnjpQlQ8qMX1qHoV/icPHaecuX1hQgosHC3nq52evRs3xSMSVFGgmj
F3LNMD7ZIW2KD51a7nG+4VyIPLT4Ue+Zl4OZKaJW4cocdaN9Rt4CwXMHVTd+/+Pu1k4Li9EG6j+X
rrQv1wh78msCIaMQqvtfOZUa4c9oQ7SSndSilJBTO+du69iLeqC0WaAddkvMXOjiS8a343uf+cFl
BghWGpnAe9KO9W4gX/Kc9xG7SB4jcmbsLXfry5VsGHUs8y8dCZKFpa8WBn57/9nwgf0/hvPwa+I0
SzY+e/9wEClA11WGkIqfX8xY1nOA8gR3VbW2JEJ8kvj5nqFLIz7gTOfpdonVLn9Qixc4tIenhsAN
hKIXnlJYuOwRynNqfdmRhYjAJQCl+niW4mS49WpO9Zs+/87lm4jWC4wPorn6G9LxZsFST1c2JJ+P
JHi3FPmCSdp5gizupEW92LXy7toPMj+ZPrwiiMuzl+FpZi7OpEVxuvb35qo2qmCUT6CCpqRAdmRQ
B3h/AJI4NeXzlaqXWKESoQ70BaXjoruiUvqGKxiFIjMVmkVEOme4RjINCOmQJsoVr3dI/18jlS9R
Q+4hJ6tFWp/1LgbS2H+TGE5sp80z3ZVooShEmrz7ZZvrjEUSVFFRgd0phFA4Lo0WFIEUp/JOFweI
vClOnde4iAUUfLF38ZMA4QQxJsDs9oP8HY7aoxKsynRcIzmK8SRbNqPQnUvWrHnGgaj+V84ViEAm
jGJ5zYcvODIm7vuFirTSJlJsM+MA6mFzEcNNscqcqy6yM63mLbux+xETB/7rNYq+mJPV0/xoBjbl
mos6abYSOnZ57RE17AlppTg4EQCwg5zJMQ1S6eA/qDVd4LbvDZCJByEf4qsDhMnUBFo2r23Y/L+F
77+REJzATzUxhlFPZt8n2G/RriDQ9E3bB0qrrfGrwxqul0eZItHT2b/LeC7fqmeyeL7ktbfXB7rV
YMWHSNa8lbjP+As4Gcas4qXorF8qI8ddswHWfspR/l9jLPe0wQK0S9n/9J6z1v1SmRe4I/cm7urP
4zdvemvaG2Z4PJlwBMs3tyya1TICOM0+6yODo5YZ9obIrJ0FU9t632qVNxMV0B1m6TEZyknAedAG
HaQoDyjweYVgMcPa7iPAHWl3QY9qJo0HStAPD3gAlsvWFToOX2QgYntCOadXQlg04zmcQkyH4DHa
PehJANjsiK30eefFyRmJJUfpfVTPDwgitc0S6NHkjeWn0qgrx/YxkBT8Vg0ldjXSeN0SfjfL0/Wg
n23AbWtLthz0dxqwCJhceNYFGDknFbliTAhoiRIsTtP0hB+0I60utUOp81JihReUH8bNmZELejFc
1M/J2Z/6uFgo8P0k/kRUKvjcpVB3E2fqA3owa4bwk6R1dC5p9TvqazLBGRom1YZdYD/HpMXbrWAk
fL3qySzn6uNfregvn7Qx4smcWoP8DSVMw6zHiXfCUs/qloQ5gr8uB9UX7cLAFDoX+cUca6xoX4CT
4DwPUfa/nqGXG9FBrPe/WUHEBWlhcddHEDARtfKAvQzbKpKsuPx/nGmqtPsj7IQSEN3nEfeiS09w
qx1O/ELIoszO/d8Z0ASLBAa5PRELhASj9kzeS4jH8HHvzVTbxovoe2411u5Cj5/1NuhiLZVdPQ6S
PJed7TJ4rMpBW6XUV2l+st8NHUli7JhDFQAiTSkyk9WNY98Pw3m+PJDsC1TtqXTth+vwrDRDF6EZ
Ee81QFuKM8IMop7QUB8/W/L16cQHuNTbzQTCJjyyKzzWger7lyo+fkt/1wCH0qYyncBaQSCz5qr4
Q31cVE19PmJHABqwz3LryzTJCMXKTFpaLlcRnihtP86lG7TZ0tgeEWg126teSLhzk0CmxvsbpjTS
XR7LLGW2hi4BdccRmK5QOTumG8YBfUKbGwWTcb9wedXP0NEysHqYoHxDiSe7FSMJT/JblG5Cckvd
lkGBa4HvodOEYirs057LPoqmhpAaTNhWx1xcKZVs2Xj/4Qpb8E/6YQKSv61AZgeTQqwge1xHf8lp
ayDm5I99KYCDGV/cMRIgeU9nmsQtgfDUL3B6xSD9LxFGLPZl2zYzbliGcQ89/xACRJwnuVm4yKeE
xRtDSEzOfNkShAmKsiYdWxXIgjgXfHYtpp/SYZjCiNiNV4o2oTBHg8jf9fr961f1A56dcm8FrIpb
PQTcaHSpUC2SCswJa5grloD/H1albn+iV4shksM2QdOl1yqfF9DmZBQpn9upyb7XmDM7d2HgN3aj
ItLJpqzOQieCasWttGSSwjorab7jP93SQ3AVh1m63IGEkMBGWupXHYfGXDQB2pjkjRlzfaURe6Y+
Rvp0cQ1Un7oCVNDWYgTtQ6wN8kRWOl86Sf9zjiuqq/E/6KgSOV2mp2YpQYBH1XYNxCmLXoLeML4O
hu9phk5c0KiURpwlPFMugu0jqzNywfaVF5s0nNJCS8OAZ+Zww2PcvOH4xNMJlAtd0xAjqAyNk9YV
3iIpFD9NOGFhMEGB+3J1BSHuyzAZtZ131IekjY12lucoqKoctB4x+rClIOXocWPZ50/++D5VIBy/
2oGgmerCtekPLokl6Ak5McLsdZANO62FyDRfEHVpTXCrLct2z38XYRlC8XJqXqYTjLewyDtSRCDE
YNYr8iD6+BLBtGaCrsDGF7js5LkXbb7eP9mTA7NS98Zw1nBVIYySOG1HNA0q5z/Z3IXrE1sM0iAU
NiRvDgw4dhPRlBuzTEYCAhQaficXxIlUEQuuokxcLnN9Nn2BWeyy5c1L2VIS9AGGY/RX22t0Qx2a
X2ovlEb0hikTVeoGYLhkOdMdG9be57Xg1zuCxh+bL7mT4kG+3S0p5FZH3Aut/XJkETtEzML11bK1
lhVX/Y1oZ3lnD79E74aVLZzBiMK3FB1BwsTB8pBiMC4wg8su67jwaZwEN5HGSNx0aqZPcPm9XP4W
CygF/Dcsw0jCqp9XFUK4dtBmFAyJQO/FZdsp3LN5Z2RZqA4cmSwA1PDvIl8uc5Au+LDlvPboFZ+w
iyIivjb0PIMeXtWsttvDCzFa9+Kna6dmu5dYzDrFm185soc9sE+Un+4mGuFQUaF7KEbhIcNQ96ab
NgDqLPUVgFJ4wNUQ1IiUM5ktAzYd2PKetjWYD82plFqhSuLqvV7Gocz91CavmLNcUXDln4itYqAM
32VJc++keIBoEZMm1AuzvagTjmpyjaI5HZtLdiLYjkQo0TW3JZRmimWgFTa5JnMZ/Yhg1/Ex3zWQ
12FDTFDFrUi7UFUVi7SanhmB+HosRaF3w7K1pg82wRNSf4n4GgA/xfl1il3+z/ik6nX8jJuSLXrf
d/dK7Y/78mQ+AVdQZYjDVNciRFSJgpAfQOLE1Rvc4XN6tg9TXZv8dJR70Kp1/KgwLRJ+EX0u0S93
nUlwMBIvwqoMcAl1blKAGPSYevIXM0tn7ODcQ0rUZQunry3HNj1ELQXdrj0CDVG52UbrCiEndvC0
JjbcHCdki4dxULsi+W1W9IhNVzHOQ6J1GGLUxwC4ArMUULfs/UTA/7/T4opvg7zPuCU2ALZWgFn7
j2b5ABLDc7HbZAY7+++vaKjQK9x/uMKZcPKIuX6WbgKsUeMA6VVbG45nQh74Nkp2upBbIVNBO2pg
1wz8zOtcbHNlpOkkrF66ZdCVWvnQKLCW7mUBBQ8Hu/HaheJDxtsoKBKO6aEf1Sc2bxVkXK9NOter
JvCZ4rJSSO50/FPtLNHX3Ro+Sx71So/iKg6v/2i9Ut7L82F+5SEuBVpSPK/Ln2HiLxn79LexdOmB
TcG8dMAm6vaFpEMIw/wuajLURlITiVUdZ2bpk7RSetJ4F7NFf/XY636YilIawzLSuTbfVSZZyMxl
4GESurqfsD59iEk20+z5WI5IqpaMYY0wOLdb86c7j270dVILWfBtNv0mnFhOqH9DJY26a0exA5P3
4CdMrPSZsFVALWZ0aH3NbNREMItvgjdmY6HlSuwYrtBR1n7FbFYF9/ro/cEZ+iF4e1wc+iz3VwQ+
2U0CUkb67WQnICprJ8sNI10U6mEs/5f9umMtSJv8S62CDQKE8lhTPwAQsgKLEEnBzZMbRWv9uhQw
BGQ0ftbtXB18v1yWnsfTTDcgmgo8GExeCMcCqwYwFLXymkhuSq4kixMTAlbg5W6LGAtNY7JtQyiC
Xud3cYbBUSuDZAf7KzStm2r7sP1RwjamNn7U2q8YkvxINimArstyE8D+09UqZcRVzmBADodKd2c4
4/4EZvlCycSLG2KMVcMQgnHb7c9WRFXubtavrOzxe9xzafSL/nluMiNm2CtL4zKzQE44bZaob1fm
DM3Alcop8W8EgMAQSrIXbdVdD48xgKe7S/ko9sl2SLjiIBJOZMSOBdrz2qSVE6ZDqV7/KZ4Y6Muz
4O1fdD95K2yl3baETb3JtTJmegy5/4haEcYK7ISW1efAIKio9cixKtAeyNdjXN6JtocIVn6FP6D9
yi5vcWuP+8K94KdWRhHM3ie01JOusgQF8LqQALDrxvqDr6GReSvg1x0jvJC6ZPkGvBZVQukcd0N1
cOpY89dVzeByoSZQe+wf/ANnI95UOKf67rbg4/o1YlHr4tAU2HmeUXQqmKjA9Qo1k2OJH6bRo7c0
zYAz0FFYuI9thcjhxQ3Nx1krjjuNdool40lOewQHmQFWanqw7T/zcmQqJ60WRI5B4m2ftybexSTl
8utagOzbH+Pq87J6Z+4SUWbzEt9ak0er1xMSCV0uiyWMrqpegPA5oJIzTlq/+a/TybQBfa/pjdb8
epkz5bU+iNLoe+4tZFdnHfT0Qtf6sQRAZgfyRKdCuMmjUuiFRuAzPYZCs4KBS1JfihRIDgq19wYQ
Jc4AThdvnc0xtTphcfgPpZFBe14Lf2tGYSftm61+HdzgVddhwV8wiTFLecsDBnWPerdMH1iB47VH
qKQN4Ln06M7+qOYkiLlxKB4/6hhdrtqGfwPjVXfWMRSc3jvgY6TkP/jt2gMfuA2v/5efAfMyBl2h
eC4uI43Vi89H67brYsJxd+Bgq0iXBj+NoAl0xHsofnoT1XxnBXBFF9aMGMf7pR5PuX+dBXsQFayQ
xkI1u+udlgyD8KIITrnHAj7HJKaZXpWy4x8+l0Bo/CVqiNrFZrJDeav5Wp8m5JuCFiHFcg+9/uZa
qvPsESAmzP8iJpvHAy1xiLhYj9QFGga24R1nzSMgidw7l8ZyoMOaTZEdQl+BP3xS9ZTt2SMjQ6dC
9/LueqOTNZhTBMnhc5pg0U5TqKYX4uXJ6sKEOHv7fXECIDLSDfRBupX+y4Wu3lB7rL9CyghnUB+Q
pNErmo6Lcr+CriGfEyxs6sDwDIw3cRZVFy5mlUh8Jsn/yB7IH8GkT9qEDZ9gvUyPmtHmmMh+ebKx
xC6X4FkLql7xtze9MxxDhc8IG/mJMQHzUh45mUul/YKfUbmKWqSmnZQysN9i1MmGvDZr+CURW4oy
L/QJJ+cFTf6rDw3HR5sYDDpUdYUrez/9t9rZ2VqBwk7UaS5NMpVprZh/qAueEKT7YaDeQLGGB14I
2TsFFZh+2k3jN8+hjQca6BFmcqe98g3nJ5DF93CkiArRXcTNRZTqXN0YSqJYvlOvxkG+9exjAZDz
dqguQTPo6zoM4/c41cmYtXW2rmP/CAALW/7MWHdEKw+ktiBrr2DbupvD/CdNGWut4+Ttkwy21PZw
8xEOZ54kJ+fOj6KsgValcBjGM2JEj+gAFQXrrxAus6iyF+6qdesFRomjZs6l9DIcTkpQEr2BJrOH
+2x1J5gioHMAWBc+vqGj7ZkCfFG46flOh5dE7Cjwmt+wGK8bIgfy/vbi+3HwdfIPbYEvpBmyNVM1
+tAzGZZev18E60R/4CzFOq+2zAdowrJEgf8yrLPdi5PRmzUXmUoFpqCsTZNlHAuqEYLh7poelnr7
xrYc/Z+sx6XvQa0N7qufxH/1slyfib8QQ55MRpN4dbz8qxd5/NG6C1Su46qqn9UpQSEQrJH0cRES
EezOVTnSDUEGsBFHu171BjXxzsg05Mpam3MpHn2BX40lSkLtqC6N9ZgKq9aYEgSFKiPXWJhoUrX/
gkH0kI4dSRCabv7EjDHdGpLjCQ3P13jblsq8mp+47IyLfSC7cK1Mm2y6/eK3NzRaDq7YYFQJHXzZ
wiUWjD5pkhYzPLprZAMcsA61O1Pm5vtyttN9RpHrnxzPdGqqJbzYV/HL7Mc6XUnIXOTBHrbx7Rer
m5bx5POwbjKmdeq2GlbM/DgxUALjw5eMcpjR7YiBalS8QFd3veyeMb0PfOtzNakFNX2EvS8ImUr+
ulsTQcTa/FZkZSJS4tU8x76tOqqGiRjcN2IpgIXShazlQ1VeBb7v080WUnfIzfy/Hara9GDDi/DD
F4J12xHQ2rEDAdv8MXuCJ99eG2LGcUMxl0sTm8RyYXboic9QRRnGT5gjc3cAG3ikJj6AtDuMF5AT
jHqFrm8hs2sWVAo3hDKhScma8PDNs7S+pmdHe0iY5KPYRagb5E8YyGYuvLsL9Ebe7LPnNydu1GLk
GBrG4dqrzZLXEaL7j1+ywhKhYEL5kDOVGj+xDEqVgmaEPNxNEk1xuLZJL6I16DBbInS//Zv4riiJ
fA2pnpQ4yOg6tzTU8X39dszZ2PbNX1J0BMuvBEGra0kU/YxQ9kEmB/tzBUeBVYMy8lO3Pb2SSYaG
gmyK0Gpn7VDUjQjbsU6UQC8mOocGCiGE4vLCgKlcWIUKaMhyJbnQUQvBNNhBYxP7GXu0L/0jNO/l
esYyhAgouMuWMRXLhqfyyY7kz/HYohQCITj4a1ZaYJ72nf9ZFrdNyTmR4HNts2PBxorDE5fSo9Oz
wPBg+o2hiEq3tnrmZ3ummhkpU14N6Nz67/sHs3X7eQcItE8mGAn9SDBfHY78cHIjK/Emc7UoHCwY
BJro/nKtrXPP2Uc2IE14NfaDYWG1aLemWRjWSCqIL/VInQ7OSrSodqWxcdrHyfqJx/HxavDCL6Dm
inZvzmsve9ejDGnPcqvFjWC0r8JzilGDf9ctQEdNOFwWQpwZ7+6vZQ3PtD78k0Pa9KSZr1GxzQl2
YxmFSg6g1GiNJlCltdeSHejtSX25ELXYbG0k3UKC29HeWu0nyWExqQYKpwZu//b0Nihq0Lyok0p+
IQHPXlnFg+4x++MSFwxiqai8mxzUH7HFdNKHN4gs9/poJtIGSayou5e7wXm+sQGSOXXnWPcM9Uf0
EWW1S5si63aFEeg+HPSbLmXt9v43/GTI09zdJDY6oup/4qySVdisbYtzBFY1UIwuSlpdfItZLKQc
BV7RVECuDczAKpsSnoX5KzwvTFCijcBhq46fb+XgCGOUhbrAH3Bd0038FvRTgIzAJtYzyPxhkyj+
YCOVQQyUQWyH0TxzffOSG6oI3PwZ2iC6rjq5yXGWKUUIHJpbvbYTg7iapRQvubOGWFy0M9KAFKz7
7pnb96+qGbxvQ1WcLj0IK+Y1uJQ6sfLQ1iNgyLqtfQs05l9/mnA7u5F7GAOG/9TlN03xCPR400Yp
oM8sBflM56biTK8GlypZDMwfbiRiRaVIGqTi1KNITs5dSIZxtLWDRMx8qIRwoWvKgo5aVGiYiHDA
YG5dPZcRE/sv/T1D9nzTYUtHHjmCk0CLAXyXkRnXe+udLwxkJU80pY9hPn+45786J7tATBU67kTr
qhxhlzswAoQGL4wxe/n/NgKQu8NKTTvpwSHbvwmG2umDoSKdMo9Iy1B1h9Vw4Nm54XzsE9Oj2qzX
CwAw3K9juVnpEDC7fETQYU4B67h1TaNpyziOejKi6HZMC/x3YS/3rrqJS76J4jvWejd5sKPAOpTp
E7wYNMKH04o7lbEkOr2RFmfEJ36FhUs5v41XmyfHea5tAHgBJLxucXBlHLT2tTQVhJYVVsDmmsc6
e4kVLRantcAAMhSa+6yv5d4w1toygdlNuwhOkPQDnRzbBcax19ia4Q2A8Glzoiyf3TRBa4RC/0TW
chs8qUNqdyrptD5eTkgLavm175Ly9kASD3qtL6jhLP56igcLKLWfHiNHPUGej3eXvnsXOWksjKHQ
pM67RNzlTsO04azh+KCwJVMMfJzzjMrQAAadRmLMKpVgAGO4+eDOvu/O6fz49NmwVHObbLdm2quf
wRilX0K+5OMTKTYVXLOzPx51q5Yfvs8ggma225FqnzODZIi3s79K/Age9xQgDeYJpH7ojAgy3EQe
L7bTkJzBa09W98HRi7TOu80T6rlBNOLwYtWwbvwwrmyG4fla8+TBcGyr81+A7ESIBPuL917WmIow
0piISSnnSl3r/O0/z6aSocl+/b+3Jg1YVWn29Tin5xWnaxiVsBipB3LIn+CLk4be72FUVkMfX2ot
8ZuUoeYdvkaAgcoB7va6GBxtN2WWImWsra4WET978HHFuqhQkxNcfTIak15hNjsYmOnG6Lyacp1S
jD3JRhFS/IBeB0XeI5rP3oLtwoG0h67i2ayMiZU09k4dWvPT/B6sx2Ixo+83+7B3ROgOAkpkxV4I
MgzpU45WpGQk7WgU/dVmJJYATd4ZA2o1hsK8vxpzo3YygXxMqZOMX5kUSo1rItg+UbSlXo3XCXwb
mNoY06ZsEJLIBDt9tCLpub05SEBPUAzintluImoKjuRIGjJvLrh4kUxLxfHP/a15zvHMDBqI8e8D
xHmz8DF2Mgs6qXdfA4dJCh9zD5phHvJ2f1p3coosIRQa1dq4MFcE8a7wgk0/dYMV8wgRiPOUMyCM
iM4lx7eszlrSrW0oJPT7L2foNjaot60AmpeajOGD0lZgw0xDsczUikkyQCxLf0Lfhx3W25I6T0b2
lmjAY/8vakiEhPxM9EfJ1ymF4auh9PKJRTKaKoyReCEgdXxEKbv0eaWII8egL8/RVep2F+nIgDkN
gPqeaiArRJAccEyrG4gtqjfSMVkw+M2EZVIbX0ixwdbxE0iqIzdOrba8IFW7oh/y1kSICLg9DiJJ
72GtHnTH6uMTs58AVkkZ38W4Bl/b+iDwZVihHKcQNXh7ltl52H7VCzfJW2FCp8muTgzq67gwJoX8
VtPNNXcTQTmj0dHDPV0iw4GpCQWlolusp7ezURdFG7zB5iXjH3y3R5wZYgtcBT/AaFxE6ij60Xzq
wIeJv76mTJKM85k3rhe+KQiGqOgR9vg63w8p48Ldjeocjmv3wIavSjHhHYmgrWQCVCEDfGU7Q2M8
bMKvwFAxSnf7g3kyllNZSHK1Nz9SsyKS3Vb/EpN6R8JNE8OV8gRjJpTFl70QKwgAy46blbUZaY8/
EZeDv0LWRX6tfSYnTmqEpqlxbhzZYQ7PBQWjBHlEG3NIN7AO66HT042UkdSlgwRJA56TLOORBjOV
ZS2OU8lkpX5YJ7A9fLw8dz1O6qOrL9WQh0SmQCd0yCW36oq5HMQLbBzSz5lW0HH9KULROGT4iny4
mz+HmKT2f2+P2IA2aoP9XDyYm0F6jexih90qOFjuNA4fDITHWoUjX9I+G5s0U15VWesJmGFC9w4J
7Zvf3hkcCDr4184Q9klOIpi8wb3/CJNCzrVvp+WCIxR24Kx7/mU1aHs7BHC2DuJB4py0BT9lRUWp
1zfUKoVDY7yfZeSa/e06Fc2joVABG0ZbX5kqOTUDGuIkvqNHrAPQgsggW0mW9VvHzybEgF6QsG6f
+d8HDH9PiSMCaSfK6/Zx9Ol/piTFA4gX6+v7BbiuFIm5xg9R7bVY8tkB+5LI58nJg5AYIF9jlhtC
nP0zGsYqpk8R7sC32T9tJNLo0LHr/T3zgmC359u8mfmwWV9wFHx0i/H69Dc6DjQ9Y8Gw4Y/7WQtz
YEx42UAtr/cmAdGHFq+J4UtUVVSmib/E1c34VCEdzcOUw7IsEVcg+UAN9G3L+icmsw9sO+VJTWa1
X1Vn8cRe5lzqe3u5fNQLv5FNbD20C0RRMdnDCmUIUvEAIF72PIclTGntQxFj2j46y0Tnpq/i1rHA
gjSWenHcgc0bNFb8TrY4zsz5znKPCYf3iypdOyfXPPdnDXNA+8FraAfK2HULu54VXoZPS1tD7PjA
sN8osd4YpVxnUUYb+LhpSqv4dvHtCXCTsD0OSjj4M7BQTKSfC5C9c1tk2u2wnrOWGrcSQXBEc3Hi
QzpBe+3PuZmzNAJ2ja83vicK+A0txEkzK6ydJ1nyNp+U68aRu1DihyAi/4U8FreRPefDtXTc/hQi
lFM1Vxh5Dw1d9jXCMcINyCuZWI3153hms/C78kN8fmeq+6BH4tT9ILO1XsPD4knCsnUGk3IIqQCb
Co9oKxUnVAhvfX75SFworPgOcns46XCnmOoENLNS0/vzaAxDWN62rQ918ZAk2aDH+k1WOPizQAWF
bLFNC4XK/hjTC/QJkdL2SD1eEDmOECYkIFez0OPYQnqHJMFHVfY9sPn4JOfDZSlUesK0CGufrT2N
lmbhglyB4YQkOZsf0JV//0+YwTqE7eaoImT8kvT0VSMrhRIr6s+//ThMlFzOmp+tYD6QXLWArb8b
YiWVpRq56oZdoVEIRSKOpDjBx4SpDCM/jppW9S04ORsA44ym5Sj6TaCUeYKTF1CNqAygxcdcR2o4
uI9xLldeJFVqnDIPCKx1x4ijF0+0WiBdddH0+/L0+FLFiuXLNsc+Nuh94fYAGcoaQgZfLGptfhv8
DYHQiL/QCSDId8gyxsy63EQVvL7ptzS0RnSyg+NzaXhVU9ylSIpoqdS0RmFJNXs/2JSJzR3lIt1+
GCf3s/pmy0A84rzpsshQYIanJDXL5dvrf9Nj7GgqdzIWklZ0LOQPYbUbR+qRxjy2eUQPiyJ9L2MM
axcu0DZnbkuvEzN9z97eLL3g0DluQAI9Ds9IRyybfCAXVRlHajPC+EsMaFW3zvjAnwrLQ56AFDeq
ISPn3dhWmB8S3Zb5mD2j/XlbBj8y2v13oaBgAI/HXx2I4t3l66tUO9xnbmUWEuPamXr+2mwE9mQq
YFId/z8QRYitG/tvqMWh8psAE3Ot5RgtC/pezB7hSYUGVbHrJ2vGTwKegqxyVj0smzimsy8UlraV
9RZOlGdM2dvFZsJq63WmSvLqk18gHWcvrlw7CJh+3x4VCvuSqMvC3DUI3GJG7ibo5e6c58eJrOBz
GTusyds97HW8vyKPR5B2gFI0d3YvY0B29zE6VytzmrTSSnhpVDHgcufAFi7kLSewp7+WNwjXKGHE
CdUqDBTnFIavSCM+6JonBsZvAwCsNji7/pwkwAY8V4X3YNdsWbu8Q+xp2OVIuRmgPW8uHQSWQTip
LeYhS7a2Ny0ps7ESnqwe9x36OC+Kb0Ib0W9+FTa6kuqXwpVA6gnjVA67XLRrRZArDPtgGA67uVkp
mVPzj9UmgwgwfLc3J3J6loPBYruGwVPsd2rfTodj3+Pa+SvTcSjJ/tyEJmRmCJw4SUlwWSFE5Abv
Mp1Da+CwZZFnlwHWvxGu6ZdcXQ6mHCUjRZzs12UM/GECvFFiypBJYXZx+yiD3JmLExgdG+zQCdhL
67oHnfPnZdsvo8pv+xuKSZIagAMY5y0AmCo3w4ahjsnLYtNAKMK3+GxxX4V7WIfb7SAxzi+YzIuA
zygtF8832P/5WIL8QecUkKa8z0cqzXNpNJt10tNEUWRU2xFRlI2WuoC9of/TniGIcs4UvHn12H/2
D0IEw1/bkXOlLsY5ALoxT/OPonyEUFQbWNwCsVFEd0G1GiID0t73IoXhAF3GTArj5tdBMQQiUbTe
/+EJyL6Af61T4x7BjtfQfI8bc+knxmnTHh5D+PCOo3q9QXWRzTWDAtggwAWlL3j3ig+4JLA53NI+
r8hhA5V7PiO3o1FhdRqwLBb0eA3s6rgWTWP0UfpFN5AJ9pVlCtwI0cClNnlGB7TqsiplgkYMoXO0
FxxFIibYcFaEN7Y9M2nIUm2YXIvrqfMNPrLGBmmnvJEvuFNN7pYIs/4CiPisyXM4RXD4nh6Nf2Pu
WNO9zAmORHeQSo0tBosDeQDTdF2wWj8sX8PuDwYI/zApQEYGzxqa5F3RlFoPiRV+nAiFzwQmFEwh
mnwqQH+Je0SoXnaMH/bkIejkuWhdBNAsQ18Lzmy8px5SCqUJhe8zCs6McVcSONElHOqfp1qpnTuX
rqb6T01FlExct0LUw1jbpcxt7zX5rutJB+d+lAiCmxCuSF2nOq3qDXMmy4u/7eMR8bbIJoeLNYRy
rAnbDxl3K7N1VOLOvrD1MWXg6OAE9gafH5UOFl2+yve8DfTm8+Syp1EYy7NlE+S6nHlXoEZ871fv
wMllDooEabtn8EwjeDVho6qkXQ0CsNPGtrlra+rVgTKfvr0wnb1BeNROfGaMRfuL11ur4VCQ81iU
kVo/MYIPF7F2WeyWAqOCECrm4UQRQkA+I84hR9DcTLrBsvI4FgkrzA4cXGA5iLXq/+2CXAKzwsFE
EOxqMyQdjnz/WCzDaKLWp4/AfznXKScJuTg9de+4O46mZStttO4KtVSf4uGh5I6zrpTSU54BENZ5
ojL9zBIXsInAHvCn99/Rk3chTlZOvCdb7rt4BVxJ6f9mJ/jRnvKdK667qscG7/NX/T+/EpGCFnAV
IA5gInFA/hhtdiQ75STS1F97Liqj22O4QMk8sBnhhPFznCUZbidp/ITsSG7hETAJvaG1yf68+gVX
AdCrWzBS+AoElHO/UQD2fk6M13TzqTioCXR8SElkMMJ+9fz5pL5A4Y8BWqDa/r4TbUxZtOC2PbgX
XCW0b0WUCDK/HuO1YivkVuNlcd5/cKr1ZKjo6NUdtvxdwHnyBt6DUYsQBbR+eObmfIK04OJ2jShw
s+FcY0J9xxLhsuFxaGHy2HHiRjXP/+KiLZcxLBWIj6TgFauwaVTZ0kifpjTLwGRvyqA2zsUv87c9
dMbSufYFW7xQ9r+MpmBaqt/Bv6rWKCceoIwiPInets0VEA1uGHI6OM1kt8Mr4yADgxfgS+oIBNql
b9KVG6lJbTGM4Y00ezlH1AkeBBoOeUFJ0bOJ8dNTEHA24A2S4TYfbgjl5Pv5chBEwEwmuZWK6UW0
H96lSqt0dB5nKpC2OuWpDYIeBu81toZ4gvMMQCOYSfe0DqMWfbKq5/WgVaLbLUCuR6RuxO6TPHuQ
D55PgrOh0gZvoqpsR1GTiDlCuW1/m6iE0jOZ6nTr5O3fHgMqpyFK+kL+dzdb4pUWljQ2htNnaciK
s1S6/xSIRBAjseZpmpItrQSxFNeOTn2jDxu8h8Oa2Nkxp7F3QG/MkZBPd9Nkaq/+bT7G0gboAqam
VGIi5iEQL/TBOr+6Emy8omDPDdQ7ZmI/r3e7jyyBAo8pvH9825KU/8qBkGAfNM2n3BxDrx1WQm+3
5R+0c/A68ZJJaePhgaALwEdxKmZgYL3sBbUOPMyvttHlcypRUr3mx6G4IMkm6AOuq30OdDIRV6QG
veBgmrKE1SXdjAvq6CdXTRW0FXdefp7164X434lk8P1V9FXHlCQYiNr2dvsesWsrGRi1T6nsVohg
EwS/a5ub/zrzpjRi/fLdV+uD4++qvitUenU6FnBfIC0fsnnW5iHAy2vex9XI6rpHnWnvd7fDNajY
G3pFxYybZZBLl9bwONYCgB5uVVXkdyPAbIYNOTn0e+2HPF8kWVLUvma08830W9v1Dp1sb0M1VtwF
SekT/rOUUiOHav4udqzDmT4MCr0fEoFCrifL99S4BPfW/KCkVtK/9ZAKVvsmV7S8JJmdUYj1nLhv
ZsGFA6nwAqS/1LwUIrRwdt8NH/ZBeiUTuZAsQ8nBZF6igBD4HnSOPkF+KDKUuFPZgJ0tunoemPa2
UYXGGVLuQMxliLDKFqGyQ4OxHiXOGdx8KHlBpbDOTUuISkE/scWsbus1MTdEHL7BHw9OKAGp9KP0
7G3vYmsYiDMfgQPqC3kVwOircdMe9dwNh25L1YW5N+QwiFiPZKt33NMxvQtUqeoP7ziGSHZsvw+R
amm16pAysgrB0f7keaPAx1gWpqZ7+elqXJ2NzGIF2VM8otgjIiL8uLBzEoSk7VEU8924XNRgQLFF
lW0zd7oNvgabnOaZitX4bBkLAtCJBxblkkO+rPM8LUGphBC7hNnTTNj2bOihURABUkilxWXhk5v/
SV2Z236LqyZ64fxDEZBoN2vdTK4pO721eB6nfi/4alroeb4EUi6DpMpoNyiq4fISN/w+rD/Al/Zg
uGmpIJiRQj9WIjmtySvZqY1inr+5PmHiAcQZ0asb4nRYi435h3sCaOuJSdsqo2zvEaRr7ZiESwsR
Cn0gDCVlK/jW49UaBtWg9IhvyFJyQGPgOHTkSUFTdRkImmaZo/fuUx4UUpHuKFE6C/lFmm/8gg51
JjQZJIUjUCO3TjzP+L3yAq9d/8PS7VsQfJ5Xv1P8AMMurZv4H8vblsehCX34kmjk01drtKtvrIv+
0RR+IRxo3Qxez+urwIgpfNrCy/n04uugU8PiWPBhu2vWIMdli1N5X2sFw16gH6k6kL1gWRLrBFxQ
qhmZH8PH58fmeeGD7elQP33nollQ1FwD3WxdA7lauHG+xAA9Oe4emyezlrn6ckFFuZbDDlcIf+sh
z+tnOIdmrzjv1QJjsNFAk2eM2j0RCBnF/c0J55DVj1a2/wbVsE9/0icEZ2Z5drHD0OZ5/GRzhvAP
V17i9ThpJVh3EoAbO8ds/EEo810jjMpl+uGBzCRjzSGpdGXaHmOhceKoPNNvpB6FXms2SN8L2frQ
KTusJTY4IuHLvkC19/kwo8GxGiUkU2GBCKKkKRL4L9ORYMsLaof9y5SB6TtktCyZ1iUWMHY1XGRI
xvvJefcn+HSOv/+YahOIRhmoc4H3bebLr3Vif6NblRiHhoYEHJyCleSIUKF7SNG0rL0AeKgVSGSO
UToISg3WT+1eZOPrR76uE21Yc/dq6MVfD4adTAxxGmLzTBlMrt9PWVF+z9MBfSqEthK98r6LvnaY
t+AIAacYPSuyOBmjY+JP4tC+C8fwPobyASY3tpCfLM0zKFKoQy9ljR5HzFmVDKvE6frIlpwpP6vG
YlE+gYav5nrsFDpHYRO7Lw8LAaIrmH+STWPe8rH97YP9fziuHHdatjoZxnqHbQl8JN6Xx0y88yvo
v9Ao/UmdRrJccU3KckOpXYNtjZheiB37SR/Mql1g9FnrhQZngOTUSM/KfHBLetTDXNJhN7PR4rmX
oLOp8brfUhsrWjdY+ynCI4+Ww3Mp4aZj9EBxvG78M+HNofrUf58PwDM+x8r+9ok4SZ5G/0z5AJdG
y22nCjRekQ79nO+s3zYZZK3iCEHep44+/G2BVDayLhXH+CLpii/sL2+nyhomWHdkOWdhcd/NlR9l
/z2QhhhW/9Ep2Qekir1q4f6CvNVU/gyF+IL79SiZ3YTPQ3JfnWWg+E3168uJvmEAL6neYXO437pu
Av81Qq3ThjoGhXzEN+GL+aJc7eY+V668bZOlD6l4EIKRIH3xYkO5UshHeMDM41uIHgJm1QYh8hCf
9gb27sNjpfs7IJK4toOwu9+jdFnMb6GcObcGXKRYiJdBV6wi0lIPNabWaJzo1klS6asXKxlORmn/
hXL8LEUMvMBorAf0+RT3HkChZUUui08Fm05zPv5E3uT8ULE8DDyxjIgiS6Jv+fJ6fXkmIZaAA+YI
le64QMBYjMuIhuu1LofAOLVKGVK7Xb/52m5tpEvaPLbCDXRbFRJ62T32kQ9qW7nhFNAbSbCT1psS
QuNKJ9nWp1pl3KIi5oEUrILUrxq7W5HvZMNcAebQuprTSP6d6JsRxShLK9hUSz0gYuqucd1OBOp+
BVY1e8IcilPyz8L2XZn2tlKlmyhIS0uN71SdsSQI0rUcyxWdH5kKit4A5mgndyCBSq42X94nO7zj
/UtyiS1J31aIsECybrXuB989YKXwmtTDqCX/cuXtGBrGSiFGFFOChKM0FvKgSkkpyIYtJxoaDvqt
1ZgUu5gCTpys0j3c+IqNi7VpGMCknpIscisYifwJlBGikcMIW3KyehoupJNjN+DNIhxbEySvXPdI
b6f7e2WAiXALGO9cMkJbOErAVVQZUeGILdAlYw7yUa3ya4uh7o1pDhK4yjUOZjDxupELDUeaLjgS
qvWL83nnFR4HAalOCy0HybNRFwKDnf5DddXAQ9X67ofkeatxWlIc6TNnTX2aD38FhygvWkROzOW5
DI6ZWtln79i/cHFUuHPrSo9hKCz9CMN1puXunsYdjXvO4kN2UvmgD8DIrGBo6iJwgtWxcp9fP8Ve
uoujhWFgW6CuHJSAlHlimJj/F5w9v9BFrGGS6LzvkHJPXgUNuHyzux2EaMwpnidWWQ2dhtvt92Ln
1bwTzMCHbFvBsT8n6LyevsRbstDIWxTkIXnrElZrzdD9xEaZhDlHl5gQlFQlXBDzgBetr5Lrf+yW
7NOhQdd53HCicBUPEdNDdvYxpGwwCKBp/BOVFOC6nMTVZh0RR7g2y0QFnqorKgRTNpcv+726blDT
+3X7mgmnkdP7RhAOSpJeH8McZvDspoy+m7ON5bu/2UfLogBfWiuLwlYCZUovcuRg8Mhb67p3lXat
HX33xaOY493lOhqzAM5TJPar1V8pzaA8UUt273ZwkZMe5eShLrkF9OHSjarfHN9g3CFRexer2NSJ
wwohhYSKKW9YKcOgZEN1E8WImW8+talQwK7Hv+/oFSUB9Oid6rmvhwUcf/k7F5ynVi9kt5BWM36B
liqMmS4gAWT5vRE7as9ZEhgLzWw6k1wLT1tMQCSy32z7qPpps7pmQR/gqceiv69I77NRVf1PI0P6
nqQjSVAHnqZpd8N0vOwYF9KggBnwVqJyShws8hKO/9IIM5wnoYDyIWX19VUOsBLWMoNvflyOrjfJ
MfIrdlnn8rLSrGj8yqHV0D47FgQJFBFTefQtcO4avBYu80D2PNIVojqTzCSZcskqzSzFNEk50fzG
VZ58ZKMuwpffqTIRV4ol/BikZfFsbQZMbBLwpROzOZ+QwguSK+N6Mh99PjE5hT/fJj4b4Dab+Nt1
oDZoIoHTOttTnFd13HC2n1U5vUeihTqdknybqFYiSHgjBXPBP66iIPE21AFrpUlOZTb2or3IJDOH
8p2PSNJ8XXnDYw6eXdA5rbt1NXNDCMbJU8PzLJ4ZYn9GMMoA1YEbYexTokfxDsvfmjBxeDmiBpYw
rQva/t4Ox+A03UF4zymK+iOuwL6Pt8Ha0qZwIzc/+UioNcbsRYA46yB6f87J1KrTPOVRdC7XoW9X
yy2+icBJAwsU99mjZ8l2L31wGiInyd+WH1GkANp3IzItONdloJl+dc6OeLMF0IuWKuQuql5TcKUD
bDBEdKyYwHm3exdyml95bAugvOnRjdJ6yEvTsBkpzdDHnPkKK1MzPfjnZQQRKMaF/d0k6WjQ/rTr
kpkO/+kdh0fTqwvjq6omTrauh9u8Wb9M60tomYtySiE99F2umaRuxZsi8cxMUCV/5zaoyQKK+UBG
iP7zEKTp33HKhgvwfbzlp/TenRWx9kiffk5azIRmkQaIQs0HESsi5Wsd3VEAo+TurtUWmGgWc/El
OLCW0K8x3o7ChxT3eo3fU0n8N3ehFNhNt2gt9W8LqtgeXvmJ1Xi5GSrujCpuPcXa7LtAGIhNsmoX
A5P16rvsNVC2scrgaW9yAp2eV5nI8OyZZJkMsTSZM4NqSI3bS57b78imf0SqocPxU4E74n7o6dyl
1xVjaNy8UF6LbSppzbpKtdV9CRz+PDK2cW7VnME0YZlRFGc6v+vkQT9H6jOmolPOWWrHNyQO6htC
T/pv0WcHoOJ1zlZcFOx7iN0kokfeMa5X0hV3vQ+vC+lTILCLM+vF+vZs+UODPD0YFZJHp3vUtVfy
GYZzvZByxEUaylQja+S2CuWhxULcfaDKiu6iULUngtiiDzejSTuVVBU/H7pwcxauORHewZ9+QzSe
9JLUKoOSarT3zJBXy1JzjI9/5EGJbk10xXoayUF4wcVWmhbUIrsrca4BEHmLd7wdBNIzRQKTD4Eu
GBJhFjMYnmUVi5mTsqUfOBeHcR30t1PsqgW4MsGe82M1Yi0IEVDpozpUE7fMB14JTwp3Me0KCID/
evp70+93FkmZpEoCERYQbfxZ5zW2HeCx72sOmXDc5x2H58tHpaPrjnRvErCOI6Nv+gAg6WwTmqeA
WG4uMjti8co5VDV47FLMhqFi3Lih0aQV3GrRMmB2hMTeWSoaUgRt1+G2hlCPZ+aNt5WgFQcmBTet
qF2K7wkEWyJB423yQ8FaRr8PVdGadp70C5SvqSAxpBrY8aTK5PmBf76kGcQA9/UW+e1WSGnC6r/o
oV6y5uOVuYgHGLRBkcmnhnKQ3hykdwTWUz8ujZL6uGkaz4HKTE+hvcJBVR6LBWiVjssbLhB/2rFZ
nqbSUNBEdVcPpoiYLY+1JJG/VcfDypFHyJmxgrFufA6ErGX+krKvH1up+cdwnps7w+DvOxxzOKm7
Az/fXnzeBOMoGlsmgyzk4tW9veIqD/mS2kxFggSg32aWKyMCMBgByKPG6f9JiODrMrlfnE7heivh
9CB1XhAFiyOsNnNGk6siwgQ3G0jKvL4Hsp0hAwO6RwZd4V1Kea7uU7D03FW8TC+RqZb2ILoQBgUg
HQ6r03v3sz4J2R3NDEBv7+o3251oPueKiRn9N7eWvAt5XvSLyFvMh2PYtxUXsGcNI1sPdgpaQaZ7
o2DHSAMEyq+zFakscUGpmC0zyuyic6Cd3kA+DYBZgG/fTZFg4azY6OURCU8KnbWZ7UF6/pn4jxQ2
wgcRLKPBNEEIqbWiDCkvF+0w4+kziAaRQAcuMk2iyngmU7LOzJy/prxSGG/HfjwXKBs1YS6khoGI
nuZ9lOdfTfoNZQqOJ+WRU45V7Iy7i8aWyqd5YEuag9levEV7hWVStv5PMscnLzZDI5oxIYVMPrVJ
YlzuqKpJkgLmEZmwO40f4agiTHtdhxvVyYeRmIrBbZCVkMsdejoffor3gIyNHnwYtOcDcsCT6rGM
cDJNVwsjvZ5DtefwfmWrCxQdVxfsT1tKT79HcWbA9lixHjNdo3danjt5cBfjMZ/j46G/xZzpo9/w
YSdCILtqb6O7VO8CxCIq7vb5ZkCLmSp1L86gzXDRc3g+djFo9GxHsChFCy9pWt1djib5GnlfIW+D
+hO6r1GZOMhO+WDaeO4KaewmRH0V0x7Ei2+zjNWbicDzbfgRjU7cfk/+Y9sHHO75f3d2ELor/YH1
zcg6nOHohVl9Vnzr9/M9um8KkMhhD+x61Y1T6ynq/bl+1DveKxd1JOKeB2eD4GPlfnvLKWG7AkPR
rPnBdUdglnU+6ezFbFJcS1cWBGtLOGG54UAdL3BKjOekAkP2plLrV5fqnt8HbXTRaK5XytHpLRZc
HL6+DBQHZSud+uLPgqt9JD2H1G7ByII+t2s3z/Mftw3g2+ZpQ/b7JqVmsxqd5cT/KoF+M1ZO2Rr9
9N+wmpqZ0caUAHKjQcbVZLDprlT2CbjvK6fh5Nfm0a00X7oxlLLa1V3WcHn9YlWYRKIJqOA8NOXH
BW+nljtMdInX2Dy0M6tgxrCZ//HaZ0cjoiki748XRItj0Jr1GncYbEu6vEWfnZ9T2cCDPXfsC6/x
dXxoAmwMYIyytqxSqA3BnbjiFalWmiAKyi2a4HRNpQezdBJ+cSSJ8Uc8+HRo/n2JaZJX/ARywwWf
bKLBnblhVT9QZuQAFXv28y+PZddoDUsJULSFLMW0FjO1L1OhIRukIOdCjTxBlVQMo+f6Y9tfSyKp
+udvPvRmaKYC9qSxqPXBX81/GxFcn0RX+fGQpA7Rj2TGISMQ+2jR5mQS/AX50s4RxcY456wo1nBB
q/s6SJWB3YZcmw2cOcMnjiP35skphgpaec123sGPb55NYctu62K1odEjSZmybK23uOjh+Bmfsc4e
E3zSfCLLjFMiZ6qSNFOY/NQi8HDslTknFBSK8O0P3AQ/Q9dTUwrvpkpcfh2ONfnB8HeIVdfcMnak
0igausN4vb0lD8g3azQjqwD5TkXlfTqSBL1avaW49cRLHFZsrN5dt1pU0Fjf6H3bujqfYdmrQGkg
kTwq15BMabPCYfPuqESRq3TfVpxgSms4H8dIpnGOXevyYCyqHMuSn61LNk8ZeJz2ucG915jHg7A6
LTBhkHbxwFOOKcC+oCS5hLKGMIYwTszHZU/br34YpCQmtgzjHIDJngSsXlTsrfQ55I7s8TXtfJdg
V3pS4AU8VN3VkyAe/r6vjZiivRK3jvlz0jJBH1VCpY1zn+lFJKqVbsMEKHQxFrZafUw/yGa2s+tx
ZuQb8uyb3Uvn8iXMmLa1gW2KrXXRo5S080FO98siEp+iCoPqTlv0LoRmFZ+9VM+jHnu8I96yuRsm
wQzRzSBGUMgxYlq4BeeewmW0OQarP3TeF6MJYSo6Se3VO2ujYPb5oDNyVNHRCt/eBaVnyrorsAve
Dpsxx/UzvFEuBjy//8b+/bI1SJhRZaiBB5kE4mfJ4VjgGYBRBDbMGQzTqGhf7SXLoguPhrWMwTfH
WEmGaa8e2LmYgvVtv0zKRYlyY5E1HnQxyOMmlGL3461nL/qxS+Vrj45EIVFHtZQ7od/sT403TCy9
31XJR7YdtlZl5cKoRWfNBxevP+P4WIgdWnpl5y5g+Y/zdGF2hjA5YXJvhDmqkJ8g8wps2yZcYuTU
zICEYVclhEb5S6TVMlioqd1bANW8CQ0AU/5mdWmQIfS67OEJW7QWF4loWgawoVHw1tn4u09o1MFH
9y6Dajbj9KjIire1HnrPRdbnMW3eQftSbpxtrO6xPi4uT901Jai5BhAYakQuOAE8qD+sznyES8wi
ATSKIsIBe8rieyqDGg7p58El/k/xJtjQp265guilNQ1eQuoqoyWuc3EWjGsNLxl3SOUpTpvYgu29
rWQrYynLWF5e5XCbwaI2o9MpIEg4GFxTBBvApLOhEkMsVqkUH1WBDSp9so5pgqUeHLgqx1BQCPrQ
g3cpHC6zft9uVPZI3hX0LZVi6awQ/+i1qB8U76jauAkFY+5gXVglwTNuCDXt5F1QKnX3i8RYYOjk
MBTFamWhQGNsCQp797FX/QBwvqDlGRpPCxuQV7nR9n8on7EfeXoSBj+HFgtbXU4CYHidvsW43Z8y
OXnQWdtmVSsVCNu/0mj+0SHS6rES8ZDb/MWsxPMYB2DRynO9tKgzXdSXz1/ArsY+wsTKVMm2QPDP
0PJvEZFQKphZrOCcn0YCQkvAvWsIPYAWIm8i1Cn7AIszLW4Bzg+mqSAU7nnafMZF2bWQcywhglt+
C/Us4EiJ8irdy1tE5cgR4H5RFaBA1KBFZQQMH5lNPMkfhfncwTcU6VXpvDe0GPRUU5VvbyICkDm9
8eFd/xmUv0olmHgQoUSSO5CfCpljHEaPB4YjIHwXwQ+BNXGWvuRWMVwRS1QNAnZZWiQX6Z4gOSMP
zSMHJaAEyIpFWHlQu5eLwBJ6qglaepjt3q1z2cPlLPgHIC5R4rbXgE5kvxQ5uEazv597wMUJ4Ecb
N2MmyT8SnVit67rTVGhmRMlyPNYDmQ8/H7P5Rq2yMDnmPVGuUj4MZ0Ui+yT7IVTXg0V8dknKxbq7
B8Pabgxe7bzpb7QEYsNgK2hkQuM0WieVWuJasDti8LTdkogTSc37KQV108kENBhzKg7TQwurVmw0
kSk1Uv3MCNiZh4sAwcoVxXqCMkxEnqDiQyvuEKTib1S2u5Qy+nEAaA2Fz1AjL2XlpsBbrWh3FbQp
TD0GfQ92IOsqFVpE7Z7JdNpgPH5jBp/N19s9GPhbx50UnJM+GYqlF4YKZCZPjNSc3WJTQsvoATFH
tD6XltMHXBNq8x6cIofXbagNlK3O/0/06fOXHzxp4+BVApviKYRCsFDvbv3f1gtwyQElZMCyMwZX
5W6H4fjQl6no22FUDwJpG2cczccCJ+yZG9tWAuJfPSMcj7GJrKCZRE65Q0z/hhhLC1CkLBTELPmE
ZWj1PaV5/4nsFvdYo7XnOqL9uqNiEWnKpKym3YFbf9ZN8Ou950Sdc/krqVaQpKt9QzjhUx+O0dL3
/U4im0cS4yptP2aSL23GY6Wh6kw8ZRUlrm8iOkP+1cC5kMB1cII9FprAmF7jPjvAtBWac4CwAb9g
oGkw0xaIy1JD9du9LgHHnRDbZwLx7ffPoEOaLEjWkdVhqMDu4P0zTKxhAe5sDcaWORnHIpQuaNHB
+iYuuMbJ+5utSuZSPcliIGZ+FQ4BRFRfy9qsW8k/xYaQiWHsm+VxZhp5M5otY9AZqNHHZzUKb307
mJIQCPGGv1CbfoK800NUBnzVH7Lw8CSx597EZLgOipJ6DxJHSYnCjL5l5elb8IJqm90XkWeFVjoq
Ef/hGjDqQ9KS+IxvIBEvutJgjZANO5n7u8dg0P+QDpucXwAtc+E7hS9lNjb/ayDcuvLxsZYdWFTh
/WqSq1zhzhoyze7kRyjRjAEWuT+Wx6bAugg4GrBSwFHgi2NjwQ1yk+sEM7Wy969WEpAfnpw5BktY
ikw4RrLPMU4jyKgAtID7xj2yCHOCvBPJ53rUJVJs9wSBTPJ/+AD2nucmFeOM2P1HepN0GHXqEnhu
VmKAlNM2GB3ZUlmdRphHm89cVoVfJHYO2NTLvREmhXvtkOJyDBF19kH3icGtXC4ltf6SDo+KzNvC
cFPHEHwOGY04R+ZguSMne8l3PcNRwHyrsVr5lPKvHoGqk/ivY/xmOKfeOTfFJ8OzI1xytzGo9jUR
XcfUp+0SWJIcMeTSUDS70gwO3CL40hHHl3sAmbvyZ0R/8l5r4TORqyux+v3YeaHkL6+J8/I3XaRv
+5R1B7UbMZZTqOyIJGeGef/SU371OHbOX1xK87RzIF2qwQOlL5cgDBpoUrLLjqBNdgKj59oIDQBV
LD+idLgagAe5858vWsTEFsh1zlxRcEXZp7+QfdCXMhIXNsyYB9/8RGoRZsq7DkClkNxK3hzPJ22o
jBEBFKJfl1H2FqiPfXlaxcU+xYSyUf5yJgv0MeY+KBAlq/SeuLcYpDarXFO9QZbz1PMzbdGGFm9k
bK/4sZymDnOxDbvTByv5HVLVVRKeUxkdlEDHG2nhFF9TVU3R2uER8r1tbkYuA7V+jwAgbQo7pdxe
weZKr5KiIEmzeZKacwLeD/ctWFX/vo9qNZLUdjLRIf3379e/d6yV3MmriVy4MThHThK+nw6rEieE
eGwXrZGmit57h5HmZdacn4SZgv/d8Nt3EwWWmAGtK9PlOcuVO8tvEakfTHLqPKmlKj7m77rd6RCv
Tz5oX1vUbec+d15M9iZTaNA3J+NfCupQZJE70/u5Wci+hnqPghd7nEtoDnZJxRt2K9pycYk5E7pY
ENdqqo0y06cnS05ZZC7B/cnAQlO7BPlvWxQqseGR1a3yjLEejMg152GDZRdqs0F4ww11jfMv7MlY
mzdfz9YxOtZhoMNpfuRQsbDFuz9liYRK8vJDB+ZvpigdSS9fC6Z7CPne//xqJFGYkgU4nPQigoPz
ptA3piLaoIbbcqYS6FHfJt/KgajYpGm5Z808mtajwvHE6wiihJZs+tmP23htNQvdHJ1ibTFEX6vO
xyVdGRfWfvJuW9lKH6YgiuIvl4rKqltQHYitTwn4MUY3ZzeERd8GpNdleqE3Av1dRS17LMKeckf5
mRBL9ME6UBHaatL++J0KYsrZjJoo88uGMvdU7yT84iOxvuepgjuTTEwOTpChTMHTNh6YRSyZuukj
WVQ9eoDs36CBIbNR3JCYfNf2T9YjdLPMxClPJmmkknmL8fuW+55od/Hi9sDI+JZIEW7gTM88cIXo
ZGU4An6E5rS0auIK4q+lUozSPtqmQD7xFuS+l3zyIDUfJMICu5WuBI6otZxGifbui48+g6ZihQyy
7/ycxKCek9apS+LzGY9V2TWCzZTf3qrWBgbbdNkQJDp+luDWcdYF4LJ3zRDjntVqBaxHfBKCUjaC
QRrHOm7rOkVYlWyIGaRcdnEhrNdaVeneuRJf1oy34AEigYjM+sTs5sRbUP6sXwXM3ySmg1QhBo+n
6Rb61sHDK+1fjCi7LMQ6/+tnl3YosV8Qavk+SJFg8uEdrHt9VdlJAYlYC2cdqVBD2m057HjYu6cN
37F+n9ekngnMsGBhZxCGOA+AyBDAUXAJpubgT85347x3i2TOYomSt/YNQZ6n6shtRLaQhUi4Z8Xh
/7ARxllW2VUnf0RGs/groInki9YFnbytqt7JtJbxa4EgrX61OlHekv4rTf4g8Y12z6Mte905ouhN
xEwZCpcjTMmibs0yh8p5PN0XreQU1qyXerWGF7tX3Kxgbc8hT6pYz4rmJ+Bdclc0V15n4lEOegfq
S8S6i+qDer113umlQ3DeWN4BwXiHQzfvGSpjjKFki5cC0AC6yZkWzvHqplIOYiLiLpl2tQS6OEsR
rHSkjwhJPV+070ydZ29jgzPfUNlQIXWg6OVf2d9s0PmWq7sX5Nu1ne3pe33GW1vyv2lxaKt95Ekc
ofSYYb39t0wdHY2tJWq8EmazOiIdppOK49AH/DJw0p/3DlSr2EDop8/qyEo5JNf4tlZ7pebzJigr
IPCTJJKEmag5aSvripQnYCp9QDEQkC6FtF1fpEYRxT5gT3YdpsLdlVhm6izSNe0U636GmZ+EfROp
pT8MiIRjwdEQ0Bf7zdAJn88L0GDj1zqSiW3zEt6nyY/kHPqRTNqQAaRX14bS8ItjG0S8wL8rEMky
MlV/GB9WQHRkc2uv3ccc1k+rCKI2Lrz2e8rLXCG8YJif0xhsj27/p68FC2D/cfFIabqM7obedJ7t
Fk/9Mn5Hat4dVtZDGPJ+YvD6//I1VQ4IhZ8W0JaBjD74k8U3hXZ+1/T8dytMfAr3zLXGNLBoFw4P
3dfY2BMpEAS37CpkCBZ+RvjhmzARe3/9vak1Qw2BqYnetgxNXZREIAZKda3+SVrUJcwTe5jUdy3u
hjC96gk9quKkPksshdW+cwOVjtuv5u+2jlID51uIRmdWUyxwGLfLglwFRLpfRxp2c4zIONjuCUYS
RiGISpWh9pXXCJN894gYmDmnrirPHcZ2gcQ6d9B+7Egzwl4a8lr7Z6XcmiuVWZ+dt07BJWpEB2Ew
uaJhpNaD2DSJlzMngyqTqf30HzQy+4KI2zTGzL0Rv8JlK6KO/dfhJQONimJ1gmQyVLrBLataZoW2
Jw9nwrq9nAiRq4epKx9uE8QsBA17v/AKYHAM2Eex2/Q+/WntvK5ux5c3DIpNK+1a1UIQjFNufiad
4Bpu6oFLyPhxTG4t8Vg3yeNAUAiffT6Ql13qQHhnrjlmBDKMcqKHY5epVmVpCCyS+Bsj7FGoL4YC
4NzchuMsv6O3ix8ezIB3rrfsUSgHbnDVjFagBextHYQdHiA2MP5FPJbHJ5LxK9d+EAkJF61Tl1sM
6iWWi7Pp+5KGg8JclQi63xFJI3+atJsFhRGdYkqKqgsVkUuSQw2XQUJNuG1HmNVMqAHCRrcprP/O
VtgN2vyNKUi6O9wnt3U608TPzVvhbz0BZzTQP9NyHQ4pHCeURNOftWYmMo9kWKcMiI50l+LMozWl
HnwIWxLuk7XY1w2/hCXrn/Do8LrvzjFSkDOxNvqeiGFJZz47KBxgAkKa9ZmsUxp8y7ey5A9mnRlj
+TDYVF57L4kGSU4GrNrqbNtK7oLDdyRkQGZ8g3lSGyiCh5UN5bpEGUSOwgoJGeYx76lStkhmgWwS
E9qRRSKDMjkmEDjM8zVsF1CVWw2B1HTrXFSznZinOs1hAM6L7E4Z6pLMcYiYje57baMuzh4RXRqq
mikImML8nSPlHw1Rgmvva8ZVpNpf+1HRn/Ts1ljV8hr7JoEn/YkPqrOdHZS6WbK+H1KoJ5AS2eUS
miRIe0AM7enAnTZS9WcuF2dNJpuIndHkyaq+wWjuIDcA+6Vfba09WTCN/QJJd+jg8A0B3nzkYseC
frQvHw8bAAEiDJ/rLyVk/12OHdFtChzoQ/F4R4LAZUte7yQPvEbaVUk14JuIHbyWnjrm6ac2PNm7
rAH8u6ACOR0GNMMus9tXvL5tO7IFMd8LR5T0kY7c0zea8E7zbaOaXnnIKx4bSii6HKu1rsuAA29J
OBA6CL84uyOAT6N6cx3pOpWonWymZYapd6l2KlyNMjXj1WUvJavDx883pPanXAfUMb1/gdAh3A+Y
OZiLJ0Nu++U41/Zn4jKWvF2Iv90IE/47nK5YyE9dVsyxfd2I6Ccr00EohDaj7L5RB46+OaJ9ifp1
0RxFvmLh7eCVSWkfCuUotA2LZoDi4nHockvhbcNw5E7niDV/JYuVHEe39cuG8ErekmMGRPGHJvHy
/t8dY9uvBRDI47+4RZzjqrLFeu+zJXNiU8wTjOV9+ihZazorCfjlELYdAT9g+XvxKO8xloHz9aJO
OZ+MvFT81dcuCrpMdxg18Ix/dR77ittWdGDJn0IHi7ZzNvVJpLfYLEtFu/JYpjvtYQsfa0Bv5SU/
bSO313oBS4EPyWn7hMf3hAhoybdRlVxEksVA3Tr3+StqqzTJYVWrg0gdfwLTFTb+PzX44UTe6ZCz
2jcP22YdVM/MOcj216+Q+fVG2ncpZIHgeJe5VTWPR7JcgGKKfto9rGM38gxeb9RcXiW9ZbeCGLns
SCy8Ss3UMAsRnw8IiL91tuSWYUNZGwTAVb4pNAz2RAjOa2MMfQW/D2YGpU5uQUeDbbjefjMyRZtJ
BJU20vrwfnom9yCgSKTdDuELqKBUyNqm725aMKH0JCiznbBcjXvhretQxnWzNpyFnlElpwLvfp7u
zXpayvrTpPL0feZdlFtOm1JCfmgTGN4kUtHRYoDSua/6X7HEykEmoBrHAe3cYxRqxTEcBmQ8bJdt
T8f4Bz3ekKE+YJdJ5t+q8Yh04whCkTO3HfQMhxPG4mIJ0u/EVw7WmKZ9T3WFWYtbSIzoVQs9xSFM
Xv7FkmkqeVhmWoRFxnhf+vbb/BNNOX4GmOzXkXMHAzQO0r52zs+Uey8tTxEVX+AXxafjTSQz3h70
Apppty6jt5Nzm0LkT0jS3gyua7S/V4WX9zSXAfjWzKyq9TduWVGMyBnQdle87nh/jvcUbPUbqPkB
Yub6ktctBfQ4mGj0fS+lcZjwaASf2l1pZ89iwiMJQ6cf9uc17nX8MPf1WA/Sm9SU8qGrd6g6ABDX
l0N4MIABn6a3fMg8ccVEOW61BhaLLP17Qrvkm8i0Xk7jOeYHiP4B5O8MzCy5Qr3gWYtH2KMRM0lJ
4S9wofVun1VqwM8LruTpuoNONEQqJjI3SHLxxtVjBbfJUAu1jUEN7Rv5kPKmilN8N1IThRRoF7M9
oSlndL0wy1C1RdF5D1UClQHq0OC7g62Mn/XONahoSAYDLKEk/0F/UspYvR5c2QfpJtK8qUFWaoA+
uiQczbf40fri/MO8iD9kx//V+FzV79YF/i3UGGE8v7bERv154QjHXK9lyLk0v3rB7i4Jynv/mRQ/
7KV8koZDI0PneX9lDr6J7Zsh4OFtUfO3XMKNLCBckWYKVrCGVgm0OE3QYVfc8NO7Bkc1eFN0YTT/
tIw4lzEGZUAW3yMEqMxCQEHXsMiwoIJJZtGvO8ivwsynbnBV80jJdPHt0CcO9Z3tg2nPRgVJxgWj
RpnFle7ExitfztjRa/DwhDvSxzfGMFjAz8qQVRkhF4B6D3efBvy02swmKjNFsoBe/uDbtzIuC05k
z4yc872Nd1iK7290jyFcBHvK9BkBhioCbOeYMensA1l/aLqcaRoINZF4lpSsjcBE/ZBf42opgQ4l
fM2vRdISVxqhsxwvGo63qmxfb1m1vd4UAHq/thMbKXLObBGnNx5OtpPLSx/62QWA0+ffT7CTjR3t
jCte9HwzF75YspvTXK/z6Atl1eBWGqQdxtzPqau5X374PeUCeLqyIejGp4+hmyIF/FXdhBGCPiRS
ONwixHcD9H5FLQ0KDa4jPvWYOr7z5plS5HYSYXUL7klbtuYvh1uxMsPhHWIuT/qrzP2q6S/otMax
iVgWhLy9tPFzfrTln60lUtxDjXFgaTTSqlIRffyR/FaZ8Ju4q/Kg2HYBN+5S8oOBWbqMWv5p/ejk
eKAi7VIW4ZCpDE+6bB7SqmYOycBqrT6xmnpt2I8fkFlCwIS+Gc7aOL6XTrLpmfHWjbYKRCccNq6b
n4kgEyFHCk1Jeka5LYijlYvtfW5zL52DqpqJ49CYH+jd3Myy8ABsCXR4mIZ0qLpeOb0uPjA6EI3D
t91Yh8F1UInOTqmn25b7aOWMnAySfawPsA778jaUMhrHcs/nGeY98XhqfykWlSXv85aKDvOKcuSM
nZGW27CnhpTDPIbELjJUqmH7rp82siNky6YmgAJHT5+eZ1zcX3j93dh0TuVWjycxIJfcZjEAaLkg
sOTgJ1JUNUpFmY5khqa5YKKCd/LXdB3tyDy2eGoJwVnfLTL2ci0TkGnC09wPWFe6FitdFPWDuwuF
s1B5pL2bL5OdPwkdfQu8X514VXnMBWzDe50/RDo93mCZ3c53F6ACOss/yd9ZQvjTjlAx9l8g6N59
9BjFvXLynOj058RS+5Pp5WzQfGo/etEG+j7CuSb9y4wt2Q57SpLWkTFBJJnQiyNtEV7xSObJPgQo
zl2j+f9qyDT/al8DSOk+bH9maXYhCUmX3bhmC3j1LERwr9gUT/rB1O8BLtK1zAgD3q8cSh/k7IOM
S/dQ/6D/Aoa4j7yOvUeCcEDfo7en3mqoJJ+EJyc8mh4T9QLqysRC9c6KdI6/Vu1jVzYgZfT/EdFR
YEQ1DxyfPdEm4HiXTcwDcZl1tjZLEQqcHg5VyoOlhuerWAcmh0fnHo08QUsBLH5umBuV/x1j5sbd
3pcLQndXvPbJNnnuYnr9YKSIhuMVWH/OBWsWe0mwRNwbJkiZ4+4y4BQvHO8acINy8XXr/xrkBoSY
lepvCOXCMtY1qYbqxkfnvJubbp9GmUxTy0iPetNCcJCMsAbfEkzr1bKp8x2FmuVrlme4WleCxO4U
HrbKPvOZsMJWIPO2NSp4hZpFGhJXNng6IdnRo0WE0JsWcSR44JQwHsq2W3TlyMJSu8RDOD2hmZSD
8LedR/+FZbUEigvT/Y0sSSPFPQ2WCuvXw6Uqe1/V0t8nzhmb1XpRg+DqFFTN3skNz4byY754m0DL
+v7ShoP8UlS2L2yzDXHz5wDgo3I/hl57fYCsvSvDulNsQM5p+sR910rNT8neg4QJlX/JkR3tIMHr
+YvdbnIuODq+mVEZfbsRPNypBAaj8+FG9h7uevoVxyQJFeKH/7fJfKJco//Wq3ecyccXcuyXatDK
wDeehAvAY1GMLmD9TIl+f82FmuJ5HThOGHi+SFfecVlHIqDpmDzHJ7lUgbQ+zcIJPVF0zVbEg6Ov
5Sl4iwiVbg69vedokWDCkdlIaKvqo2oxjD+vNyRwu/s8ILWwKiWS4umqKJ2GxjV7SEcyqWzL1Wak
LyVINQPkTHbyN9PAop3ZA33dtxQMz7RYiusbQ5vrxd0vdRb6dwpbJP1zQwQz76b2jJa7wiEwcyFi
WuyY+mD0ubMgQDxc2LD4Q8m9/03I0y1uLk4UD6L2xNA9Rr+abRybj/U+kyMG8uF4GdOuLU7dPUMV
RL1OUcW7z1bsUtxz25HfB5d35t6K4Lhq3Zk9Q2aHgeBh1R7dT46LgO/eZEzXWBROq0SvUZxQMWLw
t0qwUTjdCq8fj1vQ84/HvbIxB4x6s+LyKbluuBudCmOupC5jOjv8xRLDFxBnVJCURRsl7QxEXlj/
L3zzmQn/b/0uhrTT+Ra1AxUgTex4gthfaJoGxWZFoRFZmOmcnMZBbP6bdBxQEEO4elGGkNmViIt/
akoPG6XO+1p5RfkhuckDEs9LEkB1jbNp8edpkhrlCRg+FsdYhTzCo7fN8rHMtA7XKFJeqeSSe0Xc
FrkZS8nbhLzp3gwo6XP+uf1poK3fnndhl8/uUzmsTSqNAGP83Bbq5kwBMIO28SNDWF0iHC/eADTC
Sjm/xpZT80I7uQ5nAkHslgYDSkVrgF6IvuKSuICVOBpmMbK/r1ePt4NYi0/isV3vZfEC+mJh3GSN
QTz+8b543TlAioxKgDtb8RSW/a+MFmA70cMiWPd12mnNP2RTywpVu5akicG8kYy594IO/Xxg0L05
h5bUZY/4D6LTc5cpUDL2q/EfhVtYu4lHPz4M3efZRnNwUU6ShN2dy06pLhFawIzJTLSmrl++FdrW
ZTCwA5u24yzlTc+YGtf4Ra8whnMzGjddlo+px1AAvVmoonUrPwk4ZT+HA6YaKjrp+bqZw9gCKp2y
x4fKGIWnNKkQtdJrZZsYx3dpGBjpPz+UlrjjuinbQciCn3+qBNWbOQqDCXVCRJSwqSO9JDmKX7Ek
rg015FrcQ8pAlbonyy/RQphLCVeGmhaw7nVJF6zjvnualRUq5rdAwZvIYhEXC9mZqGIQO/402JG1
aZhXyzbonh0L0dacJ8xA4vdp5nDsm1K1GmOVTeuMit4RVwHTudoK02Oa1lcd7GCf6Q+7Hdjy0szU
J/CeLmQ0NlCm3jwzlDrgte5eagG7M+KdUF/3v/LcAlVVtPMqcAVmRAlTWX8WPM1TQWbHgnEfy573
muDDeGnxDUyI0Sv+lCW470e9lOv8ZGgsD+DuWAm9O2Qv9ZmHktCFNHAZj6dUqefNhNzrGWzvrh7N
lU67StTJIqHeoDjxPqaqDE05h37apYshj/IjOjPVFHUR5m8MSpIbrlXpPFd5z7UWSsaYV3dNfIZ1
LclV6kkZZX1ZujubLaatlVEukLZdpCaZaEmdMsSGyZ6gD24+/Rx/lJFFxoh4PXL2VK1abnmkfY3z
WwQUsBJPiWBjQrW/urLElEKFTVjL0R47i9HWzhHtkrKowAF0O3/BpiuYmKdzNwkYkxkSI6FCOYji
b/sVb/iGtxLXfdDGAXAmjpqKIu4jAGlZUZIUP952b7p5FrIJm3yx1A2tAn7lPN+wrmIatjbksVZU
7s5x94jPTD37f4mVMycMK/YoKNQzXgXJns02IDYL9QTy40/urqVc9BaZ0Kbl2R8Sd8F9vhxGNwp5
cZoCq/mLHFKDNfKmeFlsdmezSixQNbh9Qrspf0jvrS9qiCW8ZS8SPP1SdFyaEbNviRE51mrT4PdR
1S3qQ7fmmyve9A+onqMajX26uU1IgHzmaLMdZ6P6UG1UTxS+MJQZovoBSCgs7UryCiQdC1Dqw/Py
aGCo4OGBS6Xno/oe9/sUi2U0NPWlR+1H83Zrf1ncpzPvHTUmLGzR3PiAz2VCmcISRvqv/GFQGIRC
AomOiAicEcbWaxBUqHoQPlJri5QI27q4iHTmyOtF7Ew+//uBy3XjW39qt9ZqSyvv/UbipC3I8HMo
SSHt2MH6RJdd2WXWqYT2cFXVG2ykYDlDBfFQB89QXwtonrIvqjlEvp0jyzVhMNjipy24SpfQKVhA
/h5QaNigdkVRZFBXDaCzyJ7hE8Hj089KXQKA9nJpNEVqMm6fca3acXHuz3z9DXLYOXWXHAd2ssW+
K0Mo1C5yz1H+xn95Us/dIiHbDXz+hnxXxwO6sZLbZSIQgifDPafIGSABRoG2Kv95PhQfe/HsFL+t
e83qwXOxUigjpbo/k173UKu3e4XkDoEiN+pAZEP/v1sgd3jhhWZwEDq8DNlacbLu8bY8DVxbZYSC
CxiKtr0ppxT8pON1fhIvlSGcz7YyPbH8p7bUQOB4kcF6fPaVBWRp7tgQfXqGYr/qanK2XKExOi2H
INVyfTCMhwna4n1IO7FelKt05PaMe/MNP1iJ8Y6ev9A2pUbJNo4KUXw6o6+0rAguMsOTKOfuedy8
Okit5MpNLF67y38BxHasGVn0SZMBCAHwZc3AuEcLbkn24ZFOAI7hDUkWb6KPQ3ICEq8WnK4mzdbK
7eeVd2cPlQcjMiBDRNHW4Y3Y80pvKr5NpyokSSGk0EAamA7QkkLTPswq0KA8LXF6ElWaaknALEqN
vyAherbrFyDortrMmAnEnMajQnEVBt1f+BsfehTjj62BCurjCZR/dYaVO+W2LzCLbplQ7s+HH+uh
ZMAcF12Hwtkdu0CHnYFQDC4thbDIvxQ3u2WK7c4h0TkrjhMCkWML77Jvc+OKz3n7qfvKTEj8JRxd
0cg7uvn8wFsjQ2bDAYqlrOd51+olC5ySOJGHxK/WeKW/eXXgb9h5R/2srx7lBGuPd1IyuQ9chknp
O801Z4zQpJkl9ahDVeOrWY/4eEGimpDR8BDv2UXOVdBaRHEuVwmppZD+KvvgSy8qpF8VHHgPpk6K
CKkq6yVMXJcmZBAZRwuj24ohmGsg3R5kj543gx0mgjVNqc4uOWVqq1GHe/hZJd55eBbpDURAW9Ax
wQEXPtc0c4Zo3Xx2JZUQz8wQdtnB+1Bk1o2hCe4rTUEvu+bMeawSj50IgfYn5ERcfOSSqUoeCpZU
+FwNsSxDZdl7Mg791eh4ZCfawL6QmguMzEJv6pzjJvzP72ExQqrlVmUXzH9yJ3pH9ll1dc1AJuN4
JZsHVDjZ3on7VvInj8AklqMTH5T3SuIn41BgK3TiShahPHI1kXtI94hNEK0fTYoUPaa31RqgKTu6
YgpoTWw3rwXVr+2BxsLhEYS1IH073Ri5QRXPMW/raJcfHL2uFx79i9DyNapcLmarWPmJqW0zhPiA
XE7ler0j1bvi8fHh0N+jhP4uNdaIZw6x8+mjI2GpsbMWrNXtq2gV0Zbky5lJLvXtXg+bk6qsuird
LlbP537k/kk/u2v92yNtT9wrui7VC72V6U0h262IZo6sCGiiA+NnWYCYBylCj38vP8DrGaI1GaCn
ORwVGslrkiX35FMv+8ZMW/8WcbYGLgOME7J37+B7LGiVTZrcRM5/3ukgBiJIkSe1KU+Lu764xChL
NK8d1ly2Ttj3VEzgs8gcdycoLmnKOMwCmC7p2xjtCIdcEPX6EJYPOHkTyqRajuwkC2uPFB6FVikS
f6gBEtIGa5oOg6jFiRTOIu9ftfKe3fjBtLT3lcLtaDmNuCWEs3LnTOYkYQGHHuie4gLbd1rwpMJ2
ldnDQpZmcqMhMDgqjPiCIYfYqJ63dlNjpDY96xVEJNO+azvlLURnCE7AHb+Oo8UE5RyOyMYbTMUx
aVrUsI4ZmDMUAqtb/CdQl20J6b7fU79qyj4rOP70cJZbknJUAySjSEMS3X/dFUz9HbWIqK0cZk/4
PcrpwQnK7kp/lT44q1/R6kkg74fzKItYyRTcfefouZq9QyYYz2VuvNC/yqioPhCUnPw2sqQ+411e
rr8O8msQRR036xwYaYrvkI3vYId82zcCUW/n+nsRWGx4wfsv5ureh35/SeTWgNX04qHwYD21tvPN
fXON4wWyOytBEbF74VWYRQBnMU0tlSRfxuznVB7CUlEmt/OhacVLluF73EDo1FnX5jJkwSkgjD/J
MlLzY9OOB7tNHXG8Y3noAe1ddp30HG/nTzkr2XS8XJYzcoB5c01B01a7CU2B8IozqQR3Y5LMr3N1
/iPP9BxD56Vw3qiBcGv8LSOfRj/uxpWEuM9FVFsXNHoCqR7yWhioLFMnuuMeQEbDBFVbGR4Rpq+U
GZZRmlO6DdaJGvc0QDx1vBczJ8fv2s/CGPxWKgBNUfRCrYOIGFYJCZ4HEMdQeKI/LVK2+GYkLNNR
UQ1iRKXj/zs91+s+NhRtMosd5LlpNTIuOKY5KxWO6ZxiI084C8OUYTxMyr4WpP7S7hMoVPWoA2y6
971eLFuYgbYPIowuUCPaOBgV0yDtNe/RP/n+i2S5YAA9BceuKoeaamN2iIVIcZhxk/LlZWGzH5Sd
Vb4qlNmof0kj9oaawdYpBKH9DHKQSFzXhWJ3xie7wkAhRwkyE1KrXfgaDV+gIhZhKjkmdoa1lXU5
FkYF+Wmhi4NFwqWAcEYrGRYA28KGbIX8UenNqsIAXbZXfohMZ9HtBVcFyVuEM8LMkpThFMp9jhCp
Ppof6cLQ9sjc4ti84MsY9D95687WmaxGHiQmqWUMJpakc2sO1xaK2Z/2Knaf5Hk7wWjPr2XY8eWp
6zXjlyMlLOdTjMyCrPfgV2IvUxIv2TqU5qk+2Fw4IPVQXRl9EekJI9tUDb17HkartgRUhQrEV/r+
WlSsQkv8jqnmZkBhMqQ/lhSWOxP+DzFpHGDmNeAfxKMwIKQgoWXgAgROklFB1tTpf2c8a9jmd72c
FcGWCBbDIykwT3tdT2k+WpLPKkCQFOBexMSpahKrMI3z4CnuX7HTY5yOcKnhWcgnTlNYcsZK66uH
2aIoXWwhbAGWbWfQG3zcUEWQHnD1wIkZZ6QomfpocYZDgBZkVLKruFjcLiWMUJ5DF3ubNgNX4pBa
2DUhkCSIYdJJKoXH172/qvL0aCTVYF/K7A25CxKJr/aE+gOc1mbrAc+sRntF+5CGKSLY6eUfvG8F
4jWxG2cn0SrUn+JStIyDAMBM7cIcDw2kCvF8WulN5RCUae4g1WwzQXJJSH1uSnfBynn5xo0ulTzC
FbICxEQj1T6TSCreTiKbSAByQfiZWKPENbhAUqBdw0kpN3Lp+z8fnCVJX8Nkqti8UWtrQxTT4sG9
DDpHll7I3JTlHuFKja390ol8ezopPeSyUyewrKqavhTHL8ytYytlBD7kozcD83BE+VvfMjh1WI6j
tCIsj9KGXiWhTiy0x3KQOXC+gZMBOF+ncmo+WJ0iqV8cRQhcig8EZ2AjuX/EwabLDc1BHb0G+r9P
xoUJU9+Re/8XSKxFzxpVTxxOBUEYQWIyD5L4uhO+epAcpLqYpea8IUUOGzFi1Xe0rRzB4FHaKiy+
WoEefSfSOe4JyLaJqnXX1jdwQFQOBzLPUfeL5GWgh97rjo1731K0ix8G5Z2QLdni6V5AMv2zvJl/
1Cv/WOFsiw6NWI2BCYnvcSraKCASCqSt5DdllrzVr4lbYpA/z1qZZy84hRt6lkUZ6PabMde9l4VK
8vJvcV+6evADZgTHOnuO4CHBB+ZgJ9MmnzMX60ZzrhwgB3KR7NrqQ3e3k96nLRHReLzpZzkc6NxJ
AzNKDRzGHJOlAIxqSey3gESxhWnTvpiomvkFjxDBaz51BsoYIrIyvpoxpJ5kbdTBqTFpIskvDwPG
U60PXoTKN6V1sualvvLsvsz7NHzU1c39QluzvNhOu/p1na12/qRflarVEota5VMMq6gnK5qGQRgh
MqzB2eWX+xAOqm1+1xAs7Y8I72WB7hVzOozPCwTJItgYmUI77a4Dwb5mOYZVNRae/F8NJZhzA4JF
geTdna29OJLpNa+OLJw9uVUyCAzHXvGaJCq5gMTbfFXnih/5NxNOVhw+7YTo50M0+lcFMKtPVmv/
aF2m7uEBdUTM+8hAD2MR5tvpXB+ULcD+HXbZCY5L11zDmtivfGdRtzN4ynXyeZs2OcdJ1MfN9+Xf
17hjw7PokMBRPBfMBAir+2X2YQ8L+D8sLckmpMAApuJuIRwrM1mjEzqHNsOR+hNv7C0wTOfjnPk+
n39P3GX67OXYmH12ngLKOxvCYD5OuHeCTbOOZ8QUOITvoPEy7tsyfwNeOAheTYACdXnxUJwK6pRi
U6fKzoKnY5JK0gPC8JVuruEt9sb2Wp+UWstcqCBJB2nIKn8r8vTBeyDW/Mer2tss3cfEE7/Gmhyd
IUBGfMptoJ9KB3wzsA4i2Y+PkENCM0fS8tgP/aw81vSOIUO5WBA17XI4vylbFNbkzZp2+xag4ihG
nmt5+hpoeXGkf/K0mmcFTSpITBPETqMNgF2Hu91vZG/z0F/g6eS/AMU2MXSytx1BqAYwkqiFqKKX
YiAgwDBv/5AQPXlEBvJPQTIlz5Ejw/kJzHQRtvjnO1SaIffGiOLE4w8VnqIFLWi9WKzMm3C47Zfp
LHr3Ln6u1x5IE+akfVt+XmRWlMtYd5CZhYG1oPFiRmfD9M9sOaSkFbfltm38FHszlr2qgcXgUgF5
s5qvimWOw5l+h1i3ORa8MaFtZtEHxp9q/VsP6plBV7QFFbJq9dU+hA9Snmox3mpZe2YzQWYx6WaH
hk3UDO1l4XZjcUDIZO8ULK/H5Fzm5kjV/ESEgqPfdhSeleGPhTVtYau+7C3lP/kKFo5ANuLVlp5N
5cRKYsZNYv8GAErjPyBEqGFHjEyo/ilyIpqKz3f16LLD0A3PetKW+vwTkFFryLYruapIE7SG2D6M
wsgW3qMWFNW0cLBLjve3LREalMblBFQvN2L3W1tcRG8e2MpaU7v7ozJt4uknqYEZ31gDcy72akGh
k3zClepferAcTXWg3YkGndU7h6zrdGSvojuKnoUoD16KWXti+Eyde2/Y+DU2nawF0acqGgYf96hA
E6eo/sCxHJmc5qtzgim/SmMYqMsRn6BqRyJupQCx2prq7CyuDeqzQjdpVYOuh0WzR2DZobRwZplL
2jcxvZACrcAFPKB7JHMXVpxKdV/p9qCWJAKYL63V+836gtCbcMjh7Qh+g8RL4/8oXzt95mWYVsXf
6y/SnDftGxLn0mmN5K0uZLIKiQU0Mxx+Al5bNFhTn6sYFsWETRLecJh5LvmSQm1/lPLFmbJtUCJ+
fmbjWPOSiZwhYINJ5jbusQc19TfSwqHD1T+E/4mw6xod4bwIp1jSZs9/6eKocwWrFELyIh7MnM7E
Wkb1Oy0jdjbYIGx9jHyROR3m3U9CJNpul3nKluL+9AueMwGznAALE50f9SSAie7wTTtbN9MKRiU7
iAA+uzk8BLxggO8YdlB/WQzCuJFdMN2p4H1caW53TE30yFSs1WVEQEXfDaIb7hOVGPT8lbAFRGNQ
IDjkoz5Dvb1IXQouCMIk8re4KfDGtgDFfn1sT2sxU3MawwL+fU5sl8j7sOPsSgxue3BZJquiMRc9
DOkoUpw/Hl6v9+ZxVWPICKeoUeqTeey5lcNdb2S7np/H0U238UnGkTUbQxtgXsGjJNTj4l+t7hK+
Ffs/QrM15obagymJW4F6S3LbYR9QRy+DuQVxKQwxO7/uCX7+2mFCmMTnDcVt0tSGA68EqKBeleI5
zZtz/lDSSe70eEi2V1S2v8OM996Kh2o9Tn450t/mtkjj2LKxkuoxusjpcc+NzZF1QQKqXdpoBS8m
tDkSWCilJ2F6bE6iCZKhDYXb4ozq7V+UuhHpdS6aFg3EbhXFr7WkLdO08hT7x19mSLkbCAASMTZl
pjkxiZgGlE/KiWSDUnqXjWLGmfnnOOCvexCPcZp0AJHZG7vHeZHt8KxgljY5EWvzO9VwrzSwuS5a
bfZKSRt0YNiv9OFGW5wgm6QpluoECN5Xnt/fKQq6nXocpJzegAgDnL5e4C8btkpKoEYCIZkdwC5e
EzbxY8inIfQ740S/iqwG8D41aFtLFfoCnmRtnMkGAJhg+9iXaJh6lyqQ71QJUlLjvtkSaGpCS/FB
QBIBpd0u0+HSXGG/3PTvAO8uQYtiMTl88N+mmL/i84C6tURzZwagSvC4uvFa3H/GQ9asB/GvcmcU
EFyIfPTt8fEb7HgvMp+84UGBLn7Y6l6iziCNcGg0yxCYI+J9b1LQT2Krfx5/s4biDhlLgnLTwoL/
y/25FmK6U7LcnEAdc8fJiM28jSaLvtu+8YqUCWTtw4GK6zKiaqr63teibjlFC17OZS6aaqk8+MAc
GccvFqm4lqwspa7jkfmWviKnUWxZJS2jMhxO/R1VvrCU3K0xOHhjZfvfrRyXc326O6vpPddNM05s
7rUklAAr+ZLz9GRtLxBXhZHh+Zb0NLtm16f9gLyRTxwb9R7w5Fw5CFV0kqM+s5GkIANZmg0rInCp
422yHbK4IWzNO59yq7YybnU2k5rF+HAWL4cbQkOY0KiuDvag7LrgEvllHm3r/tVkTT+VtVH9Gzmk
hVV1j3a9BpUdbuqQqcdMs5Z3NzGRKDXksrcJogu2jv+C3v4RUhuuE6/dpo8z05A2jVlIp3vDCcdu
I5z80y9lVJ6kTcPtkXiwIlRB24pHiQ433P4Au4oPzQrFziMNPW8xq+XyAv1KxtZ6dyNQWxySkKj/
F5FlhduBXdc/wstcd7QI14S0BnCYFO5KIlMZG1TFb1F13U3NfiPUVYAT/ObujU6dgNRxdIXZaCzt
nuVpbkY/ybzdmn4x/WLPCqsJ8qf2kk6VSKJJLvtqMIKBHognEPSb4KPL788BCZK/h0rcpretT9Dt
KZpHxNjX2LGtRdZ2Wl1xdb9TZpB9E2THdSAXMXCwOgejaAQ5bW4W2HUoB8m4aE8ypA8zSy7wCyGN
qLz9GNMMu/DdJGrGi3H7teoHmr/G1xKEObk+GQjfetMnfwQU2zGnAwM/hVQBS1zyBEJ9qfTDTTP5
K9oSbchuHUdK6yqHJ3WSMDgpXHklIXqG0B+dKoAFZDzlFBBw9DYvd7Z8uPAxGiOrcipdrToRVkxb
xLa1TdqtfUIjEoZVJSbmcDCMOjE6VFpa0C6PXaFRL9wdoOqlHflOOxIB7+nglkJNCPtKZLhnSPPz
CWJBwXNQvHJJEd4wiB0NgWtkgN5FSn7ERiIYkaSGvnXB6ue9FpY+q7Klmspp2Uueke5isg3+XbUX
bfO6qfMMMU3tNBaBzAm3DoCqBDW5YEo4gW1Z/FghSNemakx6Bs/RR5dCrnxYTncZ1bhwjdDzwSS8
ufadhLeZB8Ri3XJjnihYh8DbiIFCm9DGUdDlIt+5cxfnqnqS4FpxQggswPBibvCnyQtFDg5sxIkf
OswpNMhX2nqCpu/dwFvsbMjuJfoE3nQPHRrz5gx7sw+6g6zQKoVawVQdWwXQjMzQHTzRToXWaABU
xQV/yPlwGPB1K82SKNvZOLyvNUd3kghMZn1zcguVPZgdhY/VQ0K9mRu5h5cBeJxRYuwZf4WzYE0X
iRiN181Ig7sJo75MXDEzQSITRIKmK4Hwj9KMsCAh2mXA2HiwWNd5ivK/FxDDM3AAFbZwWq44qegp
fncaY0eNY47JWYxsUdnBKVnK2ZRdi4xo6fkKWHeajncIpkD/bFrqIBmto910aVkNoVxDoZZ/5bAz
R287YCpQp6lT1FClpg9v2T+eoMDZ/2uD9vzcX5vpTe5podIKiiWL9eADn4n+fnTGwO6Se2BJ1T0z
KI5PsUQnIggeqYatBWBmYAmye3nxTW1TC5veCS3uBzIzcMx2tZhmuY3w4ewdvBZmtUqzRYchedUW
VglNnz4UcQ2OLLSarAiRbFS7+ILBvkr1nKK23k4bGUDIxGOSqVkAA6Iy/pP1zoylEMeysupgCvak
aIB3fZW/t/w4jDK+1UGzXRTbBXLEf8cbDaDYiq3TmWV00r8XgvrXlTyQJsrRCSvWxoIUskKFJlL4
kBnWbRxgNgtNVxxJl00wNKVmWwUDgiBc6+2GLqs9sCqdWcEyRSSNBKRIIJhy26MwnthhKLoSjZJJ
7VJenKr3CBV4oABCc+STy353RWBhx7sI3shU/KTqx+Jtn8xOVPO+lKxvExvD9y39BNUE2ZVIHn8S
rvEwXYl79y+Awc13WOR31HMZ6HOJ8a7EWbo9pEyPfMXnc2nZU6a+wculJuWiUEhL73W8rsNpyIRR
Y1h0eOj+Lwj+sxgfL3WzTg8uQi/G4Vgw70mBlo6tBoaBNtmf9gpDg8ZKRCxmsk7KbknbRlPbfmNn
HwaMwhuw50NWT9CXaNnrseijoL3M6NPHP8B/RElmFPk0gObEvIGTy6TB6K8Jm794MUEhBys5pTyv
7yQSWTwDtgzLY+iCfkSIiu7N0XwP491FFxHN/N26DpmvClpBFay4GkTKi/FklVhnvPPZr+YA1uMU
1fYNIIWr94rAoJwE0+YnawXb44Rm3laSXoXqk78ifMOvTtYltLDjZO9IyOfBIKzXv0fIjEviR7da
ddc8kFY1ZxjeJR601pWr33HX81pFbNXwUKk2WUKDgat3WjXgLgzO6ywKLGYL44dDkO4MV3hogBQw
NNfS3jAwJJ1xNA3/M4F9h/ZBFm76E+DqMDEYdPlCrC41jN/ZWD31GM6ineJHATMDjuYDnkNxhgpW
UzAfhkZ30Ar1fkOuoIt8j8vkrjLRKeW+8IuT3edkEKji7opSvL8ag613w+SOpzSuCxbBwQ6AePP5
gHuzX+3b53fYzmFSGqSggUnNdb5whXwF07eyRfOTmm+zf8HZcI7qxpDMnO7EMiywR2oWuZJYt7O+
G40aIk9Fm899T5i698sW4VCvoxgPYHws+eXynZlUF09621d+7H39yUfUAh53UNaTQBov85Mjt8AZ
/UzuqSZj1NRnneaOxzzmVwEue5AX/wKyD4LkChn+jw+yaU8LjDXnYQJqQ/wmSm80UcCnGYhno/Th
k9iOA4+jmLLedSgYot/Gn3Q8VvV9iUibzYmOA0Et0UsWhOoewEhoaEQH0GxRkMHPjJt/VKqvBqtW
U+khuEDtyHvizfXWppyrQvXYt9mtLxNy9kIq+J/D/3dZPfrcjqifTfGmrqDKLOOtgHGqbH0RqJ4R
/eDNKlzvr18Ls9kaJxPhGuDV3Nt70+4Ll7MneKT1ngWdiqdvTIySmudE+R4VbVP1DjNAhGX0Pk7S
njZ1LeX9KKD3jroaN5/PprPu+HajlJHZSbjjIsewcneb4NoZJ2v++iNNJUPokwUguF3yCYo21BRk
iENfz+VaTSseAAexVQLz0FPkNlInwoFuhTQ24GGbyGnwjGtKg/dBIP5hqO+KAZQ2TgSn50W401bX
Mwojq8HNoEUz1F/NpmIL6w+X+RBo1ZKfG5w/c5FBO9ml0etAeKTpdQB9wwIqNCehqsMtZyP7yM6b
Zt7wmyvQlfBkV4XpcMi3JO4hOVzPdxs6RqvQdWMekbVsBBqg/16wFeV6jrfH1NcF9n/BDr8nz0hm
CrFCUjjSIZ8+HtqSGJqvYim44J2yOhwmGXPpQjLB8xQ+Yl7RZNzniUF7lWDR6l0xFT6ZsdDapIvK
7CjcS3fAYhFONpI3Or1zA6aXOoQrWHsQl/EvXfy007THYnPRkVwyuUW3RNd2nBmLebqBnbLRVGvH
H9QOVqsxPa61X9CZB0hr+uCOkecH7XpmyYxxAiB2676TNrDzptGkKPBZkGrlq1km9bRD0iEbNOpu
DPseUU4Lt6MIWygXKXCaK5iDgrNUlTmd0NBwGkaLn+IB2PX1vALIcUgv4GLOHFALo3JjdBCNUdvd
TnwA/0L89sD0l9p8mMuIQ2dbkf48giufzd9PGSgQP41yw3jTP6yVxMlRN4JDE6zp7SqzB9FdzVUs
LppRbC6tJhIEkmxl5HjY+MHVJPP5WTFQim5Dmh3BY2+yMs/z1YfpormEWBuaHrtln+5lRlASXe30
MLpcB3C6Pvw59bKjPCHH9ctbZEyYwUaQYU9a/Ey3c8q2OPQdq15NLXkzbhRvI6TwNggeAAx99PqY
zIRWts2/EZR1W3DXrZT568CHLgktM67+o8cIDAvp51rZcJ+TfoLNyLNIN8KsnmCUWtiaVo798eIQ
s+eG+GkFllKdAOdz5oxjpADWk20uLo+cyKvJJDFWVxGmXzgOjEV2ZIb8wXl61S6GXD2DeJdp3QNa
sA13p42hpvYS4HDTwSCc1P6C2UpPEViw6db5JU2HdEDtbXxGFq8iKcdKEln1iYL1Z4+7A37D+Rkj
KostxJMAB0lwBW2mqf7vsH0vU15KtBhHP5HoxiekDvW3sk72PxzuFZurqJ7fnDrAhtFo+HcSP8pB
UpGKg3u+jRWRulBJH627sobbn8W3ATOjOmotxDflI2L5XmZwnb3CJLPJHa0Y68ZPQ7jfvOd9Q4eY
Wee3juKtIIO5zTdaa8lBGt+RCXrna3NHGJ+Ew8mA5IEhrXib96EX83OFvdaxvtUYXPlHZzVWigh0
K6bhvyFy1wVH3fIMHtvksKWThu8ffLh0lcsExQBGYzb/WHdd+gTGW/EO7g8lnTemYI/4te3xJ4B5
PtUROeKhfRRhS48BLhEf0HziLWDTwJ2BgKG14czPK1nSAg0nQUST/hXBvJr5hcT9YQqKehOEhrwz
YOoR7OW3eCsSPOB97+0ax0d0WfijxXK8NWQHcjHS8WkHocq29mflGYQv4jqFssDLkdt+XYUidqIq
TLKG9/zUSPoDHkX+JUMv+JgiueIFwSCqwsd0aKehMn3ltWy7o1C5R4JGkehQzcBJkrEZmFySlgrq
j7fqysHYYRPyttKacrvt1FYVFioW91WWVjAKpL082cgBk4dhOUdU9OVekP6kg1n2RmxKCXmatX1+
CCgp51DNFwERqkiBwZGUjx/3mLkE+jEMLyx+ypa6CA0q5N35hOO6HovnH5w15B5xi6l/vt9zze+i
8KHTViSK8DZuo0rXCF+Ed9jL8RTQUAr/MAQL2q1HVS9GhpuVFS8Z6y86VpsIWtp32yzlbc4FTxDi
u28+1kVMRjWKxjn43hkJdZNNdlcjBZ3s1FGfdd+hmzLOyQKA5QymAtx0oq/yEmLOPfTezc/YszVt
3uwaTe6LWU1KHkzRPGHekK3XuhfdJuG7QVhX7fWjZDehpEjG2IDHwaFjkr3r43hEJbjyz1Z9qnjv
0FSJgBEQPtwZxR3xp5asBDhODH3JJPuYEir3H7UPDv0aAzDwit8RxhB8owF20QLhhGfFCtUSZdAd
wVMQmw5ChylT+s6d97xbeKcXbqLuyrHOt/vCUFOKO/BGo0UtMkCi7Y81tTDYjq29xa7gXdt3g+UN
W9FERbIASsY2vwQOnJdbr49phxyEdVsvLrJynqwRJsscRlOU55UXKWzaNiiqxKXUlYQaFLtEZ44B
uU+1nvgxKrsa8blMS2M05vzJakaAaG9jgF8Tjka6glW3jQd79K0KdLkwqR49iaSkG6LJv+FDt0Ja
E/gPmMlgFjuFQN9y1UJTATN1RAJCBTM8lTRWA9pHsbuW3sqci9D+m7lCEpcQGAib00+9Wxm2fIpK
PvlyoBcvkwzlfooeSKAU9hqrwyjcFPAaLd4oN4l4cp0zgzpl8JYF0vTB1iqZX16PGJiPESV/geTD
af2q1YN6ZgxQMk8DEgXwGTlaRkveiZblSV2PcaZodXSVZbge+cMNsqzPB5BF/XOG+5NvGxdBmkaI
o63fZIM0S0ioVMkjZdbT28i6IaMIAcd05kWJV/JPiFrCHQHQx2hc/IYlXymmbFTi4Sn95OWQQe12
TzxrM6FIBiU/5F+nsTxT+4/I4cMqcKURLHRQyjuOnst5lK8IMv90gaQ0jU4xQA3DCUYPeAwzQD5C
PVpjauCuMuOu9YyaymA/0j2TalGVptwz/kYH9qWoyCXaWAHgIGFDumGvJ/TqNtt016OmCABXgbva
WaHdkKhu7Q+WOoSMRGiQfAJTzgpZUKjIMll1JaJtshNmoFcyN/H//RGgKL5OdqVlT2xHxECoDHYx
H4LnDr7ITPjKdF8qX3rElEa5e3+mB+ow/OOmpj8b/eZHawtE9uS+mqY7SzYSfRKB/qjz3kgGtg/H
9JCCwPg5hUOHJULkxM1kh7u7Ab3m/NXJBG530Sf5Krx6lJp1AV5qakraNKq0xb40clJxPLiviPzh
4tQZwjwMby406+cf3v0YYZUFiMeMIbU5Sso7ga429tc/hCU26XKPDRxmyPztZxygayHfjfXhU+Zj
UFr5ocjKqFLA9uMzfj595U66qrJRx/hxvjkha1/XLSsHWaHCQ0GcpdpTl5EbxJA0hexCAw6BIDVv
wW9V+Iggh2p696m0rcVElQle5fmNUVr5257PepAjacC0z54MLnligeobYhcws3iSudwnbOmeaHuR
vF1F5UErMymNdGtBDskd7Lvq92sBg/iDBPfjyN+WcEau6QjkLJbTIZ4zeErziM5kG6qY85Tb9Nr2
QcwVlMbAg7vfL67IST82/Ky2XJa/tMoqC1vVL9zOpoO0o/8TVKwZg+GR5o3oIIru/TyJR/ucEgS5
Vl97nzZiYpnylKkYUvMytNGWuC7PTRgF9AJ2qSyE/J4xxQRmj6e4naUhMxw834vm4OhEKqEeTNlo
6fR+2gIimNRArXC5i/sUoYR7kOp1Gr251UUPquSXM55DjDunKjgikfXLmB8DizY3iK5cRwGzqj+U
T+GG0OrgbcvgskEBfADx7MCm+ickt843ZrENqXjH8jJ9FFUnlEzUTRV/eZvGCVPDu9u/2/4sUV5v
284052lya4pfpo89joEpI9rslNCHo72YJNjkimgczCUL+pey27qiGiZeP8VXYh9FgIHY65ntrSBI
t9zD8vovXyxOqiMF9h3Uu5IJdb2WkcPJcVAE4gSG0MJtQc5VqrOCw11mV3FmGOMlmtNCjphf49wZ
i/0L9BytuHqDDKSoBjIuzeCFRHyKvTrdQlb9BEgwkASnhUzJm/EBsdzdz+PoIr3riMMOHpm3VUsf
B6+S0GVKJ9nrIGs15pisinhnf6UahMWIOdEL3d2fPOUdGLj8SvHwLvABhqN/SpRCQMdCk5fAfsoE
dGfrEqsZmnDYg07P4Xl6G8MuUCeR80eHTAwxRMBRgDS3oHmXwpzNfFqWbnG55I3k6fhTrIf9dISe
uKdzkQuRAxSqrhVLg1qNxcDXB1VJKU2uDjd2EpFugqI5rRVeK5nThda6NR+TFQwqxt7Hm20+jSh1
VWWyLPe81liiAfAN5VoDVWWRMjrIG04I3Mn32RTL6J2xJOJhNafdeoLDL6+QKO92DmPQF8ky7iCT
w28LpyLX1WEpCH8gfqTceZd/GjLiapqg8yMdMMTzY/rBz7J36aGZu1uGr1wsIgBIEiwuvLaudF95
XBGrvQhJPrI95Rp3ibCWNgnCORZhvHO9xjtk2blvnFRN8tnTP0pKwBgWCsKVvNV5WDuk9Lgx/8fP
jEUrNt+FtEfB417ja4QJ0sGjJ40LFc/P/S/DlX5cL0XlkW0tn/vHX6myQC/8BOJ3mhV7aSjILBMz
JPr8/oYHS5NtV67hi0oOS7NVk/z4cX3YJ13dbMigV58OtOUMQGykfWlL+0KD+Uqu9XazRI3+j2pt
3yZKoBqqWdPShIFD5R3aO7I36WsqLm4jnFHiWs/SXGchBOCa001/VQ20sM/O2/3ngmwLgwZv9P5R
JjF2tejb5ceU5kcfoUW2/lnLMlJvr83UmkJrfYyNrczR5H9KQv6cy0JD3eZ0r6L57V1ya7uNJAgw
DrJk3x6Ey9eUf4pyCqRmqnDLcQksrBOvlHW6fz5pN4huTNzeUo8kd9RD66oSxWbh9HC6uJjIn/Dr
y5OHnC6FVo6FZb3JkbJGOJI9yIlpD6wuFaKqxrAuvgWo2jt18mqTy3DhnciOCJQqBNX57aInd9ns
8VUwrWyKqFWllSnLT/wfFQ6hSqsCowoeBMzKLhGdFP+nSxCaBVs8VpqkHeHEr+R5JEwWqnj/GH/0
psN0M+22ppv2aqtBxAqJutSMK4Co7pDspuq15UXFQufSugM/rJ3Jpuo8JIs42l10uH0b7cbiOcRk
ADF479fqUKgtncOyFMbR+gs5K+MsCSt51wB0T5BSvCl1wza34JANgGZvn/YFOZKNCv7YdJiadvNy
XY08pEKkMfgQ1PComNdqWtNo5ZczDtLmJd1fk4IsAeSAIxFjKSj+1d5Pg16JhV7Nc4ckKV1wcvIv
sF8xEfFjNp6SwR4EuXHPdwQqhlJ9rfZajuHQ+hWpqTuQcvTvHui491pS8xG0xMFY7BDOSCj6FdNy
cNn758vWvmmSc26TNB5IZMmsKgK9F6gv4T4x6+7F5GQOjaIdR6YjHdLXMNo4r0N+pp1JEa++BJgj
DSkDkxufMVRNyCwzgW4bFAOO4pCIKces1KPMDsZxHZPA5OOk/g4QQZZvIt6Q9G6sEjqh6J/fmdZI
tTK/7hHDhtNl3m5xsQJAG8v7quBXyk9fVJ5JXyCi2u6U1vhThQT8MbRv9s3M49VYP7fZXuVXe9ZJ
EnVOjpMBdKIkClUP5oVmFmQgnYz3c21lgcytemnM9E0Ad58G2rQ8VSGkXGSgPFKacBpWz+dvL+Iv
6Ufm2M2wiIlNfpRr/lFGMPOUfRKhnPd9PBmxPt4XRAIm0YTyPY0mGdv4UxjpQa+SGmHW4/fmj5fk
a1xvLwcJJljSGYO1dZWjx1e9RU5C1b7DsVXxG8ozXY6oEPD2yMQWjGSwt0n9QPGJiCAkADoIFJeq
GK2tbHIYg4wbWa91s7YCebwdhvEm90eWCktjTj+HS6H/cIF2/kbPPLFf5XguL4f58LcsrKP8osdh
cxzGIp/yiUi0OFE5NPd1eu5BEKz5rjT04pqZf2WSQiXeMMRx6YWd5MWoCtlZB1qc6G8crs2EpACd
VwR5sVQRw3gTV9I2+7wzCDRkrIOxfbMyynbszwDUwS6t4FoQTXn3qRwOz6e8I2cxLJrHkqnek2YG
d6lmNPg/J1dnj0HZ4hBiOfqw2JbrPii3UmKdUVIeLalR4vMN5gSx6LGAswDoTuGnOhquIo0Z9Qhj
YWidwldzPL7WZPeqggHYLprAfqBdQb+xKrYl8AXgmOxB3eV1fRjCE3aalIVPEEhFQ7lfQnWbi5/C
AymkAso+TsIB7YgZWFpiIi09r6LwbvdNba7OaKHjsTYlhP8yfiCqXkq4139tA918/CWH3sFEto0p
p/DT2ylkF3mRRB2OKIkcixYVtMe+4MH7PYCaIJh/HJJaXlddrMontPlPSaoNmhoudb/gq2LYPZdL
dMwUMR/K0OE1IVjtTPAMoV+POiT5yb9wjBpxCPofR5O2f/L313RGZ/u3yyNlty3Copp/32k0g3++
pOnGVevCXMl5Ua3d9pvaRKzsVw99JUB6D4b9a7KE014YdmxHhWahNAd95aAwXZ4UYzf1K2GWrjxC
o+wf94xTVwhPedeE2+b2I7dFbRBdYCAf2cnaRaRJ7hONCPnUgE4oN/5JQrfM1yE+Hag75Znjebve
qmSUReqTLt1mH++1AoGAuQrdn1lZyQITfxMw5bJqoXJwFc9yo1nB9SrKgzs309gKMPBZ9n+nIgxY
dMcNE3rNz0yq3/Rp5d3xskSUcr2vr2KtJkIG+XlXivX9CdvlPlhnJQk2PySrPt4LyYi289qfZ8L1
elKfAo5KRNRzCJmLCYp6UqT5gtEnR36LmRIjboeTDvpvdSlNHptDTH8fnNSwNLl39Zc1STaKkm73
DkQtAa8YNkZO4edK00TFyey2veeQrUbVkochTavZP7xvdTdjSQr9cu6Y8IzHzoxzlDngopDn9pkc
UrFp7nvHVG7f69lPekhB2ygJBeJz0RW1oTOjcfFO4gE11INLSVkDwF6nvR4OYAZ0fEjo+FLyXQjp
mFPE7UrQH6KpQ6QMKM6rfsjdY9d0hnLlHwNKPw5GxVblUPBee4/zCpQ2AYPAdmpYzZC4CkZhak50
kLS94rjB7d3zX7ZL7MPIUfR6rrqvLOghbflWLrdqEB7rSbq4dh3c9tFIO+O5QB/3AJAGW16PJVQW
AkCurP4/UC/XVrb1tXQooTuxDG3ciuoaZiZKV/ltITzNMIBbUsbGMwMaz/zKE89p6d5kcyWtND0k
8j61XDxX6EW9PNb5Jje7+J+JaxWQeDeL/r+iRmah3t/ZuJjT8oOaB444ZDgCTzXnOzcpq+4Ky8Of
obuu2i9HihjV8SgbPcVR992PZfw4M6UdCR493x7wTik3aQuEQ5MLWqnO401gVrMjA3J9onAmezHk
mYyrpFX5JcEoXd7pDGhF3nYTmw7lsa9uEkXgaqycHbIv4MWBaOi4iGEk3AuirXboKqyyxIBc4yET
pdDZApipg9FjaSY6xGcdpFcp12lwMZFi3SiqeaSsJh2ap/PPHzAcBYxvVKn+Cvf9I2oHMWLHPyF0
PwDvHmvRQE9rH+0Y7jX92MS1tLS3W0nUbUtl96qTbyG+MOv5/EYQ39xra9ZYEGStuj6UPLZlVh9X
kXkh5X5fvjOj37ZNMaX3Xj9sCbBbMCJ1dBq9zTc9pSaMcLRxWnM4WuUgDjvpqAMvOzn+vj0csrx5
u1tvVudGrkBlXhR0+s++cHl7FKK0aBpSt6vKpqO4KgdlN4vJyVLEjdiueI9ZJOsg8b1ap+QtmS5D
PJQiRzF6fdP0TU2h7K1yTdeuiG72a17KlqasxwGUvbH7h8ix0EpNM+J7cUJVdzMQ9dDCdnlGc+rZ
WkP3juLfd0k73ZpieaHIiSS5gQwqPwsQI8N1Rz7i4/uciAPv3RxILkISClm9rPKbnkRMLoKYQf0H
cCYN7aVXc8BNZBHsXW4Ytx/DYyJ0h2n3mXk4A/5VXgOa+SSnLYSGyOhZqC3kisFKBFEcqKBC9JFo
Zj9w80UefzcBW5qSr12Xp/cCH1UQFdysjQyvhpni0vEg4S6EGP8W8/k5eAaHWRxkxgAag5JmJZz6
2FZa67FgAH9uPlykiUqjri0w9muzaUCRq/nKJAXYD33dma3VlPgRy1c5f+Hah0he0wHfYuPNebi6
vymH23tdEreAlir1T5OBTMSyVoqmhzF3wQVAeJqFejqLWWDnFiA5xiD2J9aQ5l+9v0i9fw6qGd1s
uRCNF1/4EKDgMBUTcRl4CGxpAKK8bxQv+WHEZIxKUZgS32K77/hm3hGqOlKF0hizeNZCkiZ27EkA
fOG/+FmHT3keT8xhc4x8jvl4g4iTJi3QH+1ax8Gvpi5pLqNyR3G+lfG7idNqXTGVUUy5OFKN6uy4
s0cHHJ0R8bMfRIy1L/uK2RSDQtma1j5A/2+ioZmkGHUMuvYrxYZR4jcVfQZ7Ki4ObDw/n88FKymL
fkR8gi9ZIICXEhDIyUNtv9J6UCu8yFGA/hozaYLzwZpGL50wPQD+dsfReqlJYlpdkslDbAFStV5u
Nn9rHKVsLBi7ZavCKdbFVsOf6sW1LR9g57TFq472wBGbzq3sc8HXij0HOA5R6bUC81wCYu8tC1lI
78RqQh0zYHNRw/9bBIJ7K8PEhiDYvumK/WAV/0Kl454riaHenG6SG1WXtucR9yTAI4DQ1uFyz1cf
DjNpoBvfyyiQwCjezrep+FHdp/f2RYjKOQd+j7EmKMukWIjHFrfl5+pQQ7hBIctGEHfx5VXu+nVx
h+wPROxGYsdDBD2QYbNeo5G7wcAJ9b+Q8OGf3kGUeyHSe8FZQSeWDsNcV4AbQ07S10AL/QVlzP/W
lk2kM0WPxSkvhfqdhKy4sMV0HZkptnqZI1GQE91orVAt+dVFpZVn68RoGHZiSZlvvapUpwkjri0Q
7E5qRaJYj6bWJ08pokJLji5i7yd/JlX7Ofjj6UkH9Xgmu6Lqt8mggvwKJpaWULwcSs5/Ytgb4Iak
a7ERZlzcigizzDlwjmK2Xbm1ulY+QNWRpbUECtQ+FchO8ynTx6gw1olkrDqHzlKGOhKZgdijj9Xa
6NOz7tbCyBqnaaJLg+URBrMWsbE6+YrgV5nVlB1oea+QTiBH0F3eAX5OcRp/fJvo7OhVclAiXA7D
T4FoGO7W8+WruMG0eor5WPDmUbqmS4ZwU4oRCeztPQNiTLLH19rb8Ag/si1S95np4904LwHJO4za
QC3+n7Lot3OGKL1VY84TLMOmGeFCfP7z6rT6Q3/Vt9D13FiUEQJ9g7DTPe0n2PuzRDOoLsZ764v6
pNmSc7jbm3IgbRuPTaeWPaq8SUSyXlzGAsFUIeyoIIzGVW6du2IuA6goocvHLKqQh7rQqmx2t6g3
GjL4Lv393BGQuKXOwiOyUywa89YnVlN9YXR5lRGqDgHTLI77Utl9vgCRugywu+Z9ZTc4E86muTWH
c50qaQ94Lwjt+ORtJ144CnOwLjUashMXUJUBrxyOSrbfUBBruW49gJ//hXNw7S5KqMbE9qf23/gF
1n+r4MTqR3FQ/TuAOi0aX0Eh7HnVu+t3CBGhwxuUD/WbKXedLYWUfObE5Nak989eeyo+4Y1QF5/B
LFwPE/W1+7iHovCEtygqcmzZnevB241sHvtArUtlYqoZOAf4QNNXH0aQrrla9xW65P2J0fIDiPGi
ILFfzTNU/rKvnSdKRI/FwcV+ruQm0LJMzB3WPH6/u+K3B5pUZGNQX2g7yqZeLhCjxF/QDh4kyc07
GZgRjW0mQquf/ASq21a8tjRorYk58Vgj+UpsF154nnizs+axpXML0IXO/5FdUEEnrPazzURSyNZe
FF++oBH3dsUa2+E3BR5WdjRyaFp4R/vcvP7+PqR/JxuAzJ3ZEO3S+px0fMj5iPJWp/zbjrDS898I
AEiatoo2OOxWOp6my0UHLKOGgDMpTiVH/hNxvGu6A86IkWXvqDod+lH7gipSRoW2VmXSSfx0z49W
V2VieGkcc+esF7px5Bkd31W1YXGiKTALFAfew7RhP0PjjPaD5OFdqiMeIIC8xJtXEK9WBvfeodTc
ToCYHr0GdsrF8XDQQw1hu/Gg8/dCShDEbgfIJ+gIcJPUP93bfttYy1jX0ENdLFdWZW0HTmJMxcK5
5yXT9O0c0i2LSrXERXm2B3DEjEkSMc4xBQjutkqHyOeO7P8E7J6PbLMr4RnWkaIJ1SV8D3jbvgsk
ispS7m9T3TCCwhNAMhFLzQKh8R6n+CK2TD3ifaHULBjxuyt56F+LzV1jMxxX6gDNDFCf+Ocbz9ew
ht9oMiSejxxizOxRDpNm5OFZQAZCLOUiP3SlZ36CSr1zHOQQsWfHsQbNgoQng2sHslcLdYoNjz4m
C51MtTZzoUjZwp3Gxx0PyDUM5w/BpKEHQyee0xVxXcBqlgE7+/QlDuTU+PoHl6O9g3VRWzSoLGD4
B+LfnePVqDThT4dmIzYdS6LKvbpLgVkBVV5C6dM3FRG0uYYE9qt7D7hQOx1CUt3GYttzupodrrzr
C5Ao19qd7x7AFirjyVbFmWe3F7KQoqQqsFpB7gthS4ixZpsJ+81Cjr3zaRVU7nZkRj0AM1PZJVyV
6BGZYbdMbK5jnkNURja3AH9WJdOnPEwJrEZkz+XNGYOK910ewxM1Q+9Na0NNOtXhLCneuEjgBeo6
fNzs1LQp/3dlBzBC10uqWwWUNz4br+15/TfXN9FQsRogWp3x2b10zx594X/JGlOW2ujT6kohZjvt
nqWAT38f3q9inryb9J+GPzo2jW4aBhjjkaC+1oNVjmgA9dEIo9YXLpdnLe1D4Xn/J42059r7/e6J
Yc1FScMRw6OMXkSFj/P8V/jVe0chYOIuQqCK3/i3xqHhTHw0p4xoN9mS12LehVLCJkPHLEeyJT4A
Orci6PukLc66CFFHkfw7CclRF7O4yBgSjJdL5gdlSNR6SRSu59v1BLFM7pIHh5JsFXWQnVVVw3Qa
JEEuHKazXJsaPHZdCHwqjlflfdPWzvxvtvjuB2b6eYeMTCmonbPqavrCc4kfrwIdJ/1hJFilQ4JZ
/QiCusYZTw3KdQvUvonbwtK0oM/163+YXKMOyYplvK8V34/2mA0WTVWNeXfUxSw4tFg/O9WAUYc9
d4CNIs77uq1QwCcrwQ6T+ybUAqQ9z1n+mUsQJLiEdt7rCys/W6eXf2k5DbiMLV0/aBxWVvBW/KkG
CuhHeCYdF5oR1n622tgufU5doRlqbhI8tAxDFMLFDGMemwDT9my2OAR/U5EEZcHIdvYcP6CGJ1CO
DQYWNsgr3GczUaSvFWSALLm80vxKIzMkMeH2WF7w8oIWV+zBxrw1oH1XrL28prrWYevjJU7EVqLv
JKLh/IskiYxQQgRkZ9APmAd/u39y+bjAAFLjv1XaPewyw1LDn5acw3HlwBeaZ/n2rpKmE1TLDUIz
ZT6ZimCFwz/6Jk/cy5U6EdJ+KR29ooPv85y9kbnf9zyYXll0G/fIuXv9t/BkeiP0Y9OoWyt8uxj4
7DH6FCbLWmPJMhhi2Qn0tyZdF4RVTgBX41tQwLA3EXig6dOzhYFVk9ODRGZXyu0vp5fYNDf0a5ve
+6eRVThxyQ1NCb3He/loj1z6HEQy8SgPAdHyxd2kkZuQ5slr4d4FCSirvH7+mg4gTQVFvZ7SDy4i
sJ5WEqJuulNdBiBlNdYyKfEyMs6kbhUjzHBHmFc5kgdbUR2at1+DC1s9KVDYOFF3Gi6JLXvi79zM
Xi3Ow8eYaEG7tzOEdgsnEoLncInE8UiAyjP/fnOFQupvSRCo9UMpfwrUad3+UGtvwJa0XHq8EKuU
UUyKRA7DR8U3aBPOm20tCORziV4gb/2FHch1riHUnvi3ZmK3QR93yeBvD5MyfeL8KRNk+7K4SoXi
H/TtMuJkZ8XN07fLb8GXADUHK1zjU+RRWiJw/FXQMJkDFtZbchQ9myP8LgLYsK6jRdoMKgutDNw6
3CvEq0+ldWiF0GqwXAyBebsY6koMZaqajegVjayO9QDLl1Z8qGtqafPLztN7sK0INr/RR2Zh8wh6
UH1Uzjq5MQifiJ1v3D/nZ4/KQkp6fSaoc9sSPXN7p0XJY4lcyuYlsRbnX5jucrMS841wDK17tJ+S
NreM2vahnSpg+bxqfCfdcjDO30cbJTUEEN7A1Z/ogH4bw0l86XgWsDcJ+6DiU+mCd33j7hXBe0jR
YpHPDk0MsQ0Jitb8wfDcuOBW6j82kuwJr+1RfWhOL2inVRnZDqkS70zwhUnwV6sy+ET+tAmeyTB6
E7h73gIy0z8ZcDNX8Rul/Rd25k+LK6H6vZe/J2MhhuYgGyIdSZ8I8FqNdtFsukrcdEB0rKVvYh4N
NgotXuQ8b2RfIg3fiZhM9+JX27C93w/AHfIIQ5IG6dCR0qcYx/gu60tXcI+QnXtP/b3+qvlRtrKp
3PMPHLPWg32Pe5ouVtLKQug+Xo4mOfDLE1X2D+V+S0uoIRgF/a7lBBzuYJpY5zGXv+9nu0/V8Wtk
gQgI3BFD7HPBB24CGUq0IavqBdTXQZnYfoNcTgb0CRehs8RKLIjXtQEyJ0em/y8zz9Ln5IttX3Qj
qie0wP37H9HTMNTuafgaPpHrHL22qUdMz7opf4nMGeLTaKLE6VoQaCUA1mWv5RI12AxObGwTkll+
jQLQlfV25gzHnb+JUa+VxsSC3Mumc1979SCyT6IhJMB2avTI1omQnJE0egunXL1ydvndpRinyOQV
LEK7/XfwjBKSPlt9JbnIWwQtcP573YQP6Ho+8Vac4/gKwRMDSx2b5cXuP0pM/jvPFEqeO1bC5kAk
aV+IKFIAWwq2ini8muvkU3gt+1pyVQgXPD+HQNaa4L3bKQ6BttFcrl1oVbIOUGmD6FNcxmP1xVCN
+hJXDId1zPthucyfQD9+LX9sgUYtXVGUDkLdXXaFMYmveX0f9CVnxQ+AxLmUrqhruuraqKERdLgS
BBeDswkG3dEkIfupZjnsic5SBbMdny+mqzTmU/0I5a/m/p6uWZtLeNS5XJn08F/Sy47USt2GurnM
YnvFca0NR3TUA8Blx03lDXQZelp6lGpWRhkxOBw/9cFsgvYi7MgTj7S97GHYZ4o1hFq/euSCrFqb
V/o39iol1o7NFWxn1oxlAot2Je6Pdn3GokZibXVki+hj9mZjM6zt4yzixZu+1bgJU3fKb46FHipW
nzAMJoEDimC4+vIz9UJTUq2GQe8FMbKN1NYFU6qbAAOtL20cVGJlT8reQoDaUt71Ft1XCo7XVe8B
zOW+YQwJjfObNX2ifmrNxYOkW+ablhRx0q4FMU/6J1nIxJJjJE70nlCh+VtGvWGDeJfKQE/FCdDL
0q8uC8IXPCaRoJ4po5pDTXYN0dhsNyWUkirbcuvF8PM8at2xubUAVph1Ull2zMV8qn+6zVV57cQd
CFKgP2m0XOJ12vknjmbYBLFNXt3UKPC0Q/fKV7p5Dq75Jx/McUUce6m5nhUt9p7eaFFUyU62RXk5
KAHu0NXFFZyxhQtlZyheu1NmAba5nT7JKLBI4PgP7oC/rM9dv+PJjp/lfK4GFGRrFfn/GtNceWYp
3f/vxPbZAcW8rPbXoJyGi6l6d1QDZjTZXu9B8WTZui4rleiA67X0SfYGHwj7Q45PKaTLPmB0KMAn
wO/JQIKfHmaRSbOur+ya9Hj7Erf7ZwvLaDAypQa/Ule+y8JDM8Z8P0REYZSy4l7QoSNT9DtLHj8D
BSxFLWzhz42KMs7NafvuZfDcGLPyKh24UKjYRiou42ueY1vxQno6O6gV3MxqG0EqAAfW1VyYTuAX
3cJVLAFexOTMtx4++6C1e2c3CK82lHMOx99JR8+8Wl2Cu4nT/d7ojOi4WeARUFxpIBbdkGkUp81e
avd914/0HfuoSwlXr+UiCLWmdlSZzXL2btVpv8FYQK6EKcR70e/Q4zieGt8IMDOc3D2pnSnUKrmi
c7esUtZ6VElLxGEizOaAL1KnkpLroA+uXwbo3P5HY5bZpE1gpUtwuhDf7uxJ+OterE2rC7NCwqQg
pcd/pTYTW68KbrBxGkEqG+opJau27M3BCV2AkmSlwN/LyGtAjra2OtdySy+P0EutYD1diKa1xl/e
2acHItb2W5IFfVQv24dvBLRGHNIiDLvEnsb5PpSCpYD5/5nddpjig5huElRa7OF1yHLslfwNnKJS
8vB8mQ5xhH0wdbAVO0CTuZWgss6hHj67+IQrRlACkRBXuwjTw1aXYZdpLGvDdrwL7LenMRLWIyQg
Rzy56GPedJc6i+1DlIXQvom5M3Nl/oSEUWZhx7yL9+KDKeopvw+8TBGOUGElouowCyoIA7rq8kre
l75er6CV1zSGZy8zN4eft/ukMznk3/DmFFVNG78lwiUJq10f7VYKq2A/eyeJ4aGQ94s+Rx6nBoMr
9eE/+Qx8KcDdVvYRdrYk9W6VmUI9SDnxU1dPHHk87hYqOoOtUpoxnpZZxK0Nzh0btJNxvlA8SrcR
l3a38tU+snHlO4hEjrVb3vCIzouw0ZtAm3ufutAS6Kh93dYJY4opG8RvX6Q8hNLdMeqdPX8V2hSc
74B/oMALtmTx1efZaBtuqLA6LNSN5WR/nNRst+hHGuV8iBSRzU11rc8RobV+/SSPIM3V09NhiCiK
GHoCJPFhkpZfSbAyYOYqCNNzsag3PwPLiLsVqjHA6KrXIZWoSH/l/ABHmK3vp72VD72hNsykB4S2
yMjF3wT9CzzLzqx/LILV1vze5eNhcTiuPFMStmxwAaVT8oRqcqYNfRWjC4lFmZt0Y+z8D08PD1xH
9CL92axuKO8jQM7wXwWLN1mZw2prbAC4318KLgCzc63MtJEmDtCgXHR2IMDdOTUM50XLrfmD/nC2
X4NYXWo6re6yzA50iy9XjyXuzdIhDVwZjx0L+jJByqnmbP99yeGbCfOZQ70oJVE6lpx97f0ch0Rp
/B2bz9rj00DWOV44H6rztYAW1gAOKiJlPPFt1BXa2RXT+G/HymoAlZFZz/btfk8M9HbVe5pLbQQb
vD2DxRI+QVQH7pgxIVVI5t7aSDznsQWBov0ddOa10g3kqWOPwGiP9xD5HcE4amv6DFOX4dVWdaFO
fPoSq84tEFdYlkFxXgsaAaV8gF9dwcoVL3Dn3zXrdMxVEi/pcklILgUTZsB/BKGdOvgT8KMkkoE7
R80xb2bowDiwHUp77rPyxEby1TnZVIqQeZqYHaUpX/p/5qZT37NqsF2YV7mI+gVRm6L5Zf3JF1wo
H9SPqVKu7Y33KqgXNdxe0N/6XJiu40BBpE7gU1qLFEsY64JxtlLC3kJRYWy0nsh5+yISCBeMBT1Z
JzzvybmH8N3gWi90Gq5ZOo4WL0ZsOj9AvWs5m06Hp2TK0qqNT/3znoEQdO+fsF2Y/DWnl7IlkWtU
PIQQiu1fsu0sbCs5fPsala+Ie0doBNguAuUMV3P8ZGH0d7QVNEVPvYHUoVXP+UrW4UmeDETbIyyM
su7/02UsT2adAtwm6wF2foBiqRNPmLEA6sSY6kDrExqeH9ciEycaO0oT3tAF8tKUirFJSyugJ/+p
a2sYpVvhiXKkb96wj7+K7PSkj6EoDPEtgHrqVymDiXaG+/5ABCm5OIxUnc/ToZz3Y97yMjzcEc5p
CrX4pakxdHFNju6SjUmf+D8yqV7CDD2yoDNtmclWWxSFoFponv4rTIixl2EmeAkICgTPFUJ0GLQw
Ys2Sdusi0IQHA6NAz0chIQr6DcGzl3TZfrd/skBT9vQuN5Tl3+dMMWadKmOPNOjvgbWVzSQystKE
6iyd9Rqz/eOF4ZLrNFSLqImblorARG/pi5uTyeAXFQKL6sWXaTpHqW4om3F8QH05juR6ybd5GAel
cRQ+IToUAtFodmPe02lIyyYXfzZ45Di/tZdwfeBFgVvpxsgwO107C1EPx33bpQIRFylNmcquiJu+
LsVJAcL7oeQFBqEt6EPoHyNher5+alhO6UrGbF/ikDINOCD1X3wUK366Zu+8NkuDVNsM6nSG9oux
stQGB94QNpJb1a/dygwFjxNl+t4QSWfWrynvwfRDboeg/Az9PLDxY/0yUC2CNLq8wRTcQtQi+Bkv
ZuUFDJv13R61OzRM3XXSJePTaXRSeHRr6QpLGSLwmFF5SuJgrx85sLvuJQiq+cAnA89FPEIebygy
71nXooZ6gyWWnff6dcuuJkKylua/x8QsxjAQamXM/UeUL17CmlS7Yfd3DtiZ1R1hkOaXBwlZyYPL
2mBmpOx8Q5IblT/WYsRm8tnCopmn+YbZn70utHztjfOsZ+1DAtQ5DYGtuNsiOwusQYAJ5Zju/ehR
otcgsbys6xgZabDXI5M2YzYhI0v/fYtV9L2eJgmYsXucomI3xX0qKrQaS8FRSb1uD1NS5+d4GZcB
G+OMMqyaSGqJ1mgz07lmAhxo6wFTFF0DFxN58da61fKSlElqflE//rjPq8DnhrEkE4vFVwdZLOAC
v6bURiNeECVVm2b+Gcae/ZaAVPv9A9VH4naaAYa7gx3Mc4OYsUVjjCl6BNwpQVvuBnMu4HJy24Nn
jmDr5yr020YEPgRe9oAuiaPjhp9GlM449I9RBtSg3EGOWw4hxEBzTtSDNiRORabPdw3rCeBzwNxU
ed9tn8p8fqIl/AksvNCGBIAbia6RldJbzPwWGghWnlpIxs7YiEMz7++unqi8tZeS/dyXujFHdDh7
MtT+sa9JA6O2Wb+HlZwH5Cxkvamm2B15N7YIl06iKTODwVSPtSdVV5ZMAIrYcfh1UVBvVKcWH7dK
tunl8dVBiMPrDYyzm/yStnw+dcPPLfzURH0UlljDiOETUwgRtqhLvm3fU71bCQN6yXecFRR/bx2F
rDK3GarKEuw8E3BFl/RPSmgNxtdmguApFZ4KcY/tcVlu2xLN6rzpvqt2DjWjVu29QrTQzOhZghY8
cRd9s5UFTfmkLjObhtwV3dumgkv2ttAUYp72NiZXISBjW2AgulIP6m5KfC6PBDR9D5eFVp7RE4yj
dQ5RwB7Lo9iumlY9QWSGiaVVApbfxE4VZLfcnbrAdJ0fe+sNpoeW+E6nu3tACZIybDNGudmqQRU/
NuBjCbJcR84KygODOiVD/oSVc+/yrhhtwHwri8IslfHeqycjgBn8uCXAtZLxQncOPopvipx5W4sm
YCD66K+tzo6GhvM8hRSDxMbitbPPV49T/Iu4kNwqBbHhPgJB6NjOh4hyMuv48l7bq1yoVrSchLf1
8c/mdlSGcwtxhnfQ8XZ0KvtluI/cClty7wauZhzg457i913MUDRoQwji27n03sJKEkhYf7uCLFmY
IrVFsXpar9nE4rIqIhuhGjaU8Yhpg6Oo2H8Gn5uCmprGMbjwYJFVTg5M8b7LyQWtWL6LvCYtndh2
RByshdvx3p+bydHrlI+Ggh3uvrfTbyHliAJl3F79eNV29R9tJp8tlY8cWgyT2n8349Fah8CW6x9k
ZsYu5xnDVGg15RjSYVHTwWjLEXxoVFoxi6m8IekrGSeoldBGHHz/+Aw29LMspSDHmb9WpKSp8IDH
VpTxyznG9uFLgM1ZvqwgqAcPK0OzF4dzR72HYa/+uNrMr5Lem0yaA9f0lMGwFHbyyZffwCxPfvRr
31kgmQ0CW9F0oxsx5c2QSbrNwMIAP82HaQhBBl5X8qYa6rI+rWEWJE979e1Buuk0mJb6RXw8RZuM
5gMwEttxOH+GN+U8h8zYFZDGGSepK/EWI9kMhAu3ZagJA1z151WAHt4jJZ+QklEEEbC0rC6vp+3a
JqHE0foug4WdXAGnyz3KQfHiUDxYhOLt7DAjOFtWynPr2c+5C/3NO8GW1JEA3SUUGL9or6xPS041
jtK6H8HWFqdvs0L/T68YUawNgQfardgQfOK3EXchCNXgBWo0tuPetiC0CAAjJs+vwx4juqkcFz7o
Btf96sTpJtyHwoeXjhS0q6TcNTeJ93zx7xAQ554zimeQoI41GMwEmeuCLb5HVK+BqbvRzhD+Fdcc
uZlucw/ajR7amrLuv7KpfYy75dNXTfecc0pLdxxo3W/cfzp4qFqImO7dmglXB0CBuyoTK2ZUr2hh
GX09hCJFWo4cO3AFJq8GP8yzBylfFp2sXlENFhRjtV1acaND2jEfQXrcxD1QOqQrdIiy7RgHXPF2
SD3gxVlFiG161KBu2+BfFeWdJLf80m8uq4nMawGgToksxiCfHAvaleULOX5t0919x1r3xEarja5M
HwR9zOXcwZyt1vZaAfxpK+lTlBE5U2EaE+a0XwLK6YAcI8t8MmYVy1Onqni37G5LS7orJR/hEjK2
llw+5EFl58Pu2tYeA9RSWrbuRoHCfmG4i9zFszMZd2ao7SYDlaNceZtmpLZxBQuWXs5nEShamWNQ
aompOVZb9DY36ZRD45IbdzcmrBJLLekMK5QhnPIhYrAeGsSKfAFSx7Kp7zTg+6E3CETqNrBjgMJK
iFjcOV8YC3ryrFteDUKKBa1/ow6W+7pWaD+Ti48mGzgEJNEQ6vgvgVl+45Yn561I4C4DRIRhsTAU
+XVzZZKJYNEk63vVpNM1AU7TPHK6+JPqia/2K6Yv7V3TyvBChv8MBQDJQdcmDOS7Ks5NtzjA5fyB
vHTEnSpTAoX1Az3mlzSYS1Qhw1+p7+bKR8705GDtG7sy2z+P9632DqAKG6weWKFlsPsDyJE6SpkZ
++t0e5PBh21iKO42U+6NIBSO7DjMyz1aFGfKZ8ijnYbvassqu+a5n8BGMjX+HgSrGwPt+gq21GRE
LTepEK6lw205LE4towu3IuPKxXYsV2hx1zVIKEBytPXyNn/kYvbf5Sj1QGpjm2JQEq6P+9w03+O/
KXA1vNo9Z+fR6AEY8C2Av5WDKCD85jedcGD/0+W2YR0Gaw9eXX+WWuXdWAfUXZbTH7iPLjYfJHxQ
LIdyX5JH8ZqR02pM/zXQsZpQVKck9ku87l2BifVbKnFeO8hKE8a+Jq4++ZZvnVBlq3C7r9PDkFxc
xaafKr/S3ilZ1drM7jZef9+MfQrSDwpBSpHT7ExwaBwcgwEaoHy/y7gt/Wc/n4ZsvfvWMbtY6KS/
/kt0pWs1MWEz+o85e7M9DU/z4/W4NgGg/Dx4cg/rZz/1rh/Nr9xAnTZ4nLIPoY+ST5Ki9eKRopFl
puIaVmJIkBZ8WeetazkpzGujuz1jwY1pkkfnGsIC5fyLJkE9oMgj83//AiFtYaQNY8kPd7VlgmBO
DVi/wLuWmIVh9GpJBiXzm3UwqVj8B3STVn/TE+I0IEuzSP6tGNGSkieO6/WwYELqB5tYeKlAM4Cz
A+DQPC03dTLA+aEXymMCcBWDysXd/Vk3bmImSwMPf315IUJVOShT9TobMiI+hjFX+eTIMNMtGzzn
DKa3ql37zWWX6hGZvQ8cwnlS7DoVwPsktAMVkmTNjXK5G1solN63znZrFgilageCHYw4UZlFmSkJ
YPC77eVqVGQlVmFUjyH5Hascp1APTZUOxVC2x36yi6x623R/jbixlyF8HF98ZMZ3vRDQdmhT25fA
M7zw1/iL/IE6EK5g81AtIylCVe1t5RNZgJ5rWekRynDz1MQ3kVgR6P7khlzXjyDP6abloAJpAaUm
pBwSH9WxG393ZFpLr+95+bUbZTbh8ocj7lGYqU58wJO8U4yWZn7DeYqTEVUgrUZyLa4THjGsMsIH
YbAqIHqTEMzUX+WLjDLYpZDFZTxO3K0YerAQZ2seBz+IGGURB4RD5l2UPbpR4DKvKmwFa6iPuZv0
Quavd2AJePhlubgYtnXBYXSBdVHx5iWkX3MOAyhxtsXTy0E989i6R8QUEHaYUK2nlLaeSTXh35kG
PZU96RDCUdjTsDs9wh7zdZIW+QTNE/KDjQAeKcE0Q/UD8xlb/i2ybHx36kIeWlyT+Rdc9AW0IubZ
Z+D6U16HV/WFU83TxdDAfMnxaqPKKx4/UN8ughux1OFNwM5HVHqcBlNKVxnrtf3OA4iATi1cu+bZ
+DZPa0FL1816OGaRFCn3SLGv9t5Lhv7d0FHf4y7dA0uqXB1DiLiqAQA8wKiX9aJddNpBni8ZARPS
ZnKNLHvwEtchN8zrKjF25TgMXv/bIPblzZRkMAYsPfM1/vCQmQSaVU1lqQsPt7dcO4vFhaREhfA8
5IcZOgTiIYjagZ8O04utZYU8IqbxJnXcBlqxAn+V0lI66YAqta/MaWNMM8u6rD7ifqRcwLidvsx1
lvBf5T0WbMY6KEvz5CadMYJ/yWchV5tr718DuTArTpVheaOr/IiIsO1qtTXIq8geMvqBpVvb8lLj
08Qcu7NRJVUGJCjJpbErzvOo/KNv4IZrvZIg0qeHyncqn01iQJ62c2bPHH6X4PIL4/qbpUvMa7Vy
9ys6cFDcxdNzt31K/SfFZH1GuPVdSv5eHiNmkmhvNuQ5VQLX1rY4wY/4/mS4y2Bi0Zz8P5AheywC
q2n1LG9OuLOw8LJrYjT23+ENpHDsdYLxYv4iv+IJ7r5/upo+3AMZyN8jUYS7MY1yZwsDPAkUholi
9kQQF3q3Q3CbBNS8eiMb/VKdbL+1REhTktYcQE4j+d4vZhG0FS0zP9qhcOWkcDCYDXBAPKUY0xWI
pceeFCnxONQwCNjHCyDzY2F8ix88GLUUv5foWytomcwFiL/N/MF6qLoOI7U7w5xZ60NFiIZC3b4m
9+1ThMscCbZr6PTvLGXE1FqmaoRkNlwqdkKpMs//oitNE53e6VLJ4PMK8NK/65CwKUzhnrR2En/u
2pqHXo6fEhL7U4hacekwuJHkyoToDLgi7H17UHG1+MOR3dCEgm/qpcqqCa7eAM+X3teqcAGReLxC
wef4xiH1tf9/4TdRlyVkxkm8/nskYKXcsHMmBEH/9ZkDCAwtoJIVX0RKPnkUaLg/n9kfQ/82pp9i
c2l6Mge2uQhmyaFs8oSbxbasj/iSkFkEOs+MlJkWctil0qf0B3/aPZHnMW2x1kvWaAwgTm/iX4Yb
toabVXl8J2Ml5C3fFCYMmqwO4oHCS/28p+fKNfJmk/m712K2h25gYYmEhBDqjmgM1qTCHVakifA9
XcEjfFEkRmmSeLC6+/TWWJccYNYzU3eDL/DVe30Z9Ua1y5F00XSY+vcoryeeTh/K7ET5mWPgfYYL
9cWQpJQf/DLZYTsncn6pnsuwPD7C1OBLOyBCT2abwONceIxH3mM0K5Yraxwnfpc9R8egdw7bJAs7
vP0z56+LW/DelwPyj/rgOGwTjWr+8FTFoLVCpDQLywgUuhCe6RLKfzd12XDYpIXrkcDPDfskueVR
/6OMeGLOy00FwlGK2/FcrgYNQisX5MmMJF9aHbeyK+WJHTFTGp1c1YNT0DHFp3ZT3O21SJ0ojP1m
MvZ0eeq/2ClJvp+EGyIISVGC95rwDzQdwNKI3dgzzYitdZ5AsyxPyqHSri4GCyGqaSBAbgu1Wbjz
hsmJnkfkr+h9KtlJF1virsjLRBXJphjSaRRQgs/ztRRjTpWaMgp8XogPRzTnzlvZLmnj8XAz3CTH
FBhvStAudShuD1odtv6zjlwmBQcFwJV0O6SFO2vkK5ySQM0+cJfj7kJ6dUnW5ztP8bU98TEBQxrH
CxFjQlnBB/C0K7JrOJsQDGmMIV+PRMZc0kfgah1tyhBJ/g6cplf9Vo6eEblwG/+n9p2myG4ae/cK
VIjCaGsZSiyI0lQ87e1oIde/sOXnRt+2x+nCFe4ba1ijljwuzAAvdXIHaUNcGGML0Ws+bcfOTee9
OVCGqxOFWQA4yeYaVbgCiDK6rkTknr/ZIfyk8Y9ZNb8utERi5yDbQb8gHs8nffjvMhwClXxj9yD1
y9UxWMSSgGdKIiZR2+yBCfSCPgQDhnX8kj8yA1TlNyOMW0hSPVp8sh2hBT7/uyG8qX9qwY3zDnFE
dYoCYdB9f7Q3cm4VVVDqZ+jtwRxD4Y1YMallFlyBdDmTntonHG62FntguRTFBPfKiFIf82K3IcJm
nPBaDtWP9f+1y47+oS9WSF6EAmeC6IrqZw5I/sIgGm6PfNcZJcQ+kEYnRqB1RlvxeLgDja2lfDff
aqNMF9ZcJ7K9rY72VFN2OXylLoALiRZa0KeIaErauiSM55yowckW1D1IA5XHWvDc+N0698gTmg79
Bkr71fEy1aORWBbZg0Y7pVunPVhNCsFFrQx0nT4chLTppilylgfrcnXXPuw1RAsVXzPvlYYWJoba
vlr0hOb+B/PKnDuSG6VrGPN3NmSgu+znEGK2z++0pFyWCnodlq34EIeT9AEfLWKU2eiq5lc0uj1o
Jzq4HHiXw0Dw70BbW52kyxw8QoKYEy5Tjn1VKg1+UB1I7Y75UyWk6v2fWH9ZoC0fUlAvlPvvvG9A
x9g3MX+R1LSJDsaFOaaYBPxQj8NQ4jjpKXVQ7KxNZnsK9mWoP9qFgB0rigazLkCEvf3ownvBVGcF
0461QYTdRrtGCSBbEsjj788Uu5kh4BDuvmjLBvlDgpv9pLQKApK9qTvnViMqGF5+Xk2x0wTUDAhw
sACWrW2T0b188T9gv0rXeMxzfg3zLUyOtKm0aMkYspn0CfTfqvNRPq9rytft5LdyJk1i4YLBvPM7
HrmJuc1zNiNnwFnZzT2u6JhkAomAOtExISDaLy5S5ZhWm0NPSRMGv6nbc51RcaqLRj6eET/3vj/2
M5Qmcf+pqa6A53l93L5rIO3+xXdZ1Kp3EzdrRleM86vUr4tYv+3i0g+bikyoFMBpNI3U/5cQtBhL
3FOL8N2znTJy1NOJAvAi8zWarEglP5Cz7aBBQ5KqRhIUnbPoLn3x8oYO2XPWORBR+ZI67dTpGMnF
xQAYKsioXPG8twX9eYHnNjJdTdRPa+ba5VLdZCbbfj7UokW4ui1SkFOYvJ4Q/uolpgU0TCAg48SK
EOJj84td/9anj0TWlueTtj7E74YTryUq+QWHRpynITryc+rNok4eNzvQL/BKawsaT1isLnsOa15O
EUpY2lwTPWTea7Mj19O1zluaisBm8VUBBeCObFHCzWiu8RX2X4R40G6cQ7Itj4Ga0CTC3G1NKKlP
y7qqsBYp6L0n6mv+H4zB69DPhTT3878wQMHVMrVrVvsVDyEcI6+9yj96rvsJPMubr09sEfaJ+LxT
6kH+aCpndGEV6eKJM95HDYK6gwg/7dGPO2X5GAmFbQKoz0AaNbxtLJiS1aSU9MWEF0RD5rUt0DPR
4fyeKjaubVgsE2EWGWMnbTT0ro6hL85Xva2luWh7N31itbr3hxFKixw/ZhulJcsgaB9jYspAuZwx
zytUgxzb24tLdgwEwfO8pK6mi1mTQ1JGMMl+eyQUDKqEAVAYThhaD+gyRWG5B8oNy4cVd6vqwiW7
wxt4yYqFnjDt4DevE/+YhVvjTizFEC1+WM8sP8BFhNTFLvHute4kIrZfmSxZOiLLp97wLcaYPD9m
m7WQ9+IGYAIMZYfEnoCxEh3nP/jy79MTFgwIrszBtQ0JsKgOUKpk7qqTMzhY91ofirwWyWlCroGs
Q3rHeskmrp973XPKNXNtD1eMA61AD+wHmyfxk2QrKQMdbFB7aC0aPTmkKzP9Q3q2e06VunxUx0cm
dOIXbnQJPljluK7Z7aO8R4ppoBDBvi7kmgtM0/d3Mxd6dGKgcytIGhrhck/Ko3EaLsfUG100wt4H
rqp0Wi+Bw68hQPQqM80B8IrgjIKHoUQtt0OfR5nK4EStAqk7IsRNoeNovb/y+CQ8JKwbJEcImCKY
2q3ZGU163bDIsEOy8cZWdgdTs0b7BLLVUkvrc3jD+ZDwXxrhlnCmJheXfX9FBqlSpwwgzDYFt+9B
tVxzf1vSwVXhGZt+O+zeFhSrqmHw6gq1hEEuuYlpcitznwUoJ0Umdwnsflf+e/sj5b4tAJXSU0jt
W4r4tOi/zGUbh+KgLDpusQB4pdZJ5BRQ0837wrIFl/v7NEXazLwoDFjGqj5rkp9md+oECJ07xr7z
hxSiiMEJ2ft8K/3OSWD6HhO63knJe++hx9nK/0piJ3fVaEoBb0mu1/b10Ju/i/eyCBV34sFwSPFX
VVvNPQ/VGxt7Q2EasJg1U2TXDt9mr04Ifo7Arlo+z1+/5DMwOSvSjeZdtFKRzwIca6/KXJCyxrxv
49bs4l6TDo+j7IxpSnj4ZZhvrvEhgMpSveUO+y2yiRIXHh0PGpjfL632Jn0OTyXK1oIzTfupu/Jg
zar9tJkuwq2BDoGBKpmZVWoqryL7v04Ho9zvBB1lCX44IRiFqGdyV38vvaHFu0Xpp7iKF18qQL/1
30F7V9K5yi2hxsWyMqViLKlBWHHui2k4G2iFunu+PFWCCNeCgjcufrsf2YqtOox85pg2GL1b8g8V
TtjzNTwCA8lAvOkMJvFT5lQsFKyRbSSUIst+sCrfYyrzFuQNOWi8TdqocYdA5ow7DP3jNUZBu0Ic
Pd0QVfcZJGA4DEUoiE5fB3MBobMKqPqb4WT4RJPa6WTqiZzF6Bl4c5X+CKEmi+rVzfMps5Bvbxzm
yOcRjrNKTA717e0f4+5Ww1uuyvLxZGF5CCLTowZbME3CW2yFkSlDAsayJC0SQxzJsbi8eJXXEZDD
Ck+0cB6P+tsxUgPCG3hLswlv43NZbLeK2cvwm7TPelkZdb3UxYqsDZM5XXkh+7JSGzhMn3xht6i1
2GTI/jemmSA177nJBANDkS09rM0TOF864pKVVzAjGKEWnzvJ8Iizc4yP7ilSLATbsGQDsrG73sVr
3tucM6vq60wsUBRlGUB2qvVRasf9M0o8Ia8rP4pQIsQZdRGqtTiyuy6cAR0dQ1w6K1ewT2dshztJ
VBrdbfKgY/QZu+UbKncnWECzSBbuMsiPgOJnnaE8+Ygb1lfn/Z/3BG1/Z54q610RaFuMpvZhzOII
mrvTrVmXf2PCpHv8K+u/9w2+wRUOIc/3IEhiztweZCznw9lKBaYsobNcJ7xoc76XuBZfEzdLwkob
AWjhYMn9s3ODZwq0Kt+er2j4SFEqbv+4+4dEPZL0aiZrBdAzlG5gQyiwXt1qgt1I3/5+WQrTi9io
2hUUlTANwtZElr4H8CCL8RPxjYc2zjw4qb4xvXk5jrh3UBaYD1B3hx4/BIEDvKFI0a73KBO3qlfM
5hdxY4eiWC+EagxA21q+/GqQ1WvAxg+G0OQBPwZ5ATCfxa77ZfSuz6xkOHVl6c+aiB+QtdgTubze
nPaaKHEkRp/skYrWWPokfaxYepV4ZZ1fTn8nTIy5A//q34/nBmAV+JcNyRMvx3fLPNyDIX6fosJ4
nVVd7lY3dlCot1CLD5vveLv/DayGC+5mJMwZCtb9fufkLgYIteyNHO+7M5ItnULr1dr1bqgR+ehO
dd4hTO1+XD+GkLRwwh+FaPCV8O4XZlaH6Apq9qDaiz9xgaML33OYLj7SjKg1ZRjVH0VpQil4p0er
Pee9MT6z0GYP2synTTAo8g4IbqP36pJA391p4HGQFUt0+xhk9Dk8osYpI0hM1ijUj5rexlwnyMa7
ygJXgHU+1imeEHMUZtSWIUIjHU9cHk9DabJWrsIiXU2wmrUU4vvye1UreRk8BrRAI1vGZwTlbl3n
xIoyovCPusn6hgr2cNk7N2pizxV84knuiyBD/Xe/Zycqj/p4tUnRl89tZbKP/NDnQ23gSZmiShCs
tm/4xtAxmrxWiheudSzzXG1QG8wL66WX0DG/wO5OxExu1+Cx82Xk/1gbvwveFQ5pkmJkxalZHXos
hPuFLGseuQdwbhdSS36iv4JfljjjYqMmQ4IIF7LjNnSpioaQFo2L6Ms9f3wSvF8WYC323r8okCzG
KKJV5OSfyRmJGWGCeGxSbt4LNcDCImOQrpvEMQlkZt6CID0/iDjHdg8DsLHprDG4+00vR7Pe/W+s
agMknLaTXn2UkflqiD/Slm+9nGGAU694y0m6nuTc6sxQRXr6qeKa0n0/NCE3al1OZr7n9qYkaR6J
crmZ+vqsZE78395gdBV9Z0iUR8MDt0QGf+P8Q6reR8kPHt4CyiO4H/ZvkMUMmCzS4MoBgrJwrgbC
oQN53DWhNTV8+wqWb6ZBTsTkxQG8k5jCvKvxBF5VzyemXWyqJYrqJRhJHzCBkLETnnM1ARlPmN9z
clkztLQMCpvQKf1xBKeByTOH6dhTv8cX7Z7wgQJ6N01Nm+ZEFRwnYmqmWz9t01ZzbfewOF/cxWIw
xk+eQxh+CJFQKj5Sh2uVfsVEr1cBN4XGKhY4kVKFP5b1Y/wI/5rul/4Wx5CDvXqgvWP3+k+d6ozH
21kDRNJ5iKWr8K1oumfZc4OI/eMVfFbWCWuKQXZOcQWhfJ1qroPXQ6iYwsQWPiJ7hTMMTPqlEEFi
jDFcaVqRbKQ7QRHJT3Bq66dUiGcVlMDyl/Z8zTEx6Hm62NkxQZ0CwkUCEHKEEyX7kP3Y9/Vyjm1H
LT+sgKnx6hVI30YL7mJbQcaFvtgtPDC6P5QQ05woX/8y2rZBcM9t8PDp49ctFdJs5DNcUWtqojGH
bZFsHcJoX7O8Pz7VSyvuVAJbHbbJf13MedJrAu9TAJim+HXDm96FbRYuRbi5qL5pSdUJugajaBsI
1Wy1s/qQ7Dioy5zyCuXkDPnwNBncxNZkhd7GQowzuXS6o4rnju411Er6Eg+tn7TuT32Pl6NUhiB+
h0Fd4gInkazjjZusN89Gmw18aCeRgWbTZC5qqdo6sFRW8T4lkeAX1TcLq+cKtkNevpnYaUvrBxqe
Rr6K3+l1E6S8yz3glSrZjbO3HtI5DSY+nDkEPiYQS5FyYR7wMVgjq4tuAn1gHsNiQKoiVljTcyBx
Iyh/pskbG94a5H1SW++K0uc+BS3VXWcbR4YTbhpeUEYB1m3oQy2qDxVNRg5oyOVDHQ/CBcbK/kLJ
OXqm90tO7LdpA8l8cwZx1ztERBe4es2Ffru115I9mpeUdyVEebkhNYhWALN3Gmbz5v3x8QgYxfO2
v/5qEEIPDIljLb0O9gYItaG9/yVQLneKAwPr6XilPl01KO1XNincCDeuhE2i7EHag8CsokLJ0d+h
Y8wA3hs71TAd7s4dVCtniJEbXqCyFwZWMMuyg5Fk8y6nkFqUEW+b1LG257ft/Zvuj8fIMMivU5Mg
Be6QrzaxoJrYSib3OBJnYCvp3WpCM5Ga1jaz2XmU2YE4+ukupRhoHGaT0bxebEGKluSyDeOXiwSu
o3NC0qYHAAdNsWSCGWvVEQkTGkIqxHaqFEzQM07heRAdj4Aoz8A5o+4pPjqUqd+2E1YVRKy8nPEx
yJ16u2XLKgZShaRwWWZ65gyMiwnhnecSmvvxyP5ERZT2Tf262HAY3WJ96g0+0PECFFXuERjDS4KK
Gxwy2nXc9dq+g5LxMD+/IMCFgCf6GnT/rOI277NUl/berXnZqU1AzB4NUANxRyzp1A8i5SpZzWZe
TpBFnWqK43HgLJzbrbSJjxOiVwtC6srCOVdaO1Qutteux44xmHohkg1F9eSGfRycfikTSJeEs0Ja
U8Wh3qn2fubITpYoch3oV854MC0mNmj3NKaktn6fNXNkZB5luarKoVw1PHJitRP7/XfrWyws6LfQ
rnPLLDPBpqzakzcP9iYOVkwrsRgKXpC8cXe1XLZylaVn+NwE64JBAtYSO1qTjNQ65dcFDBfZf2kM
n1W0c583C6wNyIsCiHdzOhUoP1V4IlZ+szwlu8cjvgMJfrIVXjWXQxwWq+zT27wp43QxfYkkyFqO
hi0JV4Tnr8/ym31fXPLVc27+XCrWcLs8pAae2xsrsGbxHhG7v9PurpQKs6awdl8B5YvOuu+pf8tC
xSjRq2wRX9RnAbWjX3Nrq6IRMOx1dzTNyEquO6SrycA8v9ZEMLSkrdJtNpeC7Q0PFvqed89GKzze
de/uvpaKmXHhUzaQ0R2y1TjWCbdTQKZWc46CHM6HhDfxj1iY7TW9WmGcgnWwby4drL7h34Dg6lMy
+HwqkGvrlQ+yxb29aL16TRAkMvDiJjOsEC36o81DvSsfhk/1ttl7MnBk/eiLiZZbiH1GTi4z0o3z
2wY9CekXEfSs8xqQ0JY4EFaztV3Ct5OZz+wLtA6dMHfWw2okd3nFA16gn3pmiQcU5y/xkRR2VGfl
r8R4vadx1WcqpPLUhOK3dn7UAVugupalYRPbDST0fx7ZNPlQAO+6hZ4r3yR8QHxyJTbUiBmRr5c+
+WrXH7fJRFIs8eYWxJqOPeVu+d/sdx1m0lrM8PoFtuwpx/kDLO5YJZxVpBt0EM1wZdqoBKsFkgsz
TkTnMbD2IctB5XcwfGgp/40sPAjwNx5CCXsSftdC9m6FohBeDB2X/B43B2C9w1334Wnz4SN/ovlv
0MnrMB2Ql2QX5v+639kQPYimDgj+rM16HfMhxa5EY66aXCO9fuoFg6fz8y5Bh8N1MpdC3S5Czxqr
MCSMH2Bcs4cyA4Tu6FHiQEkMfq4lB7jZQTsspowPn7uIf5346hdUNY5ZPKRdbgDmSbE41eEptG78
37iFp4vtoIxTjd+MpqjQ+7fCcV2IWZTEm3FN7gnxEhkcO/hfA5bm26+I/ZiW7Ss2REwLIwIsy2Xg
tybp2RJD7mUuAcVhEkLDHr+CnpT56QPe4nQfiJmaMoatkGVz0JMiD8nelQyGqXKlyNcKyB/APr5L
DhDe0mUaW9T/b1GU5rGEhb1VGzjR1Nt4NzE5/z2tTXg5GklLF7DObuiG354OvbnD3GV39uuL+pXs
/lh71zD/xHUsLzBt+QegMf6dU5AnFxPqrSwmlsmufwylNEC/MOeYsmvF3BmABwijOgMnWDvchEFv
sKFhwBxflw0eqqh3D04yadfNRD6QRLdt3WyYsSjOwOSw+Ys++mF1QRmV70ZrLYl6jL8cz0Zh6B7U
Cbhv/POzn9qBx6RN/HxCnNPOWP2Bwp/96S5F75nZ4pdMFuH5SOjraJEv5OFcGVn9pgwUbFm2LOaW
KMGd5O9p0XCs6PbeV4Z4A8wlzp7fOSE3vPDN0kWCXsR1J7g4r1DP0N/SfIAq/QE57N5QwCjwdk3G
Z4II3sxCPzABsR5fVWSJM/+7+N+iZA/gdVd1Xu6iG8Frb/wbkMuL73KfjXtNXqGMdFfvxjUtmLJz
xiQGCKgQ9w8hN+JV/Er+5iNrpcGJx5tnUAjjm+xHSG9mEUzKz8ms1rVmPSQI5jJPD5v7DPbq/i7n
I5TEcQF1M9LPZ95aKPWM0ZH8RubDhWLgignLYv4Gw8ZJwzK9ckO3rfcFXkZMDL+nYJhPjbd6qxL5
l6PNTMwvrUKTmJfhnhqt7dzNsXG+BnbJIZllXcaN/fkDHPE7USPExaGnvaunqyISpYLKxIMn1swI
pb5fWm6qktHZuib06wIWu66tYbZ0oziKtB/+83AGeZW4FmckiRsoaBe08tqx0PpDTwzMhyHvE6Vu
Z35q40F+PNPMtCRbvw9tooZFwQ5nFBv5C4lqIPZJ8W7RlVXfSSx9L5T2OLFxGXNsBWdHZdQst6gp
0tVpjhS17hUAB172ApEGsqSMM1aO/9QTyx3HkDJwh9CPynmb1jWGO6VvgY2s+usmpt1nIA1BXhL/
lQUZGgr0aZV7/W7hKwEKvPzFQpnL2i9WCRftMOso90vDooqoG0uvy5Pwyt/dxxg3DX9OGWwiUF6/
QijK6gIoWXGe4eijivSHHJwraMh45GR5eWhdSTTkkRPM8/l+Xj9UsgU5i6sWeRtYUBY4AJEWPeR2
QTV4fkJNJC3d+qsqqncb4FbbWdv5NPr1fIHgFPDLdsWckNK/PkMnXAQqi4d3KLsCJFCCl7n0djDP
A/Llhmepefj1wmGoEugTg/fYp9koFEYKz7Ox98oYolZm0Z08x10Sa6Hyrr6VKzlitd6mfe6lVTMH
FNYqzzQgFBkmVUki4BmEb3uqvAW6+Pco/qnUASuodM582f37zMmL0Yy+5g/FRhkNKz1KCZEgddBj
Z+HzvCULHLSnXolOB+QK5KaFRKDY2LoHnxTCm8QDuDKoam9dtd0YTdDV7uRaL3R0UB91VB+DCDiD
0367wIEdf02Q1hnCEPDqvxG/03Er6GqxEH3YkyFX8Ui/GHVZhzN1BLTSxAn0kVNCZ2qKrhmKSVVw
tYvyc3Ls8jrZ/WGJMEZOXFU2Tw68YXM0QqYEC8bCspmSCctIwyOBTCr7cnO6VxsQvTvtjqnNSU61
dSLjOp/n3eUb7lphrrlXOZBmWCJ32cF6az0NcpZPlUQJ81rG4dWSTt0eHj/6hzOAfTPfGwuD8PW1
OGVJ5c4wlNKQXabEg+RVLsyhh2vcLkhU64MYcnf67GO1L6GC9mWrhV/JMhVQjO+LsX/NdcknN2TV
nEKBdC9nI1rLuymmALGi91hRH0ngO20KgzgoffWu0CC0pnfc/h8XSAD/dah2j+RUAR4X6sa+14Re
0lACzwpY3LmypZATKfFzttPoR/+EoDs2d8YNBZoUPnUW07W0FB3Wk1Z56+dQDUZCx2mwzom9oJ2t
aFGe8o3sGFM8tP3+3Qu6Odmma7EXUudvPJ2LZ6upGDxt5HKCfcxknntA0t/XZdIspwJRcQFOXjuJ
KHAqvpBRdhIqVD246bJdP5NMrzN5Z1Wl7JWvZRM6Yq5wBv6VyqQATvQvmQq3TsuY5NWe8OpKH4U0
c92KSW1pK/HaC5ZXdyYLo3iSLumtGzuC1THXCuJM9lBbOJs7z8JoOE2Zyp/hGou3WNCxbNu2nnUO
dMFimGB4BKNJoTq4MeVwciNZqknKVnuYzjqosNtKzfm5m1Dm9nHLJ85YPyn3qPepHfWSyg4/AJYd
Wa+1S4+n80sSgeAPDcBUuClw2E699s5TuazwiR6J8r692DgtPll6mgOhRGM5L1rOocIc8rIXIF9F
4ZTXjQMeD/kDeSk9JXLt2XzuXqQYLWN+ZiObxQ1y1sGU2YTv2tnTCm8l/XGYnrTJwuh6+2zDmgLX
vrpauAnOpCeD3Ar3YOoeqmlKnaUxUvt6C0PR1U8qYXYRlvCAkSk53BUporDePs+F6aBItT1tG1fZ
G3Qi11gVBAyhooN4Thm283Syb2c8X4LU0g4SxSdProW8zop304c7tPbvtG2UIbAOvPpZDD1QWXwZ
2dUu2A2ejmRC00WrTwlulRU1J5JbAv5i8tnYM5OKPt7yBWzgvYSAfGfXkuvW7+I8SDUS5u4ytHiJ
U1CEWBK5uUTF5mnboW/nydUeq26Y1YrduL2ZlKGGJo6UBweK0DWC3onjjCWBwYOxmMfYIhdtG61d
KUZCVCpMAqzTdEJArWOfU/JMAqwdp1BKJ9a8DZ4zYRqjsFECi8DbWfjR4EnsT7zvOUPqqlplSIns
6TBtzl2mZOhZSdRfOaKvJwF7c9H3u//ie5NFg0dT+zeKx+bMmltX9iY2uzF7cseQipEIeXJghxea
veWdkvKExJFFVOsX6qT8ahnFndrk+9ebk0CYAzWDRF5t6bxMVP47/3W+dGi5GpJJPd4HXEti6M2R
b9rRq6jEHL4h3gL4Cy9wjBcMtZyyNPg/2nGp4w7ZbnaLddOovRvezRotiiYBddemQBROewuc//4a
/QiRdeetbehKSJJp2gEnkY1cGY8v6wuIz5jH57/+i8PxJRpeTSLmGOAPlUwlvBe3TjZCQ/nSXSoG
ff6qOU3wXUARoP+chLsmcJLJ4gb3wPxkHI8Tu8kIl5v4BArKGNoU6+wGlC8P1jpUronMDrsW7aO0
HgFsGGy0AkferTAC1HQRZyIHPyFUf8X3E89MICZ/gzdBmdPvrrc6ekB+m7QzCol1njS/1S/HU69T
1Yd4XTscQTmHQhoAH1aLUjhvgBWkzgl3QvCVZJ2MFtxtHPS1wEKnx72mop7c+lysukuV/uPYHt/9
9Hwel79QD/Dnf+PwebXBOwXabFsto4LvYvYmHhrnU41PacOYc4SnsExwrECrN7i2bclwcApMmPcU
Ifd54r+eAnNFiJeeXO8LGq74KiQ6EIgsp0J+YNapFj1TJpJg0yH2xwFH8ikUENx6kKCl0xQ9iuj1
a+ZEJ6MywtOkc7UGV1OPFUzA2QsYD8rKJMheFgpCDCU+lVAwB66kWU7MmH6uMqE8hHsWmlndU1FD
1+Ci/Rql+zxOBsHOE1FsdvNIFYuVMoXX68zuaId5vxoabilPeAJW3FCNjomAxAyfF9dTG+N3/IU1
PENJFgU8Tv8IJN/LaVFtYUOa1UQF8MhPeSjVmTB22exh9sTLGFpdSHyPSxdJpNmoFieCv1k1Hyii
Hc3oKu1V0GffCyKlxwqkYT5gSpf4va4XehiMdcqEIpQAGr0JenYMufSOUy+8Y9UlpOIkZedT1Ii6
QMR6ZWnKrM3QewFpnXpJpfhrMWDt3M9D2r7xq989n5M4gB5p1tEbKswUJiwJ+Zuz11fOUx7vzNjJ
UggJHcgMqAx+sK4Ag97iGY0zHIN5rCHpxORxR6xGESCHsIQ/f4eAfgCGOlLQpMXPayAL7ht6JAoe
SxhcTigtppSCOOBh7HaWMTgX1Tm49G8CGtEDBee5E03kjXVf8hETSCNQ07R2yoJqvipqwv49nbD6
MLkwAHM10FI+Q/P+tj405QjjkUN1i4M5ZDTXD3ORXhwliYbHrBD30297bVV/8VlR6VFCd+9GehcP
2Bix1ZvBrI6OPHkQe09tt5hO8OWsjZHUO7Lgr+TBsNk5PH3dYAd7W58Dcma2Pj670VvIkCNlwxuH
ugvBMngQvYPnCGggKHLBGCGDQVNs/Vwjzyz+biTuzEZbiHRYtP9SskxTZKu2xiExVRJJVJbD1xkF
PtpVINAZQA3+I7gE0O8Uql4M5P0Em5wdpRLLUT3ascp+a7qxvNoyczlK40BQZzde+xuXp2syKtjP
pcQDGnVT07OLcpZ0W/68LYjQOTf9XyIuaoPUOJm4UX6x2LoSdQFphfI0FFOdj5KwRUSPr18zYkkX
LrhyhG09h7Hy1egnjDl2XunlAQgyXysDBl0AoiLv9jqR2o7k37GYfB7c9PeOt7jWdf8fuK4SLjht
nAJlwv/im/MWshd7cMZkyU+4GSAmq62UOBV85MnvEvlFpDrodqK1bVqy/cCoPSY3/KWzIvu9z6Yx
46sn2X8tdg0wQextG+Es6DRlL/KXVge7wiCW96gSnqUo/AHq1x51CxS2PNJrnQTJf9f+rlKwJj2D
3BdycEj9zlC8CUInGlQEizq1aZg35Q8kgCv1B70f9EyT4zZt+bq7mWKJwap3F8T4AQ57zafDP+4z
Dbb/+QDUfHeSv0KI7+vJblVDa3FRcIbKeZxry2Ft+52b1bAUIzI64HIb+zGN1s4l4FkGkRUdd+Ri
EeCkwWjm0odts7rfBLptDksmsKUoYKgDvHeP7ztNGvug8Tq/GNpGcJIioXOQFfoAy9dCUkNZnGiV
TsOGSdxMkSvgzfsnPNNcEILruMBWx3k3odreNJCU7afOXiCM0oBIpDJa0t6pd8QSfsLGvJLr+lWZ
vdgTa3C9p0R1jdGAcVS4JvMTot8ZDF4zjwnJSxUhaELtxu4o+rTaeQzxSGDS5icIpMUVoOs44Oj1
rGGlNOgsifNVNiRJTXDkgl4cxe6jbLEmZSgVGXEGvDYckP2GX3gQVqFr8K3bSVPBVmwaF/b61+Hz
enfyJpcBjEeJ+VxeY7IUcZRxSpWxJQIp34vmrMvpx1PQ1nykxmkLQ2Dm8MQop2H4mRmvWM0X4TLW
tr860g3KSAnJhqMgT5XmfjgTYvb/YcIw5N35RGzXEcrtJAUeCkItg+meaIH1+w4HZUvHafnOZuNI
onmkKDthftrL/CSJXzTQxWqCqO9rqz8I8l+u2ITH9EDIvsWIY55/wTmllFWJnRus2GHXNmXsBKll
pYWLCgagcOlKjkMJQSMalDjqOYlaYkPZUGjHDF8gNpiFTt6laANe3SKSzCHzX9MnNFwxy2OaCMy/
jPqbil4yqOMVWVP4VE8FvXm42gPMSkGc3AkD3NELRm+QE9Kc+pVqulgVoMlQinqkllZd1Gv5DMse
yymTuSZEDR8ShINfZoJS5w8oIAIN/GcwnrcpeEraKPgB340dF3Ty9kQ7f0EcjSdsTFAMhrujB2KD
+64ouanIkweCu19ad8jPf6M0Q0uJ5esnjmx4iOdf2rC2v0TUrmDe85+CXefw+uis8ho/7cVjPPRw
UF6VtfXEOMlXciBgYkn004bJRO1a3NaloDeVf0tAf+vaAkduZdJbcC1Xion64fAKQpBpO5HT1lQs
OW3wOe89WV2aZ2ycgLL+fKgmsY4njKzmq04l0Uaa+XzKRu4PZog16b222y5t3d6N2MSdGFZmXCNM
/I5CCKlRwVm1GpZECtjdw4pbT4KZbzqdN4gWkfUGHJTXj4dNXFPJdBBeh5Db21LzsaWW4RL+YcK5
SQhmx54Z72C1AcU2yPJD6J8mvVYNgBOgePMtXCBuVN6gwn7AqGCggqFD2UqTdZPwSDWd7MuR73I0
YfvQf8EoYvdG6HyQZCEhOtnCuBXC+tsH7PuOgCrqg+U92bzLcaAxDphJFSstyp90UWvf1ejJWsPL
iTLNUIh+gqU42d5VA3hf9CtlDQTuS5hfgITFc5C3iHZJl59GrY7p5yqPCoUvvVZXzmFKUrhkQsHr
L89vcV4f10jHscH8nBeIOJsA9xTKmpJ2EFZ4duDWHKr/W45gXKfb+cX1maChhn/TgssE+x9mjdkV
KKvWJy/hZQyiI5JgYX+abvCGS/ldMey5e4oijyocYKZfIGFHCLCmRHFbN7zgsXrsZq/QtT2yBpyY
7P0GMkuJ/39DNQA8AAPtd2rZD7WIciIwqla30mYfmSLSN/z5pQJzKQT8YTJApQNrbc0xVXTbdMOj
RE262QSuwmCZJBWlbVz+MkQMHapPMDKpDwTUvnnK6u1xYsI5SmrVV6WZH8SY7K6yVErkQ4fGJrFZ
H8MgK4B+CVjd4fFvigigSm3IuIrtjzXK04kmN2gf/ApjdnTCNu2dHvnXxNv5CJVaGIZj0tD41TnZ
0jgnlotlQ0//Wlrf5s77l1zNhovTCdhCZjeDNIzWRyctNr0yt51+ASDg7sCv3bd0GdjveZZfxJK9
KghO8QRwB0vxE18GE9hNQtzgweVg1wQOgZnMRvyMN0mnFaODM4x5BxV5BQeH24lhxaZ2POhVRkp8
hG6C4NZjsKOal7y9dNLdDxJI3OKKE1Ph4Rx1KY2ISE9+k/re6ogH7ccE7kGWl7zBSzcvUUctR/K4
789Yn/gHSPyF7NqUPgEPRoTwTcGNNJUD4yefT0NU9T23fFrMDCp+M0HbXGT24a/+YjdLncZqu2Py
5no0k71Z06tayvOoWnFSMgc4PuMB1XaCuhMfi8zpC3zQTsWitlojbYN1zGzYKwHqfbxCg9vJqh/A
FZfQbZy4r/tCZI86zBGqc2sveVk5RfEJIq02UYvJa5baAQnE96iSDls/ZMbJd2oVy+Hs/g9bmDCm
VYwSSuzQ7GSTEDJ5j5g2xvTe9EB6zsEQFXQTF5xhT32C3lTX6ldxyjC0c5KNmdiOcDcK/TPvi38/
oTfI/CyswlFqDCkNS6VFOEQDWry8dGPIy82oVRZSLVg3i08rU+MgiznCjoZWHpw3rffKTUbv18s8
I/5x4YfadcjCDZNXU/llUmMmJcHRDqWsr8m4IEgi1tJV/QuWPfCJmSNmh0pCEIF1LLGuTFEWH96R
kpUmuWJdYEnuuWhRL+E06TfIAVal+FksDFjjVEuB8dVA7s16FlO/irVhObm33HjaqInTC1VrVN5a
2k4z16Wr8P1oGCxLl40ELCZq+uD9zqs968VuifHzVrUvwbxCE/kXT/deKgbOo1e6vQNvkzDB5Axj
lYx3a/vUkRMDeNEqasJHnGPK+QhgOrey/kjwZLfWXUMS30qwkUQZeL2gdultfAyuerep/5TnfLyo
3hT2cbCscITV4BDOvxyCwRU4iLEoUdbpbs/OvAyZiG8ldMVdvh0j0aj+ao+NZBXz8oyiSeKUJ/xe
ugFNM+Szu5vqeVREifvp9/4HDgtEyJN4diI/w6TJ0m469SebQracLyVk2lu/MdsaJZ1LMbLZ4gvh
e7BFabaJaSOX27X6NQmK5aILKTLcJdvsLuVfsF/ICN+YwwRCgnHJn0kavoCVibA8MLKgx53RYTxg
rhC/VdQFohjIXVisWVtDg77LEoPRVWdTsb/flMAnbIEYHf34LIm8xbUPlTdH5Oa35t99ZIlZFd5y
iDpxRQlHmiC6F6hUz12dwoEu/P7+YQsGRd0Ykldmr3kRM/cr5Ws57/4MN9gl4eNmNKWnyD0r31/W
+Q/FJvVE0KCzU16T6ISqrJ7e00II2RdeXG+DbT9QRynbyaQFQD0F5aSwWjHIWwYEpguufXBTaxVk
Vy8phG5LzDdVODQJU0liVkDpu8N+6kEu51c3GF+24f8mhHS6XO5zyvpUqkmpLbZHjdOupm3+NVNc
bN4G71AWG/vN8wQ+RmuyKXh7UT6b8S7EaxwAcPe/gLa2g99hF6otGnmcYihlUXGlojQPqXLx/Avt
z1eHVcj3eIeaAKx4njkNv3WYzY4PSRMp/lezbYiAIEyD4ktYms+njc7C2kyrvFfkqgNIFKWXxF6U
JN7fjq1wS9C3EPWqZ92rpLW6G4MOXSBvYb95UGNulgk8qAp+2AQYNBPZtafPfmP//1sOpmc0xopT
dAK2QfXMzZwdUzy/khVusTvwgbXfWFIxmm/Q84nXpVETHnPfXLu9eZPBSEBtzXI9veH+rpYlwzDN
E7udT/BVpaKcI1b6eOoAm12nCrt1BSgGQIzOfd5eimEfY3KFIN0OexZTODWzw4JbizWRJAGwPmcf
vGc6DQpeLJZxj7V69OBTmFXn1Ngo/f71WBbcSMcTbIsviNaSpMwfOyHCWSN/+ZFso68yJ5uSNZfv
OHqYnvqR3wZ1SOtTJXI+55PJ9Hv/+/xH3LqTS5urHiSS+yTmLJBfeCKflLSSmXbFowexnSi+kt3U
iaZxlZK8XXT8E9ohih9lcR3yeQxdBm2ylPNF5oqH3/arkZZbFJRPoTnTDNFethxHlFZ71pl6XSnN
18yVuZcW0E8e2CDr2Lor0RDii+rY5Lcxv0Xe5SKFJV11IygguYIqsScrODxXPg20U6mxm1bqepom
MZaSVHlBwJwrIgL7dXLZt0c3ZkHJYdTbZ93qcF2/u+inm74/YtwgN/TOMrpopG/A31qRQT7WZUkG
8LRt8EC8RN8d4ZwobQWEw/+l2LOGZIRelxnfqKmBAmnISRYa8vkdK83LEHYEpGXOcMZ3u1hRSbwE
PdHtVSXM0C+wLHMOeBdz7m0m9ui249p50QPc3vfA17TsmhwKKNt6ZYw7vhSuACvwWljQHFqy90fp
G+JCv4e3XOay0zI1zmC8EecZjV0O5BpD+L93dUurHw9VSoGMVyGvyNZMbzhJ2+8W19XoRt/T6YTu
lwQ4+xAZVGs6yr4TVCrEBTAovSf5IvJGF1bwEw2G4odUbjPLJm6CefYLKfwC1DJDVQ6U5x2NMwNW
KTovOUncDlr1E47G4smniZK/ckx2iTgo3IR6e2XujXxI+YWqGHkmOGk4OT/r4FVok2fnAk5ZiU9x
ocue/Rc48GSDe06t5ZCFntEwhzM6GPwl36fW15DzxrygHw1SMZuHS04PKu3sQiIpIbveZG5u9Ptm
4sOC/LrYIbn2hIsLAlFprVAHq86Jj/8UmkKaIdrMCjohROf2B0gTfRlOkXLcZCa2RSTgvOJPnLvb
feKeYp+Yf9YpmYDkZObA42NVFacz5L7Mmp6vYdqHUDwoG7SujnsRvaMKzeLjxLqzueDFO4qU5rOT
y77L4N29Un8G/ObxHe9UKbA5F7UoLZZ4R/chQmxyAN9D0EW8kHvaycK0vYOwyhFYOXgBsUjL7pQk
ov+wNkhxV1SZfcOLgCqhTX1HZub+hCVGkrBBHPI9eaonjMlGCiyXnjsqs5KoB0YAAc+bNP28GO/I
OGgG0M336yL6cn8AEcVDEk326Akl1Rhe/+9AEWGZYIL81Z6ZvBvK9pwv5zZF3fMxLUR6PGvSrFwS
BeVq806i1+ivaNvo4awOn8XsdXCK1o71mrnYMgv2LRZfCnZudJxKL2pvJaRV95c6R2LRqb/YPX6X
KH7DywMn2LaFbtH3byvsX7nmyiPeEH8EmpdUrvLxtlXE1bEcnfAAQPnVPF7oM9YqndNnuD7QHDdX
DDyDWd0OqXPVtOj35XZbgfXKw9K9uZeLCPwn1RSRUxpNorv8tDhlTGB+s+OGAxFuY0EwkaLcFFwu
WNX4lX3pXUgbSZNkLwhQMaNtHMJtb+eN86602BD4mV19BjT5cbzLKVcRNmXDwzE8+l6Ab4MBcWXQ
vK8txMNhi/Q94P//xH4H9RQrOg6ZkjEmY/E+YTA5f9XM7Y48I1NTLSuM9tSGN+xb2TL1x10xgxlX
S/efop1y7CmovNUoRjKoB/ECL3FckLi/IcnJhBwYnkUN225IXl77gRE+51nvrSopOzs65B5Y7PmY
ZjVrX4RCRhm/MHp61toF1dpLXeZfr4MDYHatyTjO058JgQxEjWDiEfMTQxGYFfAju3TrULes4N88
aSlKcu2dguLmyHX00Q6bAj6EA6Fr3FMsKY2fRldc0dIsVG52Z6+d78liw8lIFzzlnemeH+gY+7bH
ThgN87YO6gGOD30eV3400lVRTu0KY8/lNihE42L8Vf8W8rCb2qRpOYH27QixcvteaIm62N5MYHBK
tsmP+8P0hLWbihyyfd0rnjfedkjPcQUBSG2RFwfT/00MzNzkXV79K81/dBVJiKefnCP3VV/dHOjU
d0TSWA07V0rdT2QU9murTqWa+p5Z9V28CovQuynEGcNO7Rla4A1Ex9durRd/16EkF3wSbKWNdCBZ
u1t6/fj4k6AecxOY3mXvUn26RYcgNURwrpSobbO+hxICjx19YFt+wEdbrWXyz8orbs0vzbjfO2BI
26ZHHI7ry00Uq1VAGlTKzq8vUTi9W1d/8CgKuU2eGz3NoM949CV1IZtSmrykuIbuv07YJOk+NeXp
9BieRE/h1UlLjD/pT51ZliD+baAKCEHv6/fA0iOY0OQmKbPID8rDdq13GLZNhYXP4eSW0uYRpOJz
oMsYAz45WXL01+KhI3zrSSPWR1s7F/jA0gflEg+5xi1j/5F5Y30RpbKGD2vCqjzzktasZjFjkLr/
H3jKfprx5HYTYBkl/j3Y8BfKUljDiQ2B9PpF8RYs/Hno2cFNn44jfHCz3KHOGhQwirIldLauu4ZG
C7S0YO0FTDuVnKZQYe/gdWaH/GUlNCFzU16J3FXZzuqW4TIC7Nf+KUk6YOwZ7SwVBPS9lqxc52cb
bK6ZyymjzX+23Nkw83WON+v0ZVQXREN+KQzg+rRR1fmLyPghSBMtS0hMnR793SLn1ZAqEPQ7ffqt
AN//C7Y8jUvyyuxTNl3CDtadPamRGtd18UTHpYuYCyujdaddj8rok3WMvjV0elY/cOZ9a8BD9YFO
/Yu2gzzi4ODVhKah1CZl7kEUL8Tp6AzmwHmWkrIPZqmLRH4/V8sjAQsGH/nPT+A9VYeByFcLEbsa
fSnuTty3wKn9E/qHRwy0g43nkxrSjjHaseJ7KTOwgE0iNWqlU5wHXuAtVQZQqbjfIroUgsOVJHTm
7g7s7k3S3lQ4oHu+eZ3NDOSSi5mG8sMmwaGMgTDvS4YNNxWKoLKBWgX6LNYdH+/hpR5/ThoC56Z6
MkjNuFJQh6IUuPUd5ojD0egtk1KGu4x3K0SkIMHouixIp/y3fulJ5pAq/BTs3049+R1B4p0qhoyM
dh+1I9h1exqThayXiZ3tYAci5WwtPu7FgUS7bu7gZvRuAnmH4tr6f7FH5HezMDU2dJHb9hbtv5FQ
bfxd6tQZBVGQPozlS7RQxdVkjcG7kiYI3LzWwD4qhazyQyIwP/+MRCvfkVEl6Fv8ZoObGrqLW5DE
j7gucRuHrvWI1Si4esuMEGtomaQtRJiyqMawsUZ1WXVvrV1Z8//SGOqdWA4sgcjBMwOb6Hzm0jf8
k9OrNzFjePWIN1Un6G2wBXZetots8BQCA0iOpvCK3FQ7AtmE7Bz1SWNGGOE5c0Kbs2f670tEhpS9
By/2e4qB0RkTwDOO28ok1GK+RYVBt3hXE4XwViERytjn++3NPYV0iJclD2U6Is1kzK0lWM49xVkF
XA1dzWKhyOEKHiQKaP0SPNZU3LLcOW7tb8VFRccO4cWsp6ivf11UPoUP1LnImLC2JTF8S3QgcaPi
v1QgJw+poF+MS5L/HXkJsa+Y1ZstJuxSlzJaSkRko4OB8k0EAZf3GfsCZXBcev8zj3t8lC7i8oOj
UWbbzptnB7bTacbTOAnSq4jNjoy0x9s/VUlg4efT/m+ysSiq9SpF8DaIQ5wKoiPOhQOO4XxL3lQN
rVmUF3A/iGLLrjg7cSiLAtWEIsdaYvPsgXEq4oS9cICgmQq9UfwFtA3JBjYLiX/Qgrv2olJXJOtw
LOKHe4TpA1gGEs5P5H9LwKYOt51dpCgg7VOwq6krN5z4HHHRGccYW1w4X2QxyR4xBdPCbSEB9sXJ
h36O2aUUPSP3Qhqh1wa9ql2LIaLk4v5W4paAqZpWbs54sC5HYi5iWlgwaoLTnz9pEwjagq2uzBZw
A3usM81EWQJIXhkuge5eGxgxysPhwqrHg/IcS2N1hiIlnh9NzNXv4zEMpoakZrvhrEVQ9W6ZtTBp
gNWTHQqkdSsi763QOMhQ6IvLlEW7+hEenVWUJbfDjmvlTXfc22DAa5uBUXTCXCqgfEhUjh+RJ63P
0D0jI+mJ8Y7TOX87chkbG753TygdljmItooplUWlq1TdPum6mIOMsviCa5Dplrq+qiLgcamuOxBc
ixyXO0aC7M4giBu95BePNI7n9q0s2iQrlUNUWitsqWwjsg5KjFWruHoaFL2oY5Kj7MUVX7FBaSgq
fQOv5nVp0SMOxFuqEpbRI/V1lyUGR/Md4wVme3zEUxvEHmCRkCQpIsnxZqS+dARo8iPgdq1zFfN6
6ZhyhkjeaLTF5h7bTCWy+TAoAoaxriAKHky9uY7ONCIEfTM3azUMnN9DviEu7gZXL+vr0weJFySy
Pm4sOXMAygS7gc39TjiYAYFTIAtXid4jmK8bZyqbrpReRFkpf94BTDoRqvpC/0y5wffSRqC/gxn+
5iO1t1d4bXzFp8KtoQzinkWbM14CbMihVsuHvMe/v2wVCO/YuUjHUHGQvwPniswVFMlF8/bmsEbo
AJgvdIXG6CmJaVbNzlwxA7VD2v9UIUprQzEwu3IfdTr8sti0BKR6QMi258QISktMI181QWZJED4B
8j+fjcyZpTRA1j+CvTFTF881QwDhX4OktLfcJs6sQ8KYLLRINKF5gfBNOf4RP3JcFUIcBkB9XcT8
WeHUtQUqWMCa76bv4UBS4kixXYkrj6l5crmBdHQgLS/AN6tpWgJFlo4E16xmsNGpPQBT67CPf69i
BSvrKR83G8tGn7DyR3QH28iZ91tAIct2i9ttH+mTBqkBvpi2eQTWAH5r8JJqUTjOD0KY5o651W8A
H0UUyXiMInD2ZxRkE11lfLflM+QEJFAxdEqsHhkdyZv0xfkNatEZvAJGy8BJebdr/rgXQX9GFeaT
gdBmZz8yKkaxiwHSGbgo8Y/y9q0iCV8EcIVwjkak9BpkrVEJVhXdXv1vpgb2Vkf4KQChrATXk6dY
IgupGnPr9aVlcLuBiYTz93V8H0yjRDm2keYLOVSc1heHVW6WH5w1CFDvECktSroek/PRcxIhvSGt
WuFHDqsvmMbdA6fl1+s9yxF5XB3v2C9Kq7Bo5Wc0/RB7giyBKm6pTm9azAu6SbFHXqmxP0gAGl7A
a6XDN2eslfmIJJtPY9v6Mrs2FvibC8oCEISIGrik2qyOOB0gFjrb/URAcvNym/ZhZ6cWjQsTOAmU
dWnHpb0IH33RGqjRgnS8LmqooHeVGa0IhuWAp/fDhZvdpUazxpDG4+dOAtonF3XHJojLlsjDWCnK
t97315HT64CaJ/FyJT3CiwcaMoau3cNb7vi8KgJB5k8B6egNjp7sJ4k/9NiVlLRsKJjAd/tWOpJ9
S2XfSKR868jExTOZ8osJjL7K2VUftIkftlJVXB2qiXZFrGp7IVFrKJ7JEbQHedBP4zs8LrJmCfgG
2RI5up6x67PLHNx5OfJRRmaiZsug4x9wEjI4uawSfMtkR73RNDLfKFDkfHl6PI744Npeaev1fseI
YhS8Ikk2hr3UqvdySdHc5vIWXJqSQqY6HqUJjDyuGhvI8+9/bjJ5vVQVRJWYPoWj85uBAn9kZ3l9
XpPBEfZR6q3B7YiAvgCUaNDmhD2KvSC9wwa2Z4wKbsCbYLLCsIx2TKwp6h/JU3F3KLoc3HtHwDEQ
ASWZosTSxtYGf5i5MpBzoqoq2cXHpJyLbIGFDusDPT77cEvtCYjHB+MNk/lK0U0HFmJOrXLb6BPw
rcYfyXo2aCemNGuoHAhE4AQL1cwLEZWjF9pLi6woxXe/X/F1iV2U99sHT1btnhnJw0RDuKinGq+L
MZoQK5dgk2lv5BoSj7zvU2QYEaJ0Yv6MJtHjUtKFMN6BnUtxj+2Vi0eOPJD7iiQ7HNOymmg9Cif0
xA9t9Pc3o13fNpzPk/D66Kt3KhwpDHz1BF0jYrlOjWf4pLva48izv4c14FSIK91BHj6JPN0hxxCV
QzrfAXKSBifYm083LtixfKv+L0EfMthMnNi3Ttr4kTvj/9iTA+ODmenn3TUpLRBLsecHqp30/87P
CsKmF3OMU3kLK/gYcoogjZkDlF3bk7pfmqMkj8AuXpGNAzPmeMBJKaO05EpCp2Sg5OBOgC2QJ9xO
9terEX08ijzHKZWp0uWdZx2aKlYxoC27RrxxxnlZJUFS9+af17kUF1zOSo8DB05UP5Z8g6CuKEqZ
qqTMZ2VCt8AmVDXORnAbMvzn9lj77n9JFxJRxF+m0m1uQFUWRHSX5RmeniNHYUvUrWUw8Ts4YJz2
zWZPpmjTkkfbwE7hq+yOGzKWDxNXjpdA6ye4z69uAUnlFoWi2BfoHVX5uuO8Xk1SR/MdX2gb+ouf
6DTkE5gaTfx0yLy4jRPooeJWtgHBTeozzmj+bvOkz+6DTyLnoebzz9bcKuKzwEFvrkYzG8BtqQkT
xA6lP86iQY8iAzdWpWjmWZVw7QwZ7qlyN+yOgf9r3Y1KVIWzQSXyn2MNxKyKKk2p+3mBWeC0+ZjN
1/rm+cPtnWXNk6cqxO9LtX/djoqxKcYSxY8wOZlTHtgrj6jQQq44fYcoQzN8FNkL4NqgEVuLm+Ng
PeOg1PJpvTSrz5Oha/9DX3wHvsF1Oi0R6cgO6bLj9mhxq9nb3NeVirr3lNtodpQd1G5vQUb/AcqU
hyGO0DCyRFoXiRKDMKhOuWwUSGt0rXJC7u4j2UykE7h1UlCdCgqUGC40+s0tB9moGWziby73mz+Q
lfACwBZeAxK5PhDFHPmLCfjXSFApP1B4VSilfDq5pDr3CFEusXv+ioJN33oM/wlpps3DYNtsXZDr
XGXGyDr9/ISAtK+3PyvJEXFiAZGRcs66Cspt4P2uMDdfUBZbWUSGodx1pUeT6fB/12wBIOqeM4xk
yenBJtc8mmcpViKxuCWFxodNYhX/EY4jEKTy39XRmFGqH7HQuHCW/4AaDWyfQAlEbXXGK5a3jLhK
V+vajcHJF0K7ybC3LRV6Fxs5FbUO6eF8sZOLj+AJ96UonNyGN3vr7alI/PovJaKF4lSAe7tpnMn8
s7Y9WsK5BHddKUCA0/n+f+qvyfV8Y7iSfWEgVrJwLnI43C9u+hH2JP6KVpfmNXaNkGidSBM791XF
0VFxHgJmznBexrXBq4cwJhYQvnBW1y1J8f+Wr/QUQ5VfHwYFLHn5y+O06cd5qxZiANpL16UISDKx
DSuBOSX6CE3ZFNoTbrJZwoIBvT1ccjZA/JHOdO9zBERUJbJrIt85kEQrpWfToE2cFo2nCeJ6YNmT
t3P0VvSqLIs1jdKI2FY511Vs+c9mmF5yiL9AzlFnQdtU4WFIfgf+x2odvt7/dS5BH9crnb/UP7eR
PLefE9yNZiXPH/bjLRZToOkjzIyWwJyPPlfusY497TYyCa33W8GJy5jt84iPG7s4Gow+JeTT7pOz
88/uGZugyaT503dXsAJixtNkKEc4eyh+1uk4Gn4pC86iZ1nzvw9kMWCojcYVuoLHZLtUvJ07OgMd
AAD7uUf4/BGbOw1qC3zHvDmt2qrASF5b+OnJcqE3mTx4Chw0mL//TOk/or0fiwsEZemCYodG8eaO
QlYZW5cpEopO6U5dKcdemjOzEQQ4ymkjnGWyLH+5RIon+vehHK9KeAAjDo3xOpx2Nv/q818hde8u
R4CQ7UKlV/hfM6ymFadlb4fqYNS1+1/nvPb1oYL4o74JrUDyym3cmyFn1ShiL9V1Wkr/mmqWexq0
zblROgGxwXHqjw7cZT3Kc7LH5SAeT6+hkYNYdD/u6FM/ktUbmsZB3D9liVi5VrGgRxUy4lu/PGYL
egRp0fEavFi/QLJDXDS9LFcvFmIKZp7DDueJ8xw41mXDgDNZ5Tpj2Qg0ANRYiqKRYp/0zoKkhzhl
wUUHtAPHSwRrf+Tp8q0cxNFp2yU1lDjmzMBWbMzZmlrpS+dsznSUOH3FaFkBfYkikkDyPAXhf/V+
SYucXKnnPA3/Tb8QQx9aOzhecLbp10cEd3U4O7O8nWKMmv6nmETlme+qZE+JxeCrqAJeUD4OrU0l
Lu4x3putYFsD2VhPyQkLANuQXQ41vBw5eFz/riRS89fGxz/7WVri1VM5/YpnX9a89MnVlvNCgqTF
MrJp/In9LF9EYm0LgLSVfw3hAoTMeuDnH+rcaXQSSBnRaIjmFJMKR7hk+kT31qe2pQUlZwUJVO5y
SX+vWTNWEhPYvraLpQ/gSVfqO558/QiQ1bU1aYiY0cylisgP7xwu2VueO09jpv0V+geJNo9LbgXb
DSl0Y3M/3QlL2aM/P3JwTyFw0MiV7BPq/HAkv9ALzm/9M8yWywv1qoRFR9/W6PjgZrcqYB2lLBTI
qjFwHwFMPzx8PseobkQb847Q3fKQPZkfU2D/lrUJtaym6CUNCOJ8PlJxvBEfu/Kd1a2TEEGzzLOa
QjlxcC20+VQg0kX13AlVP3bHinSnr/zDPvdJ9tRnZI2KG6giz9wvTQZA4EPCBInarKjrutduiVCa
SL2CbxcCVag8b1p2G93zPQ4W9kDkusN6XzJgqJcCeQkqLbXY5fGngnFTJx235bikzUxGwGBK8Z7S
dc+VMh4bh7xWCE7LHjANukJkU4oAhmmsjqTfJ9GlXmRgBUBYd3s93dPoENelXCjXmg1nHZ8m7fxt
buzhCr3zL2QkN7KwpXGim0b0NwkkGyNnQA2aJYZimLd4n2vjlGn8YbpQWhiIHXHZJ8QG/hCjkzSz
tWqW/UCejOnY3nqF9nhNWXksejb/Tt3IMWjVQm3s3NA1epbj4TXD48o+fJPfNbcCBqwDycSknj+Z
fpuL/D+D+pAX4t+aWPvh9lrpTWyZA27shvL6MG5VocQmTgAQpcsv6DyaJHiR6AkAhN/9zTZN+QpE
22jKjYG65ObEGTOR9iyneJvBvGGzK0gjZF4ZruP2p0X7Wu8iFXmhn+k8RWpeIlOcnTKgFUa3xJ96
kSZ1ozVbUsxhITVcRx4OqMZG/8ABI8ke2m7c7QoE6zWNngCH9JNMU5ETPvg7VzKeGlwwHcPvlrH4
50HUsKyvK6uh9VAcQAYAzSOu3PFB7hlEqkVwgmu2wI2gsILdtpIJKnY00FFQxybJ+WAO+S1aMQHa
vKRIP3bzgDa7gyqth+E8Vp+SFFoy0Qe4OMrjmDiVZhv/I9tVg/PNv8d+kYi9lywiE4YrRlzNctP1
aJavEA6nZuJVSxJhkf7+FarANimrRrtGkVYhKHUj1Xq69kG0QbUgm/05L7Qb9MZVaxXda6K/4QAG
PP/vBg3anL6tbsUwlLAA+OCtk46VAriOR9D3g4ls579KduyrDFEFn8GiZTluC2MAqkQ5lFRULgDJ
v9fxTtjmp58phR3//tRlCCcbBr/3c2xWXayuXovdMzoE8i4wx+nyTs0DWS7YandzIFA/sMPjfxCc
WOdbmRfhuU0UhxKD6Be2p6tDgiL+t0oqpmp1zCN+KXGRWuPvYnv0zLX4TrewWvjc6cEF4oZ/oNRu
Pqy15iuica1agmiqvChJKMM95Q1/uK3+E3O38GdDexY0BXF8oUcofMcdWikIP/AzgAyz8mUkHwcZ
tWCruo1sBkCgSZK1Luqz6J3TF8T7RKyyPrdMD3Ahlh4C8XMlNdWRLDaOlg3YybNO9c/mEtDkis7o
+CbumyHe04us2/HAVpLHF6KCZMGpEO3JJ0UBJe95UhOVNkoqphHGmdbKEWAPMFLAvykHdNb7YNXg
QkBhDdaXvZn+GWlJ9eFuj786w97g8h0awOnYu7ND6JRUuBl8Z6DXBMdp88spBQKzpUvnr4xPVglU
L7THww4yDhzJyDgWGosdtkrnx0fk9hNb91Cey4cso7bvGlS3DucOOi4p0r/YCK2+w58jMUcZBKX0
PUl/X9ahnpN9JrR6o8N4iueZrCMdflxEUiqbyIxlpWZG1rUgIv/mC7F0S5/iS7Q8GxrsFXxBxi8c
4FsB6LU+HPG1GMCwiIH7E+gzoa7s89VY6nfeuzBMtKZbfwcXHGHdrCQlSL27SRsEFYcagConJOEM
TVy/+ibCL7Y3VFfU4cIKXZNkDgXwcvbUdC8qXc2/uvXSeta1qYg12Z4YzGpz+k3b3wC0LOyPDJg6
ECcxygSFCQfQ5yL92ahHgMBojRq/ttUeZX/rdtYqubwXAGdm9UXhBxZpJM3qy8fWAID5KEf5vru7
KUyAzs6hugMkkpIkbQpubrKFhmwAKIWyXLKend01Ht515WsRzSUtvEwXBp/pJVZxgeoS8GvahrGu
qd9aSfuTYN4ayLXff/NDgETySQXGEmGnfnR7iYlQ17PhQxBDoQ/es4MzhwWyeSfewYTC6fC8JBqG
ddUr8JrvNwjQRQZEikT4udef7vQAGYYVkBkknJeUwDsZsXPF2qdKOBTfsqcqymI7eRzcd9BnjFDP
EdZ8xicNqAGl1qRTFAcZ36HJxsiGEl8v8xgJ1DYGIKev4DjEQnRv9754+ZZdyxhgtG2ljAyLQrkx
qx9TFxlEQFOIr9fraokPyZyuVLSBbSnVTKGUgTCPUqaJLUnP9yja8amQBz11fPj6ZkYRzfd06Jiy
Bf9WlqXUKVt0vZospKBjp8khldSAXHZ2TGwk3SelDGX8TGYIHL+8Oz9ReFZbQ70YzSb/7mZn52rE
i7/MGBcWPEaEQcn4xk7XrFMxLzt0STBMD61wosIOztspTj1AxHQ5COd8leKv7Ktxcwskjqn4HbKI
5TrIs+7zqvUn2oG7ODBzXrfSDjfxVWWsVzPJa0Ergrw2FtXe4cYIjllA4dgZNst8CqprlCC0/N+c
v7oNtX/nEiOu/UQLTVfWlu4eOIMonirv84PU6f8yoZYZHX0RgE0X+hSSn3QkUPb//pBNDZYMaRRc
g6/XwDXairKqwT+FOGnSXF/v30ULCNWGDPj2YxKEBmIdLCd0G3eBqnRystB0fg5runKLIAiIxazu
TIRnGtypeyB95I1vkDH0RIaLHYBZCW+SRX1di5x2yHE7Abo8XI+31d8911P2JGVcCSr6YGnrgJJm
h01cb9vx7CzWh67IxO5j6m73zwduuNWOF3CvT0KNKU3l0ixG3cmKD/RlnZQZOf+YC+/cA7A8TTnP
wM1wNHeoTDoJuRc/pBlVo28buuAuY2xmW7FKSzELCge2OCo6RT6uK7msRu4XchvW4jOKQdssL2Hk
TUoyC91iIRDkADMTrfeuTCpiyzJL9pfgoFwr0I+tAVksF+X7RojpPS71Usx3JzE/oPBrG9Y2AO4x
xmACCshS6BinlWbXvo1CSxNvl8TCRyTZgEqfDcPVJCS+H61IoFjXocQCtWKiS+UBU8QGNjv14PyT
QKDnWvwr6An8NIAi+A2gPoNvYMq5TQvJvsBwLPqbzu77UHoSpHaWmojGvZw8wXs9P9i5mAywiwrG
BnvZpjQq8/DgG+FhTTuypsPK3IM5bNVdIDbdDNtkkpaTXZkAgtT26t6sMw5gTAZMTDXUlghaJKaJ
SRFjJybT03jvq5D85F+6kK/JDCul6t/y4AZXdPjtBQRRgVitCfeLFvMBquh75qloMBrgdeNir70O
3liCu9HmF27YFowYT7UWsFUq0yxMuHiQe1kKcZ+8/Gs5pGSHrREefeJlEr7WSENIBvwBkur6t3vE
oIXBZSIVMnIGFa1sxAXEQWbdmvL9laY7p+v07qW3CVJBFaLSC+za8upxxRyTCZYQwpxfPj9CIwlU
jXrZMHxPbj1n9s6cev1hAemueMw5NDzII83wOb4YAHH9P6woK3SRxSa+EGDBWDB+yLJRPCuIpbSg
3Z30dcI7BzbmaRfY0E9lFQDYFWKO0rIB3nZzKNJmdpknwJPXkMVKXauVOK6KJwAqI5keHWoCV+RK
ZUMzZ64IMNh//j22wHLRYBfX5PzZHddR2sOeyAtYC3BmO58WmZnoYYepXsqAzLiPQpyKCzdNkjyY
UI+Dm/WSF4mlLPjUpW28RmkpjjXBOQHlHBd8pb4E9kzd7XrLC0Iv0XNFvv1HldlSSiFWRYNl9YR/
ZXGGpD4faOagr4UgRQyWsEq5eIBB8qldOENE9mM9lL8uABjelmLZAHZo0MIV5cVDVFyGsv82xXZ4
475qwRPbo0o50muJQ8aDSfMOSlKbSTax51L46PxWfRllzvPF6CHm+CU4lJuUoPSkzbs4IjorvK+E
aHuunKkyRT4xf/cH6twrYd2BXwGcvvJ1vJ+WIBZ830ECli7dIHenyL6Zr2D8Gh7IZXWx9X6/aYuH
bNgM0HdApuMNSCDdalOj64/ENgymv/nA/VtyeJpkWRYgAeMFx8x5pyuYTWYm3LeqM5978OdzYT50
DI9PDztxaBQ9Dn5oubK2UsuYnu1Pl4MJ5WMm1329KpLEMfU3y4jzrHLfXwqGwvh189n8X/FjANDH
ow8jTA3Ge8EzeyOZjHR1Mqa24UZ6Rs3ykSz5GfsJnFkaQW/7zHWyjjLF9UlxbpCDcZ+HHU2936Oh
D71A/pKT1SKgK6XaasBB2hHecWbpw1Puxu1oud4ENsHuVSp2wuVenrqyV/QAvjpN2bKJIgmASfZv
qTAApHw+F2E63gOIZXKt54yHzg99clwXCS/4WwTWa2Ht45iqeBGdrFZagthUKD/NCcCvf+NTb/ZH
IofZjaHPmYeCHFm/VTY5lUN7X0biAbS+B556/gXcWgAh+eDtOLU5PpaxLV0oFMHcKFv+XY3T0t8g
oI7jYmjEQIO+NYHH0qU9JBL+vRbd9VP2e9bSlLpwDFGiOwj1Utmq5DgEjehu3y8vepYefrrfPE7i
vfbq6XYZkrKBksQ22wC7Ero7kO5jm0EySyKW8q7+amBLj0adE2iMGHR488fJmYGujF1ijWdqNaJa
mJkKBpzFi6wvTcEHA8a1wxG5Mpg6xZJJOsz8s0lzaMMD9DVBViOJLmrb7+0N6unexb87oCSuaYvd
xyaoMb7hJlTx2MbY5J6u4tZJSRQf6wt9lpEOsmUBHItFhVzOM2DAHZVlrMv9h36uFTcOl+Y27GpA
4uyM+ZUeEa8C8IAxl2DRlTA4rmUMHtfqRbz+Zq9mf33/6gzglakzJMSY2vIKk5Qwpv5e3OVnFEHf
Brv6sM6/uCAf7otwXtnW6cSPAsfMIbO1johk9xTzySdIlA2zTPVZEq/O8RCqH5BCTk9NMR1Pa1sC
EzAkEx0+Azb7mu4Q7Hxn9EqsUy8SmXtx0SVRcK0W427jYKzEIrmOtRS3TguJuewSUL9x7NTjcpov
ZdxGAGvIpjTBlgFG7pG7a1LhHY6JZPceJHV9Xyy5fScbNdQqtpI7jPsz5yuOAk2MOYHLu6+pnv6a
9EGDH3cJrHx1TNlv9gQRqDrtqUaueQTQI4Co4i6wNZm69XOf4FiX9IBzqXkqSB9sJLkywzOTaE2j
6mSxrFuu3fpYhlOKHlOUI3lXnSFAQrTX5fOlbHicbxyEU5aS0H0uVO7wIfZhQc2SvDfxMQjqQlH0
e8qRzJIsBtUwu3zxFQJHB95LNf079ITq6XvFOpplW4f4Q/qORs/blKtOFf8nFzzcFLBBmmaaNHGd
9Kzhsk5enLH0tL+6zPSDFJ/tIDT7qPJXyCTNiC9TbJDbrh7rdvOFjr1bmA4p2hB8wuhlRlq+HxRz
Wn+kLdpGNOKYBSqhpeAH/MyyFfXTt+QYp0roTw7g23z792qu4ercEMuPr18Mx3MlSrQvoKvbsWOT
hGqX5T56aitY9Ko7YU8ato79Jd2zay0CUhN1YEBKNFANR0VWfxWt9gDACsbEseZUQwKFyi27vj1C
NCEw916FppdcYkG1ZAs0Do/dD4ITIgIMBMFx040GIpHXcZMk0WjzwqS52S+odcHKBTveUIcaBdBF
f/ERzhRtZT0xxyygxgF4FmEv52ydpzZJx4GI/+GYiFesxqyAt++JPEQ8vY05jbcZbffjCqQxotUB
lL0CwpsRuAb/iLUePYZEtGzLNHsTijR1PZPwJ8OXMkxOoH0GsvkO/CP7ppv9Wa7W/ZByNRufVt/4
hmDw4ynIfqVgDeLAZaxC28Gm0491LGUM7eFEPYTvg2Cmzp75lPE3pB82D/V8BQRlztNvIElm5awc
WlzOGW8+76cm9n/SlhP4fR6XlWv/q8SpRm2FPhtwhUfBpmFcPRTpSZtCRFYSeLUDLZM/77zSwPaJ
6Pe7/C9vIriXMzlsoeLGLJW8QUqP/oLWcQTwQZMa0R+BxOrfTe0FGOkyVIMSentUJBqPwgNdp0j3
W1uYfadUJRfNh2pMEY0nr6ubGGtVosiXOq9axxm07AA0wk71w8Cw/4mMZv1y3HBIjwwfz2KX8en0
SlZ6NCXsULoyeuefsHq/3Ye/1xbDUEMnWfouely+5q7aXjx0AoePO8ye+F4pYPPIcVXIBVKCDS5y
58CQHeyXBAFNo2Nc3U1ZrxwCdy2V9QEBExHagSXm1wpstQ1IhEB1K3JcOvY8ylEzScTdQ3csy3uK
/Df0pYRokWXV891l3nNXsBGnnuJnNOKISnaBEKNvLgOtG/AOKeBVi8fzsHsRnv4ciXLF0OfPLUif
NIpx+50W/sTg1pAShtUSYyJZnd5nJZG9ueibc0teF052/CoAkRWGLz9aF6eTk4Gxn7YiJGaUVNU2
7g/eJFw2ntESqmSy06UanbLO6H0U+0ypF4XGp9dKH0AOSmPKO5D/yEzvDQT7Q+MfaD8+4pM4P3kK
weEv9r/Aul26bvDqkT8y/ur1XamiQTkvgmylCBEovZY//Bn+RjeO2ucH4Q8i7OYmQkCiYNaduhp+
GAeVW5x4YYALPJS8gyVsM6HpY78Ft8GPumJ1fS+g9RB7NC7xVZjaSbanpIzroPSWejPIvsB63AYI
mq4RUSYRWTtDy9vDgCHzVuhb5VFKDVgySHCVF1c2vqUDHX3EOc3I44icM/XsSVRXsnGkHGTthndx
Fog0tUUT89+SZLVHn8mLt3y6yAmpKCfH8l1VCJuWozZx+TBKffEwPKdhiAZ5Q1o8hJOpGzwvB8PT
vBxzt6alVo3AFHNcZWo7GPz1AYedF5SezCjI3vukLxDg77T6p8UfjoCtdZiXKhUjbuCEqV7ELUy9
QIB3wHg81oZwiENhHE9vqeuXG8QsDFkqDynbuKGjfvVtH3TcStwCFPXRtHx5FbArAvAYQVkHJXbf
KNYoFanQNZRfD+6Ndd6xcboHeEl/j7CaFy6NxKsMLPeyOvF+iiDmtRX7rhSKuWcvVLXuPgEKxDxB
eGlcN1qXyziR3nhCYh/LkYy3GykzHlCIibgw+k3G2WNsYDIM+n0ZbIBfLsac2g35IT4IObHKsFFK
msZeUdqNYgpb4IBXZoFEjpQ+EfHJIe5NJx64UUhtZXn5T6nLvpvj4Z5IWvjDD8bu8m021C7aoY+d
l45DDIN5y7ESjF7ke6o+3UG8dITHm3Ne7/FUWyHmREl4DQRD4F7me8rfMmbVJoPtHfoXFHOEcxUg
WhoG2rR0SR+RU1zppmiJQB4BGOxIFLCrYR402kux9jNhToeQN7Z+y9c7c58bZ64XLdoHXz80tBqw
hhGS7tJoFflGP3naqzy+14gpSPU7xQ5IlC7pj86tsCWeII3BWXG6a18wPNmkaiOMUez+846YU5bF
bkKjJRTHmW1KwbttmktYLecUpa1Ry9+62pP5l7pvcSuJj0ENC2R2EBN5/KjMYdek0+80/12X9IAP
NtSIWd3Pcsgo92aYrA/sRwJeCcT0mQPKMbV8W555t1HoMcXc9OjqobEfKBS6esyN+jSf7hQhFiQK
vgsSmqFI5Iy3RuXCo+uOJCN9LjLDsfLp5hQ42nviBE3pyDuC2XGaJNHiCAjg3x20BvNHFe9tJu8r
t8KjTQtSOvds6Dbnj1fkl94aSeBch3y1reN2OOO9sYYeZHVNoQywGvFDwF3Y9dZL7DuJnYt1/8z6
4m9polKu6NuMD5DgFjWXoGb2DnA3VQxIrfXi6awMdnX3ZSP3OWyEWYn6MlnbD6XThM0z43IIODAJ
x5oCB0KVGav/g28ot4h+6gAz5TEFnleO1GDjW+0i6SWwniK8NGPlPh2+bVbmmhpPblj2V6qDW5OE
8ZsUgDMRHtYUtiF+R+owN50hyA6KsSekCgpNwKVS05lkbKR+kFCvMzY63mc9svo9rbGRzkCs+mSh
XMElEdEa8KAhbhE3vuXQPJcb36Z+tUKoQuFLG/YfAyg51VfiqPhnn5jJPrxs+SGHWiDpdKDOo64z
8mPSW/sLN692Gwk5agDt9JXvo6xssDiPYRVCxX/POn4tmU+hy4gesoC+FPDw45sUNyB6jjlV2FYI
NVTgsPOn41HAWROXmWZVNipqbhik51qwNH8uTbCrlcJQzKTYbSRqfwuJCLMmtxUoHTcfBH+jZKuB
AEex7mPXZ60RbIbZmim5EpL9JF4LwJIpiHmCzYQjzGwWOW/9xTgV452NUQ0R1vrnvRYDhmabydFb
P9RpU0YNxZDZMzjSMCTbIYqNn10ySPsvNRNgRjV4z1yT1y/r7nHKX2HxE+3zZiGn+klHVEXpZCPF
b15ZtX/uGPCzP7KjFPZqwLPw+qn49FWvn2UzBrLNW8RubVPcqVQ1+1aKTB5EG1pIai++Dd8HRNbo
uO3TWwIfQyxUNQEJqkV2RDgMPS7VlFAcvO2Ki9FfFBQrixLQiw7UnwMogrXInvdZADbtcAL0lS8+
vvbeZNVhqlVdrrSm5Htu4Ebc9/uqIo89lkcZTGiloB3YOdL3a4YUvc1rHdT58A2ozj6PfHC5v1Du
wJ1ixizYMgHnrRn25u3W69a6eLTnqAe3CcTrJU2j/2hvrdSnb04dwfnCiDGmmmSrVXk63RybrTyJ
IRR1NCDBtObBFgxUiK6FmkQtZKcwOxGLFQFBgn/gv4L1O3YxuofuSQUj0ZFUnXhVc2xEUFAGYhTT
EFy4MYTad/KJw2ZwxB39pZZOkbN0CmNG5kOiAZPaDF6DHQpkzI3wSCJpej4EA/gXyclbuI7LMxUi
WJ9NkSyXJjIKEz8QCnrCSI1lBvvTTlcUwv7SwK/CfT4NzR4zZNiz79ZADLYdpgWJU3nc2RTrg8bv
RAzZ4oDqrY0AQ+0xtvFedhmJGkxaSejrJ74E2GANQnzfaMOP5QMtb//T8E2lK6oHqVyHds9v9oZQ
4VXWPpODMpZI0DV4QWbMOO2p8pen8iMt3Wcv2PdYxtPBq3VIefEk8TfsjUzW5baMFMla3NXdWc2h
Q1IJE0vpxgau27r6mEr+fi3rC8/LZrBDn7jZXCiDC0GODBY8AKWrIpXp2Y0gNyJ2Sj0uu43LN2+Y
eOAa/YmonNg25Md+4cP44mNliFzpzL41IEd+eMDtipuzessfQ3iCDuFaRA9/wE9j5LGzx1bTUV9Z
YIYWRQdOVbUBufWxHTpeX7duUHWYAbpHDsmjz3Zj+fLFij8jPOz/jtI7D3rbToKriYsBrwbdMeTU
UrfbyuuWuMNjBhh+sLL9DaUxXj/mYnc6JFlpfWDC/4S0E6et2OIK1cjmxOGnMaTVBNHM8re2luFb
76O/mcQVpvGCV/X7tptI9tUy9BJ9PfEHHOrpCVMHwvHJxNKTHcGOX6WnQ9jhh4UvoeT6zKPmLCYN
1nP2971TTlXWuSf3ZPY3AONHyRLkfn96v2ww0FDkPM6gTbxEhFZ56mLw+BFpT5J0Vsp8hKfH0/vE
AaX9/yWYM1+Ln14MVuvbv4mgzrzHWX5ItwAfN6hwzl3XmyozYOLnZSeMGV7ukmj8mMbKGDoG1qTD
uFSPK6qgGdiM1l5zk+o1sc4wgXy6GhZSAG3sS0jBP9vDyqmLKnQerJHLOaS89W3N/R9h+sdlJWxF
Yk/cNpu+J+lqmPZ2pUtlkYknDOj4ofJl+marcVJfzbJBBc708M1Bvneh6EXKnsDHhcNohh2zcThi
BMAl9ax89/QDhimfW+lp18cl1LGUtx+y7vDNZLuvqh9/ogf2AzLbRuoQfvzvh8ngOc3E5UhRvkFy
T9suqaJBsO5eMCnzB5Tun78Gc/VbeKTBU/AqZbpIR14XckQmZ1bOmoWw3AT6vHWqopAWfvuBDu+K
3L/wr0QnDa2n4NM3pd6ci+VzOGPncVQhXC7IEi5SUyZzdJEX1d+jOht4BtISV1FWUsLBpsM/f6/n
IeGI6QumxrA95BGshP26B6bvh4dHbaFqk/VF9RIqolK0MiN5IbB9oY/5CZUMjYrVm2nDBfoxMd6S
WKjFcgPnuqj8TCA0TL9WhSATIXlnz70p2ejJJVV8z76J6TcpNffo2l3FI5ecd9rs17gOLDc/eCu0
sDgoO1YjJaVNA1HaapB9XfW7GV43YhqIYu6BEoLa76X+N/kAGUSDDgikWD5K7T1E9s1coCN0xWvn
cFFY1pZlfyHFhaOv6V99CHUCFNWKPausJOYEvPyvKqkLOzMywCNo+jKkK/9+Tng1iV29yHRQzsk1
I8WeoSsVhsSDANg2dUprnz/fSMHYFuoQ1cUdDFhr9KVs5EItwwIe1U9F96JGQzqXHGTuV0xvVXC3
Z5gLwWZumNg+4Qil+WGr2K49CcRaP95f8ZHtJwV8cX3W4R2TlRj/iRdWtF5czwixXV3SN/Out2dp
iZRVY9qLOGGG8bcza6YC1fgGj19MCUg+kBz6BCBq7p7yf4ZiS+ldDU2hvCVae6VJC538Q94GhrRM
VG5tXmk1czvrFyUJrb4w7wnHLPqjoXr7vnjXu6uxrMxGmfSdY7KquPnY17jY8haJSX4eRhIdaSBB
wxmQBSeglvSQ1Agi1xRx0l42BY/vbALPzIXy4zLq+AEw6rJllXhfL1jjn/iViVkn9cXNw2NHCQxQ
DrwfqdGjkWaUBLHSfhMS9pK+hdaaegn65QAgxKG8Cy8Qvo4EoOynvlDLsdO5+Rgsh3pkrYzkMvwO
neBpqE8VMctcvRZ3y8hQPKSU7ob8wHt+EM7lzZbvWsjoOGSmtVusAsZC89rFAW0V7fOJB2v6BlNt
D4azCgJCXyzShdBezl8Ug/oeKX6FfAE8rqIN5LcrcUH/6iNs0RX/+Nr7nLk992OtB0y501IzF9bQ
TR4z/h46RDOL/BbbSxTvW3lLUG7BlnTIFPzn9B/TJWsDBnDH2eL16KURvkOPE5YT3pqah2TA0c23
2jKZK4b2QhYS4DXeGUDSDvhSNePM+WkfjkkoE5937hhG2y4d4FYpn+tBDuO1r5yFgxnOyQtKW2f/
C8RH0yaAeb3Q5Z6XpooBpwtGLCudRfv8Me+e6DxGjsZF9WkD4/TpaFz1l3RbNzsExd5s2nLgsBgC
bAh8N2/Jgh4V4r+lvXH20mLqHmo3h/zPn25gyRFNxWMyqbD5WGeTOtqKCJ9jXohV+5RdtLoUnIiq
p0z7sKaLXzZscYkL8Z44lkmshsv/+zaVSn7X1q6aDCcqKlMshy06vC0qyQcqrRFuSCcXU5fVCs+/
p2/BO+1h6/gjDgvatSSNtXd+9wmxjis3cqbHRQEMlNUDKGpc1sCTOncbUlVQJVSoUaXUBwlF/gzo
6+amllR34LSEeoGI5PARpMwuYZs9lunvPjnJDMc7zOont4Wo6Uvt8DSzcwCoFCcGAyOTEp87xca2
N4/PdLSBP+cIipLHhKY+zTJPnKH49n+ay3zM1kj1wQivEu+rh6i8ljMpXt8MaL4UVqYGiPwb2YfV
FGspoLNqUx6vKUJFP/oFZkJ41ihXs6+JFM+qKP7EiTJHhLVO2fLrtMNdQtzx/2m+lbaVjDmUHWHd
m1MW9xmTnOpw17KzAvswPcGQy+F9NwdkI95aRG57OClGEloSAlGjIu4VFmMSJonyY/ZVczzXFKBu
bcTnpt2r5gFxLiqRmIsHyZqc8CWXqQc+C5Ca5aA9z9nADgI8uwLu0ld4V6YMQTW9cbincQH6gzvv
bg7xB3xtrBa7chFomsGLslWLHp5F6X7tayMP/SaWEZHrJHn//2jhnClaehPbbVGdo16ySWAWuMMR
xbTHyoedkC8nVksSwUSAHHg6mGNGhdszOwcHmm8rC1+rr1B90KYLZlNLMYMD3FIkHVjVxDuaXKwO
X/JJqIm2l9lFdLTYH5EeoCOadtIDqPp4CctWAfqeIX1rzeomXWUUnevNCoBU0eFLzkYh1lkePwaW
YgL0T4RGVWdZWfE/5pmbWjDGRybNjqaAfkx7fLYd/kwtfRKueCBy0T/4EFBtwML1okWDssVnxgoG
ODy6W9Zo7GrINROMz35JC5VN6VYa4PGGS7858iqDPfj8mpEbrRdqYNAYUBn0kc9UIJgmkJh3BW/X
75o9m7+/wibbsR0944hf0r3YuVDQifhB98L0OdwAnz69TOz1eiUxhEac6SV7qCQDubOYSrnt2ZpT
Rk4tfZuvXxCrT1UT6rilleA6HEa/0sEz+swd946HmS6rbb1jDhdm78Jyd6Wkgl/LEtuz5xc60P9E
QC2uqd3jyfpiZ+XTAXFLMBZnG1hR/fBMR2jGurllLVDPAeEr+Dc9RBfjqYI21ST36o9MfNfJRcHA
KoMxezpSgvwm46VcKtTkyvToillGY6qLiNXjWSXyZUbBR68KNAmDWUey4ruEUbjw4s2/hN9hb5Dm
w9oCRrtzyQIZsvzgQseGF2A4sKHPzV66OG9QnoFxBu80jq4fK2H0I9zZrzck6IPr73PzrxCqhHNw
DAhlsesT/UCjDXRXYxgUIDCTOoXfoD6HbrqmQZLgE3oZmrgBg/hxhFJN/HN5UfKYAAlaCAz8gFCW
Bp+W0HRa+dirnVSevUeHMzanEdj2RvbVROtgIQsC4lCQ1nywZov+NQJDBExmk4KUY0an1l+1kyB5
xFX1HW2RsJPUPcPr/KreRi/KgJUzBkyCXNLvGSbWDp8oi2J1OY2iMeIaEDpIX1ucDoQplz3uYloY
HPtJahbEUawSPPAPs3N4ma/Zet/0HBbe2Yof3W1VW0Shi2ANisQxSHt7V7nF4tt5oeJeFhiIvlYO
x27wkJ+I23lGdZi4AS7mJGe6EXdq0BcWPAKQMfNCQQFfWuh+NNa+XdCYPeA3swzuzUIoT2tQmQOm
zH0Kvah1q/8VP9KTKZ2Y3VRjJgFEwRetmWwkRoHjIsmIkKsjkN67HVUOh9WqV3r1BAXOa2AiMy7b
D03uiLS3V3u7HKBkEAASe1yjb85Ks23CosYKCX6cZffP/0bFbPWkHbgD/QN2uw2iPnIpJqOv9FCB
E0Ll2ymxvhF1Atufah9FiAn/VKCWUDnw2yFSJebkVE4PFYPsVh89tGWiU+EIroNops/ORNFoMExZ
8c5CrsRjpUZFQZ4HwiPXt6lm63+krrBfkRD7ZdDP/T99xqgNn+/zV6YBEChIRGE7eyA6zFDUT7C0
lYixJrzX1n5EG91sWY2yFm1CNQlGGKRD7Zw96JWbLBNShjytPBbqecelaCqlVu/9w6huftM7X7lG
ZzJHGBboAdam6tig4eDGq9S919S0pimPYHe8agj1un40rs3O9N8dU2awio7NWwJkyx/stEwpKWXS
6Os7TNqpjTVoa/wCuxT2IsywVwoz+PHynYzf1VKYD2K1hzuHn+yJEAiZSTlHQ0oWbqezfBirVeZE
P/EHXnLr082QyPTytDmM5F7sOupIsARXKH1SfEG+ir2V+MWOj2VaCJQQgh3cUyL1UDrrkPlXPXCh
fSMN5hgsXAOcjRAidIgas9VEMsC3kU/VVYAFsQsIIHpCq2gPiRrwbw+rnecX7DA72y/xuU9ec0Wy
/KfcKSdW8aHxpGy12NfW5+YdKrES35+DVt8dQ3Pbjra9i29jsppA0yArEQ8OI2qashYINNy77YF+
SBg4IGhboS/M8yHTZJ4LaADsIgpBw/2hFCmeYKe3HgRrRGViJ/iDoXWfoom5TyrUgIF2ccSnKYYR
zs2ovjLRgmuD/rMcFUhcNGbTtGr8C/3pMvkqQ22yEjgsstkPe2Z+wqSxs0I9zTNMTseFOmd5ZsNE
JD8RJ//GKbbJUbVUiF9k1UaNIJx4OAHdzFQOhkyS0AM+0Te/MqowwkcIhWtWqGtkfyKSUYYF2dBh
Gu7e02eLObHTawxyBXq3IZ/1gXQO+43WMB0BWqwCkyul95DN1V8K7xfMwcu+B60z0A5hRmmu5TH4
4GYYE4KSbC8uVPuvqqEl0Ts+trxpmocd6ivYLhgsVM5pp3Czxb8oNa/fWGWAX9n703bfCEgTD/7g
jMZkLlE2rbGRM3QZF04/LR3uZVydpWh+uKKL3d+eAIZiIgLcDQR7q/T+EeNEtbRHu+IoYjPSNfkv
sUouoCQliTQEa51HVA78TnDprK3IOvSZkTOYPlRsTBnhYwL+90qUVwq14pMQJgAh+fETI0HfwgoU
q2QLa87fn6SZjzO7OMMdftfgK2bu7sSSeWlaxMPUF72yR/qhLniLHUsV/2B5kCcy59s96Yw8ArFO
f0uU4iV1YBM0YK2F5rmn4p5gmG7HTfq6hUPwJTGainUZMegYJTTkxFGpzqG/Ah2469GRPVdm4H5k
CisdNzAHPkl7dQYekurkBcJMTa/7/Q9i7b8BuiuflyS9PLCxsMwK+ZKg19DPt4gyhnssKqkt81Vm
MGkW96V5SKgRnxFU+rG+cO2WrhWsSBFDip76m4rbMvwPcxKiVkG+3bsP2OGEDCKQHQG0drZt4Xrl
OVtzq6nI5Hjv9WLZYfvJi87f0g7Z8NM8/+4BaSUUH1NbqP7xsRLTQFr9B8ZMbA5P4UkYYX59eXX7
rY3ELnNmyNP2atkPkjwkzvA91UHWSK8uVnQKkiGtWRJ3al7HABNpu7dnzdmnuurV22zGnp6GXh6D
rtH1ol5XSpfqWdUIsm8kdzYFc2FZVuNALYfVsl1Ia8a+92hs75NPjJ/5VY2D+XoYLs1mx8rsTN2q
Vb2L+5bLQY6SmVQFR6Ma6MmsJ1aFkeKoQgZrkLhjkXojq/hvdouAjqsHKz0FXARTdFvjnSQco5/T
WwCjFWh3njkm6XIS+QKZP7n2ZpJl8FJv/fqz+XpZKS50WTnjJLg08D0AYhqvDE0M0YHEHz7cB+iT
1J+8lu27oGc7YSG4oHlGK1Su1iXLOrzfMhGxNrda4jbxd9BwzR1de7rJMwbPb3k3ONbufP9XYgKy
tcAQlejRFHaAbH6BOTj9C/SPWLXirCengFJMLQzthqTEd+/ei0CFNmwxTcBcBN8rPmyMlMvmwLMf
5rMy8gmVhscvGbshKGRohmsKAtzI4r/X0A37rtN7pPJaM9qLdAUsN5t1uw7I6fOi7FfDxl0S0Fws
58ekdtZ6MRFzmmrxkK/jJY+s9uED132CiJhixzSrggoPp/ApB/GQ/V0DTnfTYeqnPn/uoSzgUkRj
hDgHob7q7GdA5vTA4wpiU8C5yv8Q3vmNY4BT3y8VgGWmr582KmwjJ6diqpuatVPoYr/UMOmBsA3J
uiZdpSBNY3i04ucSe6cJhdOm1VL4FU4N76qGNoZew17f6FRGEgzYt5YXemDmLf690S8TGkTVsgw+
QbUMN+j0c/nkW4jhdGZe0rVCq3xA8LzTkas4iT/sSu7DwevZIDQM8PARL880cTia+zT8jsAE1vLY
0jt6Z5iCDGhASchJ63UQssTPNSIPAAvjYdeNheBEXPSigjsE+HE7MbU05XbL2inHL9+8Tftw7aKy
j8v0iPrUXvcljFQuhh+UzC9w+tDXbDFx5cy8r4Ihub6NWbHHxrovcmShsvpiiEygf0pAk6dE4Wnr
RWZscZjC44ObCBxpCeiIVJu7bbAphcYGXY374qe2gAgFz7uji3Jn6i1fPlghmwuw7miSC9tTXI9G
8n+0UqFIEq99zrfj+7U/XSJJvnRd+GPV78oyB2Lg25shqYcxFnmr1Bxa20HRcwvGs1TnZu2nD4Eb
oKKloul4StVFrpZQ+PJChlHOJPaeSe/sU/BK461Dv3l3VaDIn7yMa/auJikaysRdnnwcgotxSLgv
u3F0QyYNi8lUHlVN41AOaDI5drL0CkX55t7ye8nKPVZujcdxo7baq41XI0e+ymR3LbTodIwfhPAb
xhJZIv2JvbF+mQuziFmTztDcy//IX0d/0NVPoDzG3yyXD2tLnbWlXga0yK0CKD4JsmtosholuMEn
qI+vlmtJdm13VprLUFExZ94o6SkPnOJBdHUIi7YuArpvAfngkmToNvU5GkAB5xGVKFMnXDhBtrHM
6lwyY7J/S/zsYwufa5MTUcqvQ/m4Olt9XlZ8t+WtZYQGUVb3wK3n4VvIKggbSTbALr7VFTdxRHBd
LB25I7kH5Zzs+ONsqVeAmfuAEe+/MkzDvxFDtSQEnk4sJssXtrcWw9K23KbpLaNP2PJ2rM2y3BJu
62Xx7Xa49dLhUK5aBHbP07wp4BQmBk0tMIkonureBXNYnIs91qJJgDatHEyuJgAFStALyP48OO0k
P3dVf1N1LelcP0Q47po1MXzH7s4innT85aISVPKQv6ujUT5wBHlAidmY9bMLu7+h6UuKyt+d7C/t
ZVH/aXZos9rfo/lB0A8zDmhv0bLGSqpZQmTShzoYYN9XKwUKG2BhIVZAZnvcavI4P1+A5SCUpU2X
lVXBA6BYc75jVVt8oDRnR4tsZ4aC/mK0kpRGjYRvHYZ0ycskNYnlmKH/T45EtS5MLBwCIXH7qOYy
Eyepq1+FTbRPp3x8SnXlbqmFDGtPI1S9SkK6NYWSbPiWJslcZh9V6kRjdk1XkAPT9C7+RGPMiEJa
AVUNi0jNoyxLUV8gQJYTwUetaC6Xk5uM+N4SPhBC1uSaORyk4hOA9tBysJ1oxiLTP6kPy1hjB+pu
0S+zvnTRxEachjPmS8hr9ltGnIyD8C7mhEO9NcWhCUnKpzgXC9g5jIvnhiGGI2t4gbfn2GqYHV1r
AGjbCdi2Meq+7n5tXPhrgF9ZahGZNbXSaE02YOsg+C78BPn4GMEXW6+4UjJcP9n/ILlJkMih1u75
/88tT/gDc7OL+pDkFI+kL0Wl6l4SV+bopI0goHaAqx+clWzKA+F88KbnYgdljvFSJSv9V5LVJqWU
q8bQ9jqdhKlLJQjLbfJP+H/0mp4PqCXnE3WUQPHyysHRl4npCwZ1FgnKsVKJ7LqjrnZ3YMG+AU9I
iZLpTD6wq0i8UBkrxy9KanQhxpgc6Rzw8fhcdw3jZCMQmVttUNmTCebPCnza37mSlvyDyg7Tza7s
wHd3Iw4Af1MkW6uxxiY95ECMHF47I51VHrN12S6xVdbuXaJoh0UycrgEo+le/WJzxPyiiM1bpXFV
U/Vi82wgBXh2hdUNE3s4fwumb2tejSayw7PY1ko/nFTY3vxoQ0JbqC2FH/ffeRM/O6alZwNuiH/o
hUsHnKidBGOaasOpTKp1Rj6bg5V+MMXLBMyL9G7SRMuPPJ1hcAMtXDugWNWfGj8ONjJMiq0Rxsbm
08xjvhNcznpjvmd1LK9L/+/UJFHKkVMH0JgFApU/XT3ldBLgYUJqBThS5ock7Nxhs5zSXl56b1Lh
/Asz43dbXOvFz929f1yYBZ81uA2HQH4FNZck/yMkWqDgSBc8NpN58gxJs2PERVYWHL55OZuDvlnb
FSnlgcp2uKL8Z8zH+2DnIpWG0DBgBi++oizjemw2SVMmgZxZPs55qog2XsyZy1E7bjuPDajdTux1
34vj3XfcUNWGcB1N0uwDlcGca9I27vFbymFxdQb4P2CMw+KAL9pHh1iO4N3qQFFsAfi3VXAhM1Er
pWYNpumiwSmKZxQ9vYlgz4l7D2NF8VfGjKI7zZI3uN/HDvLfPi/leXrss6aHjRfMktrsB/YlA4k6
NT8hwNQZUhwQ2P6lwYOxLQ9tvKcnsfZMdh7GtZWidPXbLP3Wu8rgF/orJD46oQYCJXM9tTiQ01sD
ktLTP315VoK/x+imb3QmBF6KiIOPSuPWNu1IjzQ2ip1TA6kRYfueTC/v1YyIKxgKk/JjObKXRjoa
T3in3v6U9hGlLX4FV0+DbgPO4bvoNaXJJBKLymroD19iugid9waol3mdSlBkI0M7GOB3iiSgb2T6
cGMmGCde0et+1zWhG+osPCThArKAi6OWM5GbfbSx42g4CNxXlPrwSL4kMh6IgrdsHto6M36jiNvu
vZVKE4sWju2mgq3r8mlYScNjdlbYsOv1IPa54OPj0tRphPSN9MX5DjEhpeVIzlxRQgMSWwxD83zc
JCB2gWu1Wfak38iU2tZsAhkKsxEL5DpXm2DppQ9u7qcnOq9KBZSa5f6YrdDcL7bB9SjZ3opUOKoS
Nq1SurCHeVsTszpoeAK3DSTiRFTQwSxMMuZvaRIqmFJjOrhBBLpRy5Nyp25QkOZb29MD9vq4h8Dl
Rh9WykK7nHfQkn/AGWrwWS22W9Y3GumWG6eDVnpk6+13NWNkOEb3TkdrKIxcgPoGoUIKjagsOa4i
3A6fx3uBWhuSNjwy8PIXwQGku/m8qTjUObkFWgNYhSuL1ul1f8WzhgszkXbfranVdnBRnyhk5C13
zhgmAuvCx/HRfPwTFV99/2fB3X6PsPr2Suc05OoshQJXCZ5Ofu49N4PVRBzosBNpT72es2yva5+0
MPQtVKwM6coMA6jyIJz7TpXLUs0rQyF+19DQ0Au6FrQ4xYu0aaN/If2QpXfaDFH7GkR2kmXDnfwG
2gR8w3Y0Q7TL6DSuYxYTKR3NRc27uf8RzyGED8ZTIIPU9icTFc4WBpzG9oNT8/0eJG0mvQDBgoEp
rveW9cUbeKUOnOHgczY2jgbvlLTgBpnqVzNfHL5Nhdv0569j28zrzSn7C0SkMmwhcIk+VSO06EuE
onB7GJ/N2mHrwKUuJQbQLKCORPJk9UMfCwEBayC24IVm/eYoLynCg/6DHSUcPbcUhEVSuh5zA+Pa
4sRiqgyyolAXbtb0+svsA77vRBl6TQqSjxOxywJ8HOwXjiftwrCUxQUhdIpg0EFJ5AdjEFqg/b0y
cp/3jFW8pj0ZmhwWojWQ8dPzBX6I5Uvy4AHredk7E9MzGNS1gcB6+cdGAXTwIwkCa9B96n598TNe
4JbTaWWZGDRW2hrlva/s5//Th3c0HgXRzvfPo9lhfVW+aCJ7Cy8LqrxOdnkGu7IN42aL81ijPJKz
UrzOGFUOdiOaQFbICC7ihgZF5ZPxOVq1p7hfFsRyL4RVS1MA4ShmwDiPgN8yo+usE6LPC8IXTSVM
pUg0o1PrI3pcJy8qdwm059ZuSvaLBxKkJVwsGssgJZM/aU2BuDon3e71l9HVuGbcLa11qrg3O0jH
IQsXEqEkNkvEE6DJpIGPHvSEpssDqJxrmY1+Ym017tHsfWH33TzAlRTJssG7TGGzmitHPoWO2cOQ
NmBQ1zc06hjMvbSJrD/LAlE7HwCkOMplT9tJLHUl+0RwBpr3d9FjwMNxSZ62y5HVs/PKLsvQIVrF
h/gKDRmkR0WUFJMgAnqF0pVc/xkc8Ac07nSKCgzuvxlrwcDf3CtAHgLOEsbNTi7v8LxbeVowllqE
rHUDSxB1V0uGLHOwD9rl43b01s/BgBPFZ8meuuf5xyISRaiKsYSaEj5ij51bgIPh1ilc6PhbZ99i
SVcWpLaS0J8VrhWyoFqnkt+fe7GA/LsXZ6DfUCMHL3sJKV4GsV7h0iZ0JInEfVXM5d1zOwmsDMGl
BkGxKWlFK25ihQwrTd383geM19IXexRq/DX7iKuOAKwkc7AffnBJ5v/3m+pBMRSz0GyZJhCmmFkU
ETkzA31c+fxjD3BX+6IKrcvWLUc1n/Kl4ny1CuFMxvpg4FVQiKVvtBiael7WLg/q1i5bYmQavUJB
2SayZk/3r6v0Kjw0gO5AxZD80Axt9WtrAVUmIuSTAVudwjF6nUIdCwRrsB5pwLw4AcBZr8dG7sRT
x2ygxFwV4/xhe5DsIWSxMxeTi4UisOYyb/kv+4T/7bdrvy+8ozPnZS9LcqQzJn28cUj//U0kSnxg
JrOFq+U6jrvCEH8DNtCChEsJKZ4w1TCfJiRNgxOhYZTGFJ1zUCU734YQhxmphr7CZUeXdc5cRolS
83wmv5e/esnFVEYFTzkc3rLx8mLzO4HOHeIFjJSbTNWZgDYk9MyUgaRZFyPdQJHUfpYaMdhm5jJ/
UrcO5gD/UZQIHOaGf+tzjDw6LADp/8b76c1BvKolDextIQX7SoJuUnzjuXhmbISsQv/zo3giwJgo
7WeblPeYAYDU9Cx64iGWTwELKpgqgyTWqlNHK1lwBtB0Ya8xreWxs1NB+bTBTpgr6VIOSPsUAzdD
8cTHYlpJUzqsHeBUqz/DfTLRGrp2Kdks5RGvOXzfE/W2L54mIRAOfNdTlZhDIzGOc3DJhZkiims3
QOU0kkxjIu65m7fD3TUfWh6wfZsg3sHVHHLn34XrG6x/gKxNRTx+YtiVyjMv+8VdmOd1SNG6VrfO
/tjxaEN4qcaIcwa/JcvigVPoet3Y3K0PvkMca2xioCrqdLKmATd0LabSPp/XutpHKu1SUqiLtFRk
TGj26G5zSqkl5iYW553Pg4Q2L79HexiO8K/LLrJQ0rinwHDWKntuaRzPmwiG3Ruor5WGBi2EQUlP
8JkTMZDKodyfIKUeGWYwJcCf2C/c54ce+i5qLtsuzOZNYFaSOcgT49bfy/EYMFj4AZF4kIFrF7Ju
ltxDXks4mT3A7Ju1+92lFtD8Dsf0KVuWscMYKMhzMjRcbXIz2YjaAg84K+Gj8wTQMupVHxITaeuY
Ev7Tjwrz7sleXbjzjoI3sXpMNSGhZEBELvYi1htJoc/T9QmREvxMP7oSO7P5ZcK3GLNPmvtvzYu5
MSB9SlWVlcvLwDD+z37MC6+KR6oBdUSCpXCEuiGTHUqidm9DoSyu6qijnQxRDS/ucDyJB0fh6Az1
pBR0exHiaXGKqHBhxRRNy33kXpx7gIBTYkBaK/LmLPCHmwc6Of8mbiuXSX9/R41Un4kvxAISkh8q
4xvtq7OIXj1ZG64ei2XYI3LHDdSG7BCy7sUb3cVTcBSxeOdbqD+/oBIMbgllLzofbiMd5Iqmrik+
bNkdO7cyj5YfeqWP5jPGzDH9ky3VCnwoArIZMoKxKrDqnP4B2bXresQF2cJow8xS3Lrf8rgwKG2w
2pFW7NGg8QjxKTGzVeGi5UsXJsKudS7rSAkx3qsgedNZgfVeCZCDpb37HoOLgsGBod4urbeoVPGU
YpAFHJbFCIaUHns7ZLfQ52ch0ziyRMo8jjmzzes2zrir8BNTTa2Su/UJALsDCOU3lAIrllGpIeQu
rQ/b+orEKEn4GfpLoonzgq/VezP2HId0cMe3/LURepSBFFWa+47VJe5kt5bmWS1044YnUlzPmPeR
1RoFYgDH38Oprk+z0IXhDPR4unlK3mgcqVCosP8ltFMNZh9ktBKGfJhe6OTwxCO+GIPt7nSVxs25
BsjzqP/ucQYsGnCnoSruvEXefWYr6VG1FxwBKSiTtdIhT8EUwPZY+nnvutUUoNNcDI/6SJoVb8Bn
Fk77SucT+4XhimjcNzaeh0ugv8UKhCVjXhziQxwBT8lyJ5aPshVfipTFohGnxxb+H6UFm+IY01sG
JhfQx4b05+JpCqTrEDt059WQaDuLCO5/ZbzlygnQbFvofpEOphFtVuXpll3UtVwhDp7uMrSZNTCF
bzgTDCN+k1XcTdTo4gH9Pn1vOuGXnC9yxdtlzN61hm05uLt40Dw6fOEcuf5m/LOlM0mtu+N4akcS
PtSPvkRrNrfB1UrlZbClGeXYFuNO29dvHh9rA232btW8EMqiOea6TGgEySSymlp2TxgqiCCs5NXA
3hCDl4km40VfNAo3huwN7a/EvgcE5klm8VG3yhFkqqwpf2kd1/maQAR7K1ea53osgUOR+0Cpf4wM
J7A3A723kr8GG+XvUIS2+rChwOH4DmxpKDFcDV4IJ71D47oOmy2T+RtaSHMA4/aricfRcyh2ruya
q7cUNVfFQyEJlgu7j2ZWZT2Ru4si4gDmA+p7Dn+qt97wL3T6n+DsPOnlLmkmyoSdBIkV+Ey+cT9G
DX70em/6B90f4DOBNy/M5J9UolpIUicpw2oP+6jhPDak3wJf0Zzo/1C2tMPc7UUS7DlvC7fOhnRt
eVOMrjPTiGkVmalUVzyz3Ato5FJcsHG7ScMcklSfy1wfsJLXbd1NIo0bEgyhQrniUkjFJ4owZ9Kb
ZupzTx609uYvlr5yqBeCAqKChfUJmX5v8bC3r+mnnRaqIX0VFKW+Dcrg3qBrEUqlalixHDbWZdvW
ZQagF0YmEqYqH15h6Tt93DTYSoft9cl+gbUlEbW5X5HX/evcXpQyUvSm2OZEG2xeJSVVpRfWczXK
seiAcdjMcdm3ZIdcqpxx6QasknowzGnxIuLJnHklq7YgkFyUW96+IoSXsCCewjJaiBPXzujUbBhc
LDIYZJMXiUbRJ5ME/NzXvnI6j3ay/wlltvvBzzo+j8SLyeCQZH6D+0oP34yxRNduZyJFs4LICJQq
HOJ1vQJnv3DjrVANvkae+upvs79HPOwT0iFdpjERKqouvVikFjDSS8S+jPcBw/Zs27ssPGCzlTgz
nZz6UfGgpvesHimN1gck5dwD2gL3UJ77BPdTX6mkkKheNl+VJX4HOxIGqgm901xiXq8hpIFxSj7m
KJpEITLIBT8/2Qs/lYzlq+ivPVJO3eVv2OoXQa1Gpn3MvLh+hyGkOpliMn3fS8hQFmbvX5umnr13
QBo+mnWhXuZJ6HuJwZ4M8/TkrtnM6VjmnlqEeSuxzUfdIgW/51F4kM/hyhpdQaQiAMCLJk2b+mpr
3YCbOQBU+toLbizsQURieeB9e6+aTmUfsM5VrhnSWr2oruqk8eVgxS9+I4/GeEowTe+hRCIr2hQm
7yRMXH/9ELOVFuKSvTw0MTqu1jT/8TmnoGXEwiKcxVAB0TJ8dcan1sKhtSVhWatxIvTuVsd13OPr
xIL6FHswt8y1oiA4mQTTKbzyDGiWDbO9OHiXdW9hpSKPqwA236PlO8lLV8nO5Pg7zmV974DkbMm/
C5fEx+Ry/fLnG24LA69xkqTP/EbkiQUtoGTCjcrvKyLlv8PqSuECsAEmFGCA+LSKaLmLOHtWXiUM
/Oeszni0ziBC4vQp3L6k5r3dEfyNd79EJupkb3G5f54rG59xWFH9gjv3AsUEVLVbgZdK+V7vad4X
/knX/0Od66Ym02ta3YAi2TtOWQ5mBRR2HYQw9puWTdqEazoBA73pJAHnkGwxrJ3Xn69ndbuLQCcd
34fCn6itIJjOhv7cv9afbfE+ioQVfPeb/TOdNDHbETjZF0u9XiRLMDjAazadUxTob4ArlbKpzt5Q
BV+hP5M8rLQynuoC9sz8BFtwZFmsYdLKnXs6TLxgPOiHR8Twf/2pCnomfZNDJmsGo0BYVnLjDYtI
ZHN1bEaHXCghEg83+L6Aksw9pW7hP88oq7rYbpUs/R2RIYrtzKU/i8mdLP/4D0iZkEFYjbwCdGyf
dhCMdcz6NLUxi3lVcWS5mfugHTLun0sWdbEuF92CC3UQmXF88QOue442oBZ4VmphrgmC5G+t1QOO
xO7Dm1QUOqYsVKTarBCEMgrd13HJNiNG6OYEDtmPmyXCDtDMfcp61SmM92VVqBkxa3jhgk0bJofy
NrwEMzOx6oUPPwVBEoRK1Hu2H/ws5vT1PhEEFS6eccv5Ff994f5BjvZGpB4sWeGVLPdx8HP4xP+W
EWP1koqHKZZDR/APnhvhU4XeRhdLfnas9e1SIwbFlGMhggedohQiIzsRSXv9mw81iTvdP33P+PS8
3BET+ThLBjR+AXSuMzwRDylj+x+2s3I/dvC3A/94l1o0Sx/2j3WRFPjPuipL9Vls/qo7Zq9eH2da
U3n31fTIUMQo9JFTNrFO4LjfTPOMFiGUdLrMI6RgATXQPwQxS9ynWLBl1n3xjH+ztKTkkdELowcQ
LvbNOfFRzdG/0G54+TAR474ai6Ci93imV83ZDaNqNlZPd/5naW4+ceZuZt0wyH9vWdpxnJIbO2YK
+Hx9hWebOUKSiREiSienYurr22r9wHaxFUU8Lj6zXyC+1oihGq3lD1tiagcbX6cElQnLNQypdEKC
b3io6NlmiRCBfncqVo30oxXcAadG6Sn55jZPjDG+/KeujSTdFnT4FOUZKYpkI+/VR+L5eN6Txka4
/0GrZ9aMt10O4PnnziUxnJJ4yeJJsJ+STB9trbnF6Mw9hOoNni7sS/EmWCUkEQBJpmctTL+34VsB
fWi1vFV/CCyWm/q0fk4uoAo/aCR0OoomnLWGHguC1mko+ocCDHT/p8OZzVKCA/Sq4pCed5o7ld5z
s0FvqfHzHxVloWORYwtUxruyIXNFc0stMlkBmBrqKaqSJhWebhBHSbY2eICNZU5+jlgdzZ48cnmF
E3u2LV7vb+PT+xXFOpVRzLCwcy9HlqTMgj9iN9gSjdWkIhFOV/klx+FJxMIGPYfM0UKW9Y+a1x0h
iLDbGEaVOBnkMXCWtwVKTrs7ADR7Eso554sIeewxe4h3aL5LA8mjLjVpVfCnEldectz61ugMZwJu
vxQYc9KLHhmu/cHcgG7Ks2jFFYYLQtK6252gWxKJmhZ00AZO++47rIVW4WET7DlVgt72iWxsbOb4
G7LU/FDy7kIxAYY8SuY3sN0Za7N8+3ZrzMGCcuSS6/KGzS2QlsYlNU+60WngAyrkLbGDGHO0qCM2
KW/Bx8oMXzvmBfGxNiJK9QUMq9/gRks16qTlHHPRt2PvgR90cME/1zuQMsEE4pwTAfNrAwFr6USO
0jzr5+3SYOgZ/wjFZqy6nQ9y9g2hpNrECgYHRi88MNBwntRgEXgRcpD2ctXEDzLRX0/HpJDTzoBj
dW/XOsaGfaDPqEDUC810hAEIw/HGDTJSB7ziAtsirFd3Q2qQkqbMC9K5eGc+LbSzu0q9ExDMYjX7
HGph2I1jwWf3eQPkiKEBo+nqfRIC44Uf3kDCNP2oNREbYqLvtcgr9dr+4nZiV0zO7a+ws0C9E6/C
E0k25w1BBSZXiWwT4mAMwK3w4F1Z6jlg7sD089c0or+H8Zw7Ra+UnhHujuYSgrBKniYt7bBRyVDJ
JTzCvBiBFvivqXYvrzS2eTR9vpIx0NX8rqA0odYKn7Jx23nWHTy4lJSUyQTEjOc3tCfW6CvAECz3
gVL6Hf7qaus7v9eruuc/5/W02n/gy5IeF9ER8WwykUmY9SJXtWNA64j6rPQmXjXRoEf9X3gtvm2P
05MqDhiQhAWQAkjXovuQmQM9Q+a+sBmTzH9rKW5n53HKduyOfEdp5wnmBEYpmTDhuTHSgNK7Juzs
jRj4blVyRyULzrs0lgt8COF/dC/aYCx2/z9hNUx9syeQTuQPJZgJQUTyVNmL+Y3wnMVcKAtHVUQc
fOkHNd5vOtPzv520vdvgvbw0wW04HqSfkyIZu6V77+6NJVOlcFZZep+JdCxCBsOIaUYjGsKlUy8z
hgPGsnYVpQFUBKRQ/yXzDzprtm2EcJtoM3Kd0/TW8zYPEbG9F4iQ0wqMgjALIicZsKaakoxg0sdb
mYpAImKpmlMVD4CJ+fXec9uu0t2HcBIq8/UThjgsD4/IkH2FRssuRbswwK0ptkBg/5dCF2M8U8oK
WPf45CG6iKFeOXz2L2k618HkHA+Lu4xleoZlTX2rIcm7FcLRccWtWyGMLu2+8OMvH6Ne6AyfO6H+
oiHEDouF/Yh+VI25zI4cBf25Q3BUjqEsfJQytBm07ILvo84dLQ4eJGy0rvY/wFspVsjzunYsA+HT
p+Cq8AoawBuySIAWl4hvLrHPI9LezCx6DZvbt8zF1Cca7ggw9EGvIbITp/5fKWjAmI2/Z8lbdJAQ
T0kpe8hwAYoiIaNT5OCK5WHYTHtijWlk3ZSKT3r5zoAW0WJ603CGVLE9NIoA0LokZPUUB7HAZfps
LmtcRG4iaDwaNewQCokaO3OLMvjrC8gFW5UkSDT/4zdEMysdoPxIgKpanFfBSF4QFCvrD8SPvOnK
1UZINTL/EWpyHrVgipMV/fGaWs9dfDVvSCBLYczgpor1quS19g+7A/Wp/yJJKGafIll99aQ3CFVQ
kdjdYZ6Vjr6qgctkHMbMoTmSkn0hicVBg7V8ANTrzoH2PnTvTDeOkxi2Y2ARCjhJ7sfBKn/3GZzF
+Q9hbCcbMAFiOIk8gAzKqn3QzE07WIJ5eMeYIaBHkE/LNVMMXfdMPFJjNeKUuhzpAXri8360UFct
313a2YBqZalt+jW8sSGaK++2/O7Cq5TW/nS1//vvT+S3sqzTFHVaQRaudE5rvEyfNeBBXwHsqa7X
WtUum/pjk2ZNaVcbJCOH+2A6T63H7eHndu4jN3CUphITtd1XOtFfIfoiIRXYAtQ4TEZhqacSkKPY
cH58sAqwxcyOXBg8tyBqgQkS4PcWk95t3CpHlzKG8/tny5TNw/Bhz3thjYtrPm3sj/MnRvAzteBv
AiKNDT9w6B57tku/2Pky5jaLkn2/rC21UHi6Z6bzWPQENI+qk4ndjknjPtRJzdMPC52rMXWui7xa
eN3OlGtGrBPJ9Mex0i7PyzweLeDbMm5LvPXQSg52Noc6PCTm2rupO/cox5bllaInJy2GjluovhxY
qYO9k1HQZ9g0Ttocud1cMZ6Px2XqJvJgb2B51JPHV8WyMBN9IZblD0vSrz3NI7zUn5VsXKjcOQdd
QjVvvcE2qzLmql8PKHYeI+WcT1mkiIze/kjAHXyefZZBlACATE/zf00rRxiKZ0xEsiGuNZ2HHj12
gXKFzS3Ivx+5HFQ19mexMwVY1RzxETAZgEFxcxqrXyPDsqILuGJNAcZhyqvoJaVqlzl1qtUKtAAY
0bxhzpEkL4mJseFE4fsddf70ybu+1hPK0zcyvkyqEFBFS80X3l5bcSEuLUnxuKC1C2kMDrRoRpLO
/s4SBmJdTTXv2twNfpwCrwadcIbj/aW0VDeSZyvuRIbdVBxtCCHDq4PoqxMH+awAfMYTVeq09rv8
SntIEtIWe1lD3h+ehUJ2ULg4UWYU3/JOFVkuZerfyghaMmatnvPVo5t6q7MeDxMqPZO243MhM4P4
yqpiHhgw4kIl/XEEHuZzX9TMTbVWLVtyrArSABGMKbVsr8xjNtO9l/crq4KQYyY41aTLNi6dpVv5
Z540psC2UcnnqH5VD3PAgawH2KnPZFiK4GR5bXnZRQBuG4kmQhlpG6LRuaNtMB2KjrWrtlSyCsz8
30bHL0HUNwjsMfVq3vlk4bmhNXDclvE/+GijgA047ik5LxVEnrU7cXT2yt0gwRo0TFf07SjbLWT9
gFlzoizguiBG37m4u9mZnns/piSmElF2X46/PgOJn3LriyoM0l2Ty8L7ZDB6aM5WErUu0z8FuzUx
j9xlymHeI+rBEaRTuNZhU51sLSUFiebeGW8+q6g5St7GssXZzLS0VUOzBcbwAbqlpmGUj7Fwsbga
guih3ND8Q9FDP3EVSbPS6HzjHfo3CE8XOKXvfO5yv21d1RXGoRadboRUDVgXU3a4/ZJzczpAnp6b
D0sbxCMNcknFX/NkegCRPOOkulKUflCLgCpTny776wdcc+aFFTe7b6nfpk4K3GqbIQqEZFZDkPvE
9BF3tCLvdjPP3P180Yya3e5DZ1o38C9+oOxWBrzomL2c+0BtT1tasurcFeVGvS840DfwlX2BsI9C
f6aKGS+bSU3EU8N6+EFQ5uSalRV0ocmsLfWnRLrMN3qjpSirTQ91iJZ8k/PasDnjzlr/q6R2fVn9
1h9TvQYvzQGdDz7gtGNdOJWNaXBeEg4qQqAU8CiNLOHiNw9C4wcYG+xK29OJgQVDhvwtLOQVLfhU
/lyPXPSRRbJAv1hxMm/naP2Y5kb1+wcmbE5Hv4jn/JsDXanBxCS6RdbFtCupq3D4Cp2kHokGXkxo
TPapNLLKbtr1H0g5EpveAEs35o9hnBAHjqlHX8/BpXgGd1JXMugQ08ga5BKJZuhwYsflvNVpiF7Z
RjA7M0LPSRw/I/7Aop85L3WZIWh/ApIr/pck/NwzUkQrVOtlwzCt+nVombQMrhwSyNZ88yRnSppw
mlQHP+So8JCPpg0/pfxZTAxRuU2k7hmjkkXPJ4U2zG8yqWc7F1EJ7iUjyLWUqTC0Z5GIiWQRhrCE
4mJRsw/8FHxrEqkmrvbpOaoIMlXA3RCuyHay/scjbUBQK0xjY7ubLS6QnPWFK3frkvR4Rlbtski+
utG5Sr7aqAQoSvkrRrJrWpLkLujPxPR4tAiQiB64SGlrVei0dp/vZ+s+Q6bVx8CMQhp5YThH69DM
AmcdxzqxlH8eBbvHkV1nO7BHUmUeWp2cR6g1gQtjm2aKtFHmJKWR/MfdPvgdAnKP4VojPuezb3SV
VbVqKPIMS5mn3LPwnEyrmlR00qCef/sr9GsztNObvjqTu10vbJ08EXMvB+ItOKg/DhDl4WkK/NnS
md7oSJ1HWIEk6ZlUWItJIy7wvm+Z9ca5I0mUwIlYJ03AeGW8inoBbj5RfCkTEVE7agNzi7CreIHS
s5ai+J+p8KLYAo8CikyLqMphS6cdgNQ4pfxAMopAP40P79fTFrnFGwmAebH93No8h2n/L6PoK01D
A78o04UNi61RQvA/2qTH/pqScjgx5i/js6VCrTgpxHXJY48lZydCt9xjttvb9//hYHSsJjkV8XLp
33Xw4bbbvY8uXNyR+Da3kIEV+tYLfIx8xws4xLMg1a0Iv92dcOn50x9MIEn1IxYNuabVW9d/50i/
HiBYG99ERNCK8GeYtpHK0lJlkBfBUMw+V1skxgxG32w7WyoaxAffVc/bPpFw73wjwfGVx21xSV/Y
5nT3l+f8uWgBN7oTsuytUly08VY0sKdmi3CMI0eTjTD6gBnXyt9xi3Cq/3LZpXa8yViQT9uSQV5f
0nMGgiiZCqM1hnwjIlW5Fxent/idFpWbooDNtjh/MbgA9lus6cJqyb5QVza7QIBCpJeBfxPkXmfz
EYS6fgGZtIG9UmYXgDXdFGlfbG3GSU5qWVTujT3T88kpQI736b9IvkRglxr4Cmsx3/+kRWX24Qx8
qbaefiZr/Hpa6wmoIuN3LbXnrkVgPyRmK2oKQrUoeYMqmNASitpR+wjb2SryeX/OOwMszJaMwPfR
J1BhAmq6mKL6Bpt73qbeQnS3XH/AKwBpJ00VRBbluSx7Fl3nVijhk+9gfQ3+lhWFsax2Sz8TQQ8F
59HsA+fnhDxY3Bs7VkkoOGsGiogZm1jd4tq30o7MiXR1xPCDLswIKv3C3nOunhjO5jzjB59VF5d/
PQnHHN7u00B801tohc31xdksD2aBbkZwxQ2g++bJF7w8WJhtaE/LthhgotvFJY+UQYoM+nXDWuzH
ubx04vCfiTqIT5vV0kFXUkVyEZEktaFLijnfslhgGjhVSUgul/e41vjsuc+ha/w0nxjI5jyvL9uD
58f38JFkYCOKvZtYcaxo3YstmGh8bGyFp19vzvAVRwof24waHK9uNLywo8GbWy47YxwMTYxZdilB
wDzmTMyzFvFKDRRy6P9DbhfD3S5MEIAPd2OJkSpO2LVwZma5CoGtY/fclMLmOt8Uo8I3C/bKFChi
3VDAq1akm/4d9bW8csE34A2N/KqbywXtQmDtueNcJ87ABe+YWM4/bZVFBO5dK59RtCwiqsIHhu4K
L+LjmGwk99snoRU7zdTdsZy5YSz2OAtpExjRrYNjPbl5mf6E365PILLzhXrcKqlsIeYKEPlnOU11
kakwuFg4nMqT4cxPnhCGU/3as31ciHGCUmbkM8gMLy45jRT/sCE6YSbNqhQ0RpRn8olXcYNAb0td
oKAwDXy0oI53EQylR/CoeW1Tn6+wALAvdskjOvy+cQAAaF8RD/A5HvqbxRbIQj7D0jt4OctE/zYS
j1gnLkjplc0iv9drRwyGnVgr1ICfA79/YxnDiY3Fte4UllKO2Pz8sfh665sLMADu1954gayT49+W
4Y81ka9paR9UI0TeSaCz6qoh9zENiUXwCotzGkYmX/7ZIvrv2aNYwt7CxhBiz2B9jICIPcJXGBop
takj8zuTvtgC1DURBn49xMs6eX9KDDYGoTq352sLmaCLHs5AWSfAuNHhYm9kEQjZr7AuIyCfoptv
KG6cCyA2BcNQfdbEfVxjHihO4mCKMqZzXde3yS/q1fh0OBJHALZCklrk+c/Sj2zU7Gl1OHGp2sIt
vAe6NKT2yW8FIzumFMQpYr4FNMyJxn1vOeQU75OHg/BPbr2A9zpgJMdIf0KhwjGjLqD2JKACsm9Y
YfcLqH7SK4xwNq9Ryi6DL0iliAY81pOvo56QIsBGHw/7hjNrFp28bKCSIo//4uEv2isNKnGzSgR6
EDQIA2nvfdOlqC4+LtrdktI8RbcB2LCMGO+LH6fzzwDgqRvIXFuCkNXb8qmQmBMns1GSf5KS8OwG
hTEGnL9hB4HYa7gotbmZc7MfVRZn7FOipbvNOZFuPLtUWZwFsjSGrwpajYCDBCWI7fD6lEuOgxzy
cOxnp1c0ei0VkBLvD4a9VAdGKCPlwtbdS5odnYokR6Fk/+TVpI92b/Oyb2jNU1pqPXVyA5jSYEtN
fTzr7LfNLkd+Z4NZVWiIOGgqSjHp7A6cgO5D4N8wvXYNn8GPG/hMmkOM51XcBaBj0GORAeMAFS5b
En0agsa+b3l/J94vHOSjbH4ysoPN11E0gkvYyeh+ZpG4YBZ2U7JxKonzXibiCaUKgIBcQ2tpZm9S
z1voRARhFj3QWA053Om5O01Y0atccVQR1L88K/pk29ymq24iUaPzRaf/iVDjerNKo7obVsDr6Rxs
S0SmHboZ8eLfJuAtMTj8xS5SuiGPIV9+SMB4u1aJmQMV3kyOOVC8RFTzGB+ToazLaisQM1SATR73
TzSDcxJhGABgzoxSPoI09DaJzCsFBn1N1u+KmETqFb8bGjBjvWlxivxT72kjDZyTVZ32DVmNBVK3
IE/KlVJ+OPrDssqLb0yqObCo3/VK9FCKQKHY3+1OIix2k0QGDBFKL9svpaAAkMf5Km8XbA0VlV+z
lo+7baqXUOAn0lFxNxtPyxZMG/lKzhGji2cCXZd/bpAU1LHNiq1cZheeMWPOqW9zpvKCe9zV4TsI
MaSdzxGtV2//gTaUt0qTOPd8/goCB9AW/SvWIgUXqDQh6L7T+b/GyIUnbL2EMKsTCH1ZoT7irhh6
VQRph49kf5Qp6CKSkAd/3rkUtCt7nL9GqpRCbtiBmEW2fmxYJc6g21yL75NvObhojk2cUaKZXL+9
eAJ+ulKZt0i8OrF3k/oCcSpb6jSFbduUjF1ptx+L5TBzr8XWIe47ruOtPG2boQ4+ZlEqBcKzw2BE
I7yTMgQQx9Legr7yWaEiqSDpyRLSYgLpQC2xGE06aSW/1uN5GnTrOKOnGys3Lv8RVp9Nko0TlHgs
/uwzRhtQhX0hEcP+licuOgYId/VV6VFaoOb3+MQESFTVrtDXo1nS+ys4JDZl44MGciJAMgUGdlMf
glks1NOJdPDrpwSqgJup3bi6hesH2FObpuu2ieHaD9yoRfaIs0BhUSvpGxtucpK1iXb1OJ1A8uMC
U94yARI7oxGaKoXIjhBB/KcIUXNmiinn4g1OK6gw1ECP/2FvEO+v7ijYM7psENsnkm83YK3vJCKD
qvdbmXG8GhLYZcULhtcJUKOq6NtETKg/7e05zYb3uxjSYuNCLq7a3lcqMHy+F0a3bVy5hx9eOuEk
UWoS8VKMOn2xK1b6yJdyIVgyOXqqfNZgQ/3xs0gqNK1iBLBhH6zqw1zyjrSOQygc4cF6/BYm6tET
OZ8SUJmDf9yFfaF6cfl6T8FHAg5/WWspfjBdCpMMeVfz34zDd4qzXPWsb7mjS6WNWbhZRjbNjzeH
KZ7fyOGTKherrwT+oAZ7cyxdRSGE0D/uVHGfMZ1xlWFJg5rADZqcJxaPyzWhE0nX3X37895UYGut
Slw0nNQFvbfTOBGTCnBVxmfIkSc6KfzWp6DlvkV0nsOZkzFQr71puGOdNkMdLI4EFAkzFTa+tOcA
I5JZR/eZpKxu7m8zsEI6nWYIGvZsk0JA5SYnxe/0UAcCRQsIJj2GZminjpLX3YswqJAogCd9VrAb
E0dtQy8g9/L3R8a6p+ViVukMEHJCMjkcYHZ3TAdkiV53b/i8+uizYqbJULGSHR21OWTC7yFkHJkn
9G2Q8PMDrwCURDZaQuHC4USh/TUPFyNgsQ897XWs5+GZDzujQyRUlmXGUSGsoeIkZdqvcLEgZK0M
Kht75i+yeXxhD0gKuDX37o4LgnzEv6JU1Gkohrnu6MgU83ob167EGVNK2rK3mMebsI+S35RA6RXn
ONLbLIox2s3CBCtSM036Y6gl9z4mxcHoyze5uvqwhOW/n/nhMcoLkpcG5CJVldA0r2otkSTJf2Xa
NCwwSgNgIXF95dBeEKBWKjqf/ZzEN5LhQSp1ZAnLNMpyqDjq05rNSIDOLazRohLhAfbJw5TGHm9K
ioiBYYqrNXQyAzLeScXbza8z4981vcgl7h/kUHYOLtDPJTzklzXAY87sYPa2DeTwjBLhNVODzY/P
bx1s0rtjYwKrfzxdWwRuLByGEFf7Jy1HyUb+S4umT7DHkIBH4LWw1dVeGJG4hWl/lDiWnnA9PaIR
5lth99crwcxtpW3iJb7o8VDjVVWnP8nlkFZWtSbK8abV9OnVW5B//q+6goOgNjM0RsrucgrK/hE5
ANtHssqgBCguIAJlNpxur7o2UnRWUNQx6BEK2wEytOKVAEnGW4xURXOG1LJSYWqXQK/MQyke9BzO
TQPArzxO5FfSE6KRs5AmVBIy15zEC9+g0AvKf0DV/Xrf8Ju/EM6cbRG2zRwHUuvKd7Xub00kiPgB
d87RoizAJutYNUd/75Z9GFUqBgqP8j2sbEYHYYM1hB5LPmfjY3kG7LZSJATM5jHA5APE7Q2UCVgh
u6fEbGORZ4jkIZwoP6WTT7s5SgsgciVikXccvqBU0kq/DeF/U+/xbbz919F7W6LkMZMiFup9X8zU
tKxpUMgr0dVNaPE17eGQuOB26f4/xln0nEYwoM/HhcTe6JLgIx3JI0aes4vn9itwPasls5jvNGQ/
gdJrd5+7vYTgkmQDLb7abtuRGdIPOM1SExQxtiyqZbUZ+dwSJcrSgkd4zuB/OOmseTL8VRJD7oRG
BcuRGh/trGNEk7KZOS20Lsn3Y1OgJfho5vDvPBoZr6akSPxBKtnT+Eb/xcmacNeVG4Xeh44tb5hC
aEkx3549yBZGN9ikrZUtuDBsREfwilql/Idi8EIQWIBwxWzNYvicKoCX4F1xEzYZ3pB7R+2POKuQ
QT83NaRsTjL+GThVebmftpJsSt0po8kZoZaeEnT6dHobFo5k4DpASSjDrOERDZKBBMKaTyXKj3Py
+I7wT6xY3PXzlruQJQDNuxTJU+36BxVWsu6u+d7EUJrlOk/sLCeSkLYapfaikTE8Zg6cEPxp6FSS
KWmoC9KxxS817A4C6vZHbotKMTG3J/ZDAokHdlP/MuHirau9pga6A7HLlqR5hHDHRIi5pmmNkKMg
pRwI0vcz2+K+m6SQCcpQlBmfWpJvQ8wY0S0Pc9RRluT6ePH3JMMFQEkNRCtVs2UJogg86Z6U8UfH
qOaOmtrUPW6uAZ8UJHTxDFB1PeHFCHO85H4tjDe5OqdPtVZuUbQO32avMO4zMrA20le/n7verA3L
+nH5mrbdv9Wi0C59W4X2kdE94GFPS0r5iKTAIbVcW69CPptvMD8Fz0H/LD+dRbMnapGPWI9C9Lia
+Arv+QMCxOvLP7RO3/cLITkLNvE5fJkgnbLKNZh0HwTJrwOzv8MKquCRXU0c5L35VCVWWhN5KlCt
dkXISFkmQDDErThe1pbnNjBSjvSzoZYRabutnBeELYFpSTbgaqIu/sQh/aaELnCPNnI4Ht7FauKT
fSQo5F2kIapVRyVpOahTCmIlFogd9psWShSkJlLZTh4aQDdzO+Ue4pSMhpxCcbOZbZofEwrMdXI7
FvCQEyia3UE/LL4Tz+CmTFqCOQTZHBxBfrffm+RNc+YVEe3j7clJZKzZPjQcbKkzKi0R2U/e9zzM
MXPms2X0n9pDfrIWtDZiLDXSttRfnGyibm83dJZ4d3+R3qakSAuNytP2ib+MrmtO5rWJDSGjqdkI
90wpQdhfYpPwC5PGyCPq4J9eQMjm34Uf98WkrgMhoxqadw5ENrSrwGBC8ssc6Ss5KsApTsmfOqdp
BfuN8ZpbPdXe5f1MByY6qEoFH6RkNXmmmvIudQdUCU2EypIFBNFMwaIecRjXowM2BVjmH0W/gDFC
2DnuZcJk5fV6gHNcuxthLMLpBqHGOk5JjXHpW8ygA8qy3d7byq3FroQHvJ56pbr78OsX5pRRG9N0
7pfV/l4byhcZ5bJTPMVO1kb6M+qzJfGBoRDETHk4/LLYKp+r0z8JHFAguGbSlBNoATiW/J6qnt28
rx8G6A1L8VMSVZPTq7di44V1PJPxye+Wf1xKnkK6kaQTLw+AmcQ+DofGR40qlNnD8B2aEVfvpWek
PJnPKm2btlV/k8El+3bdFlRGp40YEhGRYKsLC53yO5oxwB69IQLs6m4kVnSPxN335JnbcUoa/Noh
MikoUVc9yRw4Zpny8ptRpY//6+p+qiPAZaN5gxyDE/brIXJA099zqdvoI2Jk+4PajfCl+hzyvXqH
5MdAnhFMlqhON7tdFn6b3FatWQow+L55+F/Hno4wZNHkK6Gab7OBnZw6oVrqndHef74XLP6QXAxQ
CtI3R3yw8x1Tu7IqTx+iiSkIGGZ61McTgfeOyjpKphRFZ52qzuQiySZOAmab2u/1PlT1RsYczX0H
fEeOIqujyWylEnoSo+F36dwJGSshwUXOTlDU93F/lG0v+hFhF8K6mTgFVtyjWwYAgBEWTzQshSYh
7UEAxs35ddLTNXFosYcuV1yTHuojaNFA8UDnt64MNz6YPpCeCAfYVduI+7K2Qhr2AdW+HFvt/su6
64ICZvISXawpF0yHsKalCPtVUglJPezanewzpQK3Zt3kCfwWNuOIWdz+oC7rLP0rYAKY8+leVCWU
CqDMxJl2uBwe9UfwmTaQHd5lsKHKgagqh0OBsAQlUb3xdSo6JGIcymj4p0Gko5AZDNzPrwXbxNY0
CTz+kubixYjjgbLfnYWH5TJPQ3nQPYuRDOduPHzJKGfpoVisP0CorS10DR40Y6h+inCYzyEg02yi
DGfsxbc9a5rznhb0MlM30FnrpEgdW2j8NjP6tzuG1OF6+Pri3xl6/UC4bErNPD/sz/+3wsOWlqz6
wx3/Nt7p1fRw584UcKRyYVMv/k/FHDq2/pWaSuBawQj9k9/4dVSp+4uY6M/k/qmNDW5dQ8McA5TD
KlHdOyWPwuu2TSG4zWuLq4BwTDm4CajIDYAUpmyT18LClhUxTVY/yz/QrsQC+MaI5DUFm1VXFtAu
PDTnkUegqgISQjaly+zUzuqoIk/uEZH7sx7IaOKH0U0K/97YvRYOaMu2bV1xCURjWWd/baSI6KFl
h1U63dUzLKjnsFLmZd8w6XAl9IFhV3hsZj1t9rnwAEUQ1H/FoA4iIk13VqZ0ncAydOWNa/xwtOYT
2qYJiv3B1+7BfO5LeJ0qcek1exdrKaSt9WkeWOMpZZQ5DCmJqFM8LuVtWeebmBs1h2vE0EB+3pSi
Zbs/M4tGJSPBVHV2LwmH19gp5VoDZZ6ZTWvXchfFRB17/0gfakMXQ6NK15KARVl5J4esAoFdyI7m
Y2gJD1T5qkEx/tSWIjPtrc/1CNMJ9BWwV4IpU3V2WjoGWHsUQOe+6fhZqxgMH4lQ16efbtNFIP7S
SmWok5tiVWkQUbC8kWjAL3wFKTvlc8gT5rRdtkkEi5JDsvVCrX4F8NTonvOmHS3+2rBSTycxTLXG
FvJHf54xoS5nOhLpKuMhH4NAXcK1cl9/6RnXfREyBrtCaVUG5GBAPhHnczybWlDfvNAn5LZVVcYX
JHPL04vTINIlpiLat36fp1N2ZGTiUDIXxDf4+iM2vfecH5BXPRo4pimxcu9fiq8tXlRYTJTmex3p
WZ9h6VNh0ARbPzQM6JeE8vQgTBO9SsTo9lHIi+XpmAbdGmw+ClEkIowU8g3dce44/TtIe9v0jZtW
rlH+CK1UVI8OgTSNYcqhn6uvQrC2TAbo99NtFDFRy7FAVjOrZYyp5FifIeARa3TqT6YKRB3dyC0j
bdXwlMHxJT8qWA5PtuDMhG/JlVfgZ5h5qMXaWdrUNx+g6oNIbEpcTcgV+0UtIjl8kqpmxvSXo0MP
HZdlRe7S09hXTWBxD6iShWuWh0NmqmjrXvyVwzmejn9dZSBja4X+PqGVnMsPz9RvkgN1aH+tKSyw
MeTtUrnQOIW97fQEhcR7a3bwnc3+ON/nLv0PBUaIl0vSTwbNAVbApZ1H2MR8opAFjYlrFGOYni83
oHpByb33keloqtClCENoWk8YFzxlGU71NrXhOxHP3gTvGPIleJXfk2eMrozTI+bqvWoXha4Mo19P
rRf5J/n3L5OyNHscMiflMZ0Xqxep2NyalTLnZzH6mErV2A/AoHUoOH9RK5my+kowQk6T1C3/o/eb
uH1SCfGUoO9/pJ4dxjgp6UrEJO/68YKIBqgPnlzktTgPPL1RxsnHiiOfueuakHEMLOA5h/gZBvqq
QOIIq35rihqGKyBhzHVXCQv8tfBGaFJci+dN0P+pQOaw/xdOc4BztfKQD0J9u725TZrES4mifkIO
8Jequcb/arPGzpX/MQ2gEvC7nC4yF9k5VdaWcC0OBitj+J6MfGn2qEucwcVLaQqbWBqqrljya3ZD
J2NW/ybiqb0++04wEJTZgO51DnqgBislehHCShc8TvoL0QHEeGOcLx/8hjrGkC2DTrFAlsXRuopS
igG5L/Y/k0bMhFYG+HEWiJVI333OKvszV5L72DVSGiuQgCBcStImzyCuCO2ZNqCqv0txvSYLSN2a
8qSZSpj51MPsoAJ6TblOSdcqKbUkG4LdpjVL0qGgi39dcIXsi7QJeWQZVTY0QY1nFbbaBNDGflrD
m7YD0qQOvVRmD6t//1J7IaP7t46YYd2GDKVlEPzTvX5ymYvFDVSlUIT+5NSxRgT2+9k1wTuYaRcD
Jk3kcRQ6VOh1Jlh5voHAtMJi39za6C6CU3Lb4WKFfIJJywF/BCjGXFnKUzkyAvmREyuMbtdPbLpw
eTXDyBlh6VJP+SvxwglwuSKPCpeJ1K/IHra5udG7KKfpnuS2iCh81sp6CAdtS2UmKBwsOf3Zjz80
0oohj3gTHNGCq3SAz4qS7pc405pWqM/8WbJtzdUSRwFVhvIThgN2ejhyvsPOusXpg4CXKEfqBUyS
IRHKDXU9/FABDqb2yorkZDbNgj1qKkSjrpkhmKzCzdEB5rkCyjETKBwuqAij74H1gT718CMOS4GE
vbQ+z+esW3x03MLAFFu6FBD/xzLeosk8CeVw6D4zp0DVUqSkmUpQG4uqBxIFp/a9Q/l5GCZBOx6h
Tc9cnLFQCaPi+2ShlT/9exE2IyN2/dy8mahjh/+g4AOcjznUTuMKwCr3xRlpfnaUnXgUpLGLvTYJ
QoHJ1rn5o4CpquRW+drlcCjE+Lu1rgV2b7YyG65eROSGqAr8eR1Iu5LFVKR755oZvtlwictdhsQ+
UUs1AVZxKV8F59CxUhp+nJeeUXXcop8FOuboQRsyMq38zuDY1cD6+laJU6NgIevwCjss3s+gkg2L
ijmyYIIHWeZvX5cSuf59cdZIQ4lwsxTRhb3Ieb2yXVszB2tiFVgy0QuBQmxz1rSvxXPx4h1cX/LU
xTcXx9M4lqV6871lvpTgT8WFDNalddtrz/dwjzRv/h/xVvRhyOFoQRRnebz47/0B7zv1xRuMv7Ui
CUHhLdF9whTS6FdZDmezAprHbWhFT3nDtjrqesnEfAKxYBq4BZzsg/LFW8xc6Axi3ngXETYM6oiK
pWyt0UR3Sbz2GHBhjsqh1YpfRhwzgKlUYebKcHprdNupN/SVxOXqI79vVXyga75b4M0SC6zXvRIk
ONkPNKid/NJlV8OQ8KKYpJiInt78ML8X5eFsbfpVSgdJOEOtM59QmEawJBOBggAI9/HAecRXGCWE
QfyjMsU9Z5q22QpQn2kF47qXY9fch8u/hdHcUV1oT1KnviggA1xJKsBecTjTQYNjVvEpJtx6buWt
P+W8taMZ9JgWMbTI2e8HDlwjdzvwqdgygQJ5invgGamAD4vGmyPC2J7/5r9lDz1KCMTqQuB4G/LO
U3eWIdgQa3tzo0AVgYueUwcybDMdOBe8tMW8LXSKWaAs1PzVJjONsk96tWvU1bmXO56DF18IrOa4
z+5NlkTNsHPIgQiXkZXHHieoC/aKy06wRAT5Iwz8gK6DsxLfTMvu6aRgyYOFpOeM2REh+vUjMsxe
Y5ZPi8O/s+AKRAEp4YOAvYUOaC5IDKfrZnFKV/V1D/AOcjoPeurI4gfRnsv++wFBwkpm00kOaqAk
rew5jrKheQyLjWOZVrsWsFeco9W/ex1XeZpq8r/eQhryVO8Kjft+7mAjZR3B8lZOBAH9iufuvtPd
M4RcsmlhXLz2oDgpiwfgD3A9hwgXm1xjOh1Sm5sh4B8KOpYYL2MDqEAt5Eq5lylFz5c5Mp7SJSyw
MF9mBHxq9Jo7ZfQpbt4si6hFptPrMZpCv7mvOJFPzxlx3AF4q9fkzKWRNqa7gf7M6g2u1saHDKNv
K9AOBvWYnzn8LtK5WtKpYYfzJGFDZ+5J7OgyRl+79Kv244EyEfjlQYEF1+s1SJHZcKzaDYfN8dD3
iB+2p8b5CPSIckrPdOrwv7Rd4jOcNTDEkhlNgSQFN1yh+NV7yJc5+1DtSV0BxJN1wAbUWpmrKZo7
0eWq8D1w1KHik1soVw+6aufub0o2ExOXOeu4I+d9bMagC+yd5cMBBw6wUjXZZGb7kAEVJ4qx9ddm
yO6W7SJlaW96MQY4xH9Lk/zed9XQ0dCiWDtcp8ZQHi/iqoRqEs6pDPLOv4mbaB4T6p+CMa9gdeDn
TdGfs+ogDnGFlncx2h6izuA0JSb6d2bMXbfuH6btdEvVkhw6vfSRi8ap+Lr13jJwYBP3+LM3SX/Y
brTWKsG4pRc/Dgq8RHHSkvNvL+Se5T3HS/UYs/eAsn/Yempu3K/4Lho67zi7fyZ3bbmuRlLOT2OU
gNJB5i0XerE2PpfzC340SeNhuqcbUEld74E3SJcGCEArPbh7T+WzhfXvlcn08i0OHYmRUmW8c5LG
awuO1sA/KJJh4G1hJ0qA5wyRbaEjD404QsY5Xe6cx+Z7XamsZJtxBM9LqEDhPU/4tLlxHxna+rEl
fPn9m+308sn4MzLonhdslkvEg8KOC7fuO6IFVGFth43KCDBrrGbcMGr2N9U0hzPcpkJSxsuGv64N
1ZkdXRB0T2hbnhXXS/vGZO07xDQyHKR7aQr6QXNgJwrYh8+Z/vcD+q4TYeVRZczQY+t9VfQ7pI/+
kssQdmXs9NTBPcBW4eOoPfzltUZ27oDKIFL4hj+ePp9RMjf47BwNBHX9eUev5RLKpMDYpTeSb+80
WN8PKrSPT1LWeopRVuYqgo6rmHvsq2CSPAmgS0o1tOfLLx5pqE3GjkM7lIoVXZQRz8Neq6xgQh9Q
Qh0EfGbfPBuIcmqHyqsF6DQJhfJm6f5xpKwX3DOuF1jBsqSce8RG8r1AxiSD0l7nBWpenB87Qj0a
/CX0+F2QjJhNcreeP0ioK9+GSoUU6mFCe58XvqBT/5FC5/Vk0U8fiklgRtxiRpI8GuwQht10kIVI
h4nUix6LKTxx3xTB/Cu2lAlxdBX9PtZwAhp74FL/CRHe5WqhUNN81zl1ZfacJEQoBPtpKjxhCaM5
L5W1a67SQ5XosD/YeUXO25dNdtIpC6gfg8lDCX6bj/UtTK1XWVKOVqV/GvQIzdG+4SD0HDWvwTGa
GmMtpfUdUQwAtZ7FlzYqcT2+Hm9/wuoBA0DIOhB2bup8qK4bLDq4Mk08c5kOr1FjV+8ayW9KCRHx
LmPJUiM/BBGy5EeJ7UP+Llg/xFIWmlFh7prtMJzMEc4h+ufKr81lCr/cqFEGqGW76Omw+ohwCl6J
rus8Gu9taVVzbzUht/U8Wpf2PUWzWe7/kNisxo54wPhR2x6SvrWN3rIQccs8QGfAoxtZDKYpnqBe
1q6J22aiKkjwPdoyJyr1K1aBzNSJfQK1Ay2iGdE5DCbsN3ijUHwA3pL3w38c3HBy5qEaoiaMdcvn
jj5vWJn/rnyLKb6zEOiPerWJSfPpcSrIfVqFXgCwcXYYoN+Og1L5e9Ef3Nt321M0QTotnZvfwnIp
4fAdUjKQCxs5FmUOpsuNZTGiJCPWlmgeAICe9QCGFuXwRHhetTAbsCbbn4BVYGK7ewym2mCrzfuV
YvoBk7JeLDPc0onzDSyzH1YXHYcOljupSRiG7Owv1JbTOdPkGpfxOclaiOLEljwRPSrx+QZpb/8x
SzwgeCgGNW2wyyoJb9OBIB9sGsgIjOWZu1ctjCxPmOOoKpl369yu6QIPOcPsnKRzG5b1yMrn7wkp
z4VKQ7462+c3eGPZygDo5XkXmVZD/tCN6ja2msk+JtBJ4JBoIxCE4wft7fzfpgJ/gwMtuoyTMF4Z
83BB7s/WqiGYQeDZxNWA7XaLSOMYH8Z/pmcd30vN5B0t1U9OeIv1BO9xQmB3WD7RF3R7QvsXuugN
QHtA+GnI0a0HS0chPHM7g96U/KsRdfsb15atieM8qS9QTaee3WEb9QVOWwB1ygjqG/bYKmXZTkgK
Iy6IzfJNPo5BX70DzU1GBH/jxEy6TW79vaX4ltwy8ihZJiwgcoSEQFf7xiWKeBD1RMLKY5m5qQXS
dPJsLHAw7l6mEYWrmoV80HqtWnDnaeIqsx6t4bCQT+dvTjoCbzOIKlewnLVfn0P8R4zuRGX1aZd+
elnHqZzC+LOoy8WBriDylpLPD4s622Wp7Tj1YUEtQoVhCeV8lzkKoI2DJQ5ZodNwkeEtw2uyAIXV
i2iwoybhEQkT0mK4s3D00gOMHWXJyYO5+wsJEtn7wBVk3+qJiGmT8kANHrioFKi8E6ByQx8r0CgJ
dZwK/tPH2XnEVU9taiOSG7LSE4zZXnTUrN+vjj63qKdpoylAVpCI5Mns90YK0mY8x/9PK0P9G9B4
fwOx2nqb6niPxqQrVqC5kpb1a03fsZWwunGcsqVesHeEmzSjFWy1axS4TEpaPn1CAPGW7nmcCtSc
aN8IN1Z+dKPQmOfpNyzrEIFwR41jBMeL7R3Q+dg1ZUJtO/wT7dEPoJWpGAo2S3cYmAg4SAPOwTW7
ki8B0GyJu53ZHq1UfhmkmxLREgB44PUQ9aTd2r+rAmA8lM5Limvfautxfps0Y4EEbIPaJjo8IaKD
JNRx+AlY2O4DjHuigVNwr7zbxr8B5guXg3ofXicwz3Xyo310GkZEBU1P5PEDUrnKDGrZ1ckYafQV
Vl/PwmL0dr4cXVfyE1/ECMVPpwlfiGE0DAkJKkt+9X3ilEJnCrjxFur7BxslPIiKDAwvva8cxNCB
lE8Ezzf6EYlMQ7O4H1QFSt01GhutSf2vUXkiqVQj/BE30u1h8gInT+LcGEPMzvqKC7Oi2IrBj2fx
HdjbeIK7fh/JccdVHO93cJWhcjTisteaRvG8FRuxLzvEP8rum+v2qjccClSnxin8S/q6mWIjyy4X
fpwQgSDycsrOTbbuMaDebs5CUHeUJTQbOcq8okQE/hC1yzeveRoouNCAJZpTJG2nmy7ZnMYHp6A5
2grH0dao0buQMFAEJBnPKZ26tl60Dw1950bDCCg2XydCijAWgLNk3KBzYPDVgVBaTZWXWRpr7itM
18spEo2oPldZXu5sFHEDuu43V47eYxUXcnUUN/ey5RhxRHDkydw1RR15q8W4mg1HHZPEZQTURn8y
IxcMupQMJKdh6WIot3g3mHrvrPGa6ykPShK/TiU4ywBOuVn+/xac0uVlTpKtUEBxx/bjmLdm6ZKN
AjnAJkxE1V0paUWUioYqzDOXHg1FR9ohZfGaeGELZbYyT4OJ+OkMAEb9jUAnjp/hCMICGtHJGDOT
633Ql6w17cZv45K4fWRn5bT+HjRCltzchGQ7o+Hylz/EtXFIMkZbThwMdgRkUunj8w3grUL1jCpu
LiNJm5UlBddL/lhSTrwOgEZCS0R8V/5GdsaATQvXIoaAObkSBNOZhcUSZWfJwaK8BqthDnJO5Zsp
tWllhz7ZMII7lk952U7GNfftPTahDdmXiXngVOzH5CqHVcyaOsgzdiKq6/S/LuCdCDWM5VqT7aCz
Wh0cEr6c+aPR7ZNmgkBby4LdGTcT05HseMegAEETZj1GSoqOd5Zwad4AvOE61yuYRt/LImi9UHpQ
4gfpGV2NCTVgqO767Df0Wmju3xxl3pNbE61lTtPOntSxuCyEzcbD1TnL1c6NdXmxHVEE04s/4ARv
eBHTVP/vCaf5iZFOIgWG9Hgi59UYpCHx2P4cE1uhHUnV/ANb0lcw2NgeyaXG4/a41npU2UFexxO/
n6xFi0xPkYG6I3zIcf8RT+OC+47rTqbjAu+pKMLrRws+s3psGqCp9BXqcgHwaj4KBLCSW3j0hKT8
08iaCryvHLCk8IVExorKFitXadunrRaUa364x31u9gcQ09VfcSxbCaVjdpKFj3LQ78jJ8DkPz1r/
F6hwAODle/nEqXq5V0GesfUpup83yhvihUgNA885RTQpyHQofEwHCS216MWfXgp/RVGON2rFkhZx
TIv0Ldox4U7C1nDi3z+riW6Qi/ha884JoYDoI/x6iZ5ph/i+fHwnj1NcYr7hnccUvlZYXUX1ejyU
1FFFAL9C/Mp3wPeiDbImmVw4wIHMhcxWPbzdyGGO5plkk9aIcxso9gPJ8JU8LjAOvzkEKVMeY44b
PiyF3cVYf3uwLj/x/b+g/blCwZ2VZ9rmtwxnhv8Pfcy2p8Jk7bRUcCnBzzppTF5w4M8C6rf/4YW+
zNg6zz6CEKYrNGRPBbpVe5AVv786je+RDm0GBx1xiDi1cSrm8RRSNKpu52nyccB4TSlF9XbStLQx
b42cwR8v/5/YlxBzv4APZXwKL7Z9/JDUyuPk4EaIfFeu+PANw+z7Wp9PiYWrFMFdSmiUY4ytf39z
Ei4e9DD2BUS5RMJ/xfpAiUuy8wIepgZCTwRSRG/JsRugVefm0B09uleLqfRjBHzbjUgVmjDMkSN6
1YnVqqQfY6/eBMcSnfGZHn18da1tFToqkaLbyeDxF5wRm5qy8U/TfhYSY0pZ1oKO8Mvoq1SoljhV
bjyhk1ORfUb6IHmihfj9yQ4XjiV4aJjrivIzlMdkyxTB5ErWWRoNaYUWrw5VaXmPeKJlSa5uMkGA
gCnmvjmHLczCjfQrYe37rgJsUXwvM5+dDFLuUbiShXyBkJW0XFCqQIL4uGwpH3oKPGlKyo0jvyN9
dB7qHf6ryyGxYbnjJg/Ruxzg34pC5deqPZUK4/zPPSibRoT2sMyoVca/gPVgsggJT0NX/gaxzn/C
vBGdZRBkXCr4UaWfqjnTEnR61a1BO8TYTtDNvRZPT8NKtVBcZC5sokWR1Eekk7PXpUi1HASYV4SJ
6je/aWPD+kHITiCRXlBtPIHS+wd3Qsk5/xfokXbneKVneJ/5gK9LuzCP1LIzMQx80s8YJfHCrk+g
NXkjYBFg9YU4ZAymokUz7eUGlF8ZvRRYP3PfDCTGxOT6ftpSrUBOkK7WVZgNaKYOoiFX1tq0kBpC
M9g9kHT3TSExnjqLvfsqY1qvdnK/a1RBInCh/C3q1PFw3ETdA+o/kBDIpFoDB/CTGRO3xq3twFlT
oKBotdvaMIJjmcURqVWwC2f3ZwLfl7B+Bj2bpTShV0Vihssq8jeAIvfY1mqnSi/klPlOhxRCqpYo
SMSNpQwX6AXobRwfxr/6Q63nGuCPrJFHRLQpZhG3sK3B4XdyyEyY9mAGI2LdGX5M4pbZND5O1FM4
IZ7uvoM+kH+xYQsygZqZtlcBz2yFjvwjqqagNYoKgnmR+8UE51NDpH7dvDgQBwsupNQh36nNqUxD
/3DmTzPtFKuZ42GL4AIK4aBouqV3CW/8m7F6bmeEMQdi0X+3ubQyEb/ONmdAXlOVjvvJN0fXVlFD
5YCuNO0alvB6E5KIGqcTumrWx0iqsj02iICD3C6fiiKZH/i78EKaWuqwF10E8svMSQ83t3FJh09g
zX9yVLWlSKhunb9exKvhODzvaN4A2wJCuljicERqe33KwYqzfGGsZAFWoa/VAAW4ipD/fHV1rqow
e0Oe0ilEB6eFuBKJE8Icy/B8kiiUQuiB/JijmMnl+jJrHuUHXeABb9bqBtiJcNwdOZ4J4yqwNZw8
0IeHwsHhv4/Sl9CAykzF3rS/P5gIK5dzFE6MF6tYHvawWOxNXnGUOvPVHHdgaFz46VZ/+Reu+AP+
mi/iZEEGCImaVC5Qnri4Fv8ed7sq3udITcX9MZqw1VJPU09f6F9QPjbRsu5iQedvPVD+ndeuNikV
Pjqq3Rwkhu5pjaxda4BWkPvAbqj3vE+Ct5W1niuod8iyuC5ySn8qgJ48MyoTFLEiLdlPse1JZJ59
OMigzYOfYlHvOEr7Y7EQkmqMYaMbzjihrQI60um72r7g6zmVuh5H5uEIv3EFgA52i07a02vWTkoC
lRq7zttKmOKRP26AmqVGhP/uZ8AvPOkjRDMLfffpTnARWshYCbXqFkltl1yRn5eFCBEZmJ3hRtJ7
BKSTsrrLAYuICmsyIpyof2VyJNwOZi2IrHs5ULkkmma2ozgVygxcT7ImvLb0CV3g0cfJ2GRCxLOm
jhlBL8LLlMcay0LuejE8Arfzi+FEzVXmsHp59xVSfMGmJzUAhORv/EOT6JooTNCBsD7gZzixoFJb
cAvuXbEFupf/nnEB/R9YLItWVu6moVM6r5UO9I8fOfMRAIH4oC91Mm/l9SsMrNy3jNVoftLGIUnn
l6lfLtyTgzRyV+8Db9prC4CWbcjr1JjlJhBOjDrxlUFoyvhxygamgwKII8X4l9vJVit8NPlbqrs+
y++RQRI22PuK180AtQu0b6sySM1XusIclrNI9z+SbiJDBapfp/Gob2EMpbEAiQCnYHpdBPDRA5nW
+su6yunyT0yNE7mLJcbykQ7n6tKy4La5kzePWla/RlLA6u33qNCD3Qt5FOS6II/t/86U4ynIkuvP
Px+G5OSgTQcpZX2gFSeYAOGZH2+ubgT7nf3fYmoyLB3gxcnaW3aYReJwiF1EC5zF5mPE54cPkGda
SHcdQwOD1IyyDD3sWDqoZLp2VaYeHCIdFc0CbfLX4pcplln1/p2ScyTNweuzz8AxiXCXCWiVPiKE
KfTve/mlKcs6F8mOktpByINyc6Csnc8LiZp8oOJUUR7qcPGwUEyQlIdvOHAAIPyXoXiPkojXnuYv
Iq7hNspaqUmAJCXA2YiOfKT0Okle0BqroRGF3iG4E15OBU3HjcRWxHUNLWMQo9iP+YAKyao6sKHM
NXk5N7LC/w/9ZsVEFyIut8kIXjHNuUlgIaLLjrzEsqn6PO7t8fhzIB4f3bwtViQyBKEYWzBWLosr
J8YTniJp44wPDxydcQtXOX1S1HnTwuev1sditix+ignzCbvkLKDjUWWWB1yaKE94xFXKTEhlEZWk
bKM0sAXnASVJXcw/0+tfQBwQuN6nHipXNmlIxeUt69P4cW8ecnW2vQSohGfEIuqC0QSZV27xK9SG
Kku0+qaeS34WCuP8fpyslGeu6ew3xLSLCp9tU4fTedXIKvEEMLadYE0UVt/hnt9mnXKrazaLDF7j
KnrR4k2p1hPQ+ixRmp12ZvbbATbXezou3SsdDb7kIN2gR2skn/9zKEtSRTCJOPONaYt5vzvRjpoD
FYOx8CwdDyFilmIELMfsqLLoOXL1UlKOGLkrMuizsWVmwhIWCk59Dk45CUksaLUXJll9RQ+9Ku9e
Nw8+UmiBSW90KSfb4N7OfsSKjqVS+MLOJiA/lzUd3XKNj/jeHAEQNUC126aHqM/j/YdztU+bA2Ur
MzL9XD910tYbsG5X9XjH5si8AkrM+nNOxuHSjcrmPnM2gD6LZmgUF28dWaBebHpB7m+Um27Y+I+G
tvqt2QN+KAP+lGTb900dRwXcQMNvzpooOjEqkVCyAfjvanUbx79WTdoO9k3cr8Dh+b7UEcaprMWh
S35kugGkI3siz3qpl78+cJt7wwSB+zFavMrGJAtLhTI6pMbJYFTdnAtE9VOHzvzEpjsdBiZ5JrFE
c6G7nVwx108WOHqLKaRGSZmF5WxKjk5QZoZdWJmo1wGRyiJ4xZ3yeG6UmyavCwny/hMPezF0/31b
RGXJElbRCy7eZiizxb9Cfq7oYo41nwqe8ozYjNYLu7qqpAAJxB1op5Mr3lPWWPuzhDJqBS+fYJB/
srCTH7dMpjF4F/suCrBkT8wVuWNElyb+Oqzp50+tMjV9RA2hETZD8n2tmEa7pT/CwZC6M3vsQvrq
AvZJNaHVH1ohGwDos4wZKynnOhAtajICIvOAjUWrE3f5/Jj3h1lDniBVVB9FWqXst8XBgaGH2lGQ
FgIuVycRWeHlQ0i0/RywVuheILnGUmQbNmNA1tPsbsVhzK3XVIzlEjKsgd3gfgfCzvoB/iFUWDlg
AeOYxVI8x0xlD3J9uoxH2+LDYWkuYA9i3JF5NFFEryUZrZY7ISvJJj6PFbITwSb97B7aHIOrfnGF
SDZMHFeAs4ZqWIdcHUvXL+kxEM8alH9XTGX19dPNs3F4/31eDz9vBfGT1PwEL8AtabFdoQI9C3M+
6/W5+6GjNWmwEpyhlNBOOg2lJjvNXQMEobPahqDwygaja84zURZ9f8QB7z28iMycBwPwYbecI+gV
LPmwJET6+NlnBUsRiGXZ7ApSwZqvlYeKLK9yOIuSgxffAFYL/5ZbacMPouxoIkGah4p71nbqLFzY
cLfrPpJ11ea5Tk8+PzmXzrEcz7jsaWp8rAGSfOfl4KpvdtNkpA14La8307TZlLpo6NmM0N7kej3m
4a4ZwGo26DdFsRLzbx4uZZ0PYu23ap+YOwSQf33a00iS7ZefrfBntI6Jk6EiBW2d8s5EcQ5e0GP0
QZ6hEBYFVd0/XzlVvdcyLnPs2EiPl/nhfiVl6VWppntdvIou+6gIH0ntw0iGCeWYISZ0Yu+p9uZR
c+MVINt7bpotxWKGa6BbuxSbV0kJGjF60qmnfEQeJ/UM65hqw3F8LKyvtgsnVTjHNH4vuoBC9AQH
qODHnt1z34LKohWbGGWr0ZJ5J/fBp8LUYZMJs4yblef9ERsqLrfZAoXmOCP2z+GEJHlNwq1zL/Q0
s5WQW/FYTGSwJe7sen/SGPxgsOlMzcohLkEb5XMo6F9l6MTFobUZO/fQjI+FgLZm34eW8F3j395F
XKkZre2tRu/KlwPu8if4K2JoU5extH9MuiTFwz4N111SScBrwjeobgm43wJXEPvapKPGr9cGmyvh
3oUqzzIxP02KUSIuMABX699+SSS9Dvf/vR6WvGGaN0wZedXlYpUCDCe0aia42QzXOWFUT3lb6SRN
hWJy1tyWlkaEzgOJxpk69sIPDjoKY+SUhFKowGR30JuHaEsVt86kBAHSGMe4uAQ+zgW0eUSbJGjG
wnN5pHY8qccjr8QY4SxmsPjsby0GEBKSoJ5Ckz00XX1R5hzK8h+V8p1ZbC0kSrH7LAzSrrt/BgRH
USnaF4+OpLKw3AxrmVdvYBsDvb3gGFc+nfz3FYtrYkRQvMVtzqRtLJvGi8TlKu8gSrvUmzmacJnj
dyefew5nHLlXeJQWSrkInX5mwqgXjZ/7WO3mjgGF6jpeMbXHIv0PCw1736y1NSqIGfckGvOKDulJ
U4LTpc0MepEgVl8aFjleqVi1p1JYtFnQlK6m0Kg0bAP9m2zNRZUv7CjqP89zkCIVVhA0cORX09UN
tb6my+ftpEP2F0YreOi3ROsuxK8VOqhdPQ5e48J4Mhs8JrPwHDnCmSPlDCR7o6dtxOpqF2x1fbuK
4pcSzPVzLzi+/prmQBW1r08ey+BbCCCvUOu8VDz2Vk7idNV361Ki9elJBrUyfiVXEngkodRMO8Rj
Y0GuH69lpVPqv8Ql7rmcOWirFXkZIpqt5+mkl4fNGhr0sduzhXirbZX9YtgsQYJ0VKVF4BATNnpE
2o9/l5PJlg1N/vjo+7Ym3U1gLSwrKXe4Cym81ebmwRn7gNiKMAIsJK7rW7G/BkP+UUK3DAauCRNy
o6f3tXcKQ59XhDzB3e7vX5BL56+Qi7hs6gyB+ySd+mW8aozH1X7g7MOUb6423DwtKYUs1nEYd+Jb
kpw+QU0wqhTYNZhcuxKj+JBMiFZA37tpYF1z/+07KpDtfyLpdj8Pi2xpyGkPhQ+hLyss2CDpNm1v
nKJz4gwZeL5HwFwNmLscuEKFnKqEBBx6N9hXm9d/PHnlox7XbtJj/mFtTPWqpF8pPM/raWlch8yz
MJi7KDurWbFNfLl3PIyiIEMIygHVukE49FBGkAWVrNru3wt+9un3j1iAUfmN+yQx1FRYjFbZNB47
QYS3UgwnaXmFZbIo5Tk876Z4Uv9RRr+Xt413cdgeqVUQeJDJvWj1wcU6luRY5K1jhA1BbiaHmcKa
VZuFwl0le1ekFKuHO1ru9Kqg5oGvGJVfIeRoYllw/BrqUyIqqJRAn+DQgf6NY8vTIrUY4gpYeJhs
abhxk5wSzQetuhkeiTWbwerdQEUlDjg0h4l1AHXS2X7jTYpnRbzoC3PTjIy18FmVHxm5pEbdUQfe
+Ob0kKuyQSu3pESdBhJ0IjB1eBLasdMMrRNdsthyVs0JuCPJxSeQRAEQKpvJPc8Mdi27vrQAByWO
bKCtdUgjrJ7dyTWt+QRyl4kyDqPQwaMGxueyOaXimin3s4NqD0kdjLmB+JTPqWeOpZ/SJM9Q8qoV
rPV48XWAoCSROdir3dRk/6EcNKsU0uRxVBAoeFlRx0gsq/xDmeCPSrLmja9U1Q1sl/Iyq1qzTcpd
FllG/hB8IPM1xgN8SKXMQTehdi1ndm254z0j0XlQ2+NYnHusQqxMfz4TQD6OIIbJkP9tlf+sgCLg
vBBxrFRIGjzJXfps/NrS36wgboEeBNkEMtih0wQxOsdxGYULF8tFvpg7D78oHUWZeTWaCKwyupPR
GBwnGdny5gfCQvty+h+T+vneaB5TgN0dVondpIzoDGaaOTS1UCAUwMrFeistKc70PX/qHMqUnfz4
O8JBXsdrIBFzPT+jtGU9A/v45dOzTmGefnJKjyyHf2JP8myEntIz/BoCy+O54nIn8UWbuxuDyO8r
1lyqFTVq6FONNa3zpaAW/BIIewMCWCi/YSGDcW9WtHqc/0ZS7CCvy97e64lJ0/qTmTfIRiG8VFOq
mzMhIJRqXLc1D1SJF4OxkqQu2UDDhJbi6PajGcXHcG/j+mT8yRIYF+/wCP6HEHaBk9bdQPejd6qf
qx/cP7vUwW5EToWWkebYd2nWEOEjSh0oKmAFWINk/zfSUIm92pkOUjcO7MB61U911AxywR2A68mB
SrVmZDJUv6VzTGXca07FVqPM9D6HLFrUFkPq0j+0fXNDZbXJ6N2HMwqQTwKO3sJzjqv0rAyzDiyV
o4xrYUjNi6NC313O/vIbzpySHTB74/ZJdXrpsZYvR2261jp93pWg/2JowHv3oBTz1JLu48jxfVWC
tuhqxhO7htZZlms2kVQOljpezzErI9JAqOHU2NTz6blc0jzOz7JZzKSDyI0gJMOtKSLB95La6sLg
xBsyU7zef0jQ8VI0ux9kGqL/1aqxODJo/R2q32EbiFnDWl5+Wbr2fZUf0sl/kkpJWHf4iNvws6Mp
ymS3CRuOwqxXVXJoJioUrNZeSKUoOsD9qSQylxYUEjXocgAKr+6LTbDAOTq6hDYbP6RWX+no4CFG
CZ3LRYrgXQHIiMOfYKHZWGSuwg/d5SPrljCVwIU9vFJQsCuDtFLelLph8DAao6fXpmqZ4fBpkZJ5
qh3CmD0Csa+22+pNxUmdZ1z51DXAk45Iv94L2fmXQJ12E+gcrVR9nQdrmfLiuq0+5M1INyIRyJRs
r7ruFmX31rcHh+SyxllMLSWjZ1eq7dnA4pR9/Bap8AO9X2hb0qc8mYGkOwPrti/A/bjM6F2eCyAn
ix60LPNt6cZAAZxF0ZD7sVal5aKSOVhq0nmDaCQl9pJl0EE7P497dMT2p71CkhB9J8E40qxuTd7+
t66MKVOwL8DdK8X5z+UZhJQO9+6+6LIJ6W+FZ/wEmA+M3fl97drv5wAjwGdFG3nIMFrNXjrKIXRh
PZEke7t7MIUtYK/uGCh8UuivYG6oK6IOh1+cs8mq+ZL+9HJwTzfy2Wa0l6hHrXQjh+BLi5PgHrHK
Qp7fHUJdbhPpc6eVF6CHDcmSWnMEdD0DcbjXnYDNKrXOXZ/68gl726dfhtqYIo4KXMz6vEbNU3+k
6RARfZqKJ2ehB5FzTAlmMikCG5IIi0ZChW2FQyqbUbAr/1gwUOyto/jx2r14BciWHiAyy1FKRdee
sl50e4qpkeEQT9bbVg3U6ASM7ZcwobBpupPVwqXjK/nc21qJmw7KRF4QuaBMG+DICmN9SjMm/Li2
85TMr7iZgHJUKfU/lxkHyCiW4eVVL3lzRvQ7TieJJbD3po0oXqwxV5OWlmeqvdop9gFsavQ+6E5Z
fPyOOmLScOmeJ8Yms0ro6cMAhZEmK47lkskeQwcozmnaYwCpef952/Vuh8k0OAD7RD3tAuDIlSbL
nDeCnB7HwCGG7BAobpiw42bmV5P9eInpLzFlK0EOog6Ae+nHecDYK7DuYRpQoAaQWbrGK+PsVyLn
Bm0Wgs4DM/LF32dmNfCipz6G8zNwFhJOebyAcDkNB72TkaRsUx/IoojAeoVnLm9nIy0ndnZP155l
gsrHs+A2lD4atMsQuVaSCuhOF9OM82pB4D9I52LtIAMdMEBltAQnPeuSlsZWDqwACfPTvUtq/lBP
eK6BjjDfL/x6hdnhDkrRssIglf1aKVEiwa+UBKjMFvhijOExw6sfn495vEnGGugn47d1o70Fbzn/
ziLZ8D/1inlNBnYnPmmlGn9GcLX8+Ed/MUnKYV7VofCR4Q8VmULeGwmOjX+Z96twuAoNjlmAd+Bb
ffq3UQCayZi35J9Fam1rRkUsWrrSEWWYtKiHT+YTMkh0/UHw7rrVJCirStGKm7yXb8ZdO6PxyZM4
EBC4FUmGoi4dSJVFdjl+2BnoynNPtzOuNDwHT7vAG+7CYprLZH0YBs5SI9V/kf3xBVEohp3cHxKy
MmxQNAREsiWSp7JxBEEIrrDY6uSUC6R0zSmgfkLZsnodktf2f4EyV1TjbJ904zpo9zAXhysCZjcH
N+9d/NtrDwNlmqQqo8QvCeVcm4dQTLxYdfAwGr+BIEf2v0s/FGBbR8R9h84echEOl4u/Y7VE1iCm
uIkA3JprkByxvA47MNO4QKRfGvyxxNNwTfi9G/sV83GQmXgVqSN/aV8CjuV/HiLx49nNsyUVZAy1
o8wePgGB7N6fZn+Q6iBgUbpkhM8DyyvC9DvEs7F//cFShSjO89eSGqtUg0aE9q7sJnO3vBT8T4+4
SFtj9UlTXfnfoZd9Qrme90F2tGiDtVaW1KAZblE/1rEHFhlSv6Q/23e0Cc2mlab6yoTYOR+aO/U8
3rFY7q0rSEDxYtQrmNEapLg3Vdc1lVfNjEQrPl+ykZ9qU1s4N8STVAVMFBoRnDt0H3djQuZhaf7b
iLnGGu3B+4/Z85XI50v3JPpzdNRIDOUmy2O4pkr6jU7pj5+1t3MdF0Y5VKr8yodz97ai69wDJIXB
Pwuwf+jdow+CfH+lI718FEH8r0+aMEJjk1ILyf6Vs/HN2bIfbl6XjgKExqfvXOWrOmdUohh0IHpi
KbttXfXlOWW7QJjrKN6QINoQ/maiT6ZYu10CTf8kBfpZy4NZ+68TUyFcqFTmM3138VD3o3NddeMa
CSS1FmlNZdsCVsXbgm1o25rvHUqNOWoIFK1B5kp0Ju8O7BHNPNtUzCjhX4dnJAkVdS2zLoySFJ8N
unY4itCVqeWEbkkUlpBFRx/58JdyFIm+LMHnMsiJn3XLC0yHj/gAGWTHZJx89a+wCaGKwN7z6uPI
a0gI49QZWjEDKXkTaQ97BNWbTL7pdk27TL+oCnQX9OTfxCmyNfogSoOPdfAOppKFK+Kve7okZmhq
9rnqMkPEBDBTnVqwo+8p+vMc3sGKNXhf8/yvHYpY/+bGRxXTkwo6LESz1+nIi8sklu85r4NqZvxI
G+aZW6866CARvJHNOsNdog+d/MIOGIeP0n93Je1qOcBWO6GY0mY5akRHlfqZ7wilQ1XUw/xkhLy6
mAjTrLnLHwXZKiQiAaTPSA7JEg6cjpfchgAS1goWtkq3bM/4epiYntQNOi9bPZfoLu0XfNgTEUaE
yMMCeTVlWmTRJNWfWdAxxfW5VaVe32MJxculOY94a0ixMmM7TRyUNpJdChzXiqQASqdioY75yoyZ
+JlukGB4Oc2A8Hr2xJM7zjcJFAzLqk6EILj3gIfTiLzqi23UtZBP5otmD+/EgYQtjXbT6CGkCzXj
oZkrytIsnZoJ0jxfp8QTLWxdTk69DiVuYulUeqTozZoS8+cMM0EuwGF4Dx3VLxovPO8mpXMVuWrW
m6gYtmBU/Gw2i/fOMsbX+y3ZIb3rKESDNaRi/MIokpSh0s8+UYGWQOtigr/sGKiDlVxah9Iq2zwe
yKmydQTbov3OzGVlLllt11jTOxciUeqceId+bAq3UxLRDtHSa0+qU2PjxdqJfNmg9Enxn+01YUJW
yZ909xhpLTsVhn5mL1tC0H9sZ63Y79Y01MvT0RpuS9u94T0DLXm/lbSga1EJb9aA7hM0c9tUF4aX
WtUGFdNyp31tkMOimSi4l+WVR31LxoudM5a0yzwoWw3OztwBlhr8zrtG/vaFGbQrlBSF1bVPPCt1
4Wxz1znUQD9yNyzjPswuPJ95S1KKrsLO1WGxw9n03g2sgeJVAEm3uATTtwaHivnag4dBM50bYDrF
Z8qP+EKuTRsEW///xSc2chd5cUaUCzl6zNHXxrWiLMdxguIZfYXeuuGUUJS0A59Kco9M1H+rme1O
qReNEol3NUm1B0MxFPCfcmpKdffIlMXKSNyjddwx6G0QGeD6c5oQIF4FDDLwT9qkl5eFEVKYswfX
qtU9HvZ1pGAdsKZnccaJyIem/GPOM2b04CJR3zlHehASN6i6kEgGbfpsGYptkBXfySJgdJ+EnBoM
1nJAm3rFUlshamQK7yk5jzegj7g51zdtJnI81oRw9qWP6n0iqjBDQWaz96x3vg7mG9a9hmlvTvd1
IPmSM7l+Q6eZ56wldubba2sF0qumGwlDeHiwECbL9qfuxJ6GLo+E7IV8+94lTRd2IM0m6H1YTnxx
q316m1t5/vC3Fg5uBl8Ha+CR+dq+MoCBfYZYgE0KV/GrQEKatK9Fim2upz12o4oNIzWGuX3OlsED
d98fE//5I6SLC3hXZGFODNkKUEm/Yjc7DcVOrbD43spt3+g+Bxadp/9zDA8GoO/mtxcKLeHnBbOr
I44jhb6u1qqrZR9Ap7W3qH2Fg/EaG2q4woUJeUWZ6LlI49UXpjAKboZBVO5ZtBvh+S3dsC6U/BAO
yJHH5D/RswooMUIfi9wf9RUKMv+DXrl5F79dXCg7wRZavwToG0qem9DwRwkIIpfA09dHgdNMuCAb
smz6eE38Ie2maQ367qeG7KrHhQcnIKGdRWv7zMv8+cxo8vt7uZ6WwgKDecDTUCxHXrmTFDP9MToF
pc7M8BdHKPSHXiZwivnoui9nBouKWwZbKIFGka9KF7pW9gyiXp5pzo6tR8V7y2N3pgofSVViPr+A
47E34uZqpBjKtKcqN2NX5UYGeBshOzu/nYBroA7fFmtBZDmoX7xEkyzwGV40JfoFjouVmXJdQnXM
JC0uyZi0MHpKwLeByp964iHIWRmYi5Q9gXaWSth2D+enNlEYZg7Igc9WD0AV6Hcxme2M/V7w6aB7
ts7UxAxR+uXKgVnXmOT1xf/Fkh/GVHKA58/zYlV+EDo/nrxmcRVW/wE3CFzq0st4Lj96U4swJA4B
vbKSYorDs78ESVaD/Pk691bGvWgHkQREd+oGW6Zm43S3hrRq5Tf3ursFP2x+BedAzgpXNLoapuVZ
63MEa7KdvH+NW/WpZrAqwcYeqTwHXbkKIpT11hRygjZxt9OKbBycdZX9mMbjUl/2cHQqp1+jaBBj
FhMlZVA/U57QM60Wg4HTSWj6Y+gE59rgoMTs/sfcUY28fI4KCvImtL9n16p5IUJ/pr77k9PGA7pX
w/tk85UWnTBbNl7JgtFyeTVU9u5vCHpDH/nf0rSKT8o28KWyuTHXSoxwTQAOJB4pqqTZIuyMNltP
vxcnAbmRkmsb8bYk08jhk1WzYRhGvTVtg/2r7oE37hbbhniLpMxIQ3y+Xt99XAMbKv596RECWODn
RRSVOUE/0M/mxP/O66Yvnb1ITd1yXlW9HWAthSwoqDfexzvFXp6djbhWzKpDQjn5BRsUR6EN9UkZ
NZhMrxvIW6/1WP7t2275FO3Cslqyo4xMwQFBcJovynFYp5n2xfyCli9Q/6NnaGSIYhWloNiT+rPY
m4FrC5UMkR/d2cXphCRgt0qgSrzJDomBSbAZbXgirM9HuKnwrYjIxU+55gsblZewtmKK2zkG+yOX
1V4nyC7vR0uNgbThxr6HTvPA9Ufz20DnT7CXtDLdQoQeb909MhIFqkAtGwN6LdkZ4hK00itjf7Rd
5QlWGGEwOf6lo1+xj7lwZ2i6sOdF11c8szbL8tkOgOuFv5KwUW+hJZEerr0oaqc3mZTy1B9kSd7E
U9wOHHGMdnrtK5dFx/C0Jr/PgRiIOd5VSk/0HsgLk6q0fEBC8rjJmTVmIAwuI5h6jIs3B9eVKfXQ
NvZIZv+nn8HuIFtvnJUxiDljkkgj/KJKOmpC/OMQ1HyLnx5pn/FYCN5qjj/53W8OXKkNFoIsg+C4
yosOxuYuEzjUG/f82xYehmtP6hojEiHrfUmhvE9shmCXEAPej2Y+m5QhZuOrUOrn+jLfthNhBf38
hb9rcu9vJcO6Kr3W4nSHXbprIHPQR5p1QQiE/KdLeqbuZa3nVAxlS3EGiSwqzJKYo7k+pMkJDagA
yVKTQci99GBZF7if+4bT1MpCR9hK4kXRbmeRPnW4uJTElNCzuu1BzmC9oOypi5AI2LQ1Jj/cn2pN
lR4cKtZp0VSfL9vq2qpeC16Oma5ObRfAguKw9ZAVd7ARCYeTQ0Rn9xfijVR1aSXTCEf0CpUiM7eT
7t1WjObI4P4vVk/K8u4vpdnXtWqG7jjoF6PtrHh7AxXePT/K9slR+g9MtWd2okgFXjW1RzdNrJyM
LucQTtMgG3VW9cTUtRWCnJK8SiWZpHdPXTzxcDB3nstDVuEzggX9nWJZ6xSINcY9ZLBP5lvSPFdt
ui9ygj4lfU8JZveyTWUjYyFngRnLKCxM2Pp/GLAF0alcZqrkHFEMtN7B0VfqDhZUr49OL5QldTBh
q72khhqJjLkhbk+A/ge83tI7G3zMNVfVPLi7hZoR8yvM+E0gaRMTyGaCv3u4Kqj58pYt8MTABsvz
DpqDlTTghQj/R4fAaabUHMh+Kc+Lx+CWfMzfDKNQi7+1/hWLWD3EE97tP6msB5ttua11sScVSWWr
4FAYa3CS6ktk/SPkY33T5NUim1tZuCJbZUufh6teYrMhDUvlSVZ3Dxz+o2OjDydTreT/5Rvxke/Z
kywhBtzrE4D30m/3gVf4QfLxSPDxF3CUwPiRmaQJgeTfvc+2xFltuMbriDRmxOlC9IOiHN9HTL2s
3pFJKy2g9piytKRGlP5lSJmJ+UUHbuMKrUYiBAS+ZAjyr2ZzdpKEOdV2pfkv2vVOYVpnFEcYE0ek
fo42dIVHsX61SPiCkNsfLrALJolQL5/fGM5PAdaAhfsx0ZAz7E4DDwhpIm8/tG0uKdXdJY8HOKMk
mexKc/6vcZjDd+O4OufncxtDEDAbensCfZWDsgRLxva5Pp1cSUHXkPlffunsFfeOXjQwhFxZDOAI
CnfhI28xQ2ipXSD+regZmTwh92Gp1l+KncvchyNNp91qOQTRdtmEqeBZhaO5YIkVRy9jXqKiN4YC
7x3/nYM/JwuBvAE19qDJyOp2NHXex9yK0QMoSS2uuZ2TXpUgf3UvgK6V96bkRtn6vfuInv3oTbPs
rEoHZpAqSx0ut1PCZwFXzP1+masNkMZ4XQAbttg9b6mXRb36Ak9J7TvQa7tWndMrM/s2sOjhxADX
ThAbXnBPU4bYQfD0kcIaRRyKdUZUXuLlWpDMzhNAxBRb8GGsS1WJwLbYPgYDvOb2PVUPS3JJ5bMw
i+T4vJclREqTNe8o+aRPGJkUTkmCXFwVRjOL+qHXEPdW4x3iU0/gAoyW5h8QSdzXa64MNkBI7GdW
OXMqATtZr4VseDCx8tUnB9mxwU1Uyyaf9J5tJOlJ6zZfF6q3T3NEknLdwYhln3eQQ72VInURw8zG
M/9dFwtxRFGWD9Pk63bTLpJUYC7sZ5U1C/Q3h2WaOwfEhYPRXVU0ZGtN5mP858YNizauts+RLViW
KE/+S25DZRreGfdgZrYYkiyurlb487sTPB5pa61kJ6vN685zhv33RUgA8T2t30pJLbuT95kW52Wm
8NeRAclDdFiPAeL3jlZhZwPbxpiGmN5AJ1OAI+85Paaj4iLqScsSd0ks/DY1fchqf1KbJUzkRWos
dS5jHskbI4uiJHGNSirlaNs37HqivNCNbWnLO0iVTEPk7W8lrO089eLs+Y/CfVW+ggYl7i1Hr8Pe
ma/0dIvH4zvtzih2CMn1vLYddySbBbiN81AKsFkA2D9I0TuHD4OhzrPj1kYVBzZAax0KK/VP73Rf
xiZvGk3hMydX92tMBN0ma3H6K6AQvWh5UB6z55aDP+CzMCMHvRNYBwkN+LW5Q1eYfiCyGP59j+Oy
thXzZ6zRz7/AcFmmY/xdpmzyFsrfyMXwwweSQrc7hq1Fkn13ny8v9YiyVkMhQ5L+G+aBWfkq1/BM
7G+6EZAj0FfiSceQGfpp6fxa6pfujCRMJ9PD7F2ZYf4I5msAhDmg641tKgZivHAahjQcDFTKDF1H
p8dijejIUgXvYchFsCKS4QS5G4KqKk7kxA9u5AKKKT+rFlJHZm6mb817fbKHvxQ3IYCwJm+VpiO4
yeD82mudQtNovpTNzeQatWgF43/sC/aGcWg+iKM15UTZlA35bynGmC7n1yCKuZ13tvh6bqipeCFm
sbqtDvGajooAV5PYfIAJTERs3VbF4u8Eq6UaavZRYdKZjhzmyAyCS7nUpcjTMuQDrl2GrNIO5SaB
yQA6WqhAyDFN+aUfMgGuPDLhk3ejSqR07luqAnIMSwoT4vOZZCQoC7l0xe8QsMvyyZhKAlTR0T2Q
p34g40cuNBRh1hWuCvx1tHHcwCErua8H9MLoOQ2z1wwUrDoN/lkVkuOPddE1lvh9F9Y7EAMWi8oF
7tbMAB9cBAuBzbqflTXoUXDyqekC2j4WiqeMPFxFsDRu5lxR6d3iRTQ/91STIZfJeD794HpIi6so
RRMJ6o/adB4uJRBlZ3XOOhhzh+m8nq9isSDLmaihLenWIRyDAuIK15mF1oO5aFr9Eamsnvqtw9/n
q3R4DBhaMj7mf5RuEgAJgsUqx/2XjSV18ohWYxZSJjuNfV7hXrHNlGhJm/nB91rWIuewqHBR4IJi
DmFd3MM+HYqavHmy7APM+YhRkXvQ0q9vlRq9lXJBAzWtbutete+NHtQn3dLWfqZmBtDEsu7WrFz4
hit053kXoxgL2jC9M07rERXFymgNpLGG8Qkk2/ADa9PT+NkMvfyJ9MDgXGLeE2ABgqm+u/6+V1CX
e9j4jB4X8QCiBECWRv4kRkdipqB7LiZIfcdpZV+KLUZoAvneH3OYxDzByHVPOL0qGABZX/58jfAC
0VHiGIlC8WxIfDX6LV31fyBvYGM755CJQOoOWDXKCkDypgPkFwvbb1JljYZBOj7LaBiW3UyMkWWq
0d1Inj/YmKostsaPv44ChH/QQEHAfKDFVK1+l3/lH35j6Pirk/k2IQAsaeYsUpeaIWfgjZ9TnS2S
MQw1V1dVTFnlWD2phm72DyRbAR/xZ/hQjdBXJZ2WWAsh58Z5e+hlqrk3fSEM/F9y8X+VUgwlqytv
9Ojd1GGT4mgwIYoeo3sEHrUJ5EfPDxCbyFxpQWO4MdzF+tdmI4AiAajM4ycz36Dl6sxFqlMNwPKE
R0qkldOcpiBImKEHqxZyDYtpBWP69xKbJcxLQOdyRxSU783kCFUY58aA7hBOePu9U3NbyRC1KSM7
VHpuA3N3qZitHE3Q4+ZH6CNOn+SjBjgdTO39a/i1n+8Wjhx7TMwS1UFfdk9/6V/KhYZVUQf0gxj6
swu6PhB+XrZlM1yks3YMFlsJOvs34PSHdk2LYtW3CqB7nUriLqCKQnZbzAHOpfj+TI93kUq9TcvA
sQ4unYOuf6/LVv3YiJhGv4TjsXINcf+MSpsnpR6CDB+Qp702qn5pmDlM5PdPay8St4dMC4meT9WC
oNRPcH4bg1jlON5j/Myrzwt12x8L0+cpEJiLL0K/FQ4v/0QnxzrsW5c3oNcdd938wt6odSvCxy/t
NCqZ56TXDutGmRH5suW7WtXfouzTix2dhjzE3gRjxkes6BYPPFa1NzeeLHA6YC4nbiu5MDaFUSjg
ZS3dRwS58Ssf7fGaBOkDeoPOeQQM90YmwCBoiqDOK4bm2MfJ+iS/h24j8EcatqMjPGkH06B156k3
Bx41swk7W6NEx8uDBOXonERTxWpOfgOoGBq0ipR62O6fBf9oLwLEKjwT7Cn5BdLtDXyC9jjLYFJC
EaB6GsdAoWrDgzdL4Lot0qnG4p9cpPhrN9Vobi3e09zM4jHJvWw9fG7f8GM24r+XM8deDSYrZTkg
XkT8CTtVJKpm814dX4GTP+sJxDUrLLLTPJRSjNXp19CTQz1QUdkAW64OunzVcaQyxhuD35ahqG+f
tW7hJpO2wanvdVFST7cZGoHm93mgkft7OvtfbSC6jJcj9h8frCoBBRwSnIfjeynQmaUe5ofmmwM2
BAKukGQyb881M8IQ+3SiJa97qZCXV/SRn4fQPQ6/ryDM0I/y9k2qqkChXkMQ3+PNwxKcwXWPhEmG
1WPS2ZCCgq/A91dx4GaV/G/1cqYZifyL+oGi6aFVWhWOgUEH003Z14DmpnXIp1Ojqs7DJQT6iF36
MSOLJ2R+ofSf+faxKeaL778P6yE4NEvRTmCaEukjILzRzkEnwbnOwxRELXAXqfip4/pvwu3LGlR7
+fOnkHoCYsstA0Dj2gV5H+arABArSRjejwesf3Ifg4tQod+mWBGwUsxszZnjG31ixtjCCIf5DYwg
yfV+JSdZj9l0/jLIbg5e7+aXwBZBRSMQXKXvk9GAwsIAeoI1DvC7LkkUaa+hP837HqbRzURLewFL
k04fNfFrhoBOHPvsnxvU/bA8PR0Ia+RrEftR6knxVsKZpynYbc6+Ypl5JbykZ4rexFuK7N0NFW5J
hRmlZJV23DiVXAMgqivNgyNdzWef/w9xlTP6s9TedTRBe5sAt/yTzxFCLBa/BDVsltOyRzYBboL8
TYYBdocPnfXlQKQrLERhkVPrsiRiHKJM7qm/xoSNX2PKwWP1oYqMJdcHME+w56qxwTVazUEizFZQ
BdIzgs4ojo6qLQfkGlenzxFVzgE7csi+k+sJwnBW1R9kWpyCvAobfpQymAmFmfyx33shUehizw1U
m+L6mFSNrs1M8eFA8gbS61ot6OSiaEM0Xid/rjVQ07ByoF+J+chh56SokQNIhFhoRN7HuLIQpVBf
99A882fSneQbxbr/FcblZQySbZzlptRyqC/O3nrDCDnNSLQH7AM0b8g6VhUqH4n6U8pUTFz7w/F0
jnU1XnNs9bhm9n7aSempSG7/MNKVaUk7IHz1PJXCqD9ecUAty6SEwpyj1B42B4r8UEiP02VTbDN0
sLcmrHt/DTzNy30erIuiq0fHBUFRo2VHwv7QUt4WMhckSQsfeYTzhxEG9fuAMDKLXPTsAWJWN32c
ezXr7VH9jn3zeAIhZp66jJmMRqYY1KT06L0PKy0GcBiP2ux/EkuQhU22P5qDIFvWR+VtgR6fdIK6
0uo+TjfwJKpAiyd1bYknqovc1URg2eDf6IpABhoLUYoD9CqRHxn5BY/8GgeyJEtNwUTjcy60aneV
7groYXPZFghbNJRyMcq7JFr6qrRutBj0IYvH25fHRLy8FJHTWqZZPUiEfjnVNL9Ti9lu/aGZA3qT
X3BadzoiHAxDyFNiMdypfyHG052HU/ijP3qHCR8xIKsm+vwghg//o64QQmq3LV70tDEHvjwyrdP7
ZeEzpnxyYVREGojtTPwhybHc1iHFmUWQCQ9QtsJN4O5eyPFh3LEpXC+lGBAmDhM9DlRy3swtFOb9
ijOKenoeG8xJIDnuJA09XrFOKhOX0ZW6CdJeGPt3VzBWHhkqT/qmi+KDhBEk4xJJUtXk/xeU5/oP
VCLy+72mk7PsGZj+D+jhOQ0ZyjLfHq473awIl0++wURASIz9elYXKrFMTP+vTNckBUMKfoiDj00k
KOtfwHTmyhaySDz9yJKo7sp2pgRIECG1s0BA50EdFdR/cBGEN9tIS0T1oZBsEpmX1ktF6IK/VCpu
jvTjbAdYxh4DazUhaKUDW5du0bloZRcI1ZsfE5VLcmyE0H+HKaVjAZZ5b6YI5qWfo7YjBlzMuNc8
Bqp6UptUtP5Isss1u6wuLoJsz/Y3bO0Y7n3jQvnRWQj3t3xaZVs2V1hMsoLuPlnkPrbe3Qe3eBc+
HQGf9HDV/Hek1M7gTnVMAYNrO2gU/hpU4kSDQT5BchlE3lGY8ZG3x6ZyjwKkygw6JQNzhDfC/XGy
pEDfCEJssXo7a20NfT+bc/y34pLQaTsoAd1lZyfjcWi9towbmnDMfNdbzwYX4uTzx4v/Df56AjOZ
O9smSFx6cnm/21wef1MBkWvfFXx3zqkYK6LFuXUeiXHG4vkp+ujWGxOoLfS6TlHG+3k+YcGP6eU1
iwVA/fCat2AQHt7HD5MRCSvYUAEsv2hzJ1dvFsWaD3vNMgp/ddriDb4WebijSo8xBaEaDfsYuuTU
Dhnw9/mnfyygVuddIDmxNPey8g0SN2wC6OnWUtppu90rbdWvJny0t89WxzVpGINC/9fTrG2pfAVD
96qR2zQ7r3/N7EpCcmaP+kIYcHI6DSSB2n5WPz/3yMIV3b5gF9br7pSeGL7UC5r7hAcjE7/2jjhw
XhaQTOlJlMJ8c/3pDSEZj9ou4+8tGs2aZwrZvJzmbFkdQeUJwJweD1zSRa2XqrxfEHxbm4B/KDt9
Wd895MACyFtAdf+OUyUmzRmnIInzw6ODSmLq605XMWpxeNPrTwY2btv9Viy0gt8wbWiUXqa5xPvf
EbSlfv30uCDFXTQUvBA5Xmpgp0DPdq/xw0F8TWuNj7rpIynx4gyLyTDQRNtUmCAv/UjD5dGFdL5x
KvHzscmLvhVu6wp9CVFvo1dRkqUau5Fe10dIY59mA1hInjcdBwG1CR5sshvjqC/B4bTmPqisxxQV
g0DMm9mlFL7eauh6egV/7TWLcbEcZB79dtwWCW+CFzgZHHhD4Bwm/A8sbiUHCzBRA4dEUeW+hgF8
feUtOzk1iBuOONw53z2clEqnFKmR+TzMXFnaZ98VQwvUzlAry/z7Ci26iPDFFhqkmrqTgR174hoL
RFJlzPpXoOzWSWy9EpSf/x0Rxw5TLkH8oZ+DUPIewzm8ipjQKMs4kucmbSsbPVyz9UgpyQ/Pg+We
mu/BGIyqZdqyXOZrD6Dd2RZTzZZIWSyKDUlWEfjtCVij4+0p2FGrOIXBvDqSIkDKNcmQVzoYYu3a
u0jugqt//RjNu22XmVbNnxrQ9usaG3TrhtyU3TX398m8Zp/o/uU0e8P0tNWjEcDnTfiz3gD/LJ0v
pMy+e8hJPSpjKBlD8YRinGQzi+apyEJPgN/ZSxSyYlyP14h+Ne6W+0VC4ysLRdCUa9HBi4c2or+y
aBMgzhXfHVliZyg4/luKAW6SkARfzAgtnJLa1xqCcEFKOZiduOiFM7J7ouZXs+LTWYj9VTwI5RAG
7iodgpEiALJkVblwtewWwLHxZij9o3dHwpP4bX0dhZPEn2JfKsbIN8/n92iI2C2sEnEJVMkN2678
lnhxii5deQQKdBHj6S4QX/7z7G/j5bi0HvGX4nAC37uqRJrGurCtysJnuFMUrOt/UBjp308VHR5O
AgqGia/v6FLIkceBBH18TbVgYHI8f68ZxKySWipCDW1uVzTN4VGR8CcElyCVauN4z2KzH/5TFtm/
+lDhwBKdovOGHfcB6qXYGtEPHCgpy6c2QhiWZ0HiprdS83vGIiwqZfuCuAdr5skfgYCLE0bVj+wA
H184ai9IFqsMVAwiiV+2euPN/zuMfAYyc3zDUAU2vGqDbrSZWu2L2B7x4dDuR1ksRXEfRTxs3Si4
CRcbsw7XKQ+7cIeTtobVh1zvGOCeJkdgdXY6V0lD5yxy2doRVVa3nCMX5LTge1Kg0N9OD0PKEaJT
NhQuAyYbFFiXZapuPV5PsFyafrnUDqE11y9wzHSSePN05o+Fc8kM2PDuH7xvg8kJDnESeXhXd3dT
OLt5cVvuuOETKxw96KBSrQus+ft82+hV2c2yO6IIUuVg/hOTav0C4Tn9fV0SCZo//5lxxyQKq1Pz
4L2tPQF/0GpdFmRQ5dMOLd+aow51KRjcAW5uMCYipsWa5gkrCFO4w9Z3ZvIcTT6S9mp9TnDKKrHD
XETNxvMrR979vO3WUgbZQxrF+29GxGsNFlfFYbGgqrYKE5wLBtsI/Ew90hhfHuvT1gj4EAIpn7/h
0xaynlSdrRK5YFqiKzC82NKwAQwyK2Z9/nRZ6cvjVvPBNa8tnBMh0moWfe4Llbo7GRjrvFMGYVi0
0Qv13Xan5Fe0HB8QdbnX8iDaISNcm1LxjT4hl/Am/75b4ws69EOVDKdGM6+BUlQdd2oO7HfE2P9V
CBG2b7Au2SNUTgl/jh+S5GbCBGjxZ0ggGTRx7aellbALqGGOUxOUe5c5rf73WHW2BeA787Ql6U7+
MDABUs+/txQbGss3tr25PfAl85JkohCa2HaKZOUQBZq5RM2XA4ZWG7I19N8e6vJeIZBVmUzhgOaA
IYNmrWPf67lO7RN6P8MP87PRao39YdQSpU72iyH/wwOzBWRVuf1Mr5CSyEPIHJouDgGOmFPJUApn
2zDI94lY+G6nAaXnmTCWB8OaL9jpC6JwWX+pmEt8m104oI3SDV0vT4fBJ4xqETzKCNXDOoz0054p
7qqf563KWIgNqL7tNfzbp1y3YyWWfIKEnLVpVTnY9/hmtZdMJOaSc7wo/D0He5TGm/7tYM5X4oa+
jXvo2xWZtnP2HtwQxdHUQrnSWdjQVLAK2+eVKmkVuRhMQgpTyUGGSp/Mj2Ry+DgNJFI8HtDjZskr
xFfg8M47ZAzs3LhSfrO+K6OEppXje+NzIJD3kOd7ObwY94TH8x/t+wi9VjqDTkX5Yup5liPB/Tec
/A6Z47/wWtvtba5yyrUnzkQzwJBrcF3KhsqFVCDzPhpmAK2RNwSsZCYpcxSLWdL+4iUPEP1N0Pzq
RNBrGt7OYC+da/P8Sz/yy3CAhnJmB/Qthev++9I8ZICs6hUo4AEMNxP13k6B7AyH99ukNaKQrIOh
LnXlf0fWnXFiwwey6NyoiXu/MZ1LKMedQvfFAkh0ZwOhhVaajY+rLAVZVwImP8rRoF9GugVBXN+y
g8OACAVmHyAG2gayaqI9Xmvj8doK13T+jDGJnnddX58uDpGb8tYI3K+tBO9jlT3fhLQTIQQ+usRo
OdLN0myFO0AvwvpuhNxGezinIuD6JRM2MXv2C7NgYFkrOVYJ2YBzgsjX7V60InWfFzIEC1cBGg4V
CRKnSVJkx0UA8wsnLfW/jDWBD25WgISp67SCLHc2x2JedMr47EZVhPe+gYJoSK/iBn2t8BL+ayr/
nRn2mHJq/QWZpgcoWuPMOcrGOmtWPsCtKT+VKwD5FNAsEjsBDmne7skhLVcQNegJq78ZOZlECBnp
gXa8Dr4YQrBNxIFoTV/mnQdsci1Er5NcNkZ8oxaOg+jQGJQQeRZMQzkpvmoLhJ1Go8aMiHwfeAUo
JlNUABXfv0YdcPsdZL6yeDZnFA+S748jm7gH33jBPfKChx9m2ym237YmxWpQZUFgY524XdK7dbqj
m8DomebgVAQHH89pBb2b3UVl3bf0yOJLN+Jv2E/JSL9PWoezTG4Bo039vGrLJcUdvecmUmqmrzSr
6KQ1mADhcChXRRLA9gn1pe1h9Ou0uGHts/maBJfuBPE7pS51iAmncIqFPgLaym3xcOQ8eFQIFP9g
jwwtw6Jo3Uf2C1C7XWbjSPyTjPOYYMusmEYVLOI7nfN5Ihhp4s634yDImNJkEJgsGM1sthCCdnzq
E0mf42pGyTTZAd8Q4oFb2M2IKtPUdLZVQJIV2xOAxZkA3Cch0PcLrpQQ7SHwLuEKb3DId/fE5Tnf
1gusU/AjH3nga23YodhpNJ1Ngn7/sTUDj5hMcH4v49x94am2ijauAbPf3uBVey5Z79pI5PE1oe1B
3lvZdhJoVttPx1NtAOwDH+Fui4sIXO1jRrt1OlOgwg0/oGBcn5DcMreoHhKeKT+WrPeUYyq3cU8X
PfRtW2xGzJFwg/y6SaB0mwQbtxjhFe8X9QOlI3/fhJqOa2RxI6ADSHQrzK6aA3CeeAtdHx3GxQ++
g5jmkh67/I9ElaE1f77DYq27oh8M2/7HNPdslAakRHB0hgMJyQoyGjf3TbfkSatfRC7XI/CVduid
J+MaQYIAFonFUWR6Zi79wrARUUyKWgRN8biCZXsozXTcQCXYumFSQRecWh7RmwUYSf5N1C/wAX/O
I3x1h2pMTqXiTLQzaKZqJs6iAbXKIqU44wrMjOkNXVZ/vMuRYZ5rOZ6bLmtPnu+I3zYge43jPeYr
OQW82g4wm2Ej8kJ7q35kL11bwggY+e1EP2GXJ/E8TO+SS1xjIL3vNKtOujVJT1m33QTKXPU03XNx
O2s22qMs7jVNdjtmCQoGGR0Cjb4W0VhwXMQywyqc94fulAdyx6kzhQ33VbQfyzMFpibge1RF4/CA
IVa1+QUp95XDtL70gz+ZenOvt88p+uiqR+HAPLDAYWJ79h7r4RoEd6QlQv3TjF5yrBQT0z2HDDTc
qsQ7dP38T7hzixB8ULOeZKGuSgXL8FoJJZcaJGSc76z+XsLextztRNMpourvN6RQbXV0ERV6bBva
heI3YUGud4oktORvKJcPflov+OMtEvWCSKTPFxPUjmDkCB9WPE3GidJXJqpWtBlRseEPOzkgLMLq
gMbvx13KFs+hCa8S5lqZ8kYRykFmn+sqPoTofwuqxr2LTkbknd/iKPHOg/bZ5pVH4nGFrx5uc/t/
XnucK/SaFkCi3iz3bw3hVgKUqPLSEslINA9sYsgQk0vcPmNhG0KbKibwtifgeeQftKr0ApwxZyCT
RgTnD5DljtGna28Qfd4+k8PhmqRzfo/VmskH8264A09j3IbEOvH+tDbSuOX4UH6xpKFCRIA1reqz
VT/G3O0E1TfiI2ct0ZS717slnOjJ4EKbOXF5xZaJNU0hVfMCFc3WWuY/BlAVobe6j4Kydp6ZNA5P
+WS1HusDaXBsdejn2a7tVivYbLtXC8DVH2ikHCcWHNzKjZFtVasnJsJXGP+iHuyAjMH6XGb5JG4A
FL/W65pKN/G4zOwDK9oEMkMldCjlIvpmQ11jaB6VqWhGhrRfDTmZBlTsPnEX7eXzlZHaOLQJL/GF
pH2pb8P+mZ88a+t8PIlNRCWc/y//MD7NcaDk8VmIs2/30gX9QV9S6Z5afLD7xNaDX5BeGc0nGhYQ
3SEVF/ULO5hwuEYqJQSNi5XxxR9rLJjkKQ4TDL3nCphg34C/kxeBcOrnklpomoumxzg9gInpvoQO
BkIq45UvjedxnX9KHO1D/wQbJWYcS8rQEoXmwpLnmXfmxRoSCPCjJVnKXgvk3IkknDpY9snc5vij
7L4k4Yp8jWb6BxDCfyyAgRdHgsWgqQrjXVfuHqHOSsaaXRPuEZc3dSopdoJqdGh3aAzuMRzJR0x5
5kQ2PCf22S/LaAPlocDfmNusfIZNdYgr5l3vqouYH/yP37OL1hB4tV9TKncytUbrUjeE5JCoVFbf
dZmqUn+clif/N8+LuCiS/WkmQDoa+a0aZCzfWudwiVg4oYmsuRhTF3IazeysR9xXphmCa7MR/dVo
DIPYccE69Ke4pqNADjXIuEq7xNwQQmt/S7ZwytFmXBrqzdIL/N4R88AP02OHSc3fcYMQSF9W0yV/
T3LrJg/GsM8ujH22VvFd+H5jrTBSWH2lLbexKgNzUF+RU+oMoQKMwUS3+u3izwCgTqgVvYrZLv9J
oUhNTDyeeZEdUlB/s/hASndfgCMiCSjP701OgfSDwo4ToI4Qe6+fX1IzvHGJdg83LpXwyExzMJ9O
ugrhi5cydilRXwXPrClh6ePamDTskhJXCAqDZus6q7V1+VJQVfdQ9XBWdUXJZy7zeLU9XQNmLuKD
McmaXN9M1/y1uGeJ0lG0egHlua4Purrhy7iCfAwd7O9bhZgZHcsq9U+y+iplQ5ko7E7B/vaSAhBo
E2BeflAKiybQa71oW354fZe/k/17CFZ+BmydfY7bhkUNe3807N8fRDaYRZFS0mwilQMKNc5ZrMsZ
BLcn1V8wwXKaG5esB3Gp0t4eIDztGSwrNJwD4z4pnHGyXIUY5dcSzYGppEjhWniGwF7e06wjyf/a
293SjRXSwB9kCNzuTamgZZTcl6yUMaEv/S7xab1vb4G1MzlR5+G5g6j5j+rsOV5B9xO+1QkIvCHC
wL5maeRXmO57K/UqeXmBOTaIpHGOvcs1QTHbolHamfVaecFy9iNHPWzvg1oCDouebp3xuhwbgD3x
ztLAyCzW/ZREfEPzA7ZbXWZzo6RaHXjSmte3W4+b7kIOl3sO2MeZwiJKEn4+B8AdcCouZzkATq2G
wsrFrw19AEDm8yoRcKb2bvfiGqZBCuBOYj3nLbaZLMYZ9qhpja317dXQR14KHbIs7/QMZw4bLY9B
XxfWhdg22VEBIeuYC+kuDJYedQcRWsqE9Kf1lFZiBC1F4r9NMjJSmC7aZHXtMWrlOErzLbdCt0zP
oTglXUhdUuCtrmGYE2FAg0oWQmW7Myp7dE7UCV9f0T4hmWTcdBaC2MBSkZDLX2SlnEYpGguT0Fgd
pjMEkoxpaWljcllkXazyl6/fyY4BO4iAKZhMiQ6hVlCkhj7j63P/LzqmjutzCOtMVBIjQNRg5TWw
piwwPPpP8vlPzgrVQoMnLOJ6pxL50w2sKBBawgvUZrl8/VmxLvDFYgACAG13RvLEB7IyZ42jLU6h
eF/+nY3byrsP9CQcN10YjL/LTJLfq8fQrAvy2CkYA+Q6SbBN2f9HkkyM60/uSVajhg00oEufo/dg
WKFvUTaiiPBjm1l9EfzIlZf9E8BPxNkQpXV3zEJb7ofH+5dmGhfEftWucdQq5g2WV9gbiqvoVw4T
le7RPMXH5A8ZJ/RK9huS0+rczpBH7qvntV8uZVhgD0DHgyXTn3cHHtmA4sYLjAAoQZl8nvk1hSrK
PNZyc9MuWYdz1/KuAUH/CQSDZ5d6aEzKiz6m5DhldVR8SpXm2JEnUJQbGKHt+rKN/3DBTJUk29++
rtJ2Q/Lc7wNGkPY2ZWojvMS/vo9BuZboNN6tZR2ltwkS+/5OIIRkamukHBMWeumyeT/okKrgaq7y
3H/zO4nMdHrfQIWlj9KwGnQ7LxSdsXMAm+51CI9U0OUKMWOLLs2KcI+BjSHSnrBHzaCwBCHggzNR
rcFTixF1ozykDSL5Ov6DDKC1KUQLhfUrjckZlhh4A2TEIKNzEd2Sy1riE887wIB1QA8ZkAvBeiik
rnzDMtgY6y0EYZyvP5DkXHPbe/p6kQ1dqUIXQ0X1zbxSpJfwlaMBBtD2ZlHLYbSY5Z9tM4pmbhJG
R/1CwQf78oRNojF93+BQ0CQKxWW5lLHcS76dIAToQyYg3kJmi6k9mwbjnTDuRLqxVNLqtERnZYCE
8VkWK9QDRgcp4gAZLhfZ+4FK97GTlhnJS6raGvixodJXTo/nJJYOT2OHxTW4IzDolWZtiEKPJWfU
TqfeZdeRgH72PqH/ALBqtlrWnkPzzsKCPLNb3AfnMQzJ7p0+mfxVegqimVlMk4uFxfYmRM87PXef
7f3L6EtUaA27er306P//2AniVRCiG0naCDuVxTg0+tnPdDwaiV0QyrOZo56RWFZF6eY05nQG8DbH
ajSHZ5cbHZwU7fwgr1cI2IsMHvXVewcIalvVHGI0+J5lWnI3yKi7nw0pV5uHrPJz6keFhWtaANja
s8hRFt/dF5fzrlaQelKCM7wEu+u94vHQf8RSVsMfAOtXXmdWn0bTbfE0G810COUCSDly1DnCRdTP
1F1rlefD5JoNZGV/OgRqXRJQpNqxawrbBalXRW2MugC9Xil5ugPSUQFG4gFlMa7n0RGwGVcK5Ph0
vn+apVdJVe5FiOZLlPX7KGPO/pn+ysTs1XeKz7gb3l21FC6gAVDRrBAh4Y4J5+ZS4kiendBqmxiJ
xX6qDxSh12ICWN4i++bxaOtWQ3+YpO6EDvJ9hPBAK1ieXTkHphuuuqqezbTP/dc1sHwmoQbdHAt4
ulJTJv7ezrsYjKMHGMDJmqpiDWZJv4p3kcEHmSXViyVsfm9CIWQMPEL2AIa43p6xusotJJBBB0GA
g+zqTJfVgHmQhJ6eIIxlBG8sL1xa81Jle9BeWYd8HPjSOkGqqoHW5a6mK75mI0UQIXFg4do908h3
fYZPUnYXfUpJ68LL/P9FABjhjnpcWJSfOX5YyHzIb0BIoOUIpEpT4h0JCyANBCDZsuDK6F4WMg2o
ACKT+x8GdTIthseXv9fxmifVIVZCKQRykpViEBTugYh6WHnzXNbLBaP32mnrXECi7hkSM4iffSiC
LROkVOZ57Jpwxa9XsEtkP9pS62hmZsEBF3KcfYymU9djovSoq3l3bjTSb2QvVxV2QhkUiVHu8RMg
5TDczecuoFl1nmblql+RRbp3ULLRvdEp0EM55EenefwJisA4IoVjHSwDp1FONubHmsaaSfliaF5p
L5kHvyN8OPWkqAXv68Ygpk4Ib9ulLLNTDU4tWDgsjd9X6Ln74ISdtnYp12hGciiMDkDd60lLKuPg
+tZuGfaP+7BZ8kQUQDzGpQSJIIMvVGmjXbgDKhOCHL32s25PDP6oja6hfn7RT/Lei1+WBxa7nK5O
H/dL/BhoyElNpBO+mTZKu2h1O9Z8TB2ntdFM3DZ6gq9etYWgMG50goMAkeOuzxelokJOtAOjM+Dm
KHXf31x4V/BnRTH8g/jPafjlVFC9D9EKFY2VRV4MFmilRVh34bSvyeJe27M+MyU5Dpb9yNNylDgd
7MIpCKLTdQ8mXLTviETsbChMbsuucU7lYJZNO4OoeWVzEEGgq7qzG3EJbyBEODUZtA/Eki3vOARC
8FzAn4AWetGN359KOL8HJWF5nqugQSfFw+mfJ83dAzy5lA3lmk/2PUaIPY9ERXx7mu3EZvyXzV/5
HUmjM7sGok7ajqeagA4Q4g34Ww7krIYQCzSKOc0TA3owaoCplepi1I4/DclJ8ksDo91THWhe08SE
4hYnSCXh8GPGarRjW1vaJm3BgczXadmjaUAx7qQBQ8c4xE0vEnEHI7wM5zYx+o2IDDC+G8wy8wLW
yUkgWeWdItyouCpX3jbnHta5YSYjBcqawVRldAOLoAmIYGSM8RHQDOSPrc7iUIwUp7++0s4awjSu
mbtKWbYuOCeIKXlOSn77JLtCBtP3A2Xv9znhpB9O2R+7uSnu0TNYLLhfkjKzD4jliDomkvjHouFz
8SvpOf+hzyqvBbr0IyQFZ6c16WpLwjoBIh3A9fO/+XQ2Wr1tYBNC0MJeu7hIDCFShpGViHVJ5wuC
MUJRy6RFbiz9fRQxj9vTqdyVIBVwKnJV5KotkxJAsqbXM1Y0Y8Sp4WRqGQBVRpCXTjr3y6E9J1Am
j6Sqa3EGmqWErUfoaa/7uiexnCeoX42EJrCRjuFdRebEwdSf+T7u77Q66B7EFDNqkJ+Umqz71WC6
9J+O/7hmRK36zsLjEEGg8YSS1CnVpnzNqFeTZoXHc3tOGo+RcXHx9rRLN9705Ydma8v5z6oy1MrS
CGZ9tTk8i7nR6lOkB7fwx9+zwrMKvm9sQJMRU2LJc1adHab/7qAxlSaoRmJU6Od4VylWVfc1sfxX
oDTnS44CL6eIhEU4sOdF0IU46oTPTQceCzmHgmcaCIrdIryeeWOmeYu7gEU1aEAvphaS9+daTO2k
i1KQvOAa/HOVo2nlp1TL2kUjdajAu834K/uyVir05Ava3nYR1jqmVAK8KXi/ujSOnKdcdCRkZoCA
sfD7pxf3j2RRNVm9dpCrTFzFpSM53WgfuAqXrJzirIwNsKQ9z3KTux+hNbVbhkuk8T4gymNVBHmu
dWGjPMY5GdFTRtGU9H0Le2mfWQA/Nag1LA+N+WY2mRxfcMESef+ESU3FTIfqb6E87uEtcQ7ch7+v
cilS3rcXGqQyJxHGJrBXgyr6usRm/VsuN6Aq8VOEM6isJyl+agPrK2d8hHE3fF74NEoQujCSwXbv
4HFfOJ99F28pikstQDLQgd2G7XKKpD4lHcrn9x1cO1uJYcmcllenFXyPvGQs5Ie9GXTvA/ODc1Jv
ecTauGBS7GBvE9LLI+2ZRxpJ4G4dWgceAY/jogqCJwerqRtDsDgGE1slyuZYVwjwE+EqRRfhqU+j
rCxZgu+dWwvtWj+vJlehbs447RaTrB0h1cBykOez5qYT1DnGraHKVhS6rV4kVAXoI3Wv7/ujEF1C
iyjodYJn7xVl6Lp+C2CQCkB6gsMzE2sy/Aoo9OcV6XwRiIabo5wDUCeSB+GcfQGsanp3u30RX8/8
XU//nqYVkgC2QviTf4K/dNGjVzhnkVWhWycnxpgLtYTD/ZF0z1CaZhMkPBEFEtRyndulNxJZV+nF
h/IHmlTNxVXcBt6yRc2Vs8bw0okdXD5hppuBc07y+hHXQcWE6gwjqQHj0j82oFmuyjbzDKW6OiVR
HfsFN6S5A/zsOgs9vNvSsNbPQgjdotXPMj4lJJ6x2hhbzASYyS1Vbi2l99bx8+PmiRPyrBP506CB
adSc1PpKPvVrcFVOm8vJtO4Mmvw0/A2tDlWTZIo1SM2A9c3WJ5gvKXDuV1S0C6TDNiTKmB4jr2dJ
vWqCwdPTNgJAQZQpf4ohBYvK0AjazUCtidSM/Lc/wYRbpk+9S+zX3R+osxo3FblXbyzMAgzrrrKH
NGnskAdmS+WFpF53RYLEVj2VatRTWTVkvip98A66GluHBg+NNlgyyXO3OqABzIpHXifNiRzVDfUH
biy0tbac3R3WsOwo5jqihtRmoi3lvlcsRwj+QGA5wks3j/M4XlExwIzJ3fAa2PcP+EAr4q43jZBz
touwaOWG0l5UmbUCPWrRkBNYsqybGPPtgucYuWoofTrgCogzKRCTHTqdy7aqulc77ZcCllsqBSb1
l27NjL+goKYFkYhc7UthY8Dz3M5DHMEF9l8AJ7DkALepcQvH52kN+333FX9JwoLB880WzmJH2+GY
2+BeFin10SicpH001BQJ6xmNEJx3hOk2jMLavVXpV89FugT6GOksNH9WYmmIydl0EytZ7A2/9lid
8fZAF3m3g0+U5/XqTtXv3Gbd356RHOKVXOvUJ/CpMDOuAiBa97rpdKbFG8LXjdHQJXMWjXGFjq82
WSLC4mkA0R4doO8WhQN/4CsNdnLrbx17gKPsW8Mp6GuNHcq9xjh7AcmhxgHNcbXP7iMfj/RAzDVE
uopqVjxr6kqpDXM3TIP6TeRFX3hfrvJxRxdgj9SWnCBqHJoq+/ZqPnWDrR9DdpoI+h/5uWqtxyB5
HwDCeLjoVP9S3RBlz5HHAyallmsmvuDehtjtXYPG4iGk/l7wqfineDFcnf3LOl+m3Hs9wEj4iWZT
f1d7fUxcmPTdmFBJ4+8fti4WVOUCyMCNzcrWmKrom4ncr3niqUPhqkLeu+3ggRlXxzK4JefBkG70
aeyQ8kA55DCgMURsBxr+Tse9YgywakEZW2uQfZZ8SiN0O/nuCHg9+5y3d97teQaWjnAw8WWPEWdd
+PbAjoMzBQy2XB6hLB3vWXQezp0A8Zf7ykECTLCD704n0OuD9wsD5AuZZHv8sLD2ogMfRd+EjvyU
b97ddSRCGfvTNYisJzDhXZep1H/rlHbwHpbtenCBQ5hinUjWVYrDQsREmfA6tm4V5s2wxsqKuu2K
dz5CAyirVTBwy84LoJ+yKO91PB1hHMU19um9yO4hnqx6TcPRoXiwzqp8e/Be0SfqX9E9vMgm0Lc4
c8Dko0vHCFs5i1GNe3iboIqtvnItBL3KSvGwA03CAh7RTEJbOeN8icSwSdvKJDk3Z95Djsi3Dowe
JOpLKyv09WC7zjhhx/3nVwRkLpggdflBWS8w68oQ3U6kvgN/YYMt1S3rXLyd5iQNCfap622Jewsi
qZXSVr8WbnLLNql6l0lpfNIzT/gA+McLk773xAwWyiJ6EIBgUT4+3tvqN/Lz4kuG/wh5AdJaRRzF
PbxhvcXWIPjoYEfh+7xSJ9ZyTreNOKfr5dDT9PELj30ZJxkswv+SBQwIx3Cl9s4yaaniO1jypdoo
cx6Rss1Jo4UYDAyxEXEosRQn61C8aPO4XYJTWhdRDgNZaw78IpysgYvjp8OoRgRwvaeIhkIxvl0F
UwL08RXq/vwL7AfRhuoyhgdfgae7Z/blGhbnC21/hVY9wkS4cMm9CFJc6JWkLIMBSwHyFc9qCk72
f+51mF91gz5X50WEND3maWEj4z+FM3WQDKVL9b5IVOEMSVS3gRnq2gCJxcUvuFvoo5TfOqPoPsKx
7sRibc73+CFcHkAsiRvNs4SMF+Uujd+/1Z3+SzL9RiA1OO9SUV7TlmV/18YiDnvBJB309ENLmFt9
iGA9ZswZoBdUjj/2VOJt9XQGntEiih2pVj/5MZSHhnmmn+6GL3R2FX9S+NiYgHc76dqXVvkg2WBc
riXKn07n421pEIXaDqWpsiRRypcRQfVWH3yviNgPOe6zkBUdst3j7JRTss+PyXBRtW0NFhyutw4/
Bt1c2bZcP+Nm7tzc1SerQ28Q2/iw+12fd7jOrUBIrbwGc84wZPONAmQgZ8k69DkCrGJGTFRFM1KV
Qbl3n+WWSg4D/oDnHJt+ehTl2m/peGAlC4aH69yD+uH5BM8GRf/Dj3/Ovc+3UzmiacNu0XryqFd9
Zxsa26ppAf0jYjBMATzU7keaC4RGf3cSXnLHOlwTslFnOMCtkaQOBe41gpXmL78ysB1F4GR8s74J
mxhQ1AEAbx+KxgBPNQ4yeSENjm4JlT8ob3XCx8L8CbxwbZMWaNj+GRkGuzxr7Fg5fb/vtDsVvUdf
V+xhy5SqiPpfU+E0CqFBK7PfIPhVx2Rg0t37HXkDv941HWmlSswx63RA89qCF6RHFXWCL1hFX5DK
/StqMFq0DMXNzO6nMHe5OEIo20VAReYA9yP/36R9OBEOC2xZYW5LrvbqfV/8hi8lyltmLENNFZlN
v1sGchrKHsr+KY/OOnnXP6uq/2sagEGuOjfSQPFLPAPiDCDwtNurmxo0+EyBR67wdACr4SLu0bTT
GaYYDwwjixGNLO3oohv286HMiq+3WJNwDBhlSoAedNGSuAQIFrGq34kvZq9xeUaCDu+6juQI+6oo
waLlI7Ct6+IyOUmqDJKZEnBMWGwu5tuUvqCn03CUfrCYBrBFbWWGgHciZJ/pnR9dTYakOAbl+HRL
R3kQgMX4Ksm7+mdw/ZgGDUVgJo/zZ8jRYQDHL+9QIhCF2+AKTA+Uznb6wX/YiRkc11fIfzjXdpJ7
PoaX2CFrZDyfFW81RifC7XydHHNSZ9ebYq5SyN+Fc6hXi9tLyoTZmFp2l/3zI+rB3r1a7shC601g
hfLPMPVvNWlSHTogYpoIlszG9jf7qb8bCEhWU4w9zD5PwXL3oPI3xa9yIVknykBzt6/2Qs7xbdb9
+Pb3TKebZtn4gpU7+Lv5jxLjiut+Qz3ZSIS5ZroEzhgcRdgKEhWUd3jo7ckUDalfvaZGIgJ50tVR
hMeoY8no/gZUKzg95Njhi9EH+KO/fSFOoCMcPmVjbmTGN+qxka8BdYOpYYdlk9fjNVGlSE5VHjRk
8D5WruEQ+tkyVpHB9m4i43IRbZNYFrgohqu6wWYQbvQAto+kAKSO1gZ0rOqEp+4NWqicCqFj+Wp2
6W7d6c4YMWpTUqH+RNLbpU5UdnpQlJk2vQzNowGqXmimtG3zIuxnL4W5SY1JzvYk4j1+SpU6GwJy
v68V49PGywXLc2lju6SqpEnj8iv/9Uu58VTqIO7cDhs4KM7a1rFKw405mqRYZCn4xcBR5gz6fLhb
sA6Wn/IVe7h8jJ9ieWJRd2Y4GS7Qc0++6cmsL3a7phhE3NTuHoRQBs2BYD9nB74lja71KeWLS5Lj
l0hHGbfFwJTVBRJh+4wCg6O5UhEnDV6IjpV3ggNG9z5zCmaHdqoryySZaZbjKLV5ZNH6Z+EPgBQm
Zuf06DZppr+QleXKO1COUv+LI/gqhy6LxlCR9tlTMrb13Pk7gp4+bJCesaMtG1bpfm9I26Mq5kEg
qMWry1a3p3G1qDhZ3z7YrX1HI5gZtXtEQMPvy8f1K/iRPQQAqtrGTRx3G5jviVNmAxN2y9rhTCo7
8QurUZsQzUkrq62OguOIwOExAvUKkx5O7R5+rbs5q88ohuyr3AYfJNdnEIlY6lrqOk1J+LD8z5Ts
vkQqfJtXfczSRwR+EVKJJs+qKi4HdLZN3Sxzt7zKJpSEswudqsHGHHgdTYubDof6mUFO5crHTn3O
AFBHQwmBmZ2j5NxaBOtFcPvounW70xPydGCTNyaTribANl0Zf/qnSGY2k78jOyIRsqkHQhpsbMzB
clNlG4P0XhReYnxFgxskRv4NA4osd0mHO+9M7CDA3kB1/ZQg+NGjpP9UbafaIfZWSxWOYt5Rd1KN
FBpu3wUMFKYbSKGQ2jFTAz+EQ+XJTdfPkVHXcJU/aeeGu82jh90BSzCo/d8pvA9+3Ppgd6o3FVrP
MGTBWu61L+ks0ZROHUvEd3uHsnGV6oCoOmAWNqtj3//xaGCD6ooEN+AQ2UaP+4N7dbKKiRL3bo7G
/4AH0+F3XwJnQ3NEjMRI3fG6d1Ur/dHB4hcINygNA7WDsad6BtYFCUIdoctvHJ1sY0kYAniv0hun
bSAkXpcbcyOmYgmOpJL3z7GSkWry19oFDLaPmPEdIeki4z5QCBNBHWWAsvs6gwZH6CJw0rO3r14d
n+/5Jbas0ZT8t03bP/Fvb14gcUajQJMBB8YM1+44heLx1JvmUJfDbCTPtx3pQZxQRKOMek/2wTbU
y5BvCfMqClSfGMysWwAKyJR66M4zywYHHZUtzba0PQU6fa0HeyzlIxy846ZsQUu2K6I6fdASar8e
lfg3BGwcMwULgFgLs0iKtXWb4lNo2Gb9EmDwZbHP9sWAHBDASApqHSxmEcuiiZBiq+XYe7Ky31mS
ZCWGLkJUhwZtKcWTqOG7CD9I3TYeXRvRFgvvhKLFKl0O+q7LxoqeHgxtpcdPEQIY/F+TkQuLA7Br
f5PBsEMsMy5I8W6iwSDRCiXny8ttNRrS6qE1U+geH2xGe4FYEmtTBU9EGgSrQwoYQNesy2UuIdSW
6Vxi63VNK1ABmgETtFA2AirOq+6Luo5xc8+T7Ahn9mYfCwYZFLwazrjlQQlTKtANpAdhSo4dcVzV
yqFl4g8G1dQNQbQdp0zhw7WSsxnH70W9Uh2mb/FJEzExEdQtHc4VCdTvV70iZN5M2HrX+QMF0OPq
3j4DWWkkUD2v+Q6BX/NFVZ9oxXns3a7KDfZUwgNtg0403xcq78aZdKui4pTf0tG5SGMFWp+nXwgA
XLakenU8aYzOxd4JMjgZb0VeNX0Nm9bFXy07fm/E4WEI39CPwifdUOm2gDPQIU+oSDDb9DkRpPNs
v+nX+tH9LvIDYozaO8dfd/HwAO4P0IeJEWTrvSZ3x9lfO/3if8szY2WRH7RjxmZDgAGHlsdVy+dO
fnsaE/qk8Jdb03iQeJm6Q8ukqYqjnBv8T07RDbgI2LOEek8IOEHaY/L/vRAAJM59P/ux4+Q2rCwx
bUQuKY3DdrL0eR+FOVh5Enh3o0VAZHVIXZjfS/50fldxajVE1dp3c87vyWHHFtPHvfvdz5tCbmyr
ZrVpebR+C1bUfzk79Rzypp6MhXpgHVh6UFDZgbVSDS68nAofLRfux+3NQCecBYBJu7TBnj5n+9JC
r6ANWVcyZ3mGTN20iG5lTUIwJf2cwc/cRueemSw2sa08VpPab8U4mpa55OyiqO76MzYaLv0eQSWp
pwLxL8KnxZIK6C1Vx5vEYv6Akif4s9gzQDezEbKmyfsvRJP7musw/k8QEeL4RxMqzsaHdbZbv+c/
zaTL7IG96P1wtXLm1V7Coj3gJd3u63GCvifk03xnmY/zngtifpOXfodGWAuqK5FGiOKGZF850V8O
/y7awSa0hJeFtzJCwUFdaZcgDidVbnsG77WOv/W3XAqhns7OhjUUdFwJ7Y/BEFFJbLYvC5ED+h1v
tx4cS+0y4ZP1Nl3FvQhaSZSEh2psYSngctLJV4Q70LFhoKNghCOQpQbjLSPg0uljNCUBzEmjOkE5
zeaOsDBgrQS4lDW2MqVE7kmyw/PNNGEBpqLI2CEAesTW+vmsV3J0dId4h1TpJTfUE1xuEntpytXK
9z/T1sE0ej/w/ZbXlGsdagrOOzQTprN1+DzNMQUHxbudyASMTjx9PBX+LVoBt/qx8Jj8H0NS7bus
HCu6wLla3AoIzwlahPtsO8tjgR8YcsORMaDbewbHRa8FqumyS8l4j7roXC/uF3cXSr/TKNZVtt8d
DZaAdccK94+G0N49TcrIgrdHvTjun9NepHK2WVqR6MeA7u8yDwvDXWziLcdIVkNTzrpoweFn07kJ
F2sKZkZ4I1cGgj3QYi1pYWbDvFW/JKDdi6cNN0GCd3gyMyVsRJV490h5m+mLxD7oz05LBmLtXLz8
/mApTv3FboQghSz7wWJDhCGVLwsysKerMgz/VC4ELbMG12cN8ZMm8ILZ8H3IBS1fzas9p90E7HW1
LZrYMPTDccdW9FzY9ExBtWZuAhMbzwSwIQqmjaSTFcr3ncV16o3wbVC/KPBSgDVI+RL+CUr7aOwK
znNF/zjN+M9m50aJW0LGvUb4wZcaJx0hi1uxqyTBo4xWUBh5oKSAHoqDTdG50UvGwYnBr3EWo/xn
uHC+172XQVn1djifwRoSnaOi185BpxMCgAj8WhMnXHYewg5arsmDMww+rtsvgfCUrc/BkGJ7mAMU
Y7F5kI/T1/RqJOT4IkgKSFVgYzvMIS3UQ+syxM67OcdnYD72Rccpl3A9f3kd/jGpZ91ZgW6reQWo
hPuXBm3pYU8ue6NqR7GuceCnYXHJv8u7Zk9arSZUzMApvX3AC9Ktp9uoWVsUP8c5LfwadsZJfNFE
HoAIfJTajyEAFxhPZ5cILo4Q596AQQx6EU8chUCG8PitSIALnwLSvJWPtoP9XqQL6ZmlHHAUVyYM
wDV28CjeYmrYTFXCNWmzTvbmrBnVQotslWTW/GIQexZnbvQ3D2iRHQufgFvRNktgBtdTIdAWG3ER
oqVzbedhL/2e/CuovzJNkHYsECieFtSwI/7QuYMTz4nFKE+S7gPG/UXJtT319Bi1u3Noip0CM854
PGJU0eegsu0000LQwYlU8qh/lAqHqAWyLH5E8lZUdOjyp5CA/XrJBt2TXgm7YISjelTNx+UAoApX
YIsNNpK/dm305XPGdACOa2ikmMX1VGEPkyG1AWvskb32zDIhyTVJjU9iN87DaJIyWrHVgHPgEtSc
nNor0zCdFrbrM+8ekRjmKK87iYz+P8afC2NicVwrZJBQstCdo0BstKAQ/2b/6RKTwWG0Li1qfbbM
68pTLyaFdsFCOV2T27T1yJFHGoZuufk4QmpmBjmuW1OolrEH/+HZIg/pvJ7RJ5u45/rSo6xh8rZr
JzT82i//wyqXpkbNGGfrUcR32N+YVSbzEx8Rp+P9VULngdMuD2cmmhqgrRtYhxvQb8lnE0Q/T0X+
BlUwfO71NSy1+NJXz9hY3LYtFpzG4QwiIlzQPGHMD5IAO9MDnxW2++7d6GRQuHIFVmFSwSnISMsI
V0yOZNahHMmydLuvR7kPLuEeuSPZK6bmA543YUnHqlzMyhfpmZerCoFw9fuH8KkaphjSVoaHEUlT
ZgAXgqNy5IPgpPakdg/pvlj1JlDMYY7hBVtFFj/rMwJ5DxZpQ1mf/6V2aYJkZ3+NQELygaBdMLn5
GjWuHoeD6l9vLV87meD9gMibELIX6uKk6y3QGmSFRhQeJfY6xwLUShidHZTrdhRK5GFg1lwqcTFe
Jec4yx+nLk5DfIibD4Gn4vH0auQ0d54cx51J6NeKcmdfMtHQ7Uf5HJB4Cqadm9SnkeCcgkKjHFqv
7f4AG/CuKbTrJO3C2eEq3+4blpXEFhJQMpSvM+5B+Xev29d6jCEdoER5MVmvX+DYQ2BJWpavm82Q
O77hCgc8bK5Pt7vv4ylc17A+KefOQTOYDy0UeshwgVpnld1GspxApc1TpOG+dQIGk8M/0a5nujWR
/IcbVHGaVT1E1h/hjwBy4k9VV3tvV/mDpL/pEwK9vTrVb179cSljxmLU0eMxbkYy5RddRILeaExa
Cerq+NRA3Vqa+Ttx76dXs0aewnsxHNVURsGmYlY1x75RYRQhiutwehXqhoE+QY2fOcjMFwqNR8Dy
Lmpk2IJ6XmPomckYa/2FM2zeWGRygFmId01mXfC3gtnJDGChDo9CXq3uspOnVb1kxPyl+ntzCwX8
ksJtT0rGUNXAVHiQLJCR4ek1LsL+qOGFRIbkzCVD0JhzCOYnqxlVe2UO1k8FCK68nWv5G98DuxU0
dYFCrlyHct/7DrurbuJKbxV3ECaG2eGkRaElJ5T7oPZjOHacZFiU7RLIvJZZ1X3iKIi+1cPh+k7o
WUHERVZ8JbYoNMFC2b5/kBW3HfwdelLxO2BTpQBEgmxP5RTb3yxIa9WndUjOc4eBoeKEm0D/p1fl
I+7YotWSovAi7iwGGiFvbXg+uncFgE2kErLTrnKT6Zp8yMp/KCeNVjVGA4MeO/cQg2SyZba8VUiw
/9MLyf/GX2YA+NG8kYqA9CBHEkvE7txGg5rskmFNls5GWilu4Ltttm6mFQfu2MDQ59RXyWKb/viO
9naT9wpBC0U3js4/ZWDy0cH+iG4Tvsg+2+piUo8sqfrQhychGSkSLrfz9WayHd06yuwo44IgeJld
cNWfbZE2KRx7mQZM/E20ECm6a1bJA72K2DxD0tCw3t64kptsrs74bGCRpcr9woYcn+yOl8y+jBr8
NVP/j8YHUMmOj6NK0NqCUzthDqBBZeNM7/gK5N7+9YNxJtVCTAnHnU3xeiqcWu2KetbzInxq1nfm
ygw8BqaM7qs11KQSk3EOUK6T2xHrjlSmTkVZxg6bFvN3L/oZGvtxZnyq6ofynqZxKmoW14ZaKXMJ
BLfoYW91XlnYmedUZdsaTlqBy8t+/vYRiDppdyDmAAPOSsodk7Y6nU9uuqzZlMSU8EMoIJst7zZd
CdhE0Hoi5Q/TI/59KtML15MLYl0eAroWaM3mBeGY7BumiO3rNZKLgVKbOsp83T42sMQOTwt7GpPD
gtDnCpAdrgrce1KWsIVCYhQ72FgNvM6vxBPqlh2MokplVKUG1i27fWP6yULBdSNNDyKB93CKE92P
ySt1u/fkpYQPjTSbLMwLz2VocVHebGLRBbarxt+9S729D5eB62FKwQDyal+iXszzcIEhfTZBWad1
h71kWy4HBWS4ZbrHL+CiqknCZrOFG39iA/mfijzSzUSpzcvzEjeO/O7KsDp7VlO/NiV0AKka0bq9
s7hDjCqXMjhgOnntERuPQ9wH+2CFAa4XMQgpthg5El2K/hsxoCEaJgwY8DuCSnyENQsa8pAhoHFv
qebVHDCewfljEop9WjTaDehqz+9zDxTNha3Qt//OYXbFUVY6ZjMdE6WyNMBBMFabm33wajgedsd2
vZjefhKPXaOUvfALUBQHd+S/ECjTFzI4kdC0hEfOsaKbcjZd08OcZvNLXq3uAWMt+bqZCWzNwYrK
npjeiieCe++G4V7oP2XkouXDjXNDzqfPcTgrZhd7uKKNtC0FWd7Wq85t/kTuCqLWstaWPqgO95hb
jdK6FScN1tVAqetTov7SV4qpGK6s1+iYeJ6aRfrGp9JvJsRGaPRzW/BGCVmWJi2gvXp/vEpQ+Kcr
6pVS0ot3QT9Vq2zUKlObyjynDCP6QxJ0R8JJQAIVD0siXZQosRLcMb6mM8WvYc4lgN5b7Ym5JTSc
khekrMEhEl2eNhNtuXuFxL10dWdkEGVSzScdHPFHfgs442SqJ3SLxW3Suu6irx/YwVs7GRFOTr+t
mze29YSH4G2p86mNpgbR/4Elu2Bh7jsgTensltUwkIDqI/zd4vvl6XlcykJHjfS31SodxODBP9fs
BQ8nv9rrNaeecIE6cCtnv8HTW76J7C8+LxxC1UKUh3aTO/8id9be7/D5AOPHsNZgvTOynVExzVlb
0/IZNkyBLtW2ezi1PxpAc7gfQte1vsedODsoypZwhUBcMqtG6Un3zdAgIL5xG0j+/RvCYydLO/Fr
7c4H/7kI2YwLW4gauWnuMNjALFEiIWIQn3t3mPvPtLLTLvrTcDtKTZZuHzfoPtE8gUgq53uvByJ+
UzUbHZ/iRpjGmdlabU+AIECBo98jBSN/tq1MVU524WnG2J0QrYbjSCRFNRL/egegYp7UwyvgXAzs
qAZ7U7itZxHY0H1RejMdM7u+O01UjAMWzznQ1iDF9fJn9/c0Lrf/LhYTZmD0DwLr3SkMeNCc/6an
rq0N/pIk2vDOUMJEp7r83mME0+V1h2tgQVAlkzqmtxZjqWT/oPj2f/RlD4QyncQBNofxAIGZvuRr
7oepzdAu9NQycC3nFMkSouBl9Sog3ADXEaNsLxTL9LdilkQumOtjKnSQ2LQKdmj8BMEgIj4HVLFp
WRbrejFng0Y6X+s5NOnuqtjGzlWGR0/G7cAeZ4FvzZMmqgp+xEXGiT35G95PC06VQzCpTXpuDpIo
WS4KQbMxpQw2tWCAbAMBi0mwkri2KQf+l2PfV/217H977eg1f5iWUCn+l4Ns5tL+B/5dtlkF0N6m
f8IEPpu+vwLZsNfHF/H9rcwtktGN0zrSRxfIPssAqcDzc7Tbp0SGqGuGlts2kKkdw7UdYX+hlcA+
bda8yOqOkDY+t2zLrzYBCOT0bNxBR22/t7JIwz+wLH+xXpHCgy/kZTAOtwGuCLb8cHnGRAemu9Qa
y3UAUiSssuzA2FwxA8bxUm6hhGOB+WgV1qrdeQlHjK/6FN1hJgBga19f4wfNeoF1OrXWl9WeZQza
Y2b6qMxmSsIE/oCSrxrPUiZBaO5PuXsXRGYT0w5bttqL5O5hhFOBce+bq+46dSJTfEOJU6za05ot
NHZK/N+W9Hv5xEOIvSAeE80nS9gbHB/5afO8dlyEkNy5R4yQmcq9KjqZTY35pO0dhzDoRFF1pCrJ
rInDSAD2mhAILzAw41S0+nVT3VuFnapZ/24KAUOgIP7131uh7ZXWCRPsDfre2SLIyJpVTr2jhcDe
ZPnCL+PLBqMgziGDnVEktQj+PRxgFEVFHoizXSk3Xsmf0d7eixwPrasmhbeoVQ/JcekmrHo6F0f2
uZfvI5FMRaux+7269VEzjvG7EVA2dNC3Oo7NxrUYcW4IrKA5G4lLdLSpzpT11tRmEo8F9eNID2m3
WiqJ7lj11aVdWmsLFZmcyYs0mnuU1i1VVK2OXxCdAlIg3tJK/E0LYoH7lj6XcIeaKvyovFbiKNf4
psnKWMbDLIlhjZBATH6rtlTtzQhWVAMTN25bo79eQzdIg901Gm5taFjDRsFzkVLZnLG7U4mSSced
PA1slQnDKoyGVdMt71pRKPFV160jioJXlvRzgvPkcWJ4ERBbTqFtJeyEFcR3CgKoMOKhKy9TBWMo
9XGiRbz26ibahd7ASatFNwKwYNPTUWFAYPYRE2ameuQWjjS/f/PLAPkYsLvg5PPh4PgLk12WPnXr
OHL0reMAvaaIU06McjYOSxpmEh3gjYz98cathe12vkV1tpxJqgc5sm2p9C3AF//jtRxNhkcSeUV7
yrLcdNl79R13AYwTL2b6VwNbhwCZGpMWoiALA3c6+hUf8oR5wtGPTkZTRsjzkefHyqXT0x8Jk1mA
HV6nvZTVzRp+FXTKjwiLEzYwwoqm6a/jeiV7bZQC5mdZSHyxjXLTKWFJbGFXpUC9d2iAALVW2xX7
wg4q6forEBGPJdtYsgiHUY0VKIBX/SVnGT4kpI9fAlKaw+sswZSh9DIKBlVWJjRZ4z5K4+e9Uito
TY4nCZXqsxajmL31FqqSV0WyUsEh3pWG047puMdeIgEY6ouYNDg1cNwrtGAxx8OOSIz5qmXXiNXk
guNl8dwUfH3Awg8PCiYqnu/+WaOmzXC45FLh+b1PfLXPDX0lqyjEwI6NaJIpVjojWWkFzTc5Bva6
ByyX7/ybHmH0G7CBtcnpJ9DKtmZZjfTJVNuovJl8t7waUFrlPHipUEuYR4qhrHgrDLDCjwvKaKoV
sst37L/l+BpmzaZ+W1FDnl47z91WGTXFal+3xIJ0KNqqeKun2+mhn77YR4/GkQ2HJpXLaHpu0ZLU
DSMhJ3HMyo4/WhrddF1/TVhz4v1LG292c6aeWlW1W29wzs44Q66Q2M3TX+EGACoydjNZ2Ei1YhbB
uKcFikPqSEz+CrZvVr+lqWl5WG4QYW8w07VOYee36A/70qlM6hCBla3+7vYT9g2pQF6PfTmCrXmn
/KICLZhs2um6jfrXyRYCW2zFpBs9/Qt2GIaZagFa4wl+mWunyvdnW5qRqQ3lhBjh3uUhLCIDyLQv
QE3V9Jes3Rz5mPBJBv2UJk2IzPgfkUvgLMQLYpalePGmBpuFSY4ku+HglNignv5vi2H/tzBFlovl
ZOL7ULI+OFloWmTYaVi4AAZ6tokdjdcegwcijnwE5eY/Kf0qYqNpcUhQiHj7TwUO6WGnjAySKSm+
dM8zHEeCerS6uRbCXTJ2OlH7AzPLXVT1lpSEiY8rdsJJ5V4VRrxYTSKj3K23Ba3tjjbePhJ/jfmZ
ZEdW07JjyrpcJYvimbLowzV64C4xm8Ri3mQuqcUDGp1/5u8zxRotd2DYrjVVQBQo0rJU0KLv8IXx
qYRCq8pPpKhYpAHF6ydvFteTwCPbgce/yrkL8pKQM+jIhmzDHslcze17oKbHmc+a5l+mYMlhWGmK
phiU9yxLMymE0wS9GkL9iL+SJZtFAKdLT7nVavtin9zdKVolPjstIkl8i7zPmHZIlNyV9sS/S5Q0
5b/KpnYQG8osYx/4+9mjdhLipufxka6R9Oh2LvdG4fpeGo1FMKIhqMhGKC/u8/oRbMXlxrHXtBtK
vhT1ZY7MjfGrsSZ46Kiku2T3XAn3QGWjzyEjT8XvmcoUHSx13o0qMey+yxNuEFsDT3pujf0mq0Vg
8uyfPggXyd6jNMvJ9AQd4TQeW29F+mlhHfDn1bGtzFKq8s5zNE9XiT9qycQi829Az0TDb1MbRIqR
UCeZT3vC+mse8orXeSf4/aM9shl/e9NrPlSIOhxbLwHTQGtAkL1nJM8PDSD7pyck45ht03okbsv7
apDplZDAuunu8Nu3IPiCzmazL5c7aZ7l6aE2eMzJ5ygSB3U6tgyQYiSOgClsJdaLPe7CMgtnUg8z
TkiVrZiwG0urFjekR5pmBQtAjbYTHOuQBXJeBA2oRuComYmIKxgcVTc4IwvGMl0Oa/gAgcGvAg0Q
l5Du9AGG6G6jqN4BrCA40ZamYpWgDoqAwlaSBoNfqjUAFz/1KA2ug3Ykh/Mf7ThPXdxV051hnq2a
NoTbx3BVnSrB7MKkffqwagugl/50f3rzqeX4mInEIHGcYoPr2ScL9RolelHfkcLmyfz6IPqRPZf2
EC7d5jGD1SwrsjaNTHvnI0qM9zSqp56/ReEmbyHeySM078ZjwT3tiIJOMVtzwGII5SAltISZbV/f
7m6LEZqGIWzyw6PseZisKiMjmwbPaQfbJ24oBQUEBR9kxxqEebQVOUOtRRYezBcThmpvSxj7EZMu
HCwsz8powRvnwSxqXJsjV06+cwRp4uIHaSW/wmiSVmvkRfxx/+je0ka2ydpu+/PF2KMT/6OTRp74
aO4q5YLpYsFBKrPIiO9w5T7eBRJuW7EC+o3hmbcmCp8BRKjMc5gDgJVSy/HwQBzQXAk0S0JNmdb2
AYA/vsMFZqvkTDujGgvRtZnRyPaNaE1WB8MzogA1jnzmJ5H6fe1Fu0ofEXOFPrMz5ws1P5q454/S
4U6MywLoyWHoTIyoZKRWQGMJqKRTzlUB4dXdJGt9FFa3EuNhBNghaxXlQw/IIyYzY1vOOgZ4xi7u
TfnHQaQQpcoCv+AtkrvDE30jzUBAx8SsWIvWaeEkk79gO/Zu7+fw5lKx6RU8Rb9IXI6XdxHw6QYd
gOXcdXXVWBekE4zcrbWHPlYSW0eAiCsbcIPSZOFtQZK0K433Avnf0MruqICD5ztI+J8W8qpGxzdV
GSz3NlHHYYoL2TJfBfK0j3aqwgSGbqFsa107FDWXl8VlfNh/IDgEx0tIdC5p/6Lc8lHP5orFNMEc
xivVhFySZwRkfm6TK2WM5PA9u7TPh5QwLgCdxW4HOY0jmbTpBQ7agWbq0A7VY8Pbgiw1xB/JScsm
E7UPQlUxkx7djsNm/WfT1E5ubMB2CDbQYRNs6rpNF9Y11OoTgoNTolX/VCzQ+JuVUoQpGZDVR5fg
mDECbZQDqJp9NmoIwc9rmlaxng89Q/MIoS20e3iXx0hIzg8Y5NcOcazn3Tc+cuVHSG752LSmGwa6
qdREHm8uMwpEcXh1dt7EI7AX5oHWQp/uco85dQJ+bmmalQ6UTPD8vj1TRW/RTPLAmDWPtbgvqa66
wmskVn3m4WIRPznYsRQqOfh0h2iqL4MWStdGIDZspBJFEZXMcUvpG47qZ44X+Kd2mqkr7zMPvaEj
Z/gVT9rkLAnxpMN+Xry9waG/TZfOIUDu6qNVqvGaXSgVgqbMAT/zwroBJ/UTz14gBJym53uQaX+m
8fJPlOiNdKSpLLE05EDOxIAJ8ssLLt7qsfCZVeAH3QFo/vmNUohXXo9BkDqU3xWjJxlfhkm/HD3U
0wyuKFxUZzy4eXNKFI1n+887w+awy39Wg/HLf6VsNWErGE0rc93FMf25htOhnv+bfMqpbPI1AAkl
oiVMPPTYBoPPE6dQq/fMnAcb3XDZa+ydrZ006JG6QW4nTeYarbdTL/lY447FIqM0Twhq2xcKJZ5b
scd3fKDiyl8MfKonzhuS0nzIyRM3EPsbcYqcDAfUmER0EP549gbSurNmPV0WcB+QooO8xv74iVlB
R/7xKwD0IEAhCqVG397XuGvIkgJ8ghlZYJPl5PHIAtMjjvdtiJY8Ynm1iNJa67VzJW8qRDRxquJc
hoTMLQFUlamAwLa9Ymn24aoK0ktsUbFJB4D7yLE9NLa9+58zsBYk2ZrlHHbHKwm/5o2/d1Fa1VQZ
j+otYgtfcnC4ynIl5OABpFWFPc9iWMbJEWof9bvBgNoywYlg/MMNIGJU3Q1F9dRrxLVsCLwrBPVK
s5pmoWjNKgJDjhf3WfmUj937u/gquf8VkPbxjdBfWWiB1L02vyIpVKS7w1Ze/GALPrFpguKIBNn1
nYLufj2OyqIPoMjl/OKWTG35d/GAp1iQjLaiAp0oRsN9aBtQGfyMm5fxupLkyM2b9+6eATFM9sFJ
JNhh5RkQVOmame5fxtPc783IGZmHwlzxFWAvj7snQCQVmAj1jsbytCMA7xKn2a0HQABqcu7i3qWz
5OcDe4dJ9aC3oQGp7zqJ4t7o4+WivMeUpg3NpadKPm6Wooe1oYra8N75c+oBFP0lrpzjMR38icJ/
ySKV/rd/fOVPkE5SFkOrKLnu9Q/9dnY+P6VfnneXf+ZAaxE+4qVG3mDEXzTnvwZdYFcerfrFzIbA
CfKq/eqm64BojbahvVFffeJ4FjXik1BONwWuDhUZWy2v1NgdBXvCJ292xrHuq6fNKCryQmqBqQR1
8jj2eboFNIFHJmCQcmTcxYC2R41mG7QCqcO5wghKPw/9//z3g6pqkms9gHmZ/ZkNTJzT1baRfPUI
r9g0ExYCpopc+0O1EiRAnHb6v7PwQQXUH90HqmldK0l0LsdrXUTS/2jQcBfUXtawoXJUv/TE58bY
kk+r83csj9NyT3I39xynjMv7Yz+2HwnKnfQHzTBKTGH+4g4d7wHBtZc4pxgEKbE6htesMklf4feH
UoObFKW7AEcHgbqsYiJQZ0i/302tK77jB4nfnV9B2h4EhndnqcespafrM2tGOcdEINq4IMOEvcpM
vTv8SS+jULNr81Elt53mEw++AFbT35uN9cU185bbLEiJH+B+W2s1n4QEbdKC2JjDfO1ApjR2Oop+
M/kxpdk8PxaVJyYID76X2EJj/S9jc1kESmnoM9NzRYd2JocDnqVkQsqHWaOkRyx4fSqSrhAbivck
eBvqc5NNRZr2+hC1mu2dPOUhJb9m+c4jyRUy6NyANP7c9i+6NzO4W9YYsb94QFigr8xo/ziPwASt
41vOsQylycLVZGdurmd4N1DXHN2qWBb/Mt+kFi/Yl0Bsp96e2G1jXU7bZNK8zZZWiaMRVYa+EC8g
13agpfN3BYwIQIdx21Z3lx17RrGTGM98+erL9aXaSlMHzsr1StqjFzBArynXsXgOh3Zp5Jh7Pb1T
plnu3P//J5qto18H4cfe4T1J7tUAIiPxtCelWSttKBSqwPOFj2y0W6dRx07iXB/vDr7yi7GEpW22
o7SngpQQ4SlT8sMSCfbLiE1+Pc8upgrrLHOHQSRtkHSYbFXyJXjiqE6N4Cuyokdg40S26ej+aOxi
C/ZysG2S0ZKlTWZ7jKM+ce3TngIwa5RFlgrJfaZP+Hz5lV1JWnbJxejpaYHlLY3dU+xi5kGLcOVx
KKo/jWpz+QaH+siwmr8LNac0G12N71zMJN8TLtQUNblLtXHMi3ZiV7shJIy5AApI6Sg6hyXxnima
ASPE31IKpjjgTC9oxA95nA9NX2Q5MPPlpaJ5+b42gywQMBzhIGqxmVlSyypKyfFajQjNiJLaLZyB
iiBTMg66kP+eTKaxCBTn0RbbX1RnEsoXJMbLpH7j9M9/aC7COc1FuHRuIq75f9D8MSDZCtHkDx5a
BBvKhDhunYPrSemLiBQjE4bx1KM8JVkIQ00yI0Wuqb1Q+G4S6cR2ZiCyuVa5m3Ld+ZPn7ldTJ9qU
2CmQcT9iiFBrp/Uh6vvukGmZqWOXvxkW/nAODicZWWlRvzNjxhpW4Y05AROKF8HQSI0g0NAuxfrD
EJs9enlUZgWnZhYpep65DrMSJYR2GD0cmhkH+yK8HZc3EkhUdu2LTki/rNNqBt5xfkVS0uhOjSYD
adHM6GZBzLKMMTSxkp4a5kuD+3hGoM05tInXVldI2Xkyl9oa7/Mfd/s5AiaCuu1N7/AJkdZI62UZ
L2a4Gzyefakq104s4MEujksk6xlL04R0G9z94QtXpUN+Bm1r0ykLYsdqt1E/N0fyrUzj9jwzkiEK
kLWncJ9rf03UsAjehG5/l3+FeyORvKSFukQIsssQWWv9VmFRDqOGD3p6c0QMooKM7oySRGXXtVZV
eHvqXoDCAyrpDnK8I/+WJj/Tn/Lgl4Ua/JjTgedLlXaK5z7JgegJBQGRVQX+kg20YxDiMGfhxWob
a/FcPIMgh0tosH6E6y2VmmkL/UdNDZaCmfp+fYlZq3JicVWHRIS2IBYpgdaBkgnARoF2KoudTXVE
XJZBrx9Er53PIP1cLNDxqipJcixOLbZPr0Wa+HN0fU++C1ng+6AQgNUM5dNcKB/vVCE7V1ZwBvB3
eyHrd4sbIK9cOIGp5yxlc3BWs/8nuH6/do/hsIimS5xivFHMbheCTYkrqjhzOMEu4Wwm6jk+X8vt
+sOgNrtvLIsewSs89mEWtvpZbpQkCzjQyCEK6vyJavcjXuqC0/FsVQ+Qnz3ngkhaqic3m+GonT/P
L0kb32Ohh7EpGjXWrEZ5ZWfJx4K9cMFOK7ilqNsTcnecY6NBFTRZL2MDWUxHFX8+J2xTNwWbNEew
FY1zKP8evJl5Tu8S058vY41Z+JA8WCbDVpslg2te1RXNhMj3FdaBZgbRk06lF+Iizwx0vkS0qHjk
OwZalUKLB4oiSd9SsG9hPgzP5aaZL8fJ86fAxsLhPtW7P23hZTyz8uH06nxhJWiqpFYRJi0s/j3X
cMi6QxBLM8hn6QnA+AWm1hjBGS21fUZ9Drmv5HoLI2tdBFtYfWHMezFozMcTYYBjrsf2N6MVQI+r
8Ne30KzNo80BQ6xNH1X27exL5Oy76FAe9SOZvJrMzlOum0SUNSbr6TlV2Qm0QnfUamLUcDopndwv
yK1owBu5RdHQc3VhhHxup5cLKYV/3xvFovOaM0huvs96c0AscVtQQtHXFaH+JBh4wRHGrf4PJntk
cMa1b4tpjxjPW6/AQhYMccXLYIWaN6yvjS/bC0yCF0sip/+5vHwV+rtMPLQ09IzRkXvq6I0uvkty
5uZ/JmAOX//t61dqq67hqb1jyIbwE5KXOHVo1kC4zzYZ9MqBK8AqDJDQGI4sWRE6oDuZSq7tXBBW
r8F1QXl8dIazDQacE968D6VgtMJ8d+Xn1KjO16XQVfmKIVt1Qx1bFhPVwZFZmzC1LXVhKdpDLPYr
2gKqIiPvx2lbtyPaG2tWdcuHoJkfOJqHD1de/JeehWPBOBp9IHZ1NfIL57ATxyVnfCljZFyyqde/
iIbN/oYyn/Ck/Wpnrht17IwhUl1Fi/FPi8qj09K1my9np7SaaoZ3+LavOncZr/7R3iI4d6p2Z6GB
u+TId34Fu1X+S7Ps4YwFQlktcj/GawmVEpXXQoI9GzYVgR29ceuPRq0SFH2VjlmpkN2wopoiaOAb
udvoewZyr0k4ovtRGTnZCt8kOyAotma853LDhWVy/uVBNM/NSS7ADPGdSZ2h6PVzOntZbj/3iO/E
Mzt/Ix5aCxziCnNVHx9OaIK6MS3YNjDUUwcF+gCjFvuj+rl9MN5T9tAfc9B4AiSXqVdtre7OMzjw
GJ2E3+Pxj90FahQU89MA2U7/k9xYgmEO/TWN+hkVR7VQ5aXGsV+9z5fhk5+tt0uT6Wiw+SAAJ4Hs
WFAvAdZVSDq6KS6BmyIpBL6JhxBmjlycjEkD0r09j4NSXXltS20wTmOFZ9Z72ykz0EM54o00cQw2
/aqUl7pdbzWT5FkWY6bpn37QOMgcXJJa0jQ/uvEVZU1CtYavMgaN1K5pDzucn683ZiXRUozFfhhB
T9XxoXoihMoDhdt8196M8C+G+Z3t0EIvs/bo/2LInPeUXJy5JqXyyWiLW2XjUBobnIVMP3/J/Y2n
rsGa9ClDX3JNEiBdOM3phtyijSkgs+w5EkbcPX89vRYUI6aQfL6+Hrb+qjmwo6nohhC1QcQqBHAs
wYTNPuJGkigj5ODh4HpH3OtqL29LMDtfoUDNmMhJ7RfYebFDVio2u92LkVoQx54x2gjtUlBVaQ62
pNgT9BAAX9fwTJ0SAk/+zyiqiJz4BLjQZ/sepUPUcRVJHE7iSg4l7quqmhWOrrsEJRQTVdTwuMbG
eCdlkYoZIz/7AiqZ1+zwCbfFJ0wKaSJ/Q0g0ahDYRee6a2pJgS0A+jJGqw0gREt4CLuxJCZtzX2s
hoifoTln9mw7t/PqA2mvvjWdBkVYLn9jBDWJOick1sH2MMrHCZdCqSO62nu76TUrjNymMkcg3k7g
Y9RMpbD7ca3jxw8ghG1em+LoUjWuO12teZxLGOFz6ZQYkFu/S8gLP7lhmH+EFuCKEhA54IAI6eQh
2f4/1UTGPHJBDUUMl+BbQEjEZGtI8SMjrlLM8Cxk42/31Aw6+NB5oXoibwjNIodF0WW7mUZp51Xe
lBQ3wWnVmfCBvrwNUr6cppwmCxq1IrLXJWnzzIFogVCtFGBQXw+Yo5Slo1vXPLNn2F2AD7JuesBE
Hz3GPT9W8VPXB41s4BAajdYYeCwm24Z2MVy1nK1VIWKz4V4Bze93wfdNiKSF4EuYEKAIS7rk+bsK
EqYqPkMe/XCC+xDbeyv5BoGnC8QBHB841mgMJAx2tjLLZUO3UCmhB+FxpMTZ+DduQAm3FoX6u/o0
oFkuBBHzNhdvgtYATCl+iq5EMcmXxsy8gCc9XbpUEnVdfk9xmeEXMTLaxaZ9sbU2+BJ6TSAJ6Z2z
WG+sGWEpoow8s8d/riWlgrKgtTUyDKzmu1Yn8HMuzxauLsuB0NrMEOEDbDnkQFbxwNLzz4svgTXE
hR4zwhn7+AWmm4b7+R/X6PJltrQq4WfNRDPQplwX23fg8sVObpBWimL0Vej2IK/sBkySSyBlqCuc
NovLUH8DrtBr5XJKsTWRTZTVnWE10cvoFjA4Z3WtH4xARJeGt0xdwSJqMy0W80KkXOF9bubyHqeW
yVBqx9TTLNdWFQzIBYK+skd9sWdfNQtDFynkjsGgO+mH/l2P2Wv4lcubnedO2VP/Byj5e0M86LdO
CTuvOtvbXZjVkL/AIWY4aqNfFn0rHxh2n/9iRI9fZPWfYwJxv6MGj3N3V+v+LgY1A5t7K16+FcmZ
akTGEL/lCXZJmPOVs3o/p5DeC3CUzn1/x4UEmatjXCXXU5r9Ku+fh8pRKWV+26+d90hIeZRA8VJ1
bMTWAs/ah+PLIe0kcg5axe/MEC2ulbUiHbf931LcgC7b/nF1UqIfMNEFXvX5gs4+QTgBehKES/hS
OxML7pRZOQchIkasTaQvDsdCnx+cfChIrDsnyUhSDzGXY37yAcNQeVRtnux/9eYLpumpGvOcSBWm
MzXIn3rqZ44lK87GKyVZYan5hYvW4L4khNPKwwiAwtKbXYgsYOldA99RojjZi0eVrJQ2YBzUSbML
iskAqKS4Vab561IaApjlcwIcrgzc3IIXB7CIplBUFU7xIkMaeoSYx5ekGpXJ7DE5Jtw3PqHDXLVv
UZtr/wziDRC1ZdB18mYn6YJhy7Pm6NtjdxIF+eU8TSF0Rw7es7xTunCVa9vC/UqSwF+CKzQYPgMM
IWvidP6iqeRGAFWjFn0gQqW087l2EMDninS0PmaWlcChscYrxOkoROhKyC6WhLWgLYM0uJIzhgam
XiYdkHI0DBngKdg294k9c4j+6ewFznvwxnB7mpEJR87+Ht62E16KiVZclyz+EFuXq0eGaHIit7yR
VW0jCgKQy8s1VHQ2K94okwH7xIZSb6gnElCr9Dj6EHfpg7BUT9WtYRpkkVTFdibagzmrLSKaM94E
uAyLr0YwYkmsfUFzrn2kFsUppsln2jd8ezRZhv5T6ExQcQ+7FOfs2ENCfkWi1sVs4E4uWFQdJx1B
jtGxMTBd8DNCtMUPxhTj50S6qq4UuGoiH8AHosDBQkcwHNnoH4uyBEwbMaeiv9X7bHLoUAMUtcOm
jONJsKHuUl4pzJbXLRwb/8Z1rZfwMN+M2JkQDpqcLi1RYxVoWNbBhz9jDx0HPqs7DfYSpD6PxHXy
2UsFKARHKpXIVu2vEnpgqetWh1TkA6V6ZDENuk1Nq1m0M1drTIPmuh32KDFB2y11OxA0oYUF458A
0Ng1ck8fXo1Wm+TEqBQjSUGrAZ/BVLtRJvFwsUIh0wHK6975GhRW/huyA6m2b7RBglTt0noHIeM/
otVXN5YzE0OEHSnm/d5Tqq8PhJ+a9KEZ1yfg8A3O34b0n27sKBAT7BvumSiRTr45jjcESFBOzFjP
NMmwMjFcUSAVMfl8in8uMlPKaj1EDh+AZuqnEqsi12Yh6W8YMlwlOG91muO2tZ9vEYP35jlyEthd
J4lmyBLIq01o1dvU7iQi/BDrcjuCaR28WLnChhJeuwU1Y0XftZcGz+gx3sc6H46WX0E3PzSJmfxZ
mfkSOG1VUrvOaniel3iQbW26oAAWG5xJpLTaXhAd56eTWe8s/JN4Zk8PJVvXdo7Om5dphbk9+GIi
pGqkabzBKSIFxTMywRKiiXtmk7+2M60cKI6WXWfiqAWMUf4AC97seKXyOaddA4qX2IYwyffc0H7t
BjXoFdxxv4YJU57JORviY5+Ba8SiDdGKUuJ2Ie7MOEnI56rRv1gCMvC/Ch/dydkg5+H8KQQSxlR6
DTAERc9RHm3IccX4EsQ71+kMesyXfHvQG2PxTv27MOk4KW2GxTbaePQ3vTqolS5/WLN2ZvtvcrTO
sqBXa56BrsIfjv8shfPUNMuwPqBR7O9/SN78+SDiIWAy2MmbEzuX/GtD+hr6tRLitCBX+gXW/E2o
M1gXVmfNdYuBNgLl4jgZXZ7qoxq4NcenmQ37U6GKlgriohf1cQAdsef4tlQuN1B01FTo/LoKJYXX
tgdvX1R7nVhc6vMCU9IcIb4k1DbF5a7yM9HGmQwk6hgMJDB6edIBb3YbAvHz5omjgAxFEsf8Mujk
9IJq8IY90H+xKzc0nkiddRu4JZdbA7SBCwbLrM5q7wV5+hTd0Uy9TEUwM78EVwoa5eBsC7b3Z2t6
9DEiyxqdijKBDafoIgkfC9O0xJL3sTzdmSUe/sB551EdFJOcd83ex5PkHysZOaLsMTt4TH4AZxZJ
bGHP8sWW213U1vyJgbW8pxTB249P1/qJGDtDnEu7oOqiSipCb/63o6+NYgMD/QmsjmiSw85EyrSH
hpcvOe3z36IXpCUcSIDm5YbRZMlP6hlaoRKqbOXw1pkZJOHPEsQvxaDANE338NiuIFCoBqO609ie
ferRabF2CFj7m9TM9yDdMImWA0Dd7IZvCIjq/sD5INMm1W8X/Sl/EHeRpFn/c/ZuCHYdUDc8e5eQ
zQX9shalpc04F9PbDNCAbYsi4oEWp9cXWdzs1QS1MpR9u0H2KmtLpoaUDxAULIHV5N+EW+H2XVj3
itzBzrnPFc9Mcupw5gyZ4odZG+lYUNrd8otDcpwq9ILQ9ZSulPKVXrymOOaDBwEkaB2XaKzkWEa8
2iEvBEri6aNI4uLGl4sXqUoBB6dw5tqJue31apZFrkNOtEVRWFtN9cOl8mq6/oIvzJBzXGeEgh3a
tm6Wzlb4iNLSp2zLUaP53AWHQDXhg5vCb6KtAyGSMZx5rsTFbuFD+60i76XRkgcml/MFgK6MDSR5
yUZj8s4FVhgH7j0F86YZ6H7swURe98eEfTjCSl8NuBnpKHnaBRaLL3E5fc61w1bCO5pI4TbaNLe/
g8QiaDcfpnk2hizikbHE4QbllH178qCj9Ow0NuMReG/5QoVYPJcJ7wyE456sP8V+rVspG8YwTw20
hkmofPvZZsKowlbn/dMNfT8HFXi4x0waBQ3S6h4aFFO6VEE/Zc6x3fiDjLkPP42mFqEqFv5lQyas
qQrqKmnW+nuGE3dp4XhsaOs0LJdfwDpfkZDsGdK+EI3dA2zaK1pTdVHhFFBoBOvkJdjb/4iwGhBE
t/X+WlttTMnvXbmizoYt5swATCfuF5AyeDzD8g5IvEO4GdrwSsZxOPyzC9ZMLEZkdiWSQS5kE8fr
f3YFFpwY4mb4dYPGL6P/KGW4QGz+OzSU1KO0UVVVMknAEblzsrslvpIQXA9l5z8B28CpBB7+chSQ
aXlcTdO8DUD+is5k8L5Ew9uDUmZX5pNHTyhUKUy3BT/wes/aY8X3uuQG2F5JqsaoqG6x1zgpxhqT
xiZEwii6T9utleDEa+8l1TelG3+ImF8Tj4gkNFFgyY/LF+XcoqmTLH/ywabQhDr9L9ABSP937YA7
AZHluo5kZ3UOT22o95m8dUoPFC9yRDhmLpvdTqp9aesRvHxLUwZXlp5m+w+74/0e6Q2fDG48wp+D
h2D3EqZAo6pU0T1NJynjFri9RSCHjWNKl4FRKCGiBunryRXd3F3UISGXRfpoLGuKh4vs+Q0R/XnX
8HVXzvLKh2RJ/KJEt/1zUDhfYBMDUY74Lyrzpaw7Dyqs7ddkY0HjHHwm35dyUO/GvDfBF6Y3x12y
bWDl8m+eCDCMRQgPzaT3ELd4sIP4EojIFln0AMxWYdlHMfcgl68TzwgKq3xmaVbQZa+KnS9CHY0C
01RG1vw0ibHpKz4krDI5xLPZjQSWVpN/6oVkvL9uKwMfgPVUuBPQwSNlTKITpGSqQbEZT4ZwaSyV
l0Og2QgDyuzNCzGskk50dowLV7WTriCBGbavcL29MIRWvutJCu2Q3LL4742+y7md4sdlG6j8w46S
Y2nX30SncU29yyaTXcaChH82sLxCzRxy/1QmJJHpg3YPR0Qdjzk/D5bVtqfEIPceR6lkuZGG5UGR
mvCXDHjd1nSUYtnD+RZ2t0X/c1CcMeA1+ZXC6xlROc36s0R53bPivp3vE5inGQ2Mf/T9EuO71Xsq
X7JlUHf6UOfhoI9ZnebHahOJUdN4NjfSHmr30WIX1FKYU4x5i706qMeA9Dx3BBwqv1rnB70oxJnZ
3qZChr8g+bsiUu28xYtO+2IGxUOm0jJcj29tHZy9UlAARcAg612HuKDms0Jd1blTza2EitaLkx5O
pfYp/JdVdSAoAJNMrbYW8InVK9p8s3H8ooOI+yU+h7FJ23id4Pe+mE4sYcBslptmxkvjJqyS3iaJ
nmh+wvcddOjWgHuWzevUJGie1Ejr2u30EsnVItdMD6h2UnYTZgLQ1N9yJObdWO6aeNC5HBgJAl2S
nKdvJBh/F81V0qPw0m6rrh6lNeMoEXN3c+TujiDP+7yfq0CalYuBGvT/EMLFrnda02RbSMxUahA7
DNP4RZgcpKL/sOCn3DQEBg3qX+nk2ZD/m2e3pizncsTBq0j6/qZmC6ogpUXs++0f7SXIOv+PRuUl
HyV/5XGQioWEk2+JO0LehmIDZVQchnFYNuLUM4cb8dvBHVY3dcBafwIf2vlEuiZFnl2Ux/yGJ0Ql
BiAjI9SeSCuO17OcFJ96ZExcFQPlJ0VkSav9bKNkEop1q8lTBPcH5w3IxL/tBzqm0KOPGslchDjU
8/dStMaR4BSI+7YBU5eCN0l5AsvQ3Pv0gr+A4Gfc/QeFhtLs6tekA+Ld4/YYUndc6ej1cHwPNNNB
njXGv3O0z+sA8dLKKIgq4fi63s3TXjWnsoax6Y07Fg0oihIPMk0KzBslNWDLx4XrBZH5A6LW/NMg
bD/v80/rjOTuDBXrynAxvHmFgibgxoVDijJA4vPvAxTDNaP2S9rePDhMdCOAUnRj8BY+GXk2958/
7xZ+wGrpMRnWPtFRh985qEIWS7l7OXvvR1MFUCQ2n7Tqk0/LQl7JVEqRBieXqDVZ142/y0H6peYF
2PxSC2GGnuRLIeSasiyYLlAfMFL88fOilhmgJ2P3DevqFOnUiJmkngRvk+n27vM0PUNMFem1MBMF
Rg81qW9uzixEqKuIG6dflazGlFF2sexpYajYImt22TCq8jNIDVwb8j3+bKhacPR98+PSjufW82Sr
QA0ZB32noDQWc37FXgnlsllyfzElNeg90jghFULWed+C199EIWk2lKlxkRI2E8NwLZc9IV55A5Vk
/x9wqCftMm9fYMIfvi0BOeGJLnqMlBT4wAk2tsdQmJO50IyVzMjSk3Psu2hj4gTXClkpmUFj4XJe
xy6NUdOW66UI/7/tqdB8vVmJuZcSMYGq2SNJurgjl3yqCFAFRUdllA6420PdiUpdirBu+/oJKroO
E1edwgF1CL8/Q+IhUmt5/oS4vfqnLjCeG7r5Fi8ATNon7c6pITMcwBjfeNcoQRZ6kPmSQM0F8Avg
DpN66H+g+B5c/Kr6Lnfpt/0HAir/MxeOJjV/aLn/eklTIHLKcKry0TJzIVYgyg3OYir9smQf3Ar9
sC9Y3uGXGk45pmaWodfxpySmQbdIibtiQnCWPdPSvbGpWDacQ8hNii69VRAcB2s/3YorinoYB5Hh
zgdIVFuiz59DjsDNgo3XVp3rf/I6KXV/gQZfmR3xUUcudDKhYqtQI6XS8/yucvUFDboSrfJ92br7
FEUQhBKfIPcgA/nrNO3kPK6VPwBljCa7x7G6ASiIkG0akRqWrUIYJJMf/gqZCpEXpi1BWMF0Lm+Y
00pCcDU9t8m/6TUSTVMF5l1lZb/b1c+Y9ecoPafIqsugwVQEa1SXvpympuorTuG9wEX+k6VvHh3V
DiRAh1Prb258hs9yWw/xSbOIuvQ4WKfsGwQxcdwf2QJ3pG1OXVKLxbVSqs7GuaRVB8CrJNt4CIQ5
fCphOWXHhjnRkb3s2aryNUnJWa+ShJjx5bRdqUDRhqBD+xwOAhuzsqB7AD9RIWJ314zsHIRtRGSW
VqNW9yl25rpS/jqFuJhHFc1MHEhB3bmmhHHz0J0bpFB0t7a9F8QZ4q4pKs+FTQD+Z7hgh7AFqt9Y
dElhBotGUPhYfEytpnaM4Dpqx+iGS4po8vBRmn5n09468QTvJ4Ly1ytJtiIRjcDvPIyocNvfvMFC
2PknifzwJ3/Lo0NGKNt9LHHDiZWMHMn1IEbBofsTy1hexVXlRqNnIfu0KeGg/OgsD3DD5nk51vdu
MK8/ma9EUuDkpF+Dd64x+zYjFmReONDZn58+EOwS9fjU+lV8yAQkdDm/SdmT5Maa/lvEmKmbn5xf
16ak+Yl2DOG4JR0AXX9DWQk33SrKl5WGEt5Q/MzDDE82IVXkBaHsd8XUd8XfgFwywmCGmzWdyivo
cGLS8m29tJPm7y4N6t2aFTinCMUD1NrIGzmIsXZ/i4sTm6zX4HowLZiRs3BrHI1VldiRUPcsYrf8
exkrEGSmGXU7wwbzRIWyAVdDIWgjABYIA6POcdVEFUKY1mddSWQsjrTmsO/Gyof0beD1Vf6OsxPX
PuyYYwOnhb7aCTpHJL3MFHRvyeVxFxGwqbxx2i5Z48FtMbSjpPL7LZR326DgqV0MSOjQoOrbaMo0
Pi5DleeJVZ36qU7FPSOV9JQ9Yq/x/chJaULM3aG0UO77daEheLS5ztauCDxGC00ISoUHMcF9drvA
PFE/GN+cZZHfLzcF2RAtGV1TttREKWdtg8DbpFRDsN/z0MrkMKhpedDjcWQX4Cx4a//rWGghPURq
X7SAz6IcmL3qO/Gnj7y5epu70cX8IcO3Hc9xr/FJmGAcJOGgje0C1DEvQO6oBaXt/YrD+CHXNrpU
PxxWkQY4SVxyM/k7LUsswofF7TPabUYi7mUQK0H4ZatXTemvPkT2wRrZqjYilnf1BA7All8dEWQX
pN10wkFdNVTW2mjisavUy1n3PrXxe8GThx+zyW3C1TOc9bNOQHIMrESRljgbGpDFu9Q5Cg1UjJdg
t9ANctSwgIcK45YQjjnkVmmt1hLoq6M693FMf6m0fG44/EtwPLgEj8NsSN2BlJKf0b2gpt5/Y+OK
boiEIX4fEDw9FVS299rfDUiU7GTVKLYcb+iOhAuOTgfU+CFhqrnEtbmgqbM/X6AoD/gpVZM+dagP
kHLsTM2b2/4A3wrvBxlWSPX88nSU29mQcvzHtr445x50R+G+r0Z87k0bS6UeA8PJ8MWR/m0d7ulc
azruLE8nHxndcfRUFjHM073JozR86n1403/0iYAr7aHRImaWOlQYTtmOoCEhBjtorywx4jZVLvde
lf7CuxFMPRu80M28HJi+Pg6JTQmfu7VPZbQyx6a8lmjx7CepqoHcpYLJ4H6wMVyxfP0k7Y5AujrR
6G87j+foS32sUna7rmVWRWZNIvDjDQ26VGmLXMI1VHchHGIYa8KZOXlvBn2RmAXhHChBuWOSXIsQ
hF8ZiKeDpQtiFMG2CUZAv4q6i+Hy9TmIPEgyJKcJPbdswjogZ43mZCcVpiAOuYMlBpYL0/YkW2jK
yKHua9veJBfuLdzL2vwUAk2f5+KL6zKPaiindjlj38nQDLgZNH72D/mqxmRLyxb8wIQk6EGUQ4nA
0kUK4d0a+motpHwF0W74OzwHymMYGGquw72YLfUQlYdxG8bNjc82hbG/Ux7+xnxAn43RWemBSlfG
37p1yP9dZspolAOvJihXjbCK7AzzwOdkorGoeNIjIBSyQsTTv83aNND+N6m26YlNVoGfQbDpIXwf
7l+Z1si7tm3TRj5inLeMs6xj4tGGA7BscjYiPkxYsfiRc6y4kxuYk6MNFafZnXbyKPK7VAAN4B62
6j+46/oHn53/V7t2Iby8XxFn2bamQgZ6Mro0bNbVk1RA1Qkx6vt8rkUHcXupxD/UydAJkLY1kRIR
af4laffNKDQJxxkuuoVnBgXBNWcINL0FrU9CeikO8CyuHTEVgtKMyScMZlcTgdJKPp7OLD+bVmST
lTdYC1+ORV7FKIjy74uSjjO4cWtrrdoi7lH6KF89MkVerA4zny9HyvagKg5CAhuf17QXME6lWp/D
a1824+NnNTkegc0YnGWrMUdgm1BwBqbKe0DX/uwL+3HEVXDJAFp3howOUP9FAPfgx8G5e8hG1TyO
Tbxdkf2uEXO6CbGlShlU6014f6L1yauxdZ6vi1v4Vvj1/27VcfLDp5PRLb3CyGSTBPPvs/mFKcNQ
/6IyJfvgLF05PeMu8d2XyPIl27iuZVKyUZSqTWAq8CyMKhSdBXVsSOUGk9px410RWTfYwaxCSUZ4
lhl+A5hDYiq6rJjiQCkTQqoZ783BPXbyKC7oxve7gnI+3xdz7BHbTeYsEIPEK3rQNM6pF7fsWZgd
iAMDZ8tTfgHXTF38pqR+wN75Lk7v0uam2PBEqQ+rkErXS6VnviUf2/iGeQKOEkgbBhxs5JsgYEID
OzSlJy8Q9E/7dkHJ7Y72C7Lobu+nletBDvbTy86iLrEMG6/hgWwB6PyeA23aKynz4b04OzYhPKbV
UFKpWyT1NWWN6IgwMQLfnsAUWKpQ83BuXYCOsgcWk9+2EneZ6t1AWY3QgWMVbj22x3cWi1byiWk5
L1KsqGQOVOlIfHTXxXg2vgqNqb/KFLInkaUA2FPoN+oy6tichMiLArYOJYe/IN4PEwWNWwcYkk19
kJuPqbXcoOdQPEJmOaIMA5hhlcKW0WGVHcqa8spIdJbatcFwSa6QUeuLofzJTbCwCaRS5cgIj1RK
WJsC1rq+GAJk5HycxiJIunffFkaykKyrdPwboXRZV8B4L7ZdXTNKJwiUGGNDr9vUnR3m8MVBFZzW
HIiNMZeneO1bmvVN7M3+0RP0Upf2AzpFt67Cvra0wRkU6C566+uo+Ov70gUzTVl8nq02Br9bUKle
sJtPtypFy5B0nemHgnXlfQdOXflmMisgeHflSIbKFoVZRKAAIPJYQV1SZs+iiBVD8y4+EyXZKjpF
VUSecb8dLv58TbT4ypqAyMMijeOqmXe+XxVV4m/M1F+1M9OP1GDS/KlUQ05rsdNJYOZ/CSNcsJLg
x435xFvGqwr2a4rD4fSPdUanAcrmhX9fYBVmrohKud0fP513dafDtCX4QoNFxkYz6sIAFkfDXua+
asJMrUsII3/e0kNO7CxTTlV2lF5v3GGQ32k07NkQ50DXdhoRRLi3fJnkJS7LG1pEqcwIyXXGn3z8
AjGT18hDiF30xXDk7zlH0RQAznphanYByqFYLj/JuSgvBgQEj5HPxWCjC7mPWQfN2N9AHPF92duv
3E7twKFVsMrjAkizhvmQBWU3rLw60MM+Yl5ehr8d0unUUVsAxZrqGIFR7nZs48aMw6Do1lNAon29
cN5rXKIMV1pqe+ep4j6hFXc2y9YGKldctuTvbUf/BjVif5q1N6qBbc5WH7IwrbiCz2Bo1UrXDhms
XMxOc7o7vN4xBG6k2xMS3FrFWtBJadf64iGErhdFF4mF5Jn2foMQq6ipSykLQKEugSJwNK/32YGM
5Y2YecF2TFKczBiZil2GTRESmsjdf4pbJjAhu3CVKOVTGuTaijSLiUxY4CYlPJnzoNqp9GAJF2o7
2dHywNIeydUGuKdbk9Kj6Mh0LZMPHiHekVGcz4W/Z6C9uwQc8XVg/M6XblXCRiAkIQJUlwEHJeaC
oKxKXMJ4uwbMIegB3Ust4B308qFwzCON1r2vVd+Yg9/puNZPcRIa5WqGP7H93jwSIoqeaH6vGzQv
hfSx9HaU0j6fAg6mnZIZQAKP4APIRorLzWGMxeHNd9TQ8PL6POvCWOolhC/O7zXdfI+V/t1H7qLg
ScPVbVhos1mx/t6sb9QNREM/Jf/EkSnYv9wVqm3aToja5AA2W2Crmn27RaPHG+heDHf5rELKSzHx
vWrVQVX6WAcCkddP1TQoJKbVOK7z8ECFcT3M2z5DokIAnKJ3DBU4wZ5D89RXd4I7LzVIgDNqr31m
NvawsoHWDQUC5++GS6WtYkmsl2iDzeLZgblSFIwyjr1YZ2oKBwkXYFg1rPKy7yVO0Kf77N3bi1sn
MVibuTdiBmAfpu/TJNL/mFrvXVdGPe+zU/6O/nkk1rDd6I22QgFS6n5PW/YDX+OO5rvGOgK91Yza
J8FrMhFrpNPRPC9c+zVwCUTX+FO3BiKjszSPCjKDPy7u2JafewjRbDi9zs25GRP5dlE5fEkEedh2
vrXGNZm6x6nLr2CjJj6MPaG/BIBpuaSuaprMAR+R2rVD3HeJISpylM+G0vUEcwABjAbCUyKcDnNg
2wKIs+QzD7pQDlSEpTSA+Bs0ink7DuJ2I1J82jxbL2V7EViBbv2dUNbeaE2YVHprH3MJn+yFxyhX
VlSwdFj94p0Kwi8/q8o7y/+b7oEtiqGOV6i9cPNMxVqzCwLwj5AuugFaXvOdAaY7iuQuDUCRKiJ3
hc8pdXaKqGGg22IwkruTX5cYUmhMxkp/t/RTmVmy/Yp+I0tqF5loBRRu07fhwJ4XO9zPEAHqd9fX
ZYFqx8HmTOm9fE2lhhXwh2/EEKNBkykb+3vJVgzTb8znOLrI/q8UHmCAlVnw3UccEN1R4z6b7CBO
YrSgRXIKf5dZzUmLlxRPzv63RzlKoQZDKKesJ3QymW0RUZGjqwm1tBMhpeAmL1GUUBwOTDwU6UIb
y/r6hCrXkmwhueoFvy6roFdG6KXWzDzuiQGKxZGO5CE3Pk4PDVk379uGmgG2vj+r/z8zhds3PI++
4XopuiEJhe4PNGlWL9ZTSi7oBcNhBi3aWTZ8vMX5MDzahPWz4Rw5aqc/Wc0HCtR9DYM2+KK3wxUR
XB1Wi+VS4xRCAYTMfE7NOjJP5TAoNz6kdEa7qNMVnoyjGbb35tJyrBuJ1k5SD9F7X0Uzw4Puz5yv
eUYkMtae9eZpn2aX0kxo+nJW/xRrth5wdpinFuQz6ZlAd9XSLBYsBrh6OMbrsLj4NlPpIqDS+qF2
0RJ84ohiMW2Ow0EE8qQvNwodrdG/j7nz7dXyEoo5GZXQDaskEPOey5jfdExtMtBK+/gKjjHv/lSO
ds5syLPz0DRxebSouTVIl1AsmzIMBsmlfiHH5VrLe6uc+Nd5oQIjZtEv/jbJnLCfTz5WYd6b0GZI
sTC8sR/4+SREEIjy+DOppgFeI7DYumQZb52Z4vFflmVQu9rcNaiUOd8VSlyiU6MEmWsaKOw9CkNA
D7J/XCMeWuPb6JwUh3krkYtpAgfVE4wGJhxUOPm6WgXOdhC2keRZ58Uh7gHtUm/cQcrByeARJPH4
kHNmsDfaP5A1RPHmDMJ9X7+da+lTOhM5+bx9rZgHl2hGmTi+Bmb2IEVzaoyLVALBn4ASQia/aNiT
WpKmI6UtACfMmGx/P70pg4mWNDwQOcgW4KjULfOEiF97w08MGkcCA6J25TuqDDHmCfGZyEb1yTWM
3LH3O5KmL8vQfk2VPSyzUJ1GVmdqWoI6s4OXGxHK0qLlgbRUp6jemHWvvSMd9Amdzw1vFwFnc8/y
WYgExFoS1ItzerWsnlk+kkMD4QgtpcD7J49Td3C7fdMU0zXouoOqk/sxhMIDAEh46SPz8/s9gETq
33XBYQQWLwqh18d9QN5pRGKtotSmhnHsYTn8XBenjPfm0KLT2xwMnQCrM/2b9ScpDVkOYiMCMplr
eWtwpoUpFjyNeUfrIdA6C6EIXqZKjnAc2tvx0lTydPgT7dSkuWflC34Ty7cfpSMnI0/G5yDO1Ifb
6E3iNenYEL9p1XCg6QKWFHkGrATMnMCP61QYwp1UCwXmi1kk004cfmd4R1X+elCieE06i+m9YlEq
2GNCX1fUYC4/xN/voFSazzZi55AM3Nw0wGWKK5CUR2lFEegEuvZ8UGJaHiMnyrtfRrTpzrjdMB/1
rXnEc+r1+ROhyjWtuf2bc6j2m6Kv0QUBqcNDdR2dnK6SF/UygCzsFdeSfrd8pU5dawHbS1uF0/XS
aK5P/eymclWYfl0nn91Gfh11JFmziHxcbgRxzqY2NMqFfTDCMlNgb4BILGacFEV/JOqvkvRZydQO
WlSCpiosIzqNfece3VxgllVEUC9VpxVkV/4DhjZ83bZvabOUpHA36h0YICK0BMxT46bABKiHq10k
1CwG4O6KsMX5LBB1Zw6ptpSkqniFOL4DBMXMVSolVeNeX3o0TxnI3UyjP6JOQRWmyD5qnEdwPtOY
cZOLHzS/T6FzGIZ/Vj1WQpWLl2Y8g5iSmez7pQ/Z+YYjiuoqYWK5hc82XdA+erJbq+GdJLEKMaVD
ZeRffnu7cjjFu7Kz5C6nGpNbmWSEslATyjJ0Ve1K8u4MvMAerNKt1uU12B/sN7aP7U7LiB07sSS6
XwtutHh/ooxsnW4dGMZa/FDWjAq68boFj1tRjzAotOG3bO2xNk9h0ngQxxV79cCZW8XeEIma/NGi
uFH9xhCvTkj/zz83/OcRXeBnpMCB2PUeBAleZxn7pbbOXwpHVe+Uf+mqPR9S7P4nkEu4417APHlS
ombg2NZMqENr2R5Lx0DlWcwppGitu2h+THOfhBZjR1nCBsJJn8RERt/dd2YAGgKyCdcPzQTY2Ash
pCl7EWugewoWsltP76dK7GbuVcn6WsE/gA+N2QC6bZbkeiGIo7KSLb3LzCA1m+nsdGeR56m+UGYt
IX69CdMD3AP6QKjNTbCWNfcreniZDTQCLJu7dcHvBrENiji9KgXErd79ut5034HlchUdCz5gSx9w
X1O+SO+OUnC7INzS+7OT5+E54/AbmdtADZ2+5JgsPgaNSA/BPyV3T94iLJQFb53gYxVm80mMo6p8
liaCWBlCpmhHO1irDEmMExOrRvTv7C8eGJMZgRVzi+bfJko0YhLVd2MmJqdZfQIZ+2B4cKYgoAdl
SmXyk73aGfERkxgXkItMQxBAAlI5WmMEum9JgRenGj4x8IMHSuTGqE5ucDKc6pcg0inKIcwXPdMm
qUVzl1XnI2ozmh8Az+LdtyIuHXk5Z0XRqzqSyPL+PObkVmXR04EnfIhEsM/73wHrQDZ4MO7iFI0v
eJ/WOUFSAR+UjxnHiV1KHeFI1YuKRLxAdifGNSTZ676jOiZBVMkhdYFJbENXdUeObq+H5fcAskZs
dBeZmSOMvN4DGBEwS+tIYcs58CNP5mXJFc+goz+6rDi4XbNu9mPvEoD77k9u1wmQhu686aeP1hec
CN3jg4DFDoZ2o49ufZC7HoiVdpFWFCq24wl/sArJyTq8tm5WrRGJl5H/I72jsVEiR9H4irBL50UC
kEB9ZCiST5OmR9wI6dXvRXGqkyBZE76/uI6yz0xsA0PYjA+QAvfYyuiKML1RoNtnESLyJ3SEGUbZ
FmKR9XG5TZyoacQyWW2km/apOD3f9kCtJsEZM7umFSVg7y4lk+ivxWoQ/bT0PmmQ7VPLaYfb9P9l
P6twcQGkRlQlArnarsJN7GD39LjNM68qL6pUW7RQcn+5zJ9+JWeD/2W5Sb9fxoSNmduPHqaqjDzI
qlM4SSQaHWxWFZvpqc0G61UQQb2WFbjIMuwW2B+vAGywbeRO2J+m2gSrwxpR5dPdKL2s+iAJFOis
TDaJFnYcH+dNByrOiJK3jEbmlzNx+UPNlzwuBSTPKOcGsYQ6pNwuQryaHe5mRq3iKaj4NWZJ8FVl
5a2wMsORmKwzVU+3Z+IUL07u9o8dh77vp8Mp5xZMYx9Hbhjwe5wbcDhKqKqj5lr/DXKBnkXPNkbS
a8iwWavkQX+JDGMsXI35FidDmR7z3H7s93ydaexfKmMjj+T68dqZnqxa+yhERLX3M6dr7C7g9qzA
ijXo9H1pFNfk48k0Hq8SV3jY9tVTwqtU4UGTeLaRz5jyRFwfBq3uOsUAx4+qA2hxQb0EJA3UxKO9
bn3kHrgaj8ioE+F+LKRdDnsygWS1AJMblxD8GMRYduivx/ZA9mJTJSAluwlBY6vHHOD8c1d3gO+q
SrLWPdns8X/2pSR8oSZsY/WQEhXYCe5Oiod35q7c1JZttNF4b8DzbwE2ZsT0CIOxnyfIHa24kiin
xDha5hnazEJfoStkXjeE5HzuPHWKxa9VjV5fqcK9/VKktVX+6QQp/dNp8l6DfhasKA/mzs3dTCuD
u47NNCye71u7bWLWzWMH+Yfe/VCvCQoaolJqOcdOKPFFCa2BaVvHUrPp6goCMiODdtgE43DrBdRf
3+hb9IB6CnGGnZBSMf7ZgKjjj/3uANeeC1WabmBNxyA1vHd27iIFkxVkb+whK9ED4eCh1aG1yPqf
MjkM2Tkd81EiAACCfETR2JnfGKvMVRdYnaStNAyji/f4YT/GR7jL7Ovqx6znkTJdOdIZrb0HwCYc
4lVccuWTnsSWwaw1EjCIcbFA/FGbi/C0sCu8ASEQiNmbi8nxof19MhboPACIookpI2o22qrM+267
nZ6PxOpRZ80InPMuwvlt/bm8qOK1IXZpZAQuIDByYduSxtZ2GcNJRoiz0Z05UyUV7+XaxCSetL7e
if0jDwM5qKpljAafNcIDzweAmbNnKeWC8+mf92LgsHu01pRjWh8/Sf1bNYR/jiZ6jFSHw7diMpCE
5H5vcjtEUnPhtOQULC7Ju12u861sYVFG2fMk4WD5m17pfCQX0bIF7562D1vlBH0mGEyOxVxJs988
1KyUSltWJMXmoeYXnzISsacRdnhOnSKS9ubFEXBsQRuquZP3Tt4PVNL+8ANuNu2bCx0Yolu+lBuu
aWaRACcvyYQKOzMBnZXo6QM6mO4jvDfPuUO8Li92MqTzb2/BxlW2Uto9WhiohkwV1p05NQJM+Pwu
AD2PHjI8+fm4f69Fn++ZFzpM9VJBSNAc1MvDZzGzA6YwwydiN43PgynV0Sa5wmg0Dzq/uMH+DpHm
fVAr1jpj30Uj8EG/Qe63158RZWep/W86bx8PvRNB48PbKlDWk+1Md2ab6O8hTz2+n0fhHsSPhkLO
/X1qJL/diL6Xkmq8d3S/bcMiO4FXQEupLQ+mBWS3AvBWsaqls62l1W0va2uJFkXJSi6IKZQCOG0t
HGEtwjpwBW1M0R8p7NRNY8qxYuVDRNOqJWtwt6YvYpEb623DhI7GW5bsr5QX5IslFkdr8LpvxAOW
5xHKOvan10BQ++KtX90KV6ogGpHpZfkumvvWZAxCwP1p7XDCpoy/GA5hZoKDMGoYfAAYeXp6j7q/
aGevnF9jNd3kQDKgnKnlVBVedi+Ysv3fckGaCvkWNn6qbkz/kZwLoJ28ANRoDh0T46mAW0EczXJ/
5EG16WCpflTQiJxrcp0BU3ujW7l8+1l2qtolNxAjsGTXLEen0SaLfaSXGIERI3mfy316+V5wt9UQ
wGNk8mk8048cBlLXalCDJLAj6Sj1EHUFyjbG/u21iKJsV1sXwdK32oMa+gGK1tfyMX8WDwkuNZUA
SgXpvfmbfgrWXndrPcsNS85a0JQJLS8XsI0UmUmAtvdzOO+vyKYLnxfAH3DOxKbD+U7t0DyVR8s0
rBZz6jV2tb2LvXCbKUixVqzfg31kyqXwTh1deyUrxxmU7pvBqP+u69HfD0ZPaEXF+MwZsaStL/V0
/dkn2U3Esmfn5i0U1uq8jzTUoDFWCmxYw8e7p/rqFZiX1QeOuaUk4qzxep/TDN2WnoJO18eGcP2D
w5dYuIZWC7xBw+hfK/R/beH8X6FCCkaTzlWsRP0JA4Fvm59uG9GtRAKx+iOCKumagKRUH3cdfqjo
ME5emWjLSIXOT56L9b8ZRmNUJOA0tJyqNqhfBoBV7aAOa9QyevvtZGQoVapcyTbaRsHRD1bx+JHg
YMtAbte9fjGTfM4jWpPPqTji9ZghQKrNki4dCPUuTzAKoJro6pGesyRvLGKIbbUwKhIkv7UsBVG7
rlEJAx+Q0BbSBlKSGFAQcfH+zje+V30Rxou6MmqXcMSY1uM0K5hCJv5D0OZ6m//YrfqXapy8ULkh
5pUuVIfMOYv9f0vH0mV5/lCsrBncgBPchKokokiKjZN8CjeR16jnMScJ17tskZ8x113o5rueueDN
D6UfUtNlRhLvelbwKL5Nx7ouS0TSv/GsriXl0o9nSgwgyFcrMgj09CbnJ3ZTfCaZhAYJ673r0pZP
IA1NcqWy32JgzphwiMrV2rR6xzomznAIOLZ6tMDhtVUoPVtIxHK1lNqCwkZgSNUO5V8edKG2hUv0
wG13JL5rg08i2PQ6QSnvtCLQKWd3aEPhZQmXcgxmlK4OZeEe2juP1aR37naubUd7ha4XupTKiOix
yjthULVgg+EoJZ3oeg4w4xN0b87z+twcqtcoEE3NBKNaXBcT1Jz3whbwFeKIDKpyDQm+zFdbJszT
uRFsCt9Jb4XzcLycRUE03C4lcAXNueXztzyZQ3xnfw0JqeJRoaCpRvCIajjNz9ec/Xf+Lr+OGZxj
90i0DDW1x155/qGjt982sVRMFrKRhK8Gp4prrnzx2LyQh1zd2PjqplxrSatctfoNrcbO0U0q6+wr
yQLpyuVsa2prqkO+wgMzXU/1hIwhWKZw6z57ZuzogX/Ndb3gIiAFQQWrF5q8XkJPqYGrtrkyN79x
LGm60U4L1ROaiazB7LAGryY7X0d4wfiGTKiUQ+vpHoFcfOQXcyi5iOtPj1foURjG98XB8cv0R2+Y
II6C0dc7kjrqeNSLgHLYueXzXMDAJdHHvK6tTbNpS4San2uXC+w3v926HMKPKHsVoEA4204IThgZ
wxu5Gri2M59/sZZChJPcv4t4gS+evI/uK/XDCARxo7WRoDSL0TuAZs0ZSz0aqVKAf8rRuKU5MQ9R
kxFN2wpVtTOFMpjd6TOIjG2RZhE9fEelUG4aTH+SNvNPbFIX7te/yBR3ZkrC7+0e9iXCoSnyA4kE
wRzaNo3nl/slvlBuYOxtUzIbXZyh9QEZry8BrTeS+bCP1hP1MPc9r+fQ5/YYzuUT+6NA7zrnJilB
ZYLeqE1tbmjeX2YmClhxZ9huBt6eRtpQjdIqJNu8MYkTm8t3gOAbzgSVZVAj6MEBgEQtLRzolWUq
IEYafgPs+iuAvEfyZ+J1ImtaEtb7MidnRaDjBeT4VJqXV8Cy1HmthSVhIO9r9nbJZXeFIN+uaUXY
IdJRSiwSAMj2KzSX6guOQQUGS6RBqixIsqeZ/Mtu4vDBA14gdaqxuoKlIJn+yNbKQk2IPf9eq4/L
xAcssP4hHh9Bua2MmRHxyv3tOT6FVOS4vW+K6L/GTwTcGUoPciO1A8NcYJ0Rum3s/UUl4OqMGUmX
8NRijnQ5+aU5J8sIF9bCqlgsDiCGMH4+XS54JhVaR7tmylFuTruuXGKdOzsJ+OWiE4x/lJSooEnC
QC/2P+12w7BmZ5KjcknMbBcvBBBLYPwA18ekSPdF8+Su90nW+ItmoT84MeJoaAkbihXqAG7a6g7G
sOgaewDMuA5UCVmwkZjz4Lif+OLn3gXi8jzL0NGYmUt5OK9FvRYtRmcz2QrN3v0nFFXw88Vd5iDH
hgcqk1quFXPN/RBkqq+CRpLSQmQIo75HHlMqvCD2PLZeBUzTA92r0TGM5g+K8Jsdl51c9kkVC/7W
sinjBeP0eWvfRDnCwkkqu09+BA0O1hZ/0MqrGk783X0IhdcdM5U+20R4wq5Io4iHi5ENaVp9Djej
9hiQTAnjZ3ZDANca0+7lW0qy6VPvmaCy/1HytXCjltpzeVWtmQBWdSwMdeQFJrVe9ZIOmzFO8JMA
Y674LGJC1O+8m7EXra65I/ZGkSykpPa5d1XeaH2mSy4tu+neLofins19FqfcPITXQ2hi6nQ/R19f
etu75FzmI3RA69NJ45r/LOpWZWsqsyevkzftlGlGyQq0zvqdCFjDxcWrhY2//ybag57nFBwqy0rn
R6Eo1EX4r8Rm8pHhuTraGG1lux83XLLjps4t3aE0u9ptsX22Ss1MDhc/zzEYaYj+yxI00QrnYRyY
+iZ1fdQvA3OJFHkO1HSIVncun/ocX4D452PzaOB5dv0r9d0zJwwnadYW0lKC+RXg6Y1WySVqwc6l
NuJBaVgGrUWFwdHqHIrekIv5ljXC9WbSU7Jam+QHFECsRj3Qkr3JZvNJNriGr+jDer3O63oSZ2KY
W05B8LpZG7bVJQ1mht8fcOYJ5Yg562KpzYkT4RTF4kzBgD36zBqFOaYXOlNvpUBBub6TKIBb8whY
EnhK5G9gSzk8J63vY+5kg5+V50/pzFzhrcnVntWQLGB3Sk/KvXyKWyspKH3CSsVCrP5mXFmLaflX
TUy6uyruQVo+fnUux+9Fu3trLZU0jD8E9FQbY5X4XjxKMSNYuvN9qwzZ9KNsMI1CWw/cl5WPDP7T
TiJDEdRbMTm6MdmT954ZL6g+DF4RujMbncMp4RQlr/sseRPk6jpTZnIkG5Ivq5tB7VUGRbKFereD
WjsGrbQTsBsuCITt1hed3UqJz8o/RbJygv98pg0suqUrd7kLElQfVaFxRXaJro58CZ0O3LINnyoa
D73XO6PP+53XTvpAe1rAz5K/dnqPoWBli57+buTrf05GfK8wsA0GONyml0+TT9aDhdZLjBH+7Ry2
DRG5i327XCl2i1Ep1ZVjeBZxofa8S6HUQwfNgo3nnJ5+Fc4w0H3w+ecTxnY33Uzk2lyJyYZjihYn
v9zGyfY4ZC+y/8lvazu032xkudUqFJrP7U6B4kXjwdNDWNLCwFhB1epWIanj8+vJ5NIG8HiSkNIq
94pvR/COA5xRc5Y1QpXfE619jL40XqYWNk3LLIdzYYLKN+Mu327T9RhPahnJVRbN7G+Ott4ZhYdH
/ylpnEJRbW8aUZ9Q8G+RRWY+SMEuNZc+bxH8zP9S2LZDVhywkdhyvIgMqfTw9kNDMc0CmyW8Yr8o
XerLX9JVlgzmin965SI2WG/wQ1cyw4wVwJDgj8ahHEkUjYceOar3FoXr8xvORxjBa4Yph0628qvQ
W5M8/++jdnNJqLAnyTWtdI3DqWCr+zRm+9a3PbxCoGQlj0enbcHSAh+rU7tXRgKpU0c9AXZbjWrq
ERsRkpRvkgPIxaJ4YgldhYMefqj7pHKGNUhuCGADgQKlMoRvCxawwCEQ74idFbfCxsc1Td57+7I+
pbny7ztrL44fqTRdg7KgwCwLRhQZlDwAFrXJSeyXBjeadbgGlWUw2O4uNpoqC8wNFpkr4rPdJImk
sMUAO97JqDAYsp0XquoPtBrB7n4YjOrtH9HnSufjkjLgzQuICbGiICdDCVwcFZthocZRw3fSwZdq
cG5ZPNU/p84G6PWllkHgpJP/QDt4mNwC+VXO2X1HTdAeViC8eITq7jZ4qxnzWEVwDnk7ZaCfT/7h
2MFNlvLlsNytpM+RoreMdiFAgjKZ+s9Yzi3Ft7lJk+Ze0ISQwnQ9metle4gyuK0Cvt66WYrA6Pm7
jPWyCyxyV9TUXe1WXFutMlwUvU/u2Kl23GkHGmyB5mWYdiN2ld70wsuBvFTWlJc6UE97Dpm5j6Yh
1klm1XQEYJ2/BpALT32A9i+3/WJvyeJcVCiGaWB50DcmCRsiKNG3tjwW/a6n1byDyT53zz2oGg+m
+udbXsE3YfseH0fvxdPZnCZ42lkEljW8oKdRZcfVDktVRvFxbyb3Z4pLDPHhLe+w+7slHr6FpLcD
y05da7M1Zv5NSiinVTNkoEx3T8AonRFq7ntfnGyhN/QnCBp4PSTFRnHLB81+Erf+2FowCEJ9v50P
dkYm8e81pZxg+5v33H8HrN452KtL3dPLoOXfxEWpwbRY9WiIxwjAqRxKd0iSRbjzzGcI0NO6r34r
aX/Bwe1ev5gz6BtCEI7uGuPKcGLSbjTBHvW3K+5cEh9gTgmfOG6lL1hgHhqUqxb62N2228GeZKpN
lDmaPBCncFuBRgzaCt9wMvJQEnh14fsG7KIijDe9PW5fRLzVZbIR9s90xHTi+0C/Vgmh/SD30tTo
q4cSuCp3AVRmAAxqE+edt7G+MNugD13hiZfbqNoA41Z626FQXKWeaiNZRsPYVCmV2jK8aV0auLWz
2TakRp8NuBsVwW2jePdQsf/Sjkt3uCvOnkpQmvyrnUZzPv/Jn7Fm9wxyW+hMivc11jdPP2pknErV
NwpdlMG+PrPz+D46/GGPrTCCQUtVeUGcAuZddxffF8tTfCzom4iPiSMCPtnmqxdGg3SlLQSuEiVp
euMRrt7T4aY16WdWXzW/ZSzaTgpA7fCyRve8EUTl21UiMtJBJQS4g0Ca8e89g254u7HyiqItciZc
mfVTbusFiwENvwQCrKTjtWbDus7WpNUn6f0TRGprIPCv2hkh8Z24a7wDksorkynueBbrqFSk6E7H
O0GmwuWVzxZFIgkpieTatjgxESZFn/bepkrKnskWq+y5Z9TuviqJ/NXIu+rcAhwDPoy4FfHL++Dw
ZpRWwANmfegnKKfwYLWkULt+DrgdE6GSD15GYjPuB2rADER+ZTQwTiGuyTtpmsyk7Gd5PYltBA6E
8ffTYFwqmeAhmSAMsWP1RkOAHy+AJJOyaBkCTLsSjcmiVmHWuorFNl4eHw0WRiHRXa1DhFPHzQ47
jho+epz0vlzAeBIIIJ9eER8gJOowxtcq7nMnYwQph21larhNDaqPrEq4JNTUBoLmGa9iGPrlALMU
VSS8N0VA4s7BJfaIsNeCSmZ86dOLEKicAtiUMIXaGVRQFlyWqWBWRroMHqXn7PfCRiMDFo3q+pvZ
CybOtWhEJCP8G+FSAct1kkIUEvYWAhN/YXDA6eNbw5Z+Hr3MoDxMHV6Jj8jzby/ep8v88vmMFZJ9
5RjOCvdsSvoJytdYBxzPImgPUbRPJpKktF/U9nMF7XpYC0n/6xt6MQFmARkgOvpGtQf9uQvPO3au
7KIzI1LCAslUXTaVpdz29HUuWvkyh9uJVMK+SmDpVb4+vDK06KwmdkEpIzyiqy8Bz3R8+M1NPPWE
G3yHYO0hlH3l+zMqWyY6ih+SZ/mCCucBdvcNK0NwIwMmhX//BTL0GWdi8eXyBQgF3A8aBXA24l2T
QYXtmymf/9QLEHKRorV5WAOnz+tqnnAuyiSnFkMuWx/5PwsM91YdCz4owR+N5hMjHGpZK5Ok9zas
r6x1WkPLeRWvXiUVmDtGG+WOR0d+mDXLTv9Kho4qeJOAFTqSjtq0f0J2AJ+lVju4F2g1W56agUd+
Qvb79JiqfIb9L3U8HfHl+LBZO55Wkbf1dZccqb0U072NctHXzhYpdAqzUbYhxj+wG8vsmZSwW1BP
JAkKAbvcgJVcLDEmRtq607Vsan8IPaFFg31ujvC6ZnzNopeZeike++QzIcpW7dxJfcGy3cgJzwO5
uu8yGkS1qHsHTsSyiqkV2XUR0/NvR0qnQZKMlgoRFQj6PD5AwWAKBpAxyZVwrFR/kdoeMuqLow18
ImXaciwwtTVnP6i1R78aqq/tJp+chSqgOC8FgU+IkPp+Ki3Wm1CuJhvKTHD939EDgENK4MRPLCKa
uXW0AZNiZgEwzZlHHm4E4KpkrSbQtHuCdkqqggKgdzUzaMAn6LuCE2ef/eM+1WR0gC011mjV+COy
VlocH94eRT+9zB1TVDB+hMhNnHqdX0I6rPPsDriP7+7+9O3ax6i4KIkDbTMs9s03tgiXf+5ZF2F0
DoLbqAGbAcwpxG8+61coimdvemo/CiUnOtFtkCDRIqGYg7uy37ma45vqXXrRdY8zltGDSvwpp821
E7T6IYSe8qKG2aSzJNssYn3ifRLU5+TlmdKvuo5IpNcxo6qczuipowNgzQxenDu6oOM5bGRFwRRI
sJ/zAI/PixtF69CRrsylmX5ekDHi8itFm7w9dloVIvZkm0lUmsrbYUqveRfh1AxgV8N6S5VvqtQI
qYYx7FMKV/oJEq3oDEx5lZiPOCXKQREUMHuSiliFpXWUV9gpgE7+BXQNlh9hvENyB3ZI0D8GCFbE
ktxpj9RuFVo3Fjut/VgwTOEiRQ5+PebSujW7yrtaDbWF7yzIsXL+74RlKWq6S7AAYazB9DdWVBXh
uTVG1ZOTY2v20c3CltlbP9sGn6FhGv8xiKycQ5uKycyUlr92TikgV9c8d+3XDpL2gXlJUBf3b98D
Dj8FfAVu3fQ+wg+vDPA4KcQX9dk3GfZ3YtlpD0jkV3OSeO2BejxyAnPvgqe42a9vYVo6lFW7AviP
HKd37LRV0lb/YaV7JuX6IuIKHxOLFqBZgt3jlQMwMTwvSu6M4cJ7ylwRutYHUJxUtCHjpA6h/WTT
tByFQIWIQ+tcDARfOL6n+/NgwfxYQMSxt37XCrSz/DWxBcCL4cGwlvVxqDDwgLrbLH8oAXA2DtSm
HBJuijGBEPQPmuqCLFBFOKowSbai6GfcPWEaUdl1C+JVOMN83teb/6WhEaz2peeYkdcVCpBgVTWS
tMVRMT56yFF/OaoOQ3gT8Y+iLRuGrJRDNMocH8AjOtagrfO7D/LhuADuxD4wkKSl1/uwj0JSL/PU
5WDItxE2SKqCkCtILzB4OFYJg9e7xZhyUcRzjN2HHvC2pd4bXlObb7Cmcf64TjAlf2uxkzSvjz2n
R0y9s17furgt0lHu4R/DTocJ4SLTzljCsW2xQdib/qwvwmz7/tvjG42RmbvDPxineVgmcXO4gHsE
MFCI6X35HFF//cve7cCPY/COlpDIoxE7BDCr/PlDCl9oNDjrCKsrUl6Aq8OZnscZn30vxJF3rBWB
WCunMoYOZePjU0Q30s/o7Bza3QqZb8kQEsrTtqILqMtC0XJaWyfEJ9Tw9wLQQqYmkuG8fsuaGko3
rLWwZVM9DEt6ZBuZJsApNSJ4TM3QdSGC0uSpOMw9+0CWEvYFWF4ZPUG252921TdjBSkiSLfwnBUI
TzNpqMOt1eQnqAt2HdqgL0wt7BAAiY50zobX4uhbuEsZq+PETkp5Q+tvlTZkwtRsg+wf/EfhV7wS
CicvBNg/3q6P2FB/G0CrKuicQOCLnmuX9pcA+sXa0HPFMwZkohdnyfRN4kZJE0VCnwk8UP//L7kM
rCWXmDjMTTBZ26vqy3NbSx+yr4afi4oZsuxsqhdgQ3DCvMr4l0DHJ4eqeUnIAN3lz4AO+mJ5y4V2
1mGixEPeZbuDe7/Uc6sGc9PIwMrw6+xSwCtg695Jw1j7R3qckfDreVW+mXpQlIH/49577wcCsWRQ
pUMNh919S7GHTEBQ6hWSMib4AVq31bsBYNcSzVdAyxZEGFWre4ZexYNA4Jxv/j2oy9LF5ssTFhDd
jY1URf5gRWuu0MRd0sn5XGidNkh5sS82EYwZOZIukn0SZK7LrXrgWQCX+s3tku0l208CPxMTO2uM
4aTj/HdZa56Vj3PskKkKtKUGA12rBQjFnhpJu01TK+YOcat79C5fycqFWC8fKqswudLVSvReqRGE
53zygC1ENz6H1KGbkomEnCR+Od76VwODlurR9tA+qrVJOmaJhFpnEryUlgalnqt/YOhrfeExMBiX
UQ/lZXqhK0GryOwc2Uqa9GdBZ0T57wROcz7/fptbN9AefwTERk3Y6TZ9Aa2HOTptRJHGvV0p2XpJ
jdEIMxOXkR8MfzUag30NmsCYohX/N8ZTCfkImq2qBTU9kVmoZyhRnUMrhK3W4QbHFDIAK8DtyP/T
e1PlGL//A6uK8TSvTo7uZSacg2nJ6EvwAHdhrpklCy5cBGqldfq6b1OohDoUPoToVguxMZ4jjBS0
dkxqOBH9l6ErT1Nz0yMpWw/PjvTFrR9y2hwoQCdAm9N6zZRg0ZIvFy84eC2WJ94aCuq4yBBdmgUS
CvgyUieHKKmaZLxLiShOxPiMKjLgw0JYHML1FvpxfCPJAikFpjmbYaPugazuGslgbwEELSA/SVXA
TjGJ4Y3qpX1WcriNP3lPbnNeiUB8fu9EfXoiQ6JDZvwHNslZADKldG6VkymYY4NOCWNUEUK40htW
nHqD8CRH2EnIIcdFNrC8Ip4YhkPuIvyILpQqaKk8mbOGjQ2V7I2EvTMiTDGahKQwcJUkZiOWmUDZ
Lq3EQp9ClLmE6W0nEyhGWd6mfLJ/UtEGyUAspyNFGqDm6xD873pSJdG4Q9tYhBXXImYlsfo2FaKy
kA25s1MleeZqs5HM63uvdQUOeUp8CQZr6Hqwq6sjpCIPDy6tYkyAl2K6oMUCTLR0J1U2IC0gd+g6
ZuqCJhjipXVMJH0NyxPRTsbhhjaWNWNVoIOjNypj5eiogtwnnVxZkJnFS5S4VVYTPfterl+Q7gOR
RkNRloT5XNg+eCV6chOBgchDbfzJ5flgscSr7u3nSqrcbQhNZJ4XgSFG439Dh2HHo3zOew/9IalW
AdP0babV9QAQR0GPATf+Tjlvca3EMY2phBLqYnhr08UFXsoKknTmqAKmqXfnDJ6sXg/macuwJLoM
Da/l3LQCzCEVeuTp1NdFlRWhBiNWjZp6XpXtsxZSH2gXjKy4sOZ/IplZCRqMEI8hSRO+KTvNzH6p
0tbdzMsHlwhob98a8PPTabZh6+DzJmLSRGKzZQ/y4ST2i42bckGF6CyDkGMgBA9OJL24/OqO+GNQ
OX/SKPb9cNwm70sXl3uADRXCbt7Com1m622NsxCpjCYrYcG2SL9Qwut1UN7u/Sy3D9Fv29Fi7FxV
/JtRPOrPa5FPysURTab4/ObXuNaSj6EoSUxI5C90lG2+PlvKE2W2q61ziFVaae+8gepbDZCjJypD
Hw7vh5OO7vFLGEnBUJTjuurqrNKtfBcSOQOthhSXXjUk3SwT5BDIYrvZ3P8PsnUdaWGBssclYdWS
rN3+etsyMgdUfqR7XI0ag4tXmUa/95hwTPm5vJIdsJeRnw2O670nsS7D0fs7KMMHdfrB70MxFBEG
a61AfxgvtLLNBpkkWz+ylB4tU2q8KAj1hBBADrrj9RwRhNkqRz1UvqqmwFgSfXKHqGYDpbXS08Nx
E9GF/Tt4gL2o7ePgXp6jHLf0KxeTu5klVPEGYG6H/6VJfSB1dmavCUwlAcHsLCt3KfyEuvfVI3UT
ETPb45YYhOcsOxd898lOcOxLzj+9gbPwgqwhNhHTZIXK5ZvcqNfZTjjvHGfs/aDSbiuRGqkhxlk3
iLFblYketHE/R2j5ip2M/AhbftYAvECfSVbrZctUbHyydUQ4YZIe0OjL5mmDfSVVVJgxBBrXxbEE
W6U39uI1g0ZgyKddJPKrFlBniR3gzmfITnxkalsE3wmtQqzyZywXgQUqKIEeAZgL/xVoV71r9fk2
hWQeY+9jA2RY+9vLEGmlBA29AOWM6W5k/GzO7WaBqRyofnGE/lo0/vfpik5YbKSkRrVzTjQFqNTa
Z2bNSFJkh3RvOIFeC1jDDfpQHDyT6+YzbZcS5buN9BrIgCOUUc0a2/Hpfu7oeTtjikqtD4KlHLIl
CWi1Jq4Jg2SRbxEwBQNgjz64glvqgzHTkUO7fANRs5L+x1CP2TWbYKcCNf2jYwFe3xPiERpux/HS
xTCuLNdPV6LZyZGTC3Xn9EBY+t/u7I/9UThJ3S9/0JGKq/ll6TSk+d3Zd2yWIuq3q5XhtPqiY1oP
vZo/FdEMTotBmWJEvu+E1XjCOvM4dyRtTkoIDR7XLTogNqFnTQisDOMaiZ5qkBl63qj61KV+FWhi
G2u25Dnkk/drBNxDXj2ZKQEflH8Lxp42o75kDpPJNMjAkw91S0q5xfkULiBUfPDFXsGFUxE+/nfM
UaSF2MoeZN3vl9pa2hK+hYLkeZgE+aJNmUwwJx3QHRAI+ZCBa9GPLvFFEN1HiGASeRP6DhiAa78s
h8fF0VSHsKFOSb6UUWI3Lwx++jiLPb55ia7brdWngx7rxQt1hewjD4lAb0oxYhzJUII8VcsTVDvF
b2j2EyJmRbWyksWMXfZr+irtbbZ37oc7X3WIEKr1OagH/LF0WkVExzMC0Os3ieZqPMPc2z8yx0in
QFUjHw3gXRHV6hIx/lbV9fJFDHElkC1U9Gg9vGLV9qQojyOZHeyp+kD3SNzwgsdNhhU5EwTFMHVr
ZVIDLwj+Ua2p0orknkEQSjXFC98zcDOW9l/Pmn5wwKONu9mNZ2Pf2OSzPUtPlWDGcDqFhRQfrzi6
1BNINsn8m3tTzSZgMbFYMVFSMmXn1PEBXainjdn8+OwpsHcQcP/HN26UWRaKA31WvgJL1aNKphsa
xGOjVazsgQWdko1DQegE2/azPT6kW142BzOLB9rpqOfa0rYaHublQF6p/vQ8Y9B0Dg7SU/EmwiXP
JEmaS70RIh8SvKDhYGJtPiSilXdYep6r4TFJvVcwqGp5DCyr/76zLPAl9ff4tbnTAMHWdmzib2O/
Kshp4PClFXOZQmt60/MRAb9tznM3z+6y1Ber3oblK/oQZ7KlJOZ15sz9cuGPHF9hjwxDMzOK8qTr
tXu1mtrLCvTi37dGDTPmeYjs94ErOw8OTx/TW8KN/LraCe9kP9BgvEncnMbCIl9jmruWqlFvuSyw
UzXype3QqKsZh2+spN9faLsGM1OQINM9ZactEWTLsMjoEFoEjdYq3kVFyF8BfMS/hmpDGCWo4qPm
FwB8MaR62TEzK4AHGBsbJ/pvWwdDlH+DakiQtxfF6sdJb9z40ELCQHHTJ3JXVxrA5wFJkEKVXYiM
4pY2pLcmYg/Vbmel23raHmRNj7r0LWCjz+f5jDW2jHoA3l1z0EF4YJs30hUlewBYkV8VZUejTSoR
8kpmFjAXFPgQswZClxzjl3MY3M5e+TED0WZq+5fUC9+2zuegJc1H9KHNspUo449GLXmWguXY4RXb
1asLVU4BIZVSkUoEcwwYC/95ONQkdXHrBu13VQ3bxcf/HihmVUOTUD1cypBffszlOtsDl/MYCRYI
Zw3LNGOR2XnfKpun6Q+9KNIOP725Ai/+hcPcCKE2jkDlm48Ts4F6coLNDNNHuHjcTrCFx3C+UTK2
8TKmOzbCt2ZtmXLHKGmjuhzOV/Om8Xtumf56tDS/NexIx1ltrw/M0rMwpFwAzy9/5Db44+RP9eue
lUBfv+c2Ltgs9/ng/asiPUgHFuwpm4kEawQIXbhL16Y5y8TgE4M3skr8ZtZ0/4wULhukUPZ/reSm
QKfE8xfEQ9CoSuMPMvec4QwlIMe0c23v7YkSER1398frLCmzzNYHDadGAmfV5uMXj03rnXlA52Pu
uYZ8bw5os7MJ/xfpXiBtIcivh6J06Ct95d9zib8SHrIOSfc4nr2NEef33QnaXCQLsd9ZLH+b9F0I
V6nJn2Vxp+n2gKjCGtOK6S9z4OEkuLmjY+uwMyami8dHaXGsHMBg7sjXRZVazvDoM43K8AQM9mKA
YzRD0g8Y4CnRtD6USgAw7Ba2LooaU93IAKL642y0q952FA7OH5U+5628bDI1h8DpYEfYzFgexauI
ppg3cfsr1njaLZptXigLCrQ74mjVo/gVwb3hJXpAj3WYPuGkeR+20vFxd1qA5rb+/pSwGRphTq00
DoYY0Bola2Yv8fa8Q5Q6XG7NSf4sMlijKhInFKrTjPARhlmxuO3rka1/XAD5BqfBicsqEZesv4Di
4bt3FwkxuKqgVsQ/Kbo1Xl7mjzsh350YoOviJS1/BzfPshPYcu6tmLBXEiOx87MLR+KIZ9i0WevL
gct0GGI1QEjnS0i4/P8/iGMDFUQpYEb8m+Mcf7b51+PiNs3aGPzRhuIVAjf3DUlVaha0a114a6YN
h5sxO3EpGwFjSEECNyk4xAfmeU0KgAajiRm/RRRtlFP+/Jlao6ntpplmvasv7TKI0/GKeuu4noRZ
4sfgE31tqlpas9dXx8aG9o7oTJbp5Xhdb4Y2cOWZAE7ahZ2zD/hccvj29sDJB5s2+Q9mA80NGAgW
Sy4GnN7jsBJyAyIUxH5X3ECT4Lgk0BVSbccf+EyV+IYDOxuk7lK6X7Gic9YnrkRWJfMnDnCOOZ6d
lPw6WCIsMFymvx8/YwJt/MmuVjHKQLtiwHzHytjGb+p1G/n7xSDKkM3xDCvmhIvNNhCkLgtnLKPo
3XNlkrbmot90oPMTIDBsRPGtfEDZw3UfbNIWrB4mA7fkxteyLPIxf/nSra0+HiXRMATBLQxnOok6
Jj7rlzp3XfC2L5eYokeoMzK3XOYBLoGho7UsM1cFI6KooJwYKm/dw7cYVzm1D1++OpLZjyT7a+lD
GfJvD7X0V35I+G0sZmQFGhoWCNMtWk6NyRW3PKt//A6zs1dCHUOKyA39vIFE/pt4bGGQfPe3+lXw
uaHEQ9PzU2xhwBbR9s79RLiHTNJ9kOuqfDbbHghSqTTMNI6JblQA9tCA4KjbTz3zJKwfQC6ELk0N
fF7nP4yVVJbn4quCw5gqo/IklFeQDDr82aNFxpdxTqXoAM4vJFKxSZ72pIEHV8S9I3DGH1tFLPUv
As9S79YXuBspbYE925CUhyzKmdxMPb2MiHD2abMw3X58Q0ImisSWOqoWCaHL2Y8msnPOR+YmyLcT
Jjw8Z5TKDyDyejDTbPe+hk27nlRwZd9Gvx6spQwLTh5uAV2l41WuwQmkZIJzUjHv7fpJyCqNZQIp
v5zvBoJeU7BenuVMaA3w0scG9t3s2Q16lYovQWoGO3LyYTST4p0WUeM8WrFPIlBKzrotQMEPe1DW
rJ6Bb4TauLCSrcJYagL0m92VnOHQzAOTLARyxcMk3aALFwf86flYI7bRWqzELXVhnFK0DKI2Ia7a
2OF8LQUnxJd0rh2xX1qVtE2Xx4HKeGWMUlu1h5Du6AIvjNrF1kiJ8MA0M1ii+mtO864cXkA4EYYl
bM1XtLV+HKE/faC35s69Ia+3pDctxqPznRe+DPJ1BZmTp7QiU/nZ4CiNu5sA8YaPB1RX/bjo9R4P
RQlDebKkJc1qPE3pCN2hb3gGgexi5SIYzop451uOOFKbuei1GH3A9S31YZvKgoLpXU0ABVkXT66d
FNaY1iv7K6FvWYsy3h41qWf6jPzgu5NTM+Tcf2VtqITpJ0xkDHqVvQox9gMlpJv6pHECFBdVr7bS
RJoglZmav5TfS4LzrbRHcBL9OjUgG38Ax9GBSWjvjoZxcfqeTaKdeQhjENrR3nXZc5DyvHxA/G69
R739+bagTKUakFpgFRcy/25xCv5l+UAiIahCwYpUZl19M589rNVPqRGm3lIqLmbmEwO+Df5kiaB5
egv8GQeesLsUJqSgjtiKqeSJGMg9kMsGmNfvV7spBkXGAZYYdTfMFNZYYD9ZPS5UmhYIisw0Lh9w
X+XRDXPCc4z0YQ2tw5f9LEuAf9K4DnmE+9wYkm/eY/tWRZziCTkyXA3rcZbEW6ngWXCt21teAWQQ
ByKbQ4GYHBpU/XCnotKM3Yt1z5jWYPURomIrnDydMEUPoKq7AiyL5BMxyrP2waETkrRv/kJDiPHC
/uLjIkxBEntjrjiqtFvCn8FeCSgu9fZ3uerYrazbRFFsK3YpO0BbDunLD/nT3wr9JpnIVvEDFePc
7dvbz3ckHUQdTgZbd1m5crJmuq+Id86hxEHMLiCXE14xwsPpNwVesxQzEF0Khf7EPiFyaxc1a3sp
RsuCWQ29Bjq+KplPX9P57FgClgGrP18rETLVYwOOrkqnAhR8rsAD4DJ3ZXOQHL7edUN3EzW9MTem
iUhQEgX1B3YXGyzgXu/Z/n4j3k2k4VWasLGxeR4y6lNmBS19XhCIMZvh/EAJBebQTfXWJJ05N6Xc
fi3iwJ4M5lXfz7ZZkQliXD+HxzsnwP2mPGhsYLlbPgQNmqUz4HY0rMVRiSymj9gTcKoWaY7IiVnb
YCBMJ0QXIfQCKcM+wbFCPxsaQ2g8JB+UXF9oFmcBkHn3FtU2WX7VXjpnv+X3yx8LHtkNEj1/swoC
m4V6JjLghT7Bj+MkLf5FHmu+lodeMEgq3zkURN6lXsFQTPVAah8fnC3UAhH3JJkEE7kKkhMgVCKp
PyRPOGHDz8hjnnJJ6Ve+5nYWPTMZiKNI4EMIddGFoLOUBcB5CRmNBgj9S7j3FlQBv6EsxEOl100/
b/S2CUs7NZjcOdMyVwDMCpNNrVtBMizNeWjZjSuiRf4NKkBghZVBCVzOiyukdlaUdVELVhNZEAPs
qjhSkO+5ID5nChIAWfJOZCe+zYLjPR/fSHOWcQgD4/p5dlAB7Y26TODsSJJqp5YLa12r7VmsIdQx
Y7bQXhoam5JGrZG/f8F+7Ss5Ar0RFfXgliZJCztABjJuQIGE0pJ6eZaElZylqXtG+CyczH/vchuZ
6r3SRrnkT9Wf4rnStVUS0ha3svsI2sUFRMI3v6pcaUeTH9f5ABuzoV3NTxxJlRMTDMhQOUlOxGJV
7aRlOl1cxOkZAx3Ld0CmTqTYe2ml87TckEYOGcr4f21qtxz7ZR53OVbm6QPwqDE7xTEYWaEUfwBX
op9T6CccuOiqAUkU4YkgruyWXVkKpnpZHna4/kZ+za92njnjRaiz0YQKBLxL8nIzeXctzQJukuX0
j2sU6NY8WvJNQSIfgTCAlPQyPE1vR3Ikrcun6ER5DHMn2uJomHwBFvYYcrfUgYbbYSxIOz113UDJ
WKPK526u/hWR6QyPP1vFBSTqtXkWsB7wt5pNnoP8V4DMSTMHsgb/GbFcGm28j+ydT1TnOZFKpSF5
uPYmZTR6qNHG2cR1c7rgizJ5LK9JwbINjpx8Gd2t3XjETrF4Kmvb2v8FaIZoAW1DPV/AbPDZnaLp
3zfyCdmpNPTW3PBaL+ue+kww6DqNXd6AiexnZo500p+7X73Q90/rqvTchvPD7r7koVWkEOlyHT17
WUDtizUPLrfkuYjxx1E84M3jP6DW9Wsl/pxoXen9g/Wutel7qjbHr0ffU+VjjO2vF13xdziiqWcH
pPP11degrNBJ0t/n0xwonnmrKQlUGUaa4nrjYQuqY9M06M3DwV5dkRkQkO4hCvYSFhiBXBY36EWQ
/DGONKFBQF7NxUMDm8OD0cQvx4p3v3smPfUiSXrJYQO0+kV4DC6d1zEecLp62m3Cj4w3+TGXXzYq
Wx0sxWEIdo3DsGB2XQGiXEypBaPCrxeVKHHM/hMIwjZ9TQBks/1ymoR8C4JLArrEfZFN3+UQYehV
JtvaL4B6FfeOQDiMVGibd1dxF+SyATjB0TVDnW3DmVOV/ioojyFTf9NtOysA+o8PyjGgh+GRBOAW
R/P+z3me+LQ1zjHf4CuX+ehtEbAuwWtNnIGmr2g2qlVFriGFWiKEs2juFVwLQP0tgRGQiFEoLQL2
ogh/5EZ2MeHMzSXtyqPrDEGnIzuXeJw06H92Mghp87gQ8OJW3AVN5vMEqWWrdkM219MTI88yBhcg
PazTtjfhqzIxC214rhfNCG2m/aQvszyOCZeHnjFgYhyvqUm7peH8pWUey9OMwWlTMmgAlaEJvpyr
X08yuD1UNs37GucOtfi4ljOaspycqnKDL/AHE/4Fk9m7+dNosNAdjwmYzaW/GUpq4mnW5dTofl47
qAClJRpniWoaT9cgkO2Zhj2UL0yKyY3gb6sJl/XcpG/sHo7YeqAHFcEwvcqyXfkzZrugggnrVZRq
IWhMlba0aRS8NvI3GZx7cty/lrWWV4aN2hzICTo/ygOHEUPXGH9z/8hi/8z0TBzPDnovsit2f2eY
LjlcvevCSGIHqBgWO5nSf+LebyggSMHjHsLcncfovCA3UTpNyXWTT58w6qcn4KPvfD49zoSYh24l
e0RPcVGQqne+DTQLeYAh4/ZrSZNuXVNlxSWUY/tlLRRJKffZ34TaSXBfpOLV9i57LHYzBgCgr2IK
eoOwK5/B+RjmKucc+m7YdU0QFHZYX5WxHYe2Vb3bTzRMgqSuMDZATskrvRFGRxeMHM/0yM2o5Pbb
ftm5I++UYPhD5msvJ7+1eBRKs+oivEeODRmycJkdeRO4yTwjO8nISekwY5HZVIi06CYT38tRmSN2
DoOj01vvAC0fa1aXW+98zOIlkpiG0PyfPBOWeIDXiv5CkwvGV2FJmdRq5JCN7TlBraWA68Lpa2cg
Kq26fnnK38H6EXo19P3MUiyy62v8Ewk8BY544ZNgRzCjJsbH5hzs1oWm279JUmJ5b8kYaWMlQqwF
/99xQrsTGj2LUs56fRHrDBin1T6SQDfKVdXQok/DRG2Htn0Ersp5bwBlQkJnKrm6KNEq0nJOIe3p
rCuQf66kEi8gQVyXi6Oz5AtpgR8Y+Wdhk5IqkPIbgOo9Sc33A2cM6KNXOW8/wMfOevP64sCjr1ls
QjVrD6heKi+amDabCTfewe9r1ZkzZzkG7TczAe7xUTa/pk2csEEkqfxNhU/rkp1yOcrpw/78uMsR
zNnn9VOVdjVis/z/Mjfi2sTVqTz98d7JHL+5P45q92KBzgheWpjhcZiik+wt9Cj9DK2/Grjn7bGH
ZJh/F9ZM11Xi1WaZDelWc87zAuQyAe4oNmunbUaoMrUElWblFBpabuSLKdUCNQ+WuQTOLQ9fF+Mv
Woe6HMU14RyluvajkcyHXKsf2r4vHgrUA6Q8JKK3fakYSP2QxiqiBVD94i4xPPP9tlerJyandyS0
6wTiWpOINe8M5rbDFtIq0iGPRh6LX/55mThLb63rEvX8v/sl0WXM9p17wrVs2TCU/KgORYY0Axtz
eWjWjC0/XKH+iWutwwscY77MM7HCgcVGCAyCn6vFqqT3UZvDtszHACKfAOwejzRxV2/0eaXJIuT/
2z+3+uokbYrj7eATDkO1S0shBY4MaU/HAuGWNpUzEJ02Qgsd6c3jXV6KV1/moXCmibv0GWiwpYb2
t8xoQltUgHneouwUbuwI5cxv2LVnYf1Yj41dJSRC65uWjt5KiWMWbxclQoU9HqO9TK1X2UPHvzwS
QxXu8JMX+5alwlBv/pML7dkUEV+jDBO0Fr9xfosxRyoeJkKpzNeSMzzQkOSNfdNY1aSK8blotZvd
+dZskhmClfR2qwceMjYS4bMqxoynMirb22CRyQOK/wTSIPzTvrH3k5W/iwY/+yZsxGDpXNAIpZvg
mB9ufaH2PDXrELNpL5/WP+rDtqg4d0cL4Ay+64g6LDQcTgEp1F2pGghjSSk+j3NrSsN9d6ct/k5z
Gg/iwxbhD5RA1zJDmaEwp3Sjg+vSUybUsXqwm2ZL/jCW7gug0roo+WUsS1AlWe1BFSCqEo85Qwcz
X3LCtc3uxS5lQqsbfaxWvJWeHybBJLvPJAIDZxgVHEmtMBxUNACMJbJ9BsGdyb7hwNlkYPjLaG7A
vYz0ESwDavOqtohBAzw8WLc97OhWIpph53N8D+BC7Oi0ny4l+8owKOErcBOqWNzZJT2eOa4wzxH6
0GUXG8V2OgN7ZmLA5IeIUOaV1iL9kcG4dhix2PUAAN5tH3yZHHt5SJXuN0sxyJB8H+rN/kNV5XBO
x1aSc5G8lsB5EtHALbyk4L+UfXsk0Eq8KsfQ3sIXAxloDQPeDbXAJRdVxLJfdAoL7fVjxIMJiAyR
gxTlhdvGWFy+7Jx1c5xXBwj+Yu2g4muGhrt58KDGiPTwEQgAHCsPu+aykCbHxOf+ot/nQ8I5Z8HQ
tJ8hgz7ceyFdYb8jdqTjD0kZXxk6srTOy+lSiS5wXnGZEzqEqyXhqUzFj9qR+0XZIq2s+dFIJW7D
BZ8qQT01NYSTMqQPFVlcilfNE8RSyKSgHA66SBtRtr7mrdguCT5C4NaY3HiCZf+SW6VPXpA404Kr
ZOkjOdFyaJuI0BUDBGMBS7cCJSYtYxgGJ64Y/dlC3K4xIrpZLRxFojqdnd0FZoX/UKHLLYp+/vfe
3EmzCpW0LRpjZo1I3jhXAGgXqAKnL5IO6QKRO5GNVjFf3VcPyuqRRj/cvpv1QDPcayRWgAiehznt
QvZkFyP6CCmMWuWqDNsMAl7TsWr3QE2ECB4N5GYRCAw9VEAvpI8Jus1Zmuc/jTGS4URq3FzrvM1t
zCT8fu/4fFMMkBIgRRyWsIDAFgPr2qI9ODkDSZuHxU/9x9bstJv688K8dKd2GvgqW0aOmA5O2ZHW
2d2kNqq4mDCll02IA1RkW2Pd/ydzLZOHr02H4+yv9CWWSwtn88frntZa1U6wcsxMu/no4OCQtW82
YGWX4HtGIUfvZwP23H6vH1OEwVXp+qdpZbZ8yVjWMfgaF2FR+zX27WYNT5k1ch6ac1NQwCMV2dGO
+I7DSvScpUaJ2YVRpOn0thSrCQAWjwd85n1uU+zayXW+q3iCxOF9PS1HgL2uEvDLR0hiLVvJZcQB
rL7hluLsoWfx8Yr3qQax5jLng1WI0DJ9LMF1hw9eipUNfCiDMIuOfdR0P0mGUZxSkwYrM4WZzD6G
2pcoKScF0H9q+YPwWwYysLF7oXeiQzhwCH/SPNnAoIr3xP5m84WaLR5Zv2zl5UsoVyE6eg2DFbPk
cN+WcMlr7vuxaC6fSCVIAgKNBTuD2ak/xzhLw+Rtp4LYjgVn6QUmIjVlyOY9u6NHWppye/tLuLNW
GXFRJ3x1OY9GTZCgvKmiPyqVwahnLDug4zgzruesGPYTYB5WCzA5Tb8OH3pESVCD5vD/i2q9nJ/Z
QQDPVduwXeCgfkqvDpP0EL1y95Ri5r0KqYinFaPsJvbuxMASos8zbkWZJ9AaSR2bwhhw/rdGxcew
drHjFjyU9zpGLDjEMsuN3Sot/fB+Fa//v+EKQT+TodNZwClJqUVIfCPdrvBmpTSGNR93aw0/GDng
TCdA7qDXkUFB69GiA1BquCU6ZTyncObuqfQYmAHKGEFEn3PKJicG0IaCHQzAqzlHMX7XuToJME3z
I4bqF71J+XGeoZwliHio7G3eG4WxAa9GMiyaVkL+5j/D2XXxzisPxvjWUNXbTqfFIRpQ33hrx0i+
nzGFNlOUYd+pyjmI/akgBEOEWsdhY6uC56Z1ZylFxQJdfvIyGGXR6mm7Dx02DRvyfdVHiTNlPX5+
LK8L++FTQVlVzoq3XCCrsNSqjIMr4V2KNGI5PR2Nvch5xD6D2Sf1PoJdtWLMrrWikzk7XX8OaNMb
KVfvq8h+iAC9xTC/f9py3yAckn7pebd+5y69Nq5povUkSN7qkUUQ44Li6ysR8uIniOCYgVKU2iVX
x7T4bLEylEyWb/AToTEnbW2VP+L/vfXIwBNcijR6QsyD7Cd11X8QQ86jypUVyDskfPF9OnyXYjkh
o2VGKF61Vt/d4ezjDynira/+iDRzrcEod4uDe+s7eCYMAQjUNA0guqK8vze+zzHSmhhe4htITahz
YhA6h63Yfs7UJmzGIXZ7D6Z1LJt/rvbJshT7mdcPP3vJ7hqJoktgdfRRn8lvA2HWO3Gt5P1v+kRs
IxY6Oqp66i1bUxNinRxtr+JrXFTBNwapqJ12TlBXZVBDMEqOiMeuZ53BGrcFKMfLPUlG+OQ7gNPs
YgoLIfPhYnHpG1NK8IWkpOV2xA8W2i3NlbT9tR7S3DblW0ovGoarnTCtT42VB/fhwOdqrkwlwR2r
Ztc2WOfa0LlL65hBg5F4GHOZaZMPM/WUeLSONwl+4w7fqX+sVnmJoipBV5TFHVMV38w0vKCaO7SN
lpcH9TtoBqjhDenK96+uMkiNIyjq0eR6Meza+chB1kzmx9li7+orguZUqKvy5Xl8slz5f5b4vD0V
kk/XiKr3ipK8nMliFHyVlQrd3oHbaMCU3c7lxB0hUYcr02WWGzYOA+mRuuAz32HEG3yKxTEbkxsQ
+j7E23tev/Xpk2nvdMNpbRJbVD+wdBaZWA6gxTqlZ1NLnq9SN/tZWVPiyOYEiaSOzslIjJPie29N
D+6BZKvhjcYDVsRjNG/sQgP1MUD0Km9vsuSJy+FFG8oylzIF5SIIpwz755Um2Oehhnx3Oh0lk4r8
ZR7xhS89TW9x3RvYU2fYH9OHwJGAXQ/dPGuYy2djcDpda4xqb1/N5D3JxEyUVgIl1xEpe/AayLTc
/+ksfRUxVkhvsWl0l36gHGdzYLQNQq3KU+kR3dEb1ELXmixZRMWOFp28T/PQIzcevrbHuWEjt31I
ReKUvo1gt2Vy+uYq9E5pCbJETepVKnx+p/Ap2ymK3VudklYUJV1DWbVhc66Xgfr3EODWPBTaUpTU
zjN3O0Bshz11yaD3xhRFhUd2yxoRsJX+98e+3tDp9jzu2kCdDlV3IPVRUUNq705qokL746qnK0/Y
Do3INkYvK0XgP2zuKhTn/EXaXkp0ewrkrOXFn0UG7WpnDHuwYxwrkABxzM2draua9sHSsKblKwIq
TLjPfugYPgLCe306zxfyPYpp9STOutL+VQ3GPWFj8aewiMCH+dYaRfE6Dc1BsTEJ5LN8D3DeZzo3
NfGNRCyp4L0/YVzOKjSQUSnMQrhaXsknpo+a9M7hmjyKDZGPs+UzByf3AUFuj9AvoP5dIbGXQH/P
lIDjfgxIlHPX9riTOAHVMg8pYPEwh6W1eDS17A/+nrLvHBg/ceXMHGBmVobMxKCn6mp3j1w1rDB5
LQlBARQr0RxL/3j3P4hdsBcKh5lQRbmeSlc3vc1o8fpj/E8zcVt76ijAuTiCKXDfF0ZOnSbHO9fJ
62Cc3thmIDmjAlM/UVfy49RYwxyw/xCi03LdQoR4L/JuGGwG9M3QmHy9tJ9IvMlVGvVxzDoqP3Mb
VIfmwTEkIJNst5mQbapYF8OsJsVpd721DkSWcO2ldfA6DRy6di0GT2XQ8ds15X2Qi0Ue3ppbUEJU
8dOAFwvBHI2oPAWB9q0+y3n6c8ZvvTij5EJCYOep+zN7tnhW4Swnud9Hb0w0KNBS+oOBKjK3lWGp
6KAebF+f5B0WNcE2SCU4jpu3E9hNa7HPn8W3fEVBrtMcLK8uu5PeA49a4PkQBd9sVwI4dEv5wFpb
CMk0LrCiw9pNhumTtqKeWOCpXY+mJK9JfdKXHAhrnjsfU2/wa6jyDrl84ODtaLEAy1jTazSeD9gd
vpBmrGXqhD9clp/ynfbh08lVvnbGGuUFSeamOW+lSXJmLCCswjAPtIa9/yiO95NPgTGUlSJAmR4J
yXHJeWmUaev4puzj6lG5o/Zwr/E3OHbwegcqqsUKULDjlExo1ycPWjMryrkc8YNDpBDhJA6jFI/T
rhsyd3PVzddd5Yqbr14vE6/3WVgKSPZXDhXx9uRH/MYoxlGdT/anFtTTSNOKxS6p6604M6BQCafl
T6KviQEGgO5BrDK0X/ZBqkoL1YkbvsFKU1YA47f+axb2bYSkB1ZWZMhJLep8PVBms1/0M1ooQv+E
MbJGpaM8qcU4EM+UJQTGipFZtkYD49c0u4Q3mOPCuZxOTZYW5zEEajxLwC5Gk/PsVvG57BZWNj9y
Zdx//J/aSoBnldTM12IPPxE6DrYWUiG8aHO/u5n2B8JGSeUWdIJR3qjzCWX66AjK5OdNPXxQ0qZD
oJKs2PEbEILO3YdCHJ1KdcvFnISls85eJvDc0JAnHanLEnIw63TR6Urh4jZkRtkvwUq1/7Ndo0M7
Tah7Vv60ZW8Pz8/RYYQ6iv3ZJGcRpTuPbJxFPqq6AEFA2j5+AyESo1amYk5YksOhKAx7YAGJycsB
thG59qJh5AyV8ny6U38dQd36iIXkBlmw4TvQqtFGrZMRf3yi99zEiYQXADjIwla6qcAMBufC09kt
ZL7lwgKZ8s9phSJswtsOMXGbgsn7lDbMjWBgeaSMX8qLmJU/p3fQfVw9SzQpMzDOWFxn3llfcKnU
Dyj3cJRZXspzBD6gbBPePSgcjAh/fuWscjE5PPDNf0giC3hG+Uk6jpyZs4gYS6WHSeBd0QDzvngP
ZcBwosJX+9PQM2fDN3Bvfiica1uFSmkoMAwDneItn1LrPbA1A9wz6br2d+5IDPCOxkRWCcKF4Ka/
zff63N9rfGGt36Mg4LcdVZ7rPmBd3VP12qGpmvaOQqOHW/Wbjx0zAafFgqy2/+nUqbgPHdAL298J
5czx1rBWjsIQ/xSuren4FXC0AubfxpP8loQaSsKdopDJxHh2rlhBkGwzn0plACLw8Ep60sjoOpHf
1kMu/S6of7X+QBpYpqcqyCkavAR61R6i/SGzLoFUjwJgY/wnhNH8gx2SXVRGLDb21a+PI4M+hYHW
aPyOSUNCn2IMEGNkJcJeIG+/feBOsfR3qWhJNUgEEB0fxc/w3PMjuBuRwuqLZSLQERV1RU8fiHnk
6Y6xeb4Tl72FfKXBQsdmzEIBkb5+2Os9KR56JNx8dll6gVe8gp2Rurax9Uzm6aK1MoI3oAc+Kza+
2EMskcT8UXUvWOFC1JMTJcU1FhOWxfuhXpVYlAZR8x43oWKFZwYYjdh/8Ya8xinKxCocXprOjmPg
slWD+U2TC2M4Gf+0WT9FZcpngG+/NLhgAVAnZdwKCBHiEIQpEc+jKZYk/gPuCIoJZl/RG+0IdmC+
9HVv4nt2X2OXMwzlw/PgppxsEu+TiXgLYVBUx3rqclG2mg/grj3bHoYXWdxGFdg+o+bWcBahtYlG
28iUYilUlHv47kGVvizWQ7j4s/CzaN/PcIrztzdJ7fpjtYDN56FrsRR81+QG2Ei9KhhWf0epwYon
u8MKCK4qIFoG9qF9LztYMZ5URbnIrrucTog9yk/Dz977PNGj1vwiUiAE40balSqIcY6DtFaSmuSY
ndGZqdI+lcIePTQ16j0i08jQYSgML/TPasFzC3qyrMOUICQ9IVasDnbgQ1WxZCR0MbGWDKG0SyPZ
CMt+UqF7gzBTv5VZPzjie6lFjC3oO0YNW19jAsygQx1MfHRiA2R7lS2eBC7+k6yVG+Byh3VkwU0p
YDhc8mEhqQUU5B0KTt2Z47Y80yScqg3oaRkXkueYlb9aGh+BPpTlzooEGTRk0AtAAQIZa/vCT2uU
LeTe/xzUSIKka2Gh4tXdajI+WMBYBzx6Khnma2HauqRjiQXTR61T9PKgCs+2RV9zQ919Romncg5a
QO9r/XOGgQ1sfOmX76nSSsT89GHTH7FUzDnw5AX2uyRW3dxk9mLr9nA8uHgNMORFYcDzaNw92gpx
yXVbhXrCvV1C9o7aiUASn9qlfC02F35ScAnATqMRvhyEi6iGj4RRyfy8K0ejHZGQ6Vqd3WFUqAb8
56zbK86eaZg3L2K75bRWX9F3BtWeVILaS3x8TzGkX/WgdfjuohiJ6b50viWSEbSmn9L1+gQH2LER
2aLrfi9elT2JfhV7djgTbapvB/XK77utyhlY/pV3MSvwlfpCh8W4dsro7Hriwr42Nuw1Bt70tk/N
+a+yLL+xiqIGMdlVLekhBTM08Vo3ybFJDS2f3sDPVGAehsdSpvqwxm3Y0FjPjSbHxH4GJOqMZr9k
VD3lPmdLS4DZ83s7TUPf/7l/jyCLfA7cYSAzaZFy3bhsrTJjaIfrbLJ8Pa92phht0LjmKIWarQDY
bLuB59LkmVBvLZyGyWIcpk9P7VLwFfcD4JLUa9ev2Rz5FZ8amaOFrpnElh4I3ge6XX4z3ZREzPkV
IMJx59MHCs+3yHuIUL3zNvNbXFZgKkfbUFGfLmNC/9ejINd95YiGVsVQly1uoajQfP4gCrh/Vt1y
R2zHUB+0ekd4UEgkyFaHEzmEuxtuKglroBLMi7EXMPzb1qtZIpXlTEEawBnOjfFPqXKnFlfg7tG0
nvjEv34QTBcMwzMwMyc2ou/tMLjLy+ZeGGaxld2nl4d5i4U+NRKf/7BnPJ87KxRLk5E9lWungquk
3C5VYew8Sk0GPXwesOYhVrg09e846g0Ff7uRQbUF5diCHTuiaTL5HJGsj4JrNJVDSv2ZnMfKD2P5
AYW/P7siX19PLTJD+iKb5nfl/CUUZOuLykBtxH0kEy2FpmsYIED1HDopm5l0ptna5x4C+yMLIEOr
hIWFmPZdlmkCUlglelLRgeoxjvIXb6hfdoN0XDUyXb4EpV77OgnJacwSQ7HAfTuxt6uNcQLtcr/1
7vbxxZZr+g6cO2ZwQr0+PBfsYqJF5rw/LVvEkqV2s+kdTv32Doxp8pgFOoYktt7+vsHDi9fkhoeD
Rd0KSybYCtm6qq19VRY9VbcudK8MyeFhvHoThN/habTNzVuOnefvFalwJNWQmAUViwVTzxHEC+Z+
f6q2sM7RH7bQD7ew82aA8olLRE0Ios5JuumlEJ1XMMBThKiOngAPoDdonA8uzbfEJ5+tDkuSFNNl
GLhi9H0nSpLCUHksYbIuHvIJQqiT5Ch653IkbmSobIjumvwamnN8AgYuirLrnAqxm02sx2WZrL/4
gtf12lNJGgwq9lD9fNB0E+O8a6UzBAt8bRdFV+13YRZ5e2NluQ3g7MRRDCifcdjGABrQWquO2GQG
20TQcSM9I/RMxswkammLztjh6JaiPrR1Z9IElOfEB4nhZ1gYHjDhUmWTWhwDjzQh7psSDqbb0/Tw
jrkVUDbSeY8YDjcLZXJSB3+OGlprnTyv/igcf0uFhiJSWgrzvc52WpOGICKmeAWmXQ1hgJTwBsLt
FMRnoPQxCWJlyv3eGlqRug5scYOM9aZ2v2FbjZ7fK2c6vo+NP8mz358cVXvvI8g1Z2ycOFaVHTWN
B5jMgG3fG/QIr07NitpEnYw0sDTkq4f2+zZThMIG3JLs1avhYfzuRM3ABdfmdbm8RWsKUtkp8oPv
LaBuYWq+BFy7+17AVOjD1ozxQlWp2i3vgQ/c/A9OI2Nr9sD7ARKo6VGAkbfwCCbiETYSSD5GUm/d
lwfOajNNBA9dG8lblkFA0HYS/HgyZHwMHF/RZJp9I5boLP+j+R+YLD+GhLO553BDnfy/T6GGpO+m
vhKOqWsQZRULCQ46Sns6RPU25kedA5sQAmJvFtUd6TGOTJ2beJe0ylhkx5iAS8m5C5da1Kj8bLSZ
ol9fBTdWGgbqyQsxBBAM94EJdRI8Dt1L3z2cR8YN1fxm2WU1d5nUz3/1XSwmFkb0xVx8Z1GYvNT+
2sFCQa4ktVoNcAWgGuG5PO4u+OC8FhDbAnkGF6wZdFNSRF5JGaJPpF8GnM6WMaDFjwwjLHwMeDYn
0FnJDWdb6szn4Jq1hl9LYmnewpx6n/5PyzDTYIOTpiJAl6LXQbaDo7xLBUmxXdRFVzBFCM7f4Y+O
62NbcARuyZLL2S7+vxQKVrvb+D2msX7MNU2/3NQH+3Zvgefb1KO6yc5ANYoVRDNrYdDThq+or+m6
fKcj7JQ/vZXUTQ0lipsGEH+29EJFcksCLX+rTsN2hjWnoa8vO3n8NcB6v4aRmS9XJzsF7rAF/Nsu
fVZsi9TXZQB/MtQ0r9eJze1fHQHYeVo1iRA0n3OKdWMxudR8rcwRmKfsfglI1XimatDEd8Vj6BLg
dg7vQdSCp1JrrRDndJUnYU5mgtaD4i48DCvJaBJq0L6Q4cZD2Vislp1H4WPQc7M4MW3I/P/BtCY1
sjqPjMd7Cb6Qrr+dGnpm1EhFcynsegk6fcbSsbR4wVSx9YHodvlyWiaN+aglCOdYZNNbugfwiD2S
M058hsL5iIgedadtwXTjM7XLVwTYyB9nKV9mam7vwBEwrBuipE6f9/P35BjCALUcZsdzQcBzzQpU
0D7sgGdiizFL43vxV2I2plyHxtK2RzHIdkxx/8NSu14XEdADFe4RVPMzu1afGtonP8C+0zL9vy1a
ItdzhvYMrw4OR0dS7qmk1A9adGE3B6O+SQc5c5k3+8SkRbO/B/wMQWov5IJwbrgZgkdcaSQEasGR
p0k6xcOpTZvhL1uAwdJ0JLkwGNK2cl1c48+dmdHLLw4ARI0uXxXUm8BEkXF+kmMTSi/b7IOz9RxQ
CEndmpg33Wo0203Uip0G5c8AJD68FRtyEBCbLFpqlHTaZStGdcK8+NgSDxF2iAYCJZ8ebZzzulDQ
zsyHYS9br/SUxkcb+7tjVYq5HVncxZyvTmztGAVkZ6v+l92/HknnoAVIhT+0uKCl108ZHe6LhZ1T
8ZmtcWOhX0xIn+AdyhfeNtFVkwOQhOrpA72sOQuti7VO8tkVr8bA5zFOCLpr59h3l41zHvVHtElU
WyJIWGbMktHWGlqcUuTCODji7g8G77TwAUwk8CW/mNtsNeCwrK3sLhI7Fy4HBtdJ+z4QOGpYSbBd
wFEP7mLIDCOCU+3UxjWOOna2Ot+r32pKFyny78q/vgCH8EGpyP0D5ERp3Dil/lgYwi+2KXeTXXot
2Hh10tOisHx3c/tljdR7izOOmPKEjo+DIrkKpy8H65+p1lwraQtg4z7NViRBLBoEpzda+i2wzKtN
LExcZ39c1JcrYf85eAnUJ5t+YSs1DmLFhfj/nnnF8qoURmjJvvqJID2ouzye5M7S2eiVBQSgFZSC
RGej3dxEP46XL+STwpbxKPrk0OguivsLQkjzyC8n96zeRgSWB9Tv9TONP5ytf/rnnNkPmmM29nVu
1Si3bAdfpbnYlXrs4UuurHHJvwP04q7QnQu6m3XuTFHeTrqgRDdieUEUqX6wQy8MsXRUs++u6Nsa
cSIjffnGJ4Dre62q1p9zyDIiMYkTxYiL9PvAgF7jOJ27H8Rabg4QPUX16Wj81z4uoFVqvIffj9Fu
LPVQFHib2A1ist8j8HorHJ3+oyS4kKw7JYZSR38jEk3rDCp6yo+rSZpsyEcaemGYRuttygXmnq4B
MFKmKgEdkHcmdR/mRVfQOuP4yt3BFVuHo7XVmnpl1aH0AVwtJHSppp37lIQHynO8GfFi8SS/ODZ/
gJ0+6h13nPugJOLtFXZVuFM6u76ox1R4+tOK+E9zFeYk445Nhtw8pMRk8yCraW6hng4rPPaAEMM+
cgm97G3+IrPnwKGiPkigI7CaCUC+DC3uPjSfI28qMsWwoknzcD7V1OhtST4eUNOkeYR85t8/E7WM
ooNxC16Gv0q2eF5n/4PVRz2iUIfRaHTncRYW/9ysl33TvCC/anIr6hDDz+zWVV9oT8LaUwYSGLqQ
BqQe9L/6ReZfl5+AG/iTWfIBopzv4Ou+jLDQzodSCp8ICrgYlZXvyYqta1VrOipDKY18V3dybxK6
WUxUVn7q4Sh64HslXi2PJUolKqK9ifXnJ7IoUYtCtpX3o3WQYC/7/NTHHfG2OtxVAp2hGIUMbP0V
wxPsCzDYjm27T1qO6iFPJIX5Dv2I7Oe/UNTaMwZJqiIQspQbNoovXvQ76e/8GKf6WpesRVQmFAP8
HeyS9dOfATe5gobSE0Inw5ufL2sADosR3HWajYVsllSLjviugLXOG7aWe1KsZtMRnoJqH1AecPRF
NsAh39lkpnBkN6VoAuF6Jv/nnzcu1z+pAzHO179Dmb5V/S2EsuEUGck6GPi2d7LFBzVBu5Vrt0Ih
PdJSpE5opiW8Tybecv71xW9CeFd1kO3QUXEIAdwJzyFV/eZmF4Xt5Kfw1AP7DP4ZJ9NxUFeyr5+k
zKxF0WRXMzLinBB7zLbgXPuNLeHK1oVx4uY9ucsFPWl7AQRsHGurpeidMCKEPGlYDg1nMU2CgtI3
ANaG3+kgcTNtO+UIYJA+TzrBjTSsSS2qkd25jfn38FgYs45hlMquE6lxa7sf5Xl956C0mT5YaF8j
gmy9GA0+PJ2HBipNHb4J536hVFwA9wmqQi+BZ9nIt283RgehOwulhOujXndQKXFkyEFc1Dst1BJl
uohDb8VNoCdP+jXXeTlNRpjGtMgEBFcJ/piQCOtwzZtjhGXp1JRzlCSTH5VQmpYu1AgBb+RCdAbD
SoSPzIUnky0zCzQwoCIBRc4X9iWu/9uShEL4VdhtVripVkSVdykmhHFwfxh0czTGXAXXtEooUErx
XH80btGgAVb4AjOEeNaaxR4RJR6j9uM5luKThvJpTMX2Q5XuxtmD7XxEdfYE8/psgE9cpQduRmgH
6o5eTpFk8DODZAvrjKVuzWgwFc2Twr7mrP4pPlF2xXs7U63SCpQGp+DriDSKhBNTUjCFK+2o76K9
AK7Brb51gXESuTyqBxnG5Tj9g05vzHBDYEzdtyaBUfkMa6MH2KASl1K6/gSgkaSXyq6gvWErmIxo
RWmdXJtiyMecnSbHIzBdQNplVs4AerndY9Qr/V+BOypF3AQHIhFafA/AxpsMa6Mp8y22EAKyH7C+
so7Tzokh3ttpiT9Lb85yJEZv2ajpuAPPWzEDRwHOf6F2pVMSR4TL5lofjcQtytYcqyBGVCMxGUAn
tXHf6Nxbdm4HJ3aaK6HOoL2wQUcppUrI4SoiYM6JqfyZNVnK1Lk8BFyl6P30nv7xbM3WurvnZN0K
af9qr1ypiTMWUEypWtoO53f2jTT2dKiqNX5vQtVrLVwBihFu6v+lx8WJl0AtgMRa/Bj4BS/yEhPQ
x6v10+OGmHny8sj4WbO7DDR9VWBDVF4RXM5Y/3wvPD3PCJ3fkJ8RDXzHfXWT+ULjZlJnD/WuwEqt
W0+iJERyyJsk4OKhXyU2Fpsjj8HbU/3heQTUr0Sf5I51uSQjpST6qFKl81E+40BlSL+a4RydcKlg
WkMYB5kREatzOAqE6Gu2IFEsJS6+1qJB3nOKbVdQI9FEw8gcrUfM6eM4qd7I4D4NmELTFHJmikhB
3eg16q9IcWmPv+I9pB7bRkZxEErzP4dydKSo8B9IJxigMe35KV8vwOW4PeSmc9HwzgYzge2mB/yn
uH88ecMiermk1M1p/5PjFTe7y9YwZVq5XEE4p5jrSpsckdDKkYbLLM0rSYHHFa6wIzkLb4aStYmA
jjLB/Bn0JDXQojhylDVVbpa6ItEe8qw4+T/cE0FJDPzhGUd5Jf8nB6UzNTuv+vHMrFRtWBeKUdqU
7WKs+v8BGiTh3SoIrW7ydaPC1/vX0LKi/M0gYpiyFNX4jeWhv5oj9Fnr6RyJubrCP5SuH7Z8FfOr
ECP+YtPeGst/01p0aQ1eJW5WhQNdsEozQrbAInVc37ByZISWMmdO36vstmhxtjttROb19bgqnQSu
UAGWWNCwdc6fHnHTMNgr2zT4J7r4in++ueUWMQtCbkEl6040KBNVCntYjoO06Yqh05wLsK5L7BUh
Op+c9ZkervHVex8yEbnj7VgC63+jPI/EZWrHhFWvrW9gX/4Y0gBTK8WIQuNt31saVcYRZYRLKsWG
nNcxG5zGNqUu8wV0506ePN9SUTUi3qaNGe8yMsQI8h51pwPMtn2cvoPgKfHEZLYxcf8xnwHwToIj
Cq1aDhd6XAieKTWECqAb1GphhicK1hbTfOFK6Kq8KhaADRDEJju0zc8cwoFlDxwjfl+8Z4AHoFuf
HzNUB7KyIjxTB3kxxg9Rg2mzkOaQR2lj64PRTF3iDt2RFPIOjpTrO5B8TH2X5mh9inwh62nDzyif
A3dI5dJn2FENGYWf8tJfuJbccXbrcFAtEfvQPd+5HJJiVAe3JYfkZfUXslHGB4bR3KRY2n9Cev33
iG3klQ17xVkdRQIQ4hD5SEmHaRBIBWmZMH28YAwt4sQlOGsAlGGUk65BVh7NRuNNGRmCzqoXb7f5
SWfixEPkd8/5Kj9FSOnlQuPyfTaAvpoFxllsn79Jdjcguls4ucQo1F/ap7UEAnYnfpYcf01FqM5b
bfjSAal4kN9Ja8zjWMqG8/JtQ7i8BQW5Vitr7ZeOwXxQUroFNjt/uVEBD3ojiRkLA4qki8YDx1Bd
1DnxQVvwNqFX069yIKwxeHecDJzjs62D/sxKFKYDI+F/iPIdrGwaR1h1UDGEngao7AI5cA+OCJUl
tYQklvrusgQJxqFa5qZqAR0uvkXaznImNmW9ouwqYuPRWDZb1XPGNwcdDuAe6+Cd12OQdplbbWTQ
vSlpN30jx3FU+klfPmJb2o0nJD2B8CfOdr7kFrmjVoFJdbkQBfFMgipmlXlxX4isFbo+eed7boJt
qbQj3d7Dwzpsu6WgPOJ5p1G8BEwrj+Eq15DRpF1mZWgYnbcxfxyZiGcPlrrIbAbV62F3TGX0RAm4
p0WMmzI5UoFHC2uN0KwolVDoZ+rVKGFKhSTc+lfaHdO7wMqprmSVhlm00HSjBjLRVbXd7uKMD9b/
F0HfOHuFa9R/pkF5n0nvhnmPdZYJgwpZr6Vj2yMClX9OfoKUeEigtNqhSQ84go2+6iaO1BmAXejm
NUO6zbDLbsovewn0qETWulJyvoy7iypfsL1qr13Gxy10on7jIgpTduAXY4f0TKs1T5ePNs0uqlcK
UT4B8T7o0SwgfqL0Fc3sEbyrZqzaeC9fCbkcmpQwoQbw5854tB0N+v7PD6zTM4os1gG8n7QjP7ws
8O6QxiXBRipXs8uchX8DMQZCHg/lxSz2oSGJaEgKVUTaq4KkTSRinp5MrUYIz60OERwUglV1IZgw
bEuzSgLY9doQx1E1YR5tL1PFB84EJuIEx0W7qJ3aSZEhweFwBy68bj0KcuK5eg6tOtQwVHtqrB4r
PxNVxLdi6eCl3x3/kqeT8Jb1WyrxjwRduTfOcuUsEHFt1QxX52xjzA7XjsfKUNgZciHejNL3VO2O
L1Q/dzwqjdC++Rvk0puXR3+Q45xwxtX49EgNJHWArMymALi0SqbDTDClVOWX0E0UPOkXcA1J1QfV
xyEWUi0bJa4lmZrmCzSnzbwYT6aH1fnV/8Msho9bCeZ7n83pzPwDRhUXZkMQUSvk7eYIJZcuI+sC
R79Vn6O6l463N1fkbb+tQFhtjb4bLjnE2P1FntB0UqzuG6DfGCbmCXqC80mdbUIqUpjLoHj+O7lC
16R+k5DWik7yDchlpafslNbRPQ0E9pPGUen8+lCgcy2XrLPnZMDyK1Lbuk8WpZTiqe+vHVBfIlU8
wjBeaxHLlTkIRGbP980FhbrsUN92QbfvoUYwJcifoiDmBbLOdSIJpC+iMfEaYSnRezXKpUkK5MkS
99ABLIqLx/NNlWsNNZoxJVlYJWft7Uxrvnvuaswm/vEfyHMOOHyQukXmGdzXbgGZfHTf8LV4WHq2
eBQ8WLq2RTsL2k9ahaP1/5iWqOA0UKkxl5wYTAhCmD+1/Dblj4nAPbiX3boLMcT2S8wS4oLiESU6
fu2Y0cisa/nZ3Yu2njUsUokSXg6O6NI/beAh9cb1PpfRR15+81e2vTyAJINNTDYs2mghLdT4bP5Z
xxhKDys1d+sL/fBNW4IeKSEsf9gI0EzsiZUjopHk+rTh0pyPy0HXBsjna6krgcS0MvSLE9dt2ui1
/StBMwINXVYLLhFpBnHsTuiaW0dJ+yjSBaZNQLv93VyFnA71HZ6EPFANLtwhLPLUbGH+JQ24yQbn
bjcwVuB4yQ5lyimTD86PM68bpkNCxmX5Drx/7CokZ41AHO1YzyJgEGzVrlSvX6etjBOyxkwtIiou
LjPFG6zgeyActseAFL2INJqDnuws+3hpO1pqp5u5WAImp6gGJA8aQM9meidMlIp5Jv4zoN/St5ZV
htpi/nmTAiNwXRAhV1+pNGlXl+i57CEb4H6XN15EMs2omvcuKtndaPGGXwO+BjaTLJJNJGUPXsJ3
xacVZYVIr/09cZSJUkXc54XCV97U44wxxq7nQFXPF10ag2sWOYz7RJ/fSTPVX2qIdbs03u0Ybque
zUDa4HqyU/ko/YJ+r0C+DG5hkrvYuVg4LjcYnHnv00dUJRjwZzmdjCNxY/beWZjxMnFhdZkixfCG
iIE4NR9bJokZHHYf6GUQT6dInideHu416K/3PrTSKFmWSlAUUAGYsfkLTlXuBaT9y44uPcRWA2ov
Spn8gJd7DqyWhj+ZS9UeKNDScMvE/wwqpKeaaUrz8alq+TSlV/dafGOWjKCk31yq1gb8OhZhpKRy
Eq4mZji/jqq3Mm+R0Yu8RLQLX1z3ZlzehNMEgXJ2RmAr0LlQAE9QL+yy8rIza38En86Mfoow6R7I
f251DtE2BINXCNysdbo5PuiNqPd1oQE2oGDVQhQFjek9zUtxnFxoheqDwXhc4Mco9RqW9vJkYJnA
ixpOEBvs5qtOLE+Ksz0orquIPBER9pKqvrUAYHVIgmc/Gt4SB4uqaHPQRddylVbF2tXVR9xsZRzs
hbJZrpkN5gkXseLt8xzO5Gj5n40PSnG2y43cnxSo0drrAk9X93UQ9SXmdZPQueNV6AWlbJn36ZI9
Wo0FvmnIUdh0NopHG/rhM7t36YeQiXKphkYaUGoKZwl2yw+U8akul9wiGLo80LDsvwzqfychn12X
IS5gA/uNZEcwIX5YntmfH9UAoCAOajrlvc9pjjtHddE0bxfCX7kNxR1wPF9+DaLr5z1sNU8EGn0I
sdM5dqm7JmBNBjUU60kVk6kCV/skqV+fcG5a+jNFt7COLd3setx1L8o6TnsXgyFPxZ0fpkiOomgM
mqWI+w1MVRG6f0q2cQMrAAxqzgTaduEKGUelWakT5wVA/PLkX2hgg9Dnxx58sjainYHwLDcJnusG
gbqo8XFhg4EVZlCmnRaLNQwZwxpA29Lq+tgf7seyflyYRpfS1uodE2NdhDms2LJoyAVlCqB+yZo4
ZlUMR3K5UQjc3XWqXukvnKeI6D9CLlB8Hl2S14TL/D1GtlgU/IjUQPMmuo7neXnD/8WmHMKiFBC5
VLgBNkaF0KkYHFivtTWsSoOFXlh0dNGJilyoMR6tn3LVgUNhVLcjpOgqp4tN+Jpt2tK2HMSehQAl
VoA37OXJGcvuy8Gq4ITP+4i9DE6fbhQ4JXYE1L1MQo9YKib5/ki/qZrLShIajmGdZ1OrfqDUh1BK
2rj4iWMEJzZot7IEcte+TeQof0At21Q9oqiuwAGhCedaaBxrA54FSGpi3jTjrUgRQTe9y4o0Evds
RFKz6gNTMiQaKdl9o8aKQLVYo7SROEapOdLMqW2OJ41qNgySy38dihH4oTUZwvCAaXrnSEf3UNnp
BrhHc7jx0RYyNJSfp98Xan5TvXmibmKDKtUTiCxF/xKBr6S/Ma39jxw1Hm7WuQOjFHa/zxPoxiqs
YI+w1x8vJGVDqKuuycLl/k4jDWL9WemshuDzaRe9Ro65U/2bXw3JdemUrIOaaeY+p09KA8eOoUgB
XG6C6I/JcJTJ+LacQ2BgFs5BzQcXUOaXS4v2YOKpxC82UQr6ru3inE4AFekiQCHYZM1ULHJIUpOU
jqapc4LGsaV0WyHh/4FijpZOQqjxTcygFew2bq09E7Tus8Q0CgtCz26Rxylc6MIE+1N4Jpc3pdvU
yd+dAbtSisiAAYO0VVNygT6chIQc2ksf1+AE447AHVIY1WpVzutNgkH1Elczty8p3xK5i38PObr+
yv+VRKRXfxWTNzi9exoG0WnQ1ajJzxRMtRuWtrpRil5ly4THUmoluDfNHNdkeP51GffQ84Nu/BjS
6dlSoZK5620LH08St9Jj8m4ZhsivWfOxSIpXt193EU9Xh1ntLUlxQFEXOWxkK3rumqOoEb3I4hbR
vuNPbKrsw0Y68hOGMMdIQEdikV4v9smdAiSVRorJ3vxvtKouQLINNVQ2V9H5gQqe95YNTQMpzjiP
3d5PDTJDKWoL7iiKgl0Vz5YMfoR3vbMxNHOqFl5FrbmzLpOkII7+CiGTyX355hLLVTeYwink9VSN
Rk8rkYGJIY8iOHld0Jv/OsHK/9Vqx+4NauCHhHgX0QbYih+eK5J1Dx+/EJs7IVx/LXx4wLxdx8LU
m+PVJXNGq21hMVHhwesKuhW+L6JDp13JUmBp5R59tSsLJtB+UWupRQXoJrIMRklIBvmt7sF1azLR
DBLiZTEoFzh+i7ReDJr41j4chT7PjXLLgUCEtFD7Sgv1qU+MFPk9uDyzA3bWSbDWfKAgAc/2gsJm
s1zZWh31t7FfuWKb3x+YhkBXKobz6yfuFMrE2ONRSnJNDAmFR6EcPWMzbiCyFF42uNxFMygESKJE
hkMMvqhuVk7Ow1RsEj5IEd6DawgItpYpzcHuh5EbpgN0PlfaGzNzTHbLgpuGNwEo4Vy/ganL5CSm
RzdRGeNs8sIyyK/wpMwQhcYMFEklZVtmxEdAucFWKcRQ0agxUDEhBAAkioh8OLWSXoXyMu/GLTEZ
TnpAE32OW6YU5D1hsqwZumTIF1YXEKqyN+eZkg61KLSGP4u3RDQ+HQg64MTngca2Wb8uQ5j0H/jo
LMTycJObP9NBC2z5nZj6px5OOfVEoWC96f09mpJG8GQTJVRsyCjAhoXBC20k4fbfVDWd1Y+koHgl
mz7if1tvflHaPng69/ZzT6cjkP1qvWTHkhL+AUCXVkxVfDd1L/cBO2ChbrzY//9+rCcAJ7tnnyxw
A5NrWVO07WQtIJwI7zIz/pcb/f+MK9ERb6MQU7MUBFTtmXozOjq1pKrFivsKS8gx6u4U+6P1zqv7
7MSQXLl5i1iFsk3XYJcUSp38NBPvkojG8N1a/AEOAOktbKVtPwhbvSv4votyj5QYdx+zwSE20m6/
Q3XNNWvz5yWYUXCTW3tnupFPWunGRq2VhJt/koedOYQdTrK6oYMtWWngOJz3AOgYJ8uqGNY8q/f0
UK0YYs4urDCb2fLit9nfvczkPb5Oc2lNBG/OIJdRtiDS3GHcdcIhA5Umzr4REBUyxhYNEoKPWHDS
//lAEIaifkEonmSUnF9cuABxZSljeoQNrc2jWLQJQi0rnuUKVsTZZ1kWod4OWlG+/HdNiwVhn8C1
zT5FyzeUzoCLLbymaPtly7MXMlWIUmfKRznnDQn/095TpjHIe3DzJUI6mco7uhetDmXSw1+oGuul
KxX9BK6qqeXH1l2n9FwYVBFv3YmTKPAT5SE1sHQvErE09mLg35KPioPc/9Ktlq91c/QaSzNBoIej
ghNCH0ChdQSsEUDwXiqd7gRC9AaT2M/MDGR5Hw4y/Ui94B5AOqNO1cVE70n7iXZRRv5995DDTRY3
+2Z0/+quQYt/AXpKKMNjJy9dh6dnXRRoA7kbUygcnc9vk1OMdAxyTG8DRAd+bIPuzALGOgxu4m3d
aDkIYME7joRYMn2Dc6V+GI2R9HUYq0Ad8XLEzGscW57fQTGVaYgoWkpaukfXPA80Rmdxl2uKbgr2
H2CyIoJ1zKQqV6Hn0N/kRasSdkY09rZ40oJGC6oL+RaA34lezsdtBJjQ1YQ3QrZH2v7avkjzJWSG
NXwi9CSZ9ReGi735QFwIhOUnznCPcXw18Hs3RJ3lu+sOQ8JCW58fcNi/Uf87qKb0f7SjwcmuXNi0
mxstJmO+ORV7A9qCmAiY/9+d5n60NLfwkb86j3KDDprOamK1Tkwf04PThAAqsnd01EMcVhTUL0rL
FRYxggGWaiTDoRU/9uT3xDmOtesjidUKh3oM+tQpun8d/yyWBSCIJk+MxI9HgwMEsaiD4yLjer/X
AuDIgSpNWACc3YBgNf9g+hj8JlAmCLWRNrt0PQHh5TSIbRcGUfT+x0RpC5bdcEyhmkxcEcNnVOWd
mPXP3szinN2QrniCjnxDj3ExqjJUksgW4VTJihV7H82IHRkofvB2C59j1CU1JoEWk2IYbyPxRQY8
PXq8cOJsP9DBBYlvjre/N3jhcB67etLHjdiD1xrW8hXQ9/Dz/TvgSn+dwyP4SzonOevt288ogEcg
UH+KVbpC/VQLR7kLCy/N+LPQ5/59J/Age/2HAHOQcv5OsXKwGa7bekNa87N7iMUxq63DU1GGNTfF
Gf3hM0NdFYzmFPodEryHi4Eaqw6C5YZyENKYP8k0ovKUDVQr77Q+h/IRMCbK9ghGOnpG5arthlOt
t8rBlMuu6SEUd10ADoEC3/Rd1VdfQ1XFEGOmxNskWj+oeo0C7glq+6F/VKARwJmBG+z1u/5NtM8d
95WEcJ0bS+pzqBchgB7TLzBX6ub00EG6dePYdooKtvHhT6Q5IcyzCkshIk5NvbOyzsnlmU8I8nd9
nU2R307aGOcP9QlFuPrC4Ku/VEU4pimknQU4+eSUH892F1sLKq1nCxCDyHlslV3DohXz3oPDvHen
n2OLyLidoyWpkGwOikm/pqnHSMYx+F6mktszAZd/8rr+RZ2z6IaHXfxk7DpIXo2uSJF1LwKJ5r4k
V2h/oc4xWHWb/+cSWNl85AZtugrMljJQ1GkDo6Dn+C71T9G3vMVbqqivJE9ysGHzp6LSlqtpMf9h
yq2UVJQ5fVG4uaziyJ6ebMwChd43UN/z4Dod4CBQn6vbdzs+Vd+Ct4eUygkppwP+Ev95DaG2ZP0U
WJzLkjYZ9A+z5sJ37AmHDgnz5IEHQqThQluRmagsJEqHbUNL2XDLLXTLAL+RJok3jnor0928NJkx
PjpL3YXrVTM44bREm+oO2Byr6Qe3ZNZsmPfbYiqqC74aYtSs+QOoE+VUKrrPxW+rWxZ1mlad9eds
DYPJ142TnHxxFZHAF/yaDYmFjv8FNpIeq3nWE7mnBZNgvgw5D5L5+ERBXS0HKkqt8T3Tprl6YXIP
X7buZQS5FNKWy8mMTbPl5cKDVnXcudD0RIy/c3fJNyu0bNO9w9duti8OHDgKX1d0eXLNFZe3vSQw
m6thKgD0b9cFXjK8f+f6OpNhnun9ZfUDuCRoiyrCw1iIkZbMOwI/0hNXO3mOEPkB3yCU7VWHHDQj
lGAHeBYPlxUSKRNfQRa6n99dwzz4jgX0ZtCXscuGS8C/7ssl82CM9rGp72HuGFNxfQhsu05inLTz
Nlub/Q+GECTBgiIsMzIV0uILILuBzb3SA/8p6gXWHyhnWjoGLs+bUo7WdRvW1ilmSUzT5LeQpnMI
htT4olAHnUNjJ2Tx0s8y7uczPazF74ESKeO/7J/jI/Wt5aqrRSd3KDNUnTFIB8ZaYaZehEg+35jG
O7lO21krOlIowFUcZ5oj0U1Z3n6gDUmujJiyM9C2FN7hHNMUx4NtZACq/kV5S4n6z7V3kObZzgqu
GqiDQEd6b40fQ7yBpO4NXWd7NQk0Hf9/Arks0aUEF1s02RavDG+wth6lgWKQqNtkyjhenUMDYA06
jR6bOI9tTOU7urH8R0kmU06ojD3CWDgBd90CWwtuA/1NbWDdCuSHrcZ6IfFVZsFAumGFlCNJrB8B
czoyTC3HwMLvwu8bAOtdqM0Kgujyd8XJ/HPsc0ws1jtyZHNvJlKOTG6rW3b4M4E1xh9mU8X3df9S
MVaMR0OqkWaMERpMyImuYGhl65a1yNI+G8tujwrrU6tVxcfTJj7qUtozAmQrTPgXU93s6bv7kdOg
eeLFrg9QgVmGemmHwNonuLEm0BL1alu8TG/CqTHzzs9i3CM+IN8BHdvK08lIiEiv2HWnqZOyOByK
NrNmM5Umnz7oYYJ+UGk3p+9giF+yfafgzD9nsSbvYel+EaX9B6SjMdymTw4SGdlVpRVFH/lh4Lp5
2UptkznbSb0uE/TXkVaROFt2r6I1dmcI/7a2HuEoY+SFOZd4+FNXXoXnHPRxX/Rqc0UrQv1m5Le1
OuGueXGRgbC5Co72JhMYI+JFgTzuiLCKKawoD1cbxIFfBUZgps2eVuR4W/PKBLs5k0+ztRSe2svE
tZWCJ9a1r21UHREUbshJdXsYQsBBdVRVMAcWLJCk2AU2KZjPwXgmPVt9i9HAmUjZRI9Y1eydhJss
bcbgLhStYNmqJJYpAj/CM0MeU9XWdkm1eaCQkp0eTFDtNH40vdvXcwK8r64Zq365Cu30Czqj1jTB
/wR4hukVHWDG/KOzyLXo65aW0mxLmTlpTngf7ZSLh1PyFk2sbluiYyjeY2focYFpokt+6dVPqXS4
rWXu1EktwpwnvawjQurJe3FzM9WqLJ6BY0QMqUrD0xhjttpY38VQVn/06s9lAmeI9xM52FBQIFiy
tAYEH/vrf86B9xdhgA3jphKyi9vTUKUAe9lY+aAAown1YmcrDTtDzZ3UXyJpbu6YnO0LrmIe+XzD
Oa9cfLw99MJS8L3umh8ceCRkqfAiPjEONP9pFQnvfBZa9UfXvBzxPYYXqor4OgGZEMiFlaa7nx3x
6DUHVh8ltnIsTSB4sCpw2tm2fHD8/PeD67s1EpN65lMjCyixcydXbMam1IIsle2i2mbmq53UGVPA
dTZWAFUn2SxlUPEjgj7VZf+KibC0GjJFUqE+5P8ntS/eL81LL0mmsbuYUGhtJuhx+R6pmBB/q7+7
U476XiqUWfWaTQfzyDGiHFvHinFyQyztwvzFENv7BlJCSOUKcDa3l1pn+nWJq9FyD4bFgWBWoDyi
cCSJw8UMsjXAUZ3KUOJOax/Rj3YHHcU3ijnzQkbtPw+/tB9F9d9qmhPGpsXZFk5AAVHx+GLpA6zs
p2q71LwiFbgFYuPlCqw3s/6bt31ajArIt24EiPP+nK7QqvC5SiJAhVSCu8sDiAhsxw+ujcpwNlp8
8B+yAPXLl1uXncuOLoEH71wMkFNl5kpklkM8mMoRpnBiEP7ffJfH1WDqMv+YaxVD19MoqAoVoOtj
x8ZM8HnUGM12dmxoXCDnjas1riUm+SU3f2Fljf+8fPx78vwBhUgL+hDyetpZcWjDHh1B+JjJk+4g
oVAVctQh3Hm8bmxMW11A1V6CJz3soq85kxC0WLAjUXKfpnxa+VuFE/CHjI99hcX8A2X4UdBGwT5N
PHOY9aHnO3I+xLAaGT4HZG9x8WypPcxzu9xMc3vTHnHXD6u9XwH3n5QEhVBAQfvM3ActjxLJuZjL
hUTJUwV5qfY+h7yCsmKhhMPtnjxPsk5ze2r6mZC5SDDF0Ym0RZQ9EOuMUgDQx3/Q5hAaIB0EQFL0
eqBf3JQErtFsYrnuggYrjbr3ZHLA7JxEXha9mzFPklxFokqfD26eF+j/u+iNetr9qZRy2qjJQ9WV
prPtlIu2m4yFLuml0LlpHhlb8aMOQsHkb0Erf4iJuZkVcY3FsmelapAwZEjQfL7R6FXY+qVeg2qR
opad5doTygUzH3/iPV8R+gsE79+1Yz5YGCc1WE7oYme2Jh6N3F6kIN/AchN35A/ZkmKRAKpEbb1Q
xQZw0MDOBp8JSOa9a2Lhc1iG0LXduhkKSjEH3qwdxda4KTGHDeVo4C+3ADDwQAKv5QvRhJTGWAhm
DPbEsULe8eYz8LcxRgYT+Bu8W7oidxhkYjac2Bn0DXpSBMj4SuQp4Cv4ccIfHf8G7yXFm1tFoW9D
61UUVb1aBFzBT1ju50sUkPQvlYAIH4DvSef3RvIFZF7oQqgoO/svx74yxPGZ8UbAbTi6rX+BzUwt
jRAO9f3UUmistwCXcFcBBxM0QGBBheLTUrTybZYhzmikZp8FtuVo02XKlT2wJtECEwRYI565crFi
ghw+AQmYr0DZIXlJAYhtPB0dutE4tnm4hRDjlV/n2pWW0JKKW3ksieIwTyajWCdZ4RqVt3bNb4as
Gfkj/Rc+CV21PwaWoWm0qTxm5hbxcirQq/2J0d+gHkVkCbOdSc97ouHDG72Awzywv7+RQ07j/Dlz
I05UeGEUfYHBAu38HjCXk1mYunK4kRt9U/CafpJVssWwUET0WDOK7hKY2y9HNSO+/mt3bJ/zvH5v
+vr84F53J4Uh+RMrk44xVm+vjl9YOXTCT74Az+C56cZsG2d6Mie0ncBFwvE5VPkYvmP88/1MfNar
Dvq6GiRDiC1iemT9gNdAJaJPZNdZ4tnkXGRG0+UZkO9oVMXpLA2HQUlqXJQ9PTMSchzfp+/m6wJa
meOKdVQ3aH2HJ9l3em/QyVkgWnUdERZxtp2CDnzKFsxbkXfUu/swHTp0LLQlXWmDm5UTCdHDyNjZ
ZSr4C4PnTMQmbuSEnMJX1PoNJxA9nPYE+QXH2K+A53hBkRdUoEJwBsDEtYPD/DV36d6ndX9BLDfJ
Ix8Vr10IiNO0CKwnX5MfmABev1NC+qaK+HfPqaeO7bLMfs754Otm0KhWxwH8pkjlAooA4Sz7/+lK
bm6ZcJF3ztpgmTfnLaOt3eAHmQPpFVbAwWbg2h71Bjv7X/feD4iSF2crSBvStOa3b1ofhLYouB+i
GPdOo60Te5+XrHil29fLwI2d2DgXm6pa1lvx3yYIyBiaK4Wo/F2xJqGbQ8kI6Qb0lxN6tgoPWmtR
52uZ0bxoDTRReXTUSghxnHU8qroZjl6sNU3ZVzJ+JfbHN9BR3LPK6p8ExTgAd1hKPL0n0GdiIhtR
G9sqOT9YvuwOij7SSr6/hqYgdAmxrX846Uoq8vOBI4PuyTC/4NMOcGqvPJN2FhGWWmfFoheqe8DC
WF8KPO+yeZXZO5lpJg342IHeBBVNuOhOmTKMSw0QHrhfsHhj1ci6Gj5jl8AuHsJxTQEw3Z9ZXTIe
mC9LMUQOj66yOEmvqVDDQl2+RguRDspg50z70od9eIBCypfcIr3+WfUOqrpoo4A0ZViLHJlhVrC1
XW10a0WNFjcvVet4fVfcYIDbaUq3srZx9uC/mNwR8cJc4tufilCSM42T/xDmFW2580TxsehwbnuY
s7cIUedaJf2Usd6g/vv2ukInnmB4VHUPFED+W70gysmzpDYPlPh+pIgfR7WQgOIoqtBPjCxdcX+s
VGbjDTEyhIBscuMrvyuYiA9e1hlJymrwpIr0bMNak7tr2Fg7iHuXpcwXpDJWytSzBr/gv9fSrYIa
tR5jV0OpDLSQTk0gRa4jSqv7gU0idWvxN0BU7/rwUEIaqSo2MUECVEVbzZf9AfC64bUUQDJ/xpdX
yHjM4tDvTVQfH9M5ML3n1cYmuKI+a37uKIXrsweVk65XV+mHrQ8fbEhM0DYHdFhuziPzPGxvkPiK
AyxrFq2N7hjJsYjJtgavyq1nq+QHnjCXic4HArW4DYaMwCdl9kqldBtf6q0eRYKePovtDAJKm2nE
FOBom3Kcwchc794b+9UBLjGs47Vk0THvgekGNSj3oBaVKfhwJ0Hx3xhtis2AgkkUqO3Rnd5AEmil
fJWvdMUUIXkYBITEK8TcB7Bq4WJW9W1LTdlli2K/GIvTJ9AbYizw4RUFq7s2me+RALpIAlbVr+ru
wTqGpTCxrvKaZeClQKWExpn/PHvmvAXl+FAyEtFIYe8jjjhnin11s6D9l/ORtPSyy5wezHck/G2L
uoRfm42Zq0iVNPpe5lH0kjcxrwyivCdiSPn4a9b73UOOwqVmLJB/om0Oo+7WEz3aWXqBynI97RU3
aEGNx4slRTOi9hO6F86KncvVm+MY2ktPtudcu7dOUZGIPgYTvaOY8a/PXMvMOxWdGvvaQejQ2NCW
GtWKqGZHzZM4hCQqQegauaF28HXd273dC5K2y7csZinJ5+HlDhsO2mOw/frMJOC3xFIwBD7Mzgfj
0GL4lfBv1wx13i11tsnTXiCcNo+zGXMLm/G4MMZytfS3oT/YrbKu9Y1LvjK+bjML2KDbqDJ38bb2
S5ezRJ4u1LhA5Fam8Xq+oPLgq50LqqVmJuVTLCcKsR3ru5Ieh6NmrddWhfDbxjaVBVkmEoheRXYO
7v0XK2TnhfxF2Ds8kwlnpQ1YKasdI7Bc+/GcNAxhfjhPnRTETxHEY0x55QPFWqZB9DWkVPMYDROi
0LCFu19na+h+obIQO3/tjOaIo0eMJKZUzOTAK8eGL+sRw7RHsNiSRNbUQ5uIwgK2pv0v/gjVpUts
SunRG1oXFZqDRnTOZ9stGwQHI3/q2wujrdGl7ziab67AjJ1ZIki8yIF66K2aqxIvZPByAPKuasFm
aRavN1UDFed9oL7FiTcc4eZFcLY3Ki5mX+yW//RsxwLU9rPYgO2H/A0CIBQ2Ihgfbqx73oDqM4tg
0ThlWVS5rRS7kmXY70MKshzjrd3ffbeSEb0/sj4j3wEnpvNqb/JQ5DErzZB3fr/vaBGS4DHn14XF
ZiTTRyReGOhpb9S05n5boi3zfyMh4KCXpuJM1OGWblszrPQ84BFzc5/q/OZPXBkcCePogtwvqZXP
ES2c1HWU4S5jeAZBVxo4CUTqbz8Dtq0Syl74g2pZqIiEX/FlylB2eKP/cx43ZNmdpX0pLBJhkqcB
arh9JGRYkKdx7t94rAFRuQkHmA6Cbd/uVOlKAi0CNQAjIRlJVA8Uogu/dafgpz/8BC/M0GDxJxrn
dUkgy5QT5WJICWGCAyaM+dac+gWizvf8xQRQm1D47lTzY3UCNkjQWKmzbU9PVzq0iiUshhiKNfYO
d+8FfjVXvjLmRDZ7MPXCXqsd3hal36uxz4xZ+I/TouEkWgumcTlmDYxwV/2EGUSk+s2WQYQOb3l8
J7FQ65sl4XHAbb/92hGpggyjMjarZNOxMjp5k4Q9WMiqNJa72e54I5x1oMDVYlM0BBdOC9ITB3GS
Sde3y7hBZtOaI24VwaFlc9YJrsz76qJG7ibB/9etVEzcm4OHT+klmm+UaeRbjxZObfLaNHliejhy
dy2J6j/JOWgY3PGr3+nAdAzurZf/GQQWfCgdDGxAT83CEvxQ2/wWbV7dgyfuGsZa5pPAVDU7L1Q4
aDJBEPOtyHN43y5QoMqwOim2VuZOUfbV8+Y6VPH/8+4Qj0EmjEIIj6gP+A0vAJIL+yJbc9MX1i77
zTqW76zoIx/21fQuEvjKNmvVmaaLDGMblJRhp6cRoQs5l3V7QJH5NkMwMFaFR1Ga+SuYincZQLlv
d9MKa7/6H94gqg1d0KZSsitHYY5Q0pzKgoP2PIamCNTrxdOiMBBgjAq6eiIeGqYYWAMQDn4KcsVT
3QVh2MS2gmBjkHWVRGJD0TUe0pci/j51CFqwhokHGEFqnXUBklYbjIKec48anhozd8t4u2fgCRld
wXhf0CIp61NSM7Ljj3Y62aGKS6H12mQoDjVmCfwtGc01+U5E8FkwgIzoQJxslurCbfQpCgl5r+ty
6h+KclW14u11zXiH03QP7GjiCwgYPaeqWrFvy38+ze/EfP96H92j6SL2oWWVkMsY6KaekiYS4yT8
vXa4x7KUAevBUZg2y6onuG1lxb6rnjFpEFP+fBZw8/Xhxrx/dnaMNf1Dvi6ALpKVP3/bsuQ3cIGY
7QDf7XQE4U21vMLHx0QVnwgUiVsSOnWi90qoZTO4upRAC6PoSRED0apU1XLM6/+awVwSr8b28dvf
q0bbP7zb+3R7Ovn0uCrBfV/cvlIecUq6T1oasnEuyZx7fMYZdGX3cKwjH8G+BdoTkIlGNTzdv988
4Xfk8qq1UZm9WXW1qki+pHifgHdxYy3pj891mAgqsjZc3Zk4oL69g8HOw39E9XVO9LjzPvcqtgeq
INPKIwlxacW+7JrlVFsGN8z8/WgAkEyGwKcMLI9ibZmRzyCGAZRoGnDoMx2wUonqicKhsjwT+mCp
Q47TLxgNbxJaBiJyx6VUzs04RJZbG+xrR5IBsSXSDPOpS+ZzcwnByYl+ZDtJYh91YWLTws1hskVp
aVRBoeby39+k1LSHBjC9m7a3Bw+aBBS6nMpOBEvCGNO/N0f+BgIKJFJTXWas0Y52QXcxmgbtQSbl
G+zkxZ29uYiTiX+Bk9T6cajashetgBU7OtWZKo+VoqoQVwGrxPsYrlQPdx2cekhtu2nujisXxjzN
rWfAoCx4mBEU0Mzdhkvtnj/XN7ivRuCvqY+1AOod72JpVKyevaRQDIPJ5DktvfaJsskUEszIErNJ
WaMbo9VTmkC+WAXnumWwuBDOiibGHjmgqZKZRTIVk/U72e5zEDLiar6hIkv4dtEHMIcIyxJtShR4
1c4TkArhIV/3bxqWGNP656Y7thnBfoK9YRi55MSNwdycs+XQBbqQOFo1zlOoeow9Z0KtGLT3RoqU
o/f9bE9XA2oRGrSRLc7Z8hDm45VsYNhgtS4YlRbjhKp9Ndc7hl9eVEd23+C5PqX3/CHONWcxYLRP
1bN7+NyvmIt348fm3Bj3TmNAS79FxjNba63Q7SPJZ4KPN35awMOoKKyPpVsvdinYCdtRpui0N7zu
ep5XqrqFSMHLEyjGhMn4KKGYNlYUkPeo6k44moINzcKeZ7D1NZjVLVdsujaoeiz9lwGekshtYVVs
SdRzzQrkHE4fDLIkonsMIHcpezKfldW7KcI0Mk4vNSiPYzRHgHIH6MlufShXFO4AXupZciZIzGJV
yb1If73vOY6oCeNVeX6i8y3035XDV5J/KqKZj6F58l1dmDsZO3fhoD8+Q7kgK76AzNPkVO7AO14b
igT2GO/2qJ85JmOBZqP8JAJdY2LF+yGgCzucvQXN48THBvOte5YmcW2caL2I1CU5M/YQZS3syovf
CdNiQ8yhKLvt9CAQhkwZ8xhhsjSMW9WkhEYZ5tV5+vAAhyFm8aF3FS0BV4BuGIpvuoW3eBlrGWEI
HJ+ofd8Ymb0awP/4rNmlIw/gbwaeTVwVWDZWyATU0yy6boYJlOtX5K7FBxSFPbt0tnDM7y3UMOEs
NMDgFf105U6xUOzTh1I6APpi4qpIGFP7qKTG6MavBrbD5nLMr+3uFmBy+tbOp3bMJe+OotL+uadh
EA+na7JsZNc5Sf0EcHfIv33bFqUxQDd2/XDHJxpBwgZSjXtV8FCG6XKva2bTe2AQx+7lhpy6o1rD
mHmZ8KzKyvpmpm1GyyMwRpkIex7NP/X3YwWzv0uZL36zzkYx7YM8pHE1R3niu7OzVniYVBowzLDe
52hIGR+pJfofOdZwZsdRG3xdBTZ/wtHlXoN57W7sEeyMGOgsEbolMoNHzzcpzgZ0HBKuq83ZW/xs
LuQeA11riPTT5L7Wvu/zI8APpkeA2FuoUNZemHfifKhBbbGlWkEqkBvkgbCQx7GTZJ4pX8jMi4GU
C4Clf4C/Yx7G9LS47oE4ybx8HVcZDk7hpbmFo41Rn+vqR1/k24y1qsr4Zx/9G5yqEuxAOS8HFWWR
UwSwP44IgMMC/XIgkedtS/qZAWUiwFqOSukFlKSWziZjfdeZtIwp7IINqhx2G15KiXY4LH+WIeSS
MyL2uAKY4wuGD6vN+kI1zFzeyLVPQan/HhajIZbtikFcSf2TV8x2HsPPn65Phpu3Cih7IemVl+lt
7/BfFlwfT+oGaaHOkF6wee6cnCR/Q80mQhbnqBorE0zEVHAcZCJK5aGmIbijQVEo2B9wOaIcmZyk
lOqZyi9nDTYbatOFt42IQuMnht9EZk4rLmS4ZH0bIxRoeSDaeBUurLzn3QEb93oBnTkVpCxeXSF2
sD3UlnNIqzbprrDXYoRBwe7RJDJlRbHAfxNVrwjcQb9zBOXYGnc5MqIUg5M9Qj73De1jL4KD94Mh
njDdNI4Tcj8/NjJH0ehwUdk2indHx9Rcqqqobb1sToKwIO8RVRqrIJM89J7WD9aSBrG9+zd6mqGs
Q4wAf1MrXf8GqrNEgdG7sYxXIXHgDiNXtqfwD5IW0HIgR/1WxPOb05G7r5TOi2uo9Um3K6q+J5t6
hEeZcx/EJraz+MZxS8kvUleynPlhXLFhpKD0kgkhyyQwYULyW7t0cYwh5zVgGtLQ6f8Z7UCxN2yU
e9NY6vJ0D0WtYEHE0NesNqnRMtxsmoWbWSchALrguABq1YBKTEl7av6H+ezaHcuko7g5F5dczMCr
UCAx5g6FtDFs3BGCc3F/jTI+Nk3aGclYTngiKmoH255QUl59iblZb4iWBBtJRYQrxORshHZ9J20V
RwiqktCv1IHfkdYd2yflDdjSg/h4c3rLQQDjQiGC++33xxkf8O2tLGO57+rVPlGTQAQwdHvfZStN
SqC1TCb5rXgqjI6Rs03JPpaVJq6AXEswjJLsTODWPpimA8fF2owOTYGd9lchLvemGCFPoayDxdbH
OaVao775iyp/hl5bdZ39sp9u8M1zqOSdgbN/e/PeWJEYcWYgaX0OPW637LOO0qpUZC8jUzZVA8Aq
smd1r/nNqBoe04XyEh1JCjwPPrdEqkwE5qjq0l51HdSymcgQLzT0uz3hKBSNAkEomO/EB3aZydxh
83A8l9X7kH2ysaSzdqO0GS7PD985548Da1whZe12a+fHYU3i23aGi4WA54CX4VS4g9epIFSKpabf
28dCtBfWJT/sLnoQMtlxDyFzY4wfGTTVHhQT8KqFd2ljcOdhCNDILXd65Bgwd7JgH+IWymKS2yQZ
OqHVL3x03j5vXFZx9BTavmP9fG56u3p4t1KttNGfluho8+mcltz6b3kOKdrSJUWQUqcq0FJ/23GV
17xApoOZy1bNcM/5f0227gSVgg1QdPz1S57MmBdbV/PX+Aecic3/bDgFILR+i4nJXorkFHvZ/Dne
hnaK2NVbbn7fLk/FTNJmCEI6bossoRY6E9g+14UoROvTXv91apXPIhyfxdysdW+//JN+WjJ7iE7b
yGZ10SkKgwO5TeWXcE5sBsW0wsVZt+ZLMBTKIlBveyEXB/1lYTuOIkO/ynfV6+xucQ2hjyEUZTlI
ppsRkqTklufZ/HtFissGgVlwhRKjqx7B24iIqwX5AhJTR0CFsYNEaQAUXd6AjaqdbUb+w81VZkIK
sOBePfDlLhKD4qobNaafflcVkCutIsUi493aYmJRwQF3E0ecbidkzEAAY2i5oBASwm6yFxCNAix1
SaqDRtxFqgIuKw3SOLroTq6LaEIgIWuWxOUte584LS+dM0UOAZmCWmsFI9KV+d24k3qCBgo0gmUf
RcZplxtVULiFSVFmqBXBlyE6nsO/hkHXmLHWSagfds+Fs3X3ooBaus35pu203LTjGuY7nUVXvdQz
Xk+UJ4LHXw+wPgVzJ3qo+IsO5syq2t/1BzRH4Z6jByOy8llTRb0+JvbcRIpRXuAOQk0XoXJL6zrx
HECI8bzzC/KL83Mn2Nzom6FDFnM+OMP4XsWmPTrubTfjYFLUR0MuLudU/pwXk/6G1E7hBf0iqg3C
vAITdzQmv/aczMuLcyZgZDLWS2nXYBDc/wikyAOeMEthadahEVPGASWDAZ2qinra/z27KbSJPxG8
GeIRgVd+C+E5Rds4AnMeHO59A+J8QKFitbHtl+JOUKIqVXlAUj0IQdRRqUvhr0oAAyZYZD9BOEy9
5GJTFVVBii6Spaar4ELvJmrrnC1BMkzjgDFFruhKsVMqspvdYbUCFGPfRc00eP/9H/LyJK7Dklwg
9TH2piOfBlEl7wzU72L2UsGgPi9LqkWMtXCncKS326VIMU4/+tA7fwCmU+NvuOC+WEZP7sqvHVTO
5DDOUOZB+IZFgCuZFkadQ/qnsx0/q+8ddwpyuos4kRuJStnzh/TtDVgbitDAD4Cy31fApcgDnXpF
BaGvXKMQGYoRuqECrg9LjdDDrwdMC3YTHhpFwy1rN9vgfxIi3wmbSeLWKSzMp4DxoaJmtH1SXwOf
0GbWkhRNDNB9LSVrtuNiTpf9t3qkbZCT+1WwN+vvTx4yqZB+XrLlIdbI0i+2+h9j/wP7uievj1F1
iHlrF0/89n33T59PNEiqBuv6LwKJKDoy/iB17+Z7dIXlfM/Kl2YC1NMBvm06W5JYruEPjXKcJUce
qsQhPrs7BAK4szVuJ7PJhJrGTIuSKVUHLN2AF2PMpVmvudgOuJ2HHKDEPQ9j88vpjlIgDolxnMlu
Fs+TslT1Ana4Cip/7WLd5M890euR6v5/xdl50cRhZIRioeOh4nSSeWUADxFFWo8igjprq7I4ctNo
oTP2232PoByxBKGoTFTBeayxFSMa06D2+Ggq/YqQk6UKZBvDarsv0ivY0zGxEbNwvxDUAOspmlg8
AVkrxHelsOV3mDiGUfzLdHRWb9jg/SMwepuyMbzfsus/s/ZZG0/L+YkPMYHvBQxJdJ/6NDtt/NwD
EVvGpU0Wh3xkfsPo8528w+CYqgoNvwG5TZ4nQGZkqvizPKNAUcMpWzZg1YeS3kmIfDWqqlAGxSvl
T+yb9ozgcMoovExPi3FclEcmMllQQfnoiIuqSMh7igQ87Bd4AfE0JvjVxSj4ulYR02mDv3MHOPqu
BqYRZL7H5J07RoAoKxblUieauPa1G51Q06/1rTVsoA+bLJIsleXpVmvKFvi/+wmtrU7QAoObG4Vy
OjubtE7y1jU0WLZgpj+zk6UMgYDVqHfRxYLZluS8JIYnnCOAKXYT2iTDNGkGI+re+Tc1gCpewHuH
/3wtfpToaV/UR10+HfpcJh5p/+u+Da+RcOF/03cKdYb5Tdy2R+mOIBcf47ujHIyViL6M6aB7TuEh
yuTNRUd0NTfGY2P/USV4vuGgcOHI4W+mZv6znXuKSpjmkcuPS28aM/8giQFXT3BSaos3quGub8dG
SQNxa6U10grQe+14VvGJZ8KzgJn2IqzVnWF0EheN9+QTHKioGnVSqcJuDjzbCD3h4FxGaXh0JZ8o
FTE956pzv/Xdx2i0m4vA+vUgHGwSbUrv+U1UgYHQO02fHMcsGRvoT56CI/TPbKBPZT5MwHbzMubm
pYxsxgFz8qh1Xv1fN6N8llWPZzyCyazfo1l/I07wXbsEATCBe6eBNIH1Q2uaOpYJjCHvGOkTYlN9
YANtcF+dP9GB+vbKIJp9zb90uBrFnGhQ60C3hyjL0rT8oiA2slfpkknUGJWQIFLmgA5VnzeeOkDa
Ib2NNc2qgR18ua9oz4H1cyYoiAF0Irz6B+H4f3ojROO8xiQEzllAn2TGiIcjyvQ1srNxbEGTezya
1JVL6h1wl3sXA7v8XSZCv3ntcIRxEZPPVG/haZ+wwGwXXPoTWe0mcn4MAlCSXovgn+2ULJCtp5/j
gHJA2eeSC7v4L3MGPyhdgyWiMvdcEcelLK54lpkDgUzDKOksh7SQUhiNubh6jQhCw0RensyNjThv
79AMOb6cS5toSk0PfyycAvENE0iKpmR9EDUNyEJfqDBGvx5i1RG5cQQ3kH5LrTyhNdabV3QoygTg
2GGCS4ykTWZwEKkQy6blb+aN1X6+OmpQZmfK+/DmZFhV03BTBj5ROLIRQxl35gs5eKronhZ3hxC2
r+GLXZrGkAViJ13WQNshKgMy+BUmr+J3GgoXdj0YWfPXlR0hPmRrkGLDqDaEJeC6FVWnZ0R/RkwF
1CI/4rPtTwAZXHlont3LcMDOur5U1QSrlU2rvFU9QCnw1TC8ECMTgBtK7bOCIe02mheyOD98sHRP
2nyIbH0+YqNpq7/1DQ1gzCCTMgTnpWUxac7MKn+MGoOKfzVgxaZ4I+3ohbn10zejiRe+E7ULfb9q
SiTKG8VeknocdRipvdWiOK4mKt/Ll2CewiCT5mcn75XVFMHwqWsZxXoqF/mPXzbDIlQov7qivlbZ
X8v0fP7TeU1c+lRGfe0DeADAG6Laspqt0Whg74PUriPzPewQuNgF+4o4l/s0X6ZC6og7zo1TqmRY
So7pgHmIunqevg8UA65ia4E4capYq1+lEZJFVljVAjKMpx+5zv8Bx2ijh45o3AXKc34dqqkZUUQU
1A8+GACJ/eGew5Wh3x57hNxZRfVVqjMNT9J9QBmrNH92f4C0jy7098AnCTce3xrp1VKUdZsrMg8Y
+DE69XYOA5mEvJqZZx7Lkj6t0034OjWHgHhEwN+nXspR9iQUw8SykhxqRR8GNMdH05nDGKqCVGgE
Y0xl/xj2yt77yDmk7LifeaQpAkQuniGwmvf2FaIHB+gNje6pb4gIGg2NBiS6Ehb8R2VhUKa4JuI5
eDUVTK2HmKgfzxFANU77OD2CY1Ii38/HRfRbJUt2dscsDgu5ovZ5ZHwi3baiX3O2kZa5rNw/97rr
AovRE5cqvTi2wGxNmxdeI+5YSYgUaxLKDzb6JghJm4Zc4EaxswYSdYQ8NYcidsovIydn290nqaKn
wrYNBXIrX7ywcRp6yZ8WiYTJHa6uuLLP0zNjOM2LOMninE1RLU6Biqq/yv2bGPXxeJFVmmsdaqF1
+IaP2pazheRtZXVIkqBOHwv8zorI3bkZbUICB3SVKO9kIBjpbJygoOeu5378lbeHeGG8+7a9N3Ix
75VJvWjOeiCDCiL6xEJV7ttyjZnsKT8ts8hMIQX0PlpSyg5VFANr8OzejSpxk4sO75W9kw0/jv8Z
V0GvGtVUmgcKfs1BLtbCxTmnFFdhJuEgS9+bK/ZtF/Wu3zEG1dKj6FrOtsidViTdPwefbvaKbe7V
6SY6tMVQ7hlxJre6RXhznTNpWUEG/PcOP3g1pBncqiE87o0myC46Qyc09eoJW4CSohwZXvE2ULzv
AykzeYX7IZgnBWDIWYthQ3/+YQqLPTnsCgCgZwtPSQA51hd3eJclXH9jvfZUYBMzhwfmOykZ+omm
CjA3Lri/tLhG5xgiVCYte+jiUgkc6ztvTddxiOuwCKNJk585s5pr4fRQv4bT94i9uYtsNpl7zaU8
08us7gxdtdn178LA0iO67KouUJGHv+KSy4CFsA1WD+6rqenXMuSHpHn2UoOW2hdRi3KvEnzCvMQ9
tobBDS6KIloQ/XTqRgXHxH4rCOVSYyhtxcxT9xIuQ7A1yS8ujRG1mzKpbc4/2jvBVm19YPG3WijO
PfnKqyQ8k7pChbwTYD4z51oGqPgVYTR0V4eg02feN4zA9EVEr3oQDxMWkMx0Lhmw9ITzbfvyKzix
NRUZgp/W2ghPP7X6at+qt6UWBX2Z88fPCAP1V6wgqfadEDjGhsxu/fXO1u0P14XyE18HZHlU9ofw
xsGjo7iMIHcQxLVC+b1jPUDEQ3CJ/FFTL1eXufv1U863+ICJnoPMdRc1eUQtnoQN1aV2Dh3Mp2lW
+hRm8tmEJslJpox38LC49dppnLUsuH+DkXvi3FHFGmed8zcMPmZ0Zl1gDdsBJ19yMSIuwdjOLf2y
YrrX8hIAn/5c7nnr6MBDAbe5vtbIaoS9Dys8tA8CjOCTZFV+SRpywE/Qa5H5y8GINQbJXWjw43D/
9n9Av5j4S92swNcc/Zo4+XZhS520yy2mrQKcedwivUDaoBlv1qM4Sn+3Utdin9wbNg+Qqr9Sev+V
7MbxdUqgZdbCSf0oIQP4nIob75XhkLcj91Mutz170LHVb6q5vcBAX82KqRnPRfLNU5CJEM2PQwZN
Cbu2gK9bLcK0G8FOBdMN/l9r5MF9dxFr53d+VTtZ6+izmWxBL2QwPAKCrEN1ucHHkbjwkmeoxry9
E/227AcLijRl9ZF5d3eUjMwzGMSrShqwV8RF7+Jr/DhVka+gQKa/EHp/ueFN392XobjMYc+QjzLU
1OJrtre4pULqlw6cOLpnj/5gg9MLtVOdetbmfWOH/MMRcIoYkApQEst/aSMliuzBQN3BQsbUWThe
Sl8Z1uknMFkC/ai8bAQRhMFI1LduNhBuv0qW05FG92w+fNvjPQCaYgyzbjFLbnAen9DIgx+uKuuH
9D6f+AWmZPWWCWkEe56zPskhW+xyJqSnC73e++AzZb+PRnBZi0G6s7GQxwNLm0ag2XmIaQBUw3/8
zTyo6LN3vipdNv9U7hATqohiaRCxD5BiBPJxxvg5CzYXtIp1bD/M4jOE2BrH3rTzK+Ki4hBcpabZ
qY3jUKl5P3GrPZB724QNqVco+i8htrXLuY4lquWhbkoxayYAtOWjIFoXPSrTxRfXWJnYLy8Qjzmr
KIax/TLozL+Sxja6G7SAPn1a6u+AFLDP+DO8FUiYpk/NDPFcbr2tUt4Athnj5HwsKM1bvcQQ4KtU
s8p3xw+gVpnj1UCZFT1RLFUFR58M2NDsc0Os5cwVMB6402aTMsS1DhbNLs91eNhL8Le3CVtwcjSi
VYqq+pp9e1BZwca+AWYic8Syh5KKNGQDrg3Q7G4Ar4fo126G3USlMpZTFeCBee5mUOwUib4cthJp
ktCVWGpdc3L8hLYzfoPUhYmY7Uu8xaGlV017lVtR4Eisu/epoDPPBK6gABms5Q9J5JyJiyS7Zvnk
2nq/Au6J+FHRGdyRkJyHaRvLaheGooAUv7DIIxul6ATeGyFcUuF7ZL3ngTrClNWc3tzlDWLIC8Wj
J0hqmKC5jpJx7jxUlinCB6aYkqJqVPldx34LQ91NJPkNL2QXWOLbu58soMnLNjXGtdga0pZ3mwfs
OVkr/Z4mqS2z5IyVO86kW6rONlmmNdBubKxlNu8qy55YNj3uGSkU86nKrGoWSFy2a8KZUN1Cdc3M
RHM06+qWETJYlJZlvcB/kHH1qfufOKOptSKcR8F1Fmp543ZhoaROasSw7tKOxTfnOU1pETNJ5/T4
Lj48Mwvwnv5HDjmNB60jNfH92n+SOg08KlMtszTqunmHl5ZUHTh9+oTxHzpLXTl16PqWMkMm37Fu
V8Mp5A52CqrhEKpRUU2p3hR3ygeYcwfBphuzsY2j190AovEVxZNCtUYG28vFuUoRv6/Z8OUtPwq0
cqTUthCMAxDOKNR0vp3I8JEMu6Sn9ED5+Z/1bhNr5PzPsrC+JpxyScCuiC1te6pwLvwwrT986O2V
bhDh5DEaZU6vRnd99NZsEYwDKh9cYuANv9jy2mQO6Dhy/uUbJDvI9g8SztpUSikGScvGlqDpPl1q
lELLRSSgOgvcvNceSpSZBmSSmjEEmUXE1D4VE1Jv7x92PZ8USljBzfv7Tbw93nWqmSk3z33i3DcH
X4svWSEHBt7JiD6cjgRSxUEHIQI5syzJCf2Rz9B9KouA6s34+q6x9pzq1ZikaSRKHFjfekAyurCW
XX97gU16DAXiQHFtdf/JwI36QIDG4ZbdeeE3AVpRHqDJYWvMaMHhPkOPtwDPH23y3dRUBwuBZJXW
fRxUO1vL4D6krxuVW4tQcoVEQreYQE5XhSFKFcwFXQuC8ngEbaxg9G+SIIU4u7tytHQ3O82eIwc1
eCQDLOsiOduMbQ2fco/BF6ugreXiBDBqwDKM9mhpOGclEgDa5FaZlinCAZuk8SkXc9mqPeX34MYU
ljH1suXforCKYpzIT2ML/g/APn1mQl0zh2lheoB/y564ELyZT+K7Z6RQI2ThJJTXf9s/r9x8WXSL
lmIlWEEg7bs5txB8QohmT12jKHgqnvPkrR8XrkK5lRmIOCNt/XXgoE/cpZWliRWUQAQtdEVk4QJl
niKmwT8VyKHFbSWIYYtQu8p4rlXTWvvUQu6iPMSjuB+QSN2doDyEsqJ5khJB4tkSlVy7ZDQM0jsh
Jr+Y2QcB9UCl+bKXUZ4hwynr5she6tKuUllYWRE55mOju4p5Pmht/Tx1T09bR8TozsdBYHKSDINT
Lg0JlA9drxY3c1DhNZDoKz52ifu0QjiIo6cd8l9JfuDSj5NJmzftQ4Kau9WnqJLDjGHX5Z6t9uxK
WV7yOgWC/UNxU9D6XcXunz07X+bCZZkAAUSgq2wLo9L2QOMKlWJhSu947e2LXGe0uDJIsT4IBj++
5sYigh4XNXaSS+xQfdoGba93GYeIckh89mG1jpYthaE+HrXmlDbY0J1yYbVit6OJIhgokOu5ajUu
OBQVu+92JqeYnxstZ9oy4u78p9WZIH9Uyw2ZiW7FRl12PhqLt8D7ENzStAhr87edzAx1O0VYjY6o
QNOZ2g/89HvQgQW58g/9MPm7yYw+diOrAIJtfb1wrLsgCjc4MUxZXVAoDd//D9ejbap/qgldPChF
6vev+E7zCXC2pOjd+bLOsVgTtkN2zjMounmGfMsFAz3uKW6rPgx+/g4hYNfNI3MynIpvmOGOrxtj
e88rVTSdFDHthnrlyB5K8p+zR124DaMKgdD81ukzKq76BRCVG71B/89r2DNwRnZ5CXnrS38r0W7V
s2cgC6BkEYy/CbRTVD4p9tVubplIoUNmKOUkdEGKnclOAc07y9H9ay7Q/xKMfTeXcb93dJOSNTz7
YVbdnPYojcKVtBtiRWk29XoxkAK9mnIWdB/SeD/0b7SRqfn8SzQzNNBpkdR9oBrESeNGp24Glf/O
MnKAPNLjmX2lihyGfsF6B1O+gdkOurWApo82g8aOaCqELo2dx6S2qUfIZJU/z9TLrDlTaA1g+/vZ
+fz7vg1rDvqZOAnpxWjvgx4P/0D7sBLH8zMO7jg0SBdWYrFOCHi35CEP4SH+H+XhBNNEa5wyt3hg
ZtOWnS6fXOq32dkH4R61wlUd8kuxZAjxFm8G+eFAsQQijFot6yQOUFLPyk3MFitoAcKmqo2S6Mag
42WivwqnHRjUZGY7UrLZpsjjAsDmSFFUxJ2+VQpKp7as+kr4n0M6wncWNKBPjXKL+YdYl6YfLLCv
Ps5eaitx0I6GZK1B6YX9SnxkLE5SgKa9b5ejMfM7P3ORYt9iFB076T4Jq9q4DhOkOyT8iQxK82ZW
NPnEFrQy6u+sy9OwIeO7BfyuWB0BCzxIUC5/oehoFF0rIETDlvKQ8qMzAPs1pTG37UnMMvyLiZp+
t/hWFz2DBqQOoYp3F01lHxhokYchtbLWBzhVwIl6b1BBWauFO/v7GGh1TtRe2VjDJhKVPPxt1uzu
a0Hq7jxQtKgFMPW9OvxQGNZsayq2XSuhTEiPk4N8QQjVmdWzmfOW3wljpkqB1XKwhZrRoDgh3kHf
y9LvUl0RkelgT5YQ5Edo7/kxGX+NerRXzXTr5x5T22yRGNoyDvbS25vGetdVYaV0OpzkAsHHk49b
GY3i3i5mxamzvWmJhyZIbDP96427fU0lPIYi3t3dQ8TC4McLOIHQRTKPJe68saNZwgiZH7mboqK4
16GJQO0ni0HAFx3UrCQuLNaI0nP1OjviPxTCFvBvsENF36ikQGJT3C7tti+rWoNWsGlXk4dQLTLS
wyS6qi3gsvLK0X91sNGY1pWxOuf5RUA08TwPrkR2fua/ihW5x4bQDL5qlhGhSA1TuWqjU6CkDvY7
0kvaf18oM/ldYaHvn/7Mp4cqH0F0P2769Nr7e8QjZZI3KVkBPM0ymQd323XCxZ2XuyUEI3w1qS8p
t2hW12t8o6b5ZHf/TPYFXjm8vzAxv4wnt10rw/ymwX3IMoRuTQlDRWHMpPZwVk3vmkfbfLNJ65V8
Yd2rm9rbTVg3uWFw4JTjcUH6j081qVHZ6o0OwdreptwmcMUrd8Z4Mg6vUIl/1JGPnGiAK1RBjrGj
let+bmXmuzT2tESJK1Z19HwMu9bgCFP3oI+5a16O2t++d8GT8EWhMta/aTrxubImbmv6otwmXQwz
QUQWjKKw5hWqkzJOAGCm7qx2GMi6vanhy/pSsDP5wvm3lKh/TIwvRvSg45AoJlrUt79pEnOT21uc
tYESGfLyfe16kmZ2EgIcxZ9RfNT7BYJZvO0qYjHp3T5dcTzggKdffktIOjbM/6ulVll+SPE6On4A
4f4UAcfUAA3+KDgqo1OEz4NkaUvnWLqzCgD9z3GGLDCxhAg5cSjuAUCIduR/gstYT4jrL5yZZWSh
B9KLHYgwePUI4XkE5eGeQUBlk0oeS2vqper0BPacLb3Dfmi6nrfOj1VKKs21XkPG1hr+V33Rwbis
sHCwsogJoySTymVraRn+miyfkOl0VGRuV/uzX22+55NoWud97mobn1j3eaBW1x3ZDcE6TFJ1wuDW
YURP8L49TCvsnrWKWoIFKzdihsplyT7OMcYmNGV4zVroQYUl1TdXm7JZRx5GJX+Ds8+5ZoqquOJN
Fj3KDPSJ3B2cTBdxsz8nB61pBu4klEtN1+T+E6tQfOk2c8qBrFDS8oy8N1iyJKFJUolDNES7lLq3
W1HftsvITxGaVkN2fy1r5q/8rlHBxVf6KgzgVE8R3h0HRbSNAMm5u7S8B9saI4AqguisPNpWsiLO
e0cU0kCI0ZNJt/5S7+4BVBaDMv0yos9f5V8hoa4hmRvp/I/pWW/g390HmyhaixH2vLTdt7YRkC+T
lnif1OEMuqJnyTjOtNnFrLWy4YvCc36/fu6vjfzA7k/MoSjnYeQ4XBGfwQTL/JO7BKu5UXZKiv5O
6ltHSkViE8XQJfLwqZlavP0Q5BjmNopSW2Mjj6qYcTuSChQd6zCNEc1ZgUITVCzUrZuHv/iUdN3g
SpiRwALkysoag8wckaWTFPOizf7XjJi9a/Cet9KE1aeZfoxlZij58If1VL2otjhOGE4B73wyloDV
UhYa+Fv7JIhT4fhJAkl50fTp0tV4tQ98RvW+FP1mwvn5OHp1e+gJKdMK/RforqXivNYpu7wcsfTu
bMTTK5pTZIW1wdsDtjqyxIbNQIvHAYi6DPKnHaRWNXh/MiI85bTC1bEU20Gd7vqczTxQ1RdldmnW
JZXgJAHNRBPIjh0M9l+Su1EI9SJzwb94/O5J9d1js7BaZUNCt5sAJntmc0+/Atq/EphnstZJMmuN
8ifPcV8WXxzK2/gfmlAcwfq5hgsNdM0bp/6bPSggz/EKWRaOsR8/zEhGY0nz7MlH9/9QdyBOs3zQ
xa1KKkc8t2/XDQ6i8IYyZWthq49vfROEKp7UuVEBbE9R1RBwhVu2Rp5v6boIf4695ns1/aLFMTmF
62BMSBU0g215EsQbe9b4N8DIJC0MTHiM6w/JKGNEE54/51jROL2lm17WStFaO2nVYI/Tyas5qQ87
/omlOrwlpHJcs6HQRx3Mmr2dPGYBXqKvJ1Ay9HXOt4b5nQUzHFFEA5/pl6Tq0J6WV1ApDiL9wRRu
cLcfGwnmIl6ckNOQlthUoLscQSRfZ4XiRHtXel8GHHGtZuKIITJOi2M4CS7Np5wr+OkvWfkmLy8/
IYocA2FH8gkXW0wy/3Y0vjoDDa9HNxYLFakkfVFpkeikc4LT2uYHHsmg/gA1qe0+5UZpb7WQJ4PX
Q+2XrdX73QLNDkZb8A7094W1E/f4mrZYCZnOz36jZFWTjPuXBiH9ArQmCDrYXSWs2pWyWf8TFDLU
+1/x9mvZiyoCkAooJDVk6ZJ8wg60MVe1MIfzxDfGr4lmzmyD0PcYFsOm/VNauEmJsbW3Tqrsmpue
UCGVXbCBOoWtODqxhAaRtB6ynUj257hP95qSdRsGpXOs2wulKgG8PJlM81gPfXfkONZ3/tWzmLIh
DYLi5QtjWcCZFRexGBfKId0Fw+XbBF/GfPhMmXJHrSe7iylXLVtT2KqrHe6Fz9IfWSmJRVlIAYu5
bpvjJvzZ/cJoWQNExcMoU3DSSnjPASBHfV5ZuyjhsMq3r+tQ5F2cMZWm7ledOrJKnAwBhGS0jz+O
rBEZ0MgiVYkCh35HNtLIjw7ONqIJfo4i/ztovYnBd3pRtoTMYpT5JLrOu6MRjPsJmi4Mn4/V8s1X
0FiJbe814l2466sNIB6V3t+bTXlxYZKgig3oIx3DcKBTJfyGah8A44l3/MOYmP3zuf/ePmbrOiHi
et4KFAZ5CaFLOuLmp9l4qTWffhjj1SFTfgIH07wG1UGaMXewnDb2ZEcTVH1ItWkdIvAF9QQ3wy0f
QUC549dpsg640+bRJcYJESyKFTj+NX9BVsSGaOer+OKQ1Xgw2AW5oLW3V21hCQd/sUifNXTQ1+lb
GR8oSHOotzEwzGadn5TsnP28OG+5tCUAq5hqmVfrrBbjta+JtkI21hcAZ0m+Nt2hJPOIvJHTjtVK
PTW8MileNOyXgG8zH1YhZ85XNH034zlUkitJCBQoT8Il2tKTec4Kkmbhb1dIO2hD9X41MnBFFZeP
Cjxu33x6zAjqWGx0Eyv9OvnK7GdHmwOY6NbmydOyL8mxxoamrq1ZomkH7dtCemTJB56/3xMfGDSD
Yoo1zoQmRSd/z0eKAkfI6+2tbDlZbH+I6MOlgaIrPaocIL36czlMFyaOmRA3Oty2Llnl1DeKC/D4
jo/bqN0frBNoarm2T6hg3/z7NkIEiHapFkwJoBQOVpY8t3sdUgvMuZqF7MpybZwEtsJRSMp7+v0/
2owJlG3pFzECwHB+Fofmv3/hfXBpGeK5ZcsJ1Xk8IbOoB3iPWBsaM9KpiCdJ8Wv+54Yt8Eu/KX1t
/Xt275yDs+SfItoelH73xObIPC5lINJo22bL2HQwrwvRetJJtINZy7DLYGEdtCBir2jdyA2WDnM4
X4btlxh39hUxrG5i7wzSwH5c0fqF/XHS2Rm8ByG7q8AsZfrc7p32LLj1i5dfmhSDn72xVkKPetda
OYHFzr5YIsntiuJyl6YG/rFf3cFKVr5rStvZtoV5YGKyb4BrMbjDdKlQfPvGOYoiE8RulW3IGBpp
X+K5wTfLbLjon4KD/4yTPCDgMQVxOkJ3JJGiftyHBE/3DgXEiU0+rkSqExFXxO4Nmo14jzu6cPbK
vzV64ZO07Dbd8j2K2fn3OIslNv6vJusPJw43G9Vrz2lhYYtw8YxSkGBgx4UmHwTENB4sNY9KB65n
SXSk/sjkgDlEkde2EdXJJr96Qxnt+uTCe+AHf5skpJAQb8glYoWVcD0KcBxbAW6qqdCyYUAaHeU6
xgGmAwDbMOnOjNzozm34cGe6eW8vmNfkjIo9z9leHUZfLcVuYCBffzaDhi6HHH+mT2muAoM5OE5s
FxBCQNU6bPjURU0MyfFvm2DU4OOcalKCkYG1FTgPLGLQRzFwVzyrwtZEAFvG/xYiNuDDJtxgG9SG
BnILBODblO1scnHM7mJHsLVZDNqIbf6oXaznKfQRcdko97u51LUBvFFKf3sFFtLAbJ1OuX9pE/Wj
09j6U97FguU2sCpHMCa4SMXZswxPzm6gXwpErTFWxGOY0B0edWosTd+Cvt3UonTD9VIJG5x0sj/B
iEBbnRHg9RhLtvcW4zw3FSBjAM6drbX+Lnan3E0a7mFs3LZjwogCN/eFvZgivslbakpxcOcdUbFt
EYo6/OwO4gaSBrX2Z0liw2I0thwn1RVo7rz/91nGh+vXEkdjtnPZOVBx2g/fJXy90i0VegJ0fRnW
PDVZ18OQbi1bdkbhkPTZcdUDqz5XhwVUj1wuzEuLl+DvYvfuJ9O1si9hoWR2bNFu+p6oPyJ3Fu8p
Ogrl/R6D6U+iFyuqIcgPjzw1LusLqTxWyVcCD22ExwI6yl6yXshPbNGuySqrEi3S3Fcgmc2N6vCP
aVwJ2iL5moxIkLKezVY4q8mjNoVoXh9S5Aff8tiofWpkj/lUr/luTNTzjj9whocanNXr0vr+mEOr
Cgo+3oLIFy+u4NYpoadIYSslBXDfs5mp32KZdZm+g1FHQ0rA/W4BcJ89SV2eAdBF9cZSZqmK6B6D
9s7sSnQC0HKMKgh2dcYv7xJ80pLNCr9gCqyezCiO1IBzhugtOrcB94SDUD31fBFIWHZ7wgIG92fz
E6bpPwGFLP5nqnr2D5aO3eKAmJd1gypT6cS+z3Oltt86ehZmgpXs72HNRIUewWMTwKR7p0DzHNb+
F5bWKXfjKPwPql6Ccg1zQ8GcE3FVuRUQ7OHsEO6J7pI6mJcc9Udpqx+osZ96tglro/y9474Nnemj
/9I/eUXPPARx8i1nWYQ97SsvrrYQhCvPVhhpmj/L8ivA2U89n2qEuHkptfPuBLAS8OSgxNIC1vmn
o1sw8pMvYP2fGFKp82DtwpRNVxaABvv/Lg3HNdY2ycy4pzOS7/R7j/jyjSJjc/0RLYGPc5+bXDIM
19VXh5tw+MutS9kiM1M/IyXtqQN+/Hwy96HFw3H48OauN/t6jgOMUf678LxnNklBMHLZIVg9ESjz
J364IMwrVMB4nQHEXH4fX/1vT/InzmHUxWEjFs5kfcociXGAbuJWVaJJ8XwGG4PVXDBsza3EdIET
biMKIRS1Jy9G9xytrVKJh/m1+ao2w/ezzyPrjabR6S2f+EjFuhd5IilY0B4m3t9Jwp8Mid39/Cg9
MwOYP1QmJ9ZoRd2NV6I/4nrLGJSXAoTRjoDozPPHbC2wYVAcrWvMKDHNuB+yOxdSlpVgoNrGuenK
eBk0I6f9VUuJeOh7SwToHbf/4sgr2bd/TtEdU4MYbl+q4fSja+tXEjDdoM85EYfcAhPpvu0SUVDC
TKc9hZ1dRpyx7AwzgxyoWUBVlNB4v8MZ7rCRNsZZpl3lIl6EM80hX01y/3ACssYGzLvcwMyaS++q
KgDHHfyYBJY2hpPI/CKKLgWASwfsTl/aFWv6ceHEaUabGjcB4VVrUObUEvLGA/6zUe0lzUs6/sno
pzCUVcYJf6M+ZnX+M4Cxa1VFQKreP+ReUs3DGO+E2o+Hu4y9OjBi2rRni0YSVVp0Iu1AXxj6DXWJ
ss+fJzUaaiJkwsFqwi5kqw4F0/s9SalWP6JRmH3dPa2VcI219JVVmWdr0Oyj1GwzcDocorsvJUz7
bfsNjhyjOpIbnz/kTIF+7/o2QtdEwb9P8mKh51JyFSgUwq2SArOndBxXr87P1iXCrCmxfzpCmQ2k
hLJYRQLHcbFFL+Lcm30LZ5bxzRwZXemkbfLL/uwFmZrBlh3HEFiKEuObwkDLNBfNF8l7by0rrBVw
eknAClkmR3Ff/Ab+ZahJbHTzvPgSgHliGlPXZ36Ou7f7rMWPhn88JBof5Jw/KbDhgOsBPj4BaE67
7WyyUwRGIIeL/EC0vWPmyxAsWXVhjusLe8AOUYrvOofnLzhVzsmOfXxZGogmQ69QJa9vzibSbu3R
Bl/e7i0MmAbH42ndgfVvgj3eBpmoYplRWNa4BVYA/YS1Gn+z9RApebkd+2VJkhgAtm/4KUfTQ4n3
xZ8b7Mb48NhH/raeeNVcj8WbBu4x2SI25gDImqJjCWb6tg2YabrtFku/qWfZb3L22J3F555tfBSS
OKo3e6rtZYAhrg+My9MvrVsdLgnJY4w2x9yM8quKvVbPGqVdRh+e3JeAvSCFAYABCBu/DWO4Wn9B
FElXQ07Q3fAC3A4gw7ysRS7dtIrhuLKhZP0i8dq1XBAkbnAZwnkOCq7LSpvVBw6lRcTnsz9eXsHG
Ew1M45HNbP/FbMTcQVqutUopFHNQiszywCu3J/4sP74FYehalcY0jiygp+KXEUcBcOpxnI7EBAuF
3QG7+GaQs8FcfRkDM0DtQFCIh/KlcLEKez4aMja3WryB/dZXdvkjQsb/7/gCWi9yttTyJ6s9QdVW
wMqj982gcBZVTnRxd7ZZEXJLOYMn4EML6poQ3GzxLYlOcD6xfiPA3p8G+IGjPNKsiBY1E8nPMWmJ
eWgrBqwoEc4mcmWP6vEDuQqKRcxNvAo6f9skKtz2Q3sOMXyJ6xYCOxd6M7piMCr7wwLKFBmhshRY
pZTtfqC8w3wIuqrlubJahhCZYfQte30gbCr1pL36EbBJdxjJwPmTUZ8qk5FEXSxQ6zuxsU720biV
33RIliLSeeoM7TOLyuO28T+2sDz6bWIrIoqeLytfo5hYl7pSb27q4Y4jF2VV5/DD4zqxvmqbsh3G
x0FLW96V5A7SdlM91czue5XfNhz6Hm/fD18TteQrThdvlJw8beSC9z0WdW2Xn2BduXzI686bABiV
KX9JDGnTl1gH3VEmRg8rIZpVZSe4RIiq1c/mnFqjlQla/B1qGgUY0ws5DcNp4kUlBhvknk/lTU+5
o5JfwYeWQliibBf/rWBrfbdA+9UrajE0Cp3S/vPR7dnk5LFzwc9yT1Be8Uu6Brg8o6+sQ5B420ik
E0Q8a0tIL2WmMdmLrZAUc45lFQ7GCxQCEHbyxk85FnIjbsGXtkKx8/TC1v0gpyHmN8Ttq8OauvaP
emsfkJBhnzc5du0s3i2DrmWx6siYxsgQn1i87lN4MUME3qXC+XVkIpcWxjkk1ClEi1hNBbqvOY4j
iTA5dwKhE/jX0erBK7fYt5cPs6+8NpMr6yQ6HPV7NJGzqnDDthg/802ZOkK7I/+Qix0DGDtE2tIE
BGG0ISgAV1FHUTLn6FISwrSLkB+xWUSWBM7WDvZ3nqrziHipm4+BOO8xU3PeP42xPmH3ZComYK1w
//pMGQWObWoCTZOGeRTzXo2w0SGhMkrrLNQp8orx705Qwc4Qhu0IStdvTJgIB7kg6ozN/Vwj5+TP
N9BUVfSNSqNWWAiG3op0dAfJTeUf/iN5qaYvL1h+oCEI16R81GGkjxGEb9AAiVYZEQsSfoHWfH71
XOOSUPGnwZTqp0FcQ9FOV3LOSHgB+RM/5j3em5TqCqVEnERVRKEIzB3RiBIepSJ9i0314NUhJsOg
i7e5wLHzthQ3uyJeqIc9YiA2BdPTBIr0qvBYDdD7sErcSj6BWP5ysrQT1bnfyDEwvd2hgN5Iu1qO
KIwPu2e+yycl4k+WXfhhDvQQl/F921nuynPh9PYu2BD7o2nwTdxFq2GbbeywkI8MJpqotE1euOu9
zCyVQvRNtq4r+wZzzppiydm3lxZtev/A/t0hbkaXwz7aRiv9fgZ09TddHhLve/F7/8Uc1ZDSltLy
c2yBVJ8KRZtavMiUG09uPfbegak5Li1XdTYNK9cJdzA+TGrKI778yCfNObZEIEhiweyNzZ6Pu1BL
eUP4eKsjhlFmxy+RH9p9YABLHOtvB0ZSpoXEV0MFO4yflQnWV9FzhuoWHPRNGWwIcDSmI1UQdJ0N
StNmr79+waydFGQo4RNn99TcdSOPLDrlSeffTJ+Xw2IkI0WlWoLj4MyLLipv5ifGTscEJ90XDdv8
PJPC6dTiOQUFzPnge1wKkhLNp4GCdMorntWPRysHFTZDAdJyimacx9xUzaPYxQRD5TTLsJ5xrwqC
t8xLLNVba9mB+pAtnCptTcDTC0gs8nJeFyDzgBWJzPLajTdNCh7kBhW/CISbtwacx/TCSEsZp+py
L9CGIbI0kGDnmzrOkltg7oYt04M4tgAnqJlXJ7VwoLiJV56FSUz5byADOZ3oCOO4NpSr70JTSNWZ
2FzubmL4UIRDVBThuaxdIOCBdClaoQ1XHirEaKxf78QXPMI6aCCbyyRQcFrPs68AVxXIKKZuOD6F
/M0ERMyE7dxjHg/fIUUVH3H1E+WjYbMlyx0wgJh+WMcvuo/1X6BxXatKZA3dEwjHhclprQFylEON
FjQ/koSPreHlRudapkNBDLaO38FfEBlQzEkUjEAcrqLH9CYC3DVgLAQiC86nEhGBgFY9gXowVkKf
yybFqRopyaVAvpGtlL9naJkEK5szO3oHmMIUexjGRTq0e8OgUWZfsyRukhT57ijSHdnMwKYNTKu9
QlSx98mM32111mz+iZHcs3xYgB4T9Pb8w/SPt3Qw+yGJ1tOFfc3qbcM2zY5baUfUPPJbVX4l1wdX
/8YgAfjXa3qmDgU2HyhDpoTbhO9mkGWmTMR8QDFMZSI6/9eq62dsljsh1HV5zsTaVnXK58Am8s+m
OSoQKkTT7pEmeDa7xCy44vTHKUXdOAwqWBwgp06pf4wt3t8TgZhYNL+f43rMEL/7EhqjWJojgWKw
/PjFRsnV+ScCJA7iyCSW9n7XxH1e9jnIP/qUdzQau+IppkxQ5AxF3O4jhU1FHHdN242oLuByDerm
9R6qBjvgG/AOQFu/wCL/4QLArdMrtqRzGfRgnHJbqfvW9qUp+qI58pYoIkgzM5DPyhXl9DE6Z9Ui
+EZx6Z5sEqJQZF2D15Pf8efNLEtD26bTOE/ZWcbHhf9tvGtj9onSbalqWY4pvg3W15Q+lTI2YEzF
aRlZ9vdJ3DeOs6Xs45zMFDSsKzTQ9etfl7oeTkdGz08r67GxVB9l9jxJ69STTU0KpARTvUUX64Yu
8gtvRWIbZysNtfdH/Aqy8NqNfSTHXYlHwkQYrvHTnphuOmluELLFos49LlAvC75OkNM/7CNgVHGI
lP9sM11YV/z8zgjmlLWDR6FYo3oWLDjayMKnyjPXW1ozciQ8bRYB1VNs6phhGYRAuqJe14PTBQ3Q
Vyf5tYxSKJU8341oTJCf6vkG2x1JlZKWjAL1XWvWsSmDg+8yI2JgPJOag8EC+z0k/DOfy5C7CKDR
KAk9vy/b1z1t8fQSckDHp6546JeO79NcEf2rLY/5uzTIJdyG7Y89uKOLt2Ql3nUlf39YX+D+Umnr
1BcEIcwJl6AVWDT2dP3U2RL0DL+oIF5NX8/8X1gMpgbBBpisvTWoInSwoqORT95qGNOVgvDAA8NU
30zd2a28bSTygoP0COXgw6L/csTi8Wjx2FPihfn1MkiZE/weXGpolkXwhV9qtqgsXpiZMUv2MObh
oOle9MlKNdxr9wfmsjwPcy9aykoHrmgHd51AYcynjiZULvitwx/bJyTwOHqhvasK/yndNSzotLEp
MZPQ0mObPiyY0GJpdDXhVCeakKqChiMGX5dwIwvMnyTpKJnZs3DxaD0pF3BET9HQDSddPSzM4YbT
tazzycSTJAGho2pw4/joJCoPCe/G4eWY/zQwnpq4ZQLUt6+Hy8CARII6Oipxcs9FlMuLJvWLC8xq
3T9u4+uDEvMWIKBFjPue0/ineuWeh5PfFNnq29He1b+a/S0Fbqx1t3f6uQO+yMbP/2nGCu3MBE3S
ZcaJls8nRNemSbS25Sgav2+OsZXUy9/Urk7qJvdkVJetpLE9GPvyBFAMows3YR/t+LZ7AeBO/Zoe
SS7zAnBRLYgELgM+BJNMW6BO0ksUI444AlJO4JA1xowllqxXqw1BIxUPuQbh6KBjV73riOezdGdh
niMWKUAy4rlwODdjQie3DBfwqhNnm2gfOEndDkO71+SZ45FMQo78X/Ophz+B8jyIpTfXEgFLRfAX
QaGmMWB3X6HgHn/CjaDSkEIDTG9MKuOTRv+Kpzc7eotM7zEugkKrDaDwtadeW8wYh17SXdPBzjmP
9LNPyHfztJQZ3LF/Ze0vi30RiJXz/4dOYCi8gh9jCs6Zy1u7ZCS5P9/lvhv+gM4uCGTDmi79OkPc
KJsx0rxdrnWnDImAhpvvhQ17Cg9OjeBmMyKH4J5gO8jJEEJo0CSgp/yy0NbnwdJFQC80IdmbRhnl
Om8uT/NxlVP4y9Sjtnq0mLItrV8kwUB28Uu6vlRZDIORkXmbFbV9fsfTTh1JBwY5V08vcD5MnNg+
ccObss3xUl9w0lCAzBk5RyRhJ4aonykneTI45Rde2mSnBYTJo+aKNVfjgpJi/x87ij/Fb7zlpLcD
LWZ3E27eUFDmVnFe+lw4fTzdGwT31A4PaVQi9reAej5yxP19C+rFPvalyfTfRNLkjPb5hepb2yGn
kX3e3MT8KVpfLx95cw7gQbzoR3x+hqjTKQIWwHgOq2ojj6ph9EOSksgiAwhDOcFeVMYTTHyPVzKs
YnGNiUxfGYrytY+VxoP2esACJyB8UbemQSn7PdeEVlczFOHGnBoOsOTjvR7unN5OGFSXmouqNVx6
kR60MIJMWVoFslDl69FEVmROlwebn5ka+Rys0bsibRGJCSY7TCsPx5C+0YXIAR9JKgRv+xk16Vf1
R1amUu/5mzQWly3fP+iNLB+bRuBekqgwoqs5uZvFKXG38EpMdgAAA//MUYrrmSxOYpHi0qVyoR9c
T92teNGOIoUXduEYiBTLBbOfjp7Q/qwa0Of/cJ8NxgpeGl006MMoOCx5DdXorVPNIKBMW27UEBLj
hPsnX7CkPEks/qJ2kH4TNBN0Em6Afz/p2JG/fuGaWcmjzXrmjogWLrSbYugFMCofrEYh/+jEbx1v
7U29t3IJS4I2rjaljN+10UsvtHiwbLMNHC8NYpD5XiVNx+YZYR34yM7BV8kNG31/Dy4fHuSd+8Gz
VIDnKdh59iTc5PLIncXwOPfXAAyrn2T32seswJp8r5wDkmJSKe9Y0DI9F9VyZuKhgSNTW6D9v5zc
ElVB+2bbidAHlPwnA2KV56/VmkZXuJmLCtLy0tB4+qFdqAMa5So9BR1tEGgEcjaHMqNxEU35rRpn
LZKv02+rcDrS1etYhSf5Jiq6DSm5uzaDbfN/YW+BHsBJB21MBnt7TjrrxxEMELGTFXCKbJljCaph
0ZG29DptrVqWLfC329XpkUGQnL2m6V6Qg8Ncck/ZzuXxAGOFGCPhkIIIIvjNJ/Tg7tuj4Cmu0N1O
V38NlXiRJD1zH/z09iUUadBOqKcPnJRkbcKRZQPT2/bxO2bfTCfD+kKp/mg8Oysfu9BJoocNZRrV
reKYflfzNXDOCxGHMLULBVkAbq/Rqzig5w+imrOQ9DQKO70+bVUE5LWdn1H7H64G+OBrvWWqNIcI
ER4tuqd8rPfhRTKDymkY6ymi9ZNq8504KxaIx0ZJwfLcyXEj83Fwd2S2lxEdQNuaxdgRJw6dL+LV
EblrA2OyE/t6jD1g+4zy4OF/Mbad0aXSL2CsuTPeeK6UFMp1RcFMLqQbPFtAvJv/EZYIxP7t/ITi
Ex1WDbEShx6C37Uw24+/f2Hou+f4O4WrndE7k73RXfycs5duvlMySneOgwEAuuqf6aZlhwBJ4bPg
1kBiy87scTiZcCMiW2QiFTPPits2ASvg+eF6dgaxmtbvXTSO3Ycr7qAT9S8ZW3XWqwSIObT1MrXo
rQCtGcyRjlO3Ad5yoDmCv4nTbx2twPiSIqSovPl+7sexmvBUqfAm7YCdsdtVvls5XBr1Ry/MrABY
ky1S73ppPDqQJ0At968YbROovYczywJ5sHy63C6l1p0Lly5D5Yvce9bR5tcg4yaugB2XIrk2c7We
ee5NoWbsV/dR20JMXhCiDFKKE8akSkEfDDdNdasCPcIcfwZyByhuK9fVzHMZmTMVtDeT7yQFxdRb
gmYhT9xR0Lq9chOD4x6M0MaWVO0WYXzH8hgxnWNPcWHKWgzVcT4h4kSuvKM0KDp5RlugaGuYsBAJ
XbYv2EAvJhB9k9GuIYRY/hniu19ML+lk0uxUmjtTUXABN86WPs+1WPs5JlEtkQqfbBA8W0EkWvUe
qdwycc+NFrchG7dUdRjRHLeUTU7/Tz2i1B5+oAICkJTKe+8CR4rZp6JPWqS6NhwXjpbFVpaj1/OF
BfWcsWfgAuuXFhzxIyRBIwZiX1VhzwhThPuYykZaDSf4x2gcQFbfuOJ9GzyiHm65nkcJrBmVQd8H
00hLaMPrFiFLp+IWZQ5MFncCmXBvLId06Ysn7+q4Fu5BN2Dy7fMRQt9ZQTvJLq9zaX6XhA6i5BQV
OB0rihrPWASQG+31fsakfOUH/YbsMGQRbfDwCCEu8qmKKrFMkk6gpuvf94cZijM+MHPUnklfjTGu
Nuj6aLU1q4bg2lHXEuNtkRRe8Wl44ZSG+GMAHqTmtnCkK4tEee0mwYgtGgzg0TQemdj683HYVte1
avntyWv7Kitqtynmcyhc2f+BUwH/KMK+ffcSnCmlx5G+9tPb3ynsMiGwlcW9HhudEJ4TLBL1XS/a
aj0Cu/DKgc4sLnSryHbcbhMAE59g6d8zXnyK+sHHpbj6MqP2MnqLDl+ARGEHu96n5M47U4tqHDjt
TSRqIo3qf2NL31+SxgBGhwK0s/GcCPtfHWQZeXHFEDo3qmJrIIYZE5GfVJGOKvYJIFdaXuTzUl2A
2lItgLeYeaDQHwSZktX+D4oOIWO1J2ITk2OINq3dzt66pGJLZkvNPkUJlDYbSe8FDyjOwE6cls/9
H5L/EooOgRQhy5oyD18DyhVsQZ+91ai5XUxd2XKbC70Qxtd+DSIXlcSrnHVNLyHG4zloXpc8f/b7
YEqZ4nU9oyPo8Il7Q1+3ynPeCyH+8zxTvDS8CmMmaNGqqoyiv4MSopdaBia7DDvURHoeAeY6rq+b
8QCBcHDWeGyu83LI7H3KyC78lXafUtcPVNphlYEsY68Ft7ParRLip/X1GtBTO2h/TdPohY3PgUKs
pvo/ptubVmmmx3WVg0Y4ZlSwdvX1Jw+gVv3Wd7h8MqTHdi7VnzYRgtkG2lKG3aSbMKretZiZ2blO
zE94W42FsIgt9Q65+ob6l5JyVyDzBfZZc8Pd9plG2YAIJcmp+rqgHzR4wzv38WiPKdjlOqzu08g6
S+r1J2/jvIKK39WLCtaFINMBbG0307W3KDaHXSH8GV/qBx9W9T6m5p+RpNx77Z6S+C56jZijT24D
Puhj5sqIlEk2T2+nTY3vLKcGSSHabiueoG/Ud6UVF99pen4wZlNe8ZoVR65tLU7Oufqp49QGzvr5
uWfaky4yza76Yw6jx385QNyWNF5cZEYmJewWTSP08CDdmf8AE/Unvw7xHNL+EAgORBTepsBZIofg
C+tDncIdypg/c4+1UFNJhOwxrNDXniWC99cuhTqCOZiA1MTSHDH+Q7RHd//S+fTmt8q/g4LOpQTC
zQS8XaredSgvRZQ5SDsL2SJxgZlpkdoJb/UT0VUX0AYylpnvdqRZ+MpaPGxLHkpEjmMdk4JCvFN/
F5RS7GsaVI4Cu/IXT1OgmzOH/jM+ug+3Sm+cG2u0QKhQjnPZjtBLoVagga+UcNwV5j9XRJqaZkxP
wrIFO8Qx1d/BZlXVTATllDcJsEr74PxBGe7i1mWLyaSWEj7rjnZ17RjE4EpJchiGofvBeuOIg27o
8xJBqq9I+KBe318YOS54OGn4tMMGaOikMSU7Sm5B8sZl44Wb8Bx88CfGDA5Knw6a9PsC8ixwIk/C
i0vG5pckJxLlMBkU2BQeoI4DPtmHfvMvXWKP5ZKFwELfZT92F36JkzskLe8FAIFWP3pn6OrpF56p
moH+o5puiwD/A6ERw1Wk/lRUi2BZjGbxnMioEeXzW9doDc8FlPq11frDjo3qkwyGuzRx/2TRG4PA
spJ9SYK61k5lH3xExMlFGqoIvPr8Dsf7JYupTh+brnfpMHMyBizr1prmRhxKBKziJsd+i23h1Z6Z
2cZex6xiq3Ay3AaHG+NPqprf8OweVxH+NIjIqVWQQv5O9Q4oglCWHHd6hHaqFawaLuZKMU7b3LEP
nie8TmSB52aTQso0xfVokrPhHo7E6nIYdiHhNCbNIDL7vMyhoaDg9G+xr68JIA5SdytCsOmwsh/V
vAYcs7PoXLT4DRzXRO9gbXLB0oBOCK7Zp5tAaVdu264WwWOikT+OWrcGG0tWjJIVRlwSETN1E7Ir
K900L0L/pYQcSin0CKiFc7u5mpuQYZHl7vWblAZUV3FryhmxyVNywQn8GJ65DGU8ekMT+oARgLnM
up1LfdC0aZ+B9w5lvgGyrHDp12GXIGe7Tm8rlfnpy7ZbfNbLv7/k+CyuGiTPmBL2HuX/19VjFCzY
pBJV8YU7tK9xoBHmiLs2SkxAzCmWpdbtoK1NcyMNfT3vvvEmQPtT7gN6LpRdzQkTH+bVx9aG7uKx
dnnIBnoEGr/dHL6A4Jh7/SVvTgpozS8dlj89QlSBo0FeswrlAdlO3dgoeHWQ3lEYlO1b1BD+Wfp0
vfkrBgwyUNeAyAfgqwHH4xweq6NqrPxCAPlF7+RY5eDs6k0BFY73HZgEvVR6s9B/tvjsCfENseTb
8apCP98A7JF52Jqlexg80dylquxQ28zkWE4mbSpwbEpKnKohe6i1uzw+0VvU7ZBoDdKEGKn5mwRQ
P+WP5octFpl1FRtpyyZ/LKIBXmy7KITTX2cy2wnShaLHY+P1QIlSG49w7KYDfNxh/GKQqumLez5r
6zNb8SiUzimeIAO+b8VSsKue4NgHKsT1hYzGm8fFiz0pGcIPVLNjUIFJdstXHPX8OPIsVgdSlhYy
vCKq4eLJLUv0qsfSk1S8vH+UCo7C1w56VDd/m+n3dJmROqw/7l5qmv+FrwgwoRwSlzK2tGubdqSF
sx4qgVeZXy5Lg4va/LpgO2TTsdfTXR0w7CbADf1TMVFwHTsQY2wxUgdYoe5PS+Nf1Qlna3mDQ5UD
Dz1bGDCNyX6quOGqQ4bNiXRLBQQaRZdeXuUgM8hL4HAu/CNvjNf5Vvr+WDTdG8judaRZ+1EZvZsv
24YC0M5LGimi9HqIiEdKowlRhZLkLAwQ0N8b98zsInY60B3t1nYNpGMIqxGoCgGwLJXFoNQEU2aB
JHcxarT2++N4l5Sg11NExL0FVooCB3xVnUqSZGAVR+hwhSCJk3GHTDMCA1Aj/c9sPApqiEQylZJq
oPM98oHWhxUDW54WMYukEo6/igoktNOa2thnZNJ0scQbouKRx7OOhiXmfpttQkAPGilCvPoNXUVU
BxEhpFoQe11i3T6jAfL/AkeVz2Ed+5qEQ8yCn2FlT9/HNfbXQHPWVDu6Y41DamcqVWiKdo30FXdb
8PUFLFyKVafSo8ZRbwLGfwtLo2AF3iDYne+yo2XMEH6yE+hSdtmlNgphxRG7tmPYwl0q4ZMBYbi3
1LoYGJ4Muu5Dt1+j57xHOVxgPk9z3HGnFC5rKFC5XUF1FmCYW9Nhdhj52GZSerdcy+eFgbscEPaZ
hc8YlaCKvoNSwSXOssnYHI05mM0C8bwT2YhhJqMgTbAFWF90VSZRE8CemXvDJ/Iep7P3SAMkMNZc
Ti0rGDSI/5B94mDseILPn5NIs2VSQ5fv4EJvauxKB4+dm59RlnAaYrXSYoau17Z2TNEYS73euLdU
KbY6AvBFHtY7rNkyUD7zrWpdCiEe5umI1yoxqUdMHZpPhb55fR4X+Ff36lHePkBSqkSiSCLMdxbT
Aig7O7NgKVy24yK0fd4/bB+B3Dxe0cj3oy+uIGXliYSD0jc4MK3u95mWys6V+jziH4gYeXgBXsPk
i4JoLWheCHXF16IQ4IjktoSRyETMRybzldARFCKKqXW1ytCxrF/VDGJYN0VkjMJZ/xLYT8PMQ7SA
31Z3RowggJBcJZgZknuyuKTcRJNLTh1ZZUFZeyHiM+lyAxGOqTylX3Qo/eXgpwF7ksp/wdQ4MSwC
UBOEkT0W4K44GwRNCdDWZFW5pHYoXGJHamuGRQr7ybKkd5fu2NmaXg7O15IdfcviKOm4rYhx4M0j
bQ8op4zSybcjqfiNXFyFv/eqEVXt4UNVZpBK0moDTnRvtwM2oUQa+zVr700JBqLA2sARRhluDMlb
h6wQAhMN9Klsd4hc8gBQcjPYtX1fpXd/4ioK59YvOwUBv+IyHSGcLBzrBdGoZUmY/2xZfmM7KFgd
WCod1fzSmTYCgXADogF8z3T2PMvnGTUZr760vwShWmyqp92GPbiCNJbsjPiu2TthKJOYOT4j3mFn
qzI+lEtQUVquXURQGwRyAhfwmkBZAyIbuwZuoqoSXFVxYpEDAoNIMOG3M9ZDIIUcsdjgDriZ9uEb
+fXJk8Cm92jykgrbcf7SpDEL/nH4k8eOmSOhG9NJZW8qCY6lvaCGEfbzCs44IbQRYlpijWSzKocq
r1NF/0Py9/VuIsvpFgMnncmiN9VuEEyFljuKOHpPrgbBxO0EnRiANf/5vb89m9inOj4nVPP6wUO8
jTct4xEH71glo92oDJqWRDQFToVyd/ZFtaJoxZKEOXjzTsIBBjTX9kO9Sk58Y8D0n3g3J3I1tgfP
oZfsoPxid5OUXxXqx8AXV+3HJTX340TF2sxN5jW/tf7OKDNXKMBvl80pnM+t49V+dSbPZARVL2bg
mRyqfqUaqq413ovgvF+BRA+XeRNYu2ULnYTAA4cMh+vN4HnFE0i2/P5qo4nCAf7g8ejEg5UR/Z8E
l6C/uXkkMpim4Ev9GUX6QgeMnhM3FTdSeblMj5INVS73Eii5AeNvYeAxc0ruUVilwx8QpyTgdMPH
CpPtTxL//2MwODTh39JLgJdDLGSOo3lahZ7pzybZ2m2cRYCw5rV+EjuGjpFBPTJW36K+LnWMw5Yj
A9dDnrPmmTVWKNSng5eSnIYThUTSI0RXNUWnx3DFFXaSJJfMfy9x3EjAFWWk1oSdihJrZ7BnkvY4
7k82lRvSx/PCMaUu5GFL4oIC7DfqEesiwupRvbjsLmuolp4CgYHstaU1gn254u5ovFKEwJU2Qxov
xbu7SLXxs/5cU6rrGasIQc3C149FL+qFiASRFghSantV4hLIYLX+FYZmgwo2o8VIOW62e5ha9Bz0
ZT6Yl+Wa/xfinyihF936qSHnjAUUdpZhaBVPGu9bXc84Nb2J9h3a6ayCfeV5uZXM82MaLzTyjZ7d
XQzJ9Ua1gs5czPqXc+iKtCQv1dvuc0oxL7F/tuD5ObDx7SRpIycNwh7pBQeG8lzkUR4tMiz9mJtD
LYSF9y/sEYNvTUXzLTGmdpHqSU+ETWlPnUexwZ0RcNs1cfBIGLaLNl7GU6QCs/KOlCTK24S7QJWV
xJxbbMwhYU/va6iY0BTPy7Hwbzmk3p4BNS4Hf66ZmDo7ZUhJi+KP5gw2Xy+/pe7OVxeiT2w3pNgn
0bGZgu8q+66d0Zpwg0029uEYT5AjbHaTDgPKSbMAyTc1V3FX0B8vpXSS6JrqR6VhnLSZkdACMsh4
5tYCX0DeDVjrZDb7JB5l03hCJkShVUe7MeThSGwLBObfLE0TvGNhs8dXf2CpqxYRL4RW4UrOXjHF
iJJSI1APAc38kXWEr+YXQikERw4D/f7EROXxSji8O7cvmN+57UeeP+AJkyXx41HAO2HteuuEYIjw
79gH5ZsYZfcGwNwmNYOXmyQgw+89mfSmIL88e1BYtUtMyrZsEbpjQrsNtz+Q+QdNWdDPEkRyPmo1
4HjupdVsNC12QivMr5az8mBuqBBHdnq9zpAlK2ukCZmNt55/tCk5EvmTOMrqZ6VK97KCVYJuUfbH
M84FFFuaM749U1YGXVkpkGBZUqh9XkaXMs9NqvC2v4Za/aHeqHv8OKjrCdsw8MYsMVffVRmWtKHp
GO17gj/GlxOkr+RCz/hi20iz/owUzrw0gflAZKL1BHo2m1kuQPD6h5rb538i+D1kqarkrMvaCIj1
xxnEi6OrFa17AncTAnAydBj9MPb/wevGXAgOLc+nYPcS7GJ8QC6vosF4w6EYPXFC25ZGRq1qw9Cn
ye6OOaENs1Sh9BXNe1fclGIaBaZCNJMZ2eCJPD5OGou8up5XkbVZgY+YOMvzRGgR4Yj0s2JXkmhR
NXdoVG5g78S6Co/AKbWz/SiMbn9djKIxaGS7va/+efB0icpdoF8Q1H6guz3xN/OP7kosZqc2qhir
8Jo0228tRDUcVL9StI9Sp/TRHU+fmPSkcagI4nhGfQ/gOqswq3rW3VHAjSloD4kgeIc53WtwZ+fV
KxGh0EI/WbeMWc4oc+ldegnXYx6AeX2iwWytJtqeS1IeCidu1gM/Ovv7DC9vvmTv0iLs23lxvkPg
2Fhb2Ip+mt8hJ2U2oNaFvkHpHgSIMOTWJheiRibWx5cOYXKOs4jo2dqnPbGfTA1fZIInF42Hdcyp
vYZSeFkztQFJeMMmNEaNlS/mFFnPyXqeRTKbPRWWj1q3nOnKYHrABfOti1O6bqcyYfaXEPYH2H02
ZaYLBWhjE9ixtVd+8LkUG0RySGr0mq8Jdf+TdNKGy6zA0OFzkFz6kEWWYa3bOA+g5HsXX4cm3q5i
5IQzr8TVRLScATgNaUbEF+cytFe0K5c0sZukVkbP9358K3N2F/SRzp5Qtd6FuGfU0yy++o6Qv67e
/CP3C/I+y1MQahulkQ/m06KWLbW8ekQ9yxpjARZZ+56nGimEU3YYtTKrDmj/SK6Aa5E9fbbHLXMs
qfzuhiSkn6xo5UC0mNpA3J09g5j6AXBhZ/4YTurO47LouhnVoY6J0b9KkefB1g4d7SlhkyGXxeka
IKgS7u8ccd7OFh7NYZlNM/uF24aZeBaF6adiuY9ku6jqIlDSBT8YfVGOdtS//Hs+eiE/zR1b4k1R
2wMdjLxR3DhHfrdiD8a08BlwOINaCOmUBswhK2quTM9Bi16g9PGyZgLKAqF4MM0LoD28lLr8IAU8
g54NHcGaQOAop/WybfNtxU9/ipWvkxCnoWhRE2pEcbtlFYJI6O1TOlU3fH/pwDVl5rpuBT89DCe5
OHaPXddtnGwR+gHU/5RL8xJNdxUl2vJEULhWH2oH0Aere5oz4oTKmp1U37FzHAQFkPVJKsrgmHgq
JTkgJGF2W/R+iVzOBmUXXREt4qwh4WjPZfyOQijiM2rbZCfgqZU1hqq6TEP6ptj58FBboFYfnxyI
vJ0NrZc/YLL1JxH7o/xSso0iM/CmB+msGm4NtKNB7/jN0vezMfDKexvnQnrmQL4gE6RitCTCuwTW
itiWvlGO4Wqt5xliTvKWgEUpgQglnB+7n++pTPyIP+y3clcPdk6AuGqsh4KAkLI/LjBbG3RhPn6H
0+zt5hs5cuKZhN3IBQ3K/+7rSB2RwZJBRtTpp6B9cN/X0b0qwx5LszsBhD3mSiL38JHd7MIfDsA3
+Au+rKZ9zG7r571KvoRCppsJebR9zUu1z3E7kYXV1LGiy9TrJPgNcw4cofI7qnjf7SG2T+qlfnBk
FEqD8ZmtAQg8a6CwPsJTJGf1jU92DvToFRTlQFdFnlakM2zyhVrAamdmsA711tkexEWPD0LcdS2F
+2H1JtaEs79wNUdf4AAJpkAmNAtcaiJmrrbkrvcdsT67fR14tnocA9ZLf5oumM10YzV2Y84tJhP8
6/Kdresgmp7hL45zyCVyFNxinqTg2IHT3oRLTBqDAjHnNcno8MRZI6xisyz0xstUvQj+64SAXrRZ
O4Zc2jZioyjLyznwKXPdNlTBgPC0ADO7VGvhrPo4U4sSRpaKcwSFBpum7L0c1ru9s0zp+nHJdI10
wQy3AGhEqS2hz/VDTS6O83oXeFCEFiSw9sifm8EAq08INi/aandt0apvyigHLjfOGhalyCPGj2RO
+5oQuQhk9MHo5956D2oNfywwTkY9gaPAPnTfD1DvgCrBNf6/pQ8PaFI2a0leqgIkkGC3UqQWjfxD
FfLCrVekaMVYNJSDHtmZvJ2zPoOG7oz/5t9T9GcRfYXsj9Iq4Ghwhc24nGCq1y+28BI8xhmXBIDb
uaD/jpJ7O0XFiZeLRvMksHH1p1YgT87R2ei6vvaBa7uY/DNinmgepLS9Ds22sf+auP2IqsqPquRv
VYUFLO6RkU6qF0UMTJgSODiLRy4QTh6Dt0EIeLkpI6FQTyezO0E+ktnNV7NP7foaMQN2ls3WfoSz
uQCy8OSzDOBB73G09cu6uoSeKS3Hc3X/RTptFsu7zMOi9R8f2LTVSdDcJ9FeZ2d5o4Lg3rXFLqSS
c24LR1Y80WylXgqfSW7sD89ausUKc092bGNHED4GUVt0yvfvwoBod611L1CnE8qtk2bqUl1/Xx2L
gPA8v7xCqYkzK6yFxFeSa5G6Q5s/4y9tJNtWINU39e0ZYA9kdxoRccx4Ys18LdIsXll9wTxVKcn/
oue/sHr5JrWEdtSFFi0wiE0v8/BCqxVfr9XULMosxtyE6rT4oax/4r8qj7BN6lC95qpRc8GPJmaQ
/fI6UKG9x39W7dqgjFeKfAg955nYXdDSSkHI3g/fUjpKU0W7vCbHlxKX3qGYRAftkKvS9pierhoN
tLPfZwfI92JUxrvhK5DA2hSaAQ1UTPd4wyNuHxKf/XyNSNHlSoAUEUtZcGdRnps9L5Qm218D9MnI
/eVJNIZfeOsIW8Ww1dZoBUkTfxVSIUqFhPSWvuY6V6wBLV0wruCVb6Mzc35+vGSGA1v3j/czBw8f
iAU7W4Fj0GOgNxYidEg+cMsGAtxZokIu1L2boXr86vtLxb4oCfhwGmv78blaa3qN/MFVPdvtefMr
qoFeHXnwGTOMBIOWTddYMa7xWUM024M3HnM1Ury/ycSWvYpI3uxIk1x5Fip+JbTeSPkm9Do37d17
gvUGcOV5WCAVF/pFiAzDHtAamMJx5PNvYvezBELe5aQ0L8ypebW3RWkEhncCrAMqS3M3pE0sy9DJ
AHrkP17FYr4bf/1D8hEUWx3clH1KF/eOr/CNvkmi6lKaehGWG1q51CgPDoCjWR6+cUTJjcWsnnkX
ak3H0ZZeK3LqTRVo4oB6Letel6RECBcBx1WWXm3HUzN4R1zZBUhSyfBpkKQbYVG8p1UzgmLq5jpF
UGoaS46/sfax9q/Fsq66omiRrp33UqgyqN5z5oLziTyD40iUI4YPXuzflqqd2mEp2N978Qh8dDGU
dNirwJNZaGuG9ChaswZtY3/hqp8CG60nFInsCgzS3m7gYabdv6WMZO0rnfViQ9cPgHZ66ada3+wV
l8bp0TUBMbNZRncaIEAQfQNuhnuq5I4zUkT/iTgM4dR3uF1cWLCqHgNGvhLsbvoezRPjZvRmSuBY
G3pxqedYHJecnFZhuHSdYs3SAKbnKKROqCSRFPKEWCP6u4BN/rWgQElJFFL8DgL3AgoMs1ZW+dm6
6q/yA3VNkhhL4yrt+NM3D7yVNWsNwN0rv2wMmOtAyRw3qnm9VtVpDW8QapdlKDEs19rj6IIG3+LB
SRV2EUOpcXC7n/MKaAAcmSd3zytU4lr2dcd77Sn2Ks5pTS5CzLoaURzUoHwLN8CCGCmaYhIrBnbv
qJQ67NBIDY6I0rVKg9jg2tMWSPamAcgwm3Y2z/ozLc/SHK0/quv3K5M6InxH108eJxp7lj6pamTc
02woDEjULQAFIKZofo7+hWtatNRI4JOvvfyfWUIzxoV9Dym9PJHMKoO81mUYmIlSMYJ2fBrLhlAx
m0nItCZVNM25D7E8I20Z1vBN+Hi5MKcEZCLjaG5Qe8toUb/RA2UiFKHTY+LXGUdgyjeHkUgpEjnc
eXfvyqkkjh9BoMus/RVD4MPb//15dkxv5H+TVhKPLOOdRbXzkK6kllsarot4y/nqGayQj9VVaQTH
S9lJFWeiaslRTsCIfvLf6rJQBSuNepFm8jkQsV5GJ3XgdE4/1/w621Tc/ZaUyOKJlmxC8MnVtHkD
ICNKioG6GoJb0E6fnFKTrjFVCF1kPQ2flo0sl7H04lkTeOnkZLxOFqhGBaDU34yQN8Kh2pXncGKE
19j1eGV2WM/N5ryIOIvz0ra8MgCiwalwB+BI/9DUsEDMAJsQUt0GrOCJLz2ZAiSbaX6C/J1o7+TC
vWJQjTW8aUaIascBbBA3aJ67hGjAX4ApiRKMlR4wom6uTp7vkm1rgKRrHxvyaokkTCepOF5TkCgH
jjmx9SVzCyS5UXBKvOc1fnSk8xwOTsXZxmKT7ugrFQNnkv9CIhy9iP4u71CdUXxSAU+E2ubMeGaL
uKAk/I03eEvyEXax4cLCrlppI+1t6NmZly05HLYElRIzpojDH+qILbekeS9VeG/9OreHsP9GYvZK
EcG5x0uKW2ct7Kzr6PtXQ7Rd4elULcUSGvjhxf3pPf5g2gPYK5GnAplFAa2T5qM71bTdQW2aWFjT
omoSq3HX6glsbycsogaRKiIsF2Uj5o4PlWOmIaRZhcKTIOjypaBmv32n+aZrjkSLkP5nzQWvv54X
ASJhIswXN+rYxeMvXE71zrsieURjvzoZETmJolAaG7X8uRRxPVF/GecuVlYwgTOlItWu415ODqo+
mc2dEdLyBvmuWTgOPy56bbjXE34vgbsasKAvFTDUzpsQjpjwdR8XZPN1OWnuM6sxvUPQXFG3L/0t
yLKG4QtvH1cP6JjjPLWc2cC3WqwuNUFgsodj4DE3JMC9wYnHqQcyf1TPruO1VVkqWV6IceAQX4Id
xmzspCopQdXXhIuNfG5riywh6KST/3qc2DTnlQrMZ8hjFJ7cofbVbk5qAvbLKvYB+FjOei/ecpQe
f2rFyqaKyz2p4QN1YgpxKwL5iaoG+ol7/IXiAgipjHzdsDz1gIrqDB8LzYwZPTVHH9XlwJ0elnAf
M3O3vArYcj19da598oQNQcEt52R0ewY34tqA88sW3XJsGfL5McJLc6Q7hWVC51x6Ok87Pr52nA4E
PpBElRF61nrPHm5gJvNekBR7pY/bRQ8XTLqgNuGS0kmc9FfCi3zCos6isNBmG87U32mEnO1mSaSY
wRpUwcoAZFZjJgDj9ACyl7ixg267zb0dMWFarfV5EgfU22VoMnKulfuQuzzsE79oDUDSCfADOXsA
8L3TR+O+Q0KRJEHq2fmyXFPjBjvcEuu8/gRqnK9mHAAUuCg0to4qITRqkyxUOyx2+9L38THC0jYa
Fbjt/RxbBmsqyFmWpNk4gEiNhPFNWdtB35dz3KNKfsXKRBxEhdlJxRS2SVgT07mwgv9VEBB7ucxR
05LjfRN+Tq5hLi92LQAd6B+xVgj8LZPL3CV2Qp62NZfqhRaTvXW3F2yLUUGEhieZByuCZfO0/Ppy
3B9sOYgj789knk5KaMQfRuPNjkid4J6V5Qnd+HNrkQFBnGQRLkI21RaRQP6yPAScSS1cRMvDQnaD
3a+5jP9G3x3xvVp3vJVQrYbn+XRGZa7kv6oiQ9EpqdGU8amGUxu4BY1V0aJ+IfIKTAfk3CbFhay+
/CG5b0p4MbvLLp4L5pILpmzsTvi6vLjOwo/G4hitC8xVmZP2cr4MOoCFY8k01fQo3XD904S8OD1Q
fjoeyosHZ3MV6nAVrd5KCZWame5f79Eqy4AdniFJ+ZLyUnDWBznX3OZqGL2tfKaAimjx9bDGtRet
esIq1EiNOY86R1bEpMhLTDLcGJ0q4i+KtmTZmvRBXlAKwPeG12qA/8V09+QmK/OoMaDDs/veK2l1
1Nvop3do6kgdNJMWijK6GrONQsMBjCU5ZqVIrXlxf5JirTeH2e/QMDtg94ysLx/8KmmYKLWUyTxw
ZwKLOozUOKLXW0b1C/RlLEk0AIWMKsZO6GAB7G/07286sm6edjiwdc4DCRp/z96rnEIO72JdFbce
YehxmgaLv85mYrOta9vxtbKuVTtEIBfiq+/DcgP11tYb6XSbgEW55CpsjcjwSatMpPlEkdmlnL1m
5wGvwpC3PbipHHHL4d04QcsTlNH1FPBQjgVKiPw824dLa81npmZeoCyqUtiacLlpaUGXmeyheyTH
3l7VKvcGb2kBr0XyX/g9UEZzz7k5oBSFgsyiBlwHNrPlWtBnEQcc2Dz4TKGaqvlE7JiNl3AmqkZM
7K17kZaRo5+vwXfBLDw0nZ5x77q9sOozsnFXqEzl//VdMNCN9J7Kw+FkT5DQCichC2bhw8a/MyAJ
otEqJNevO92wp97Vri85ahXVPvfmoNDbhS5jflItQKx0/5uC7PL938GBMRpxZl6izYoh5y3ZRC+k
ZGQSQPYP11MhjspH9Mv3HIYiK6qWclP2nEwqs/nqGOcUnuc2dtyaBtkuT7PRXwPhpVscIVCNuFEz
i7XekaLlQKdxfmxqBJBlPYHJDp0NG3EvUE43xY9BobIUZBarQPO173bJ7k0dXCxxxhxVleYlB8BX
E9skrRmVo88jpNbDcWBffrYANjoBjvbfkNLTbobl/e3vqGppRtQ/qCtyYn8FIUbMZ3chZNSv9Uxg
n4T/ThEA87uWie/XsFjCuiVdQdEIgyQy7rKwVsHdd0HhXJxSVkILv/k46zWAzrnYZOFtLAWByRTW
EfzRLHPEgQz35VSip3duHzXHmGsEn2wX/1PKW+d5FIpFAnvYgN6St0Vx89YLJqeR4KyH4tA2aDYL
7Drk9lOvHJ/VN8yTqadtrjLGADcZVSiReWNcfWJlbekjNCvTEkGr31uBCX/KuA5NVEosFSBlptSo
v/p7HavQ59s6JRYLq0pikBMtxersCoZkDABZuzmVnaRhGgKjgmbDAlqWPWg64KiTJxMyksIxGLhO
W65iq5zt0safDKhTkpKdLqzIp3YAY+cdP8lLHfMHB/vz53sjRXZ1odnbBCJmsoJbsc0SLL+Zq/xr
yCHZVfP3PKQCQNTSGeaf56aes9cwXFHR/WQS8Rp45xXoffC5qvK7nZ0MeHg0HUwG4uG+xOvFezZ7
CUO/AD62BTuwG16TiCt3B7QuCNS+33CZUM3+B+x6e9noH/iPiQUKkkV4PvbIT++q++5e2OuF9N04
vUo4RlzdC07L3IU7qV0SpByQ+1+vphnE1b+UupHFZmPFR3yFlfANjCBOhIlw1BTaSQuR4Fl8Jr1G
763Wkn1xAkk0LTLzbnSoxkFR+jhRv5g1QZplx/c9hf4kBHGp7Lt9cysDeqoYfmpu8JWwo/0Y9bnE
HDNCAo44IBWuTkGrn6h+rvDKSRFUrkkiJE1gqxGd8m+QrAd406v39egLH/YkOlvrrhyfO3YcX84g
pfL0AgmzmK+9UJ394nznew86nr3Gmd7qp15H4+lgYYDpgfZXB2zdVeqjZ0V2JEPMQNAMfTat+lr+
wLxwPpYLqa7106lvL4BH7tCsWim+hAJkG+UCvIQMQR9aba2B2zNO9mY3EkUMIPzaNGe32R6F+h7S
2lUuPZzzi5VS1BP+JxfxIdP7TbMamBnCjR2GVtQWD/rIs2a0RTFGSfymvF+KCcgoi7480od5lVdm
jhSIwyyQtIsUJthacM/jjYPfGP4+lRnO3NwU23GWxQM4l3kinXfCQKOMWj60o9+RCmMxyWII/3Fw
aHd9SK8ZMSyQrMed1L+bg/GCPAz+DkzTPoTM2661q78l/d8Ow/cR/8koP7lUyUZvbpsGwS4FAv3k
poRgAGggmVt7wVHpNFyp7j+6jbxqydJuvmiNJ+EkdsxNlkqwsIBtTlj63ChIc3Qol5D858Z0HV0K
+P4gKo5EJJePeNAAl/ydZugWX+tUjbFxS76g7RtJOgrpFUDX+RdCxxMf0BjwjuJlGZFLejspdLps
5Qcj1x35SGoflOobuGoYCqKhTZDEZioP/s2bzxyCYOKx9X+BcIsCzh6eYoWuwP+0Af029t9LAkDI
FI5eL7Cjd6GLt8DCEzxA5o8HuXbyl9QTZc4iGFJ05FL5QAUJz0+ZDo4Uo/SbSd6Nd1fdlOx0nrwZ
zWrae93IM7qdxw2ay19sg71eqAjL7oWtYvSkHpf+8bHnwbl9WTYbTARI0iwEw78tTY6/jPgaS8jq
i3Bvg7k9qKjXLcSoHgKqdfAqGQsgjeDgd74WAhilIzFrW2pkI+c6yDu+HP18nG5q0mr+ttBlmeoX
aNI1JFNuCoXoSOBuGIaWRs285oEw1RrERkXy2PQDnaX6B6iYliI8uSPYzZq7/kSolU8V1t9TTnhG
seNSRSjnPWGpSdvKJxRQkgnMqxGIm3GtNTnolW8WWsm7ko8444JZ4FurGdeIb9VRZkozRD9qQQ1Y
+j5D51urql7UWFNFhoNg4/PUB7AfPf0UNbQxPKvHS84mXYOFxZC+KKfpfGmPk5FeNaxuh0WfkIcN
PDOIPQauWLCqB8c7buxCbjm261iKQz5pY67sN1XUGoLRfnr4jaRlldW7KTd5swYd8LmlDTwhunTN
Gq1+l9PDS1EY/fzBxzHG948UXtOSUCvvl4jLZhpesj2OivCH1txUahqayiLJzQ4pBW5EbZkjykpR
VTTqvygsSRnKwG8Sex+FQltyp6nI3UfJFBEWYef6ZpmETzV9QCxMItt59CqC3Pj44Otf7YnGzbX6
K65nfxOfg30SUTY1uqprlK7BRYC0+XlDnYU9feTOuxNutOuHsThpLazvhNUv7JhizLI14LskoLs9
DYRUf6VcnBiAyEdIcr6f1SgJfmjmEnihU+MbemNElDbrJCthLSZzW+suGlXI3L50M4Lksv6FRQJ5
1vZx3UZ+ph0U6Ssq0crMYLBxIyRwj0WQp5c7pXLHFGzzJTlo26uQbZI2GownNNZOPhpqez4LzVul
EDXNdKQIs2/GB+TLML53aQxN4s4MxDUAZJXeTag5fCY1AJ/+Xc96EVyFgDzlQsCryoVMUkl/gK+f
G1SQ9IZXpiMiWFcxrjLuqriWyhTyavhtp6YqLLVwTLg2mW7xd3fpWgqNvLrTnJLmDSXamvHzYCcs
R500gBDbRzLMhiWj6rYdYO7QcC3utOVTUUzXJdUqrcd2fTtiTGQB0b/B1LUqIQLiQbnNeOA7YS/t
rpTiHomx+jGP9LDLtAGZEyXZ42ySFSqtWLSVFdJWJ1/2b0OyfzN2V44vLcmndbO34JcdSVPL/8CG
eyqhifqwgLKW1qb6ts+mmCDb27b+tddlLxquk1jO5FkcFA00nQMO70MNRoxF7qeH+RACIxmBc45F
zvlqM0zQX5Zfpc9PRGzE5GE2qOvkBcVIGNkgChoc8Ig6Qzt86fZJ6Gg5NiQw/P7VPO8nkyIjmjuG
5gCSWRSdvkqxLBlQMy1Gf4CgBvfhxPvZKAbCJWLz8At2UCE21j+izfATHY9ZG7BLCA577xGZWgzJ
cf5KgalO7ye5A2q0FZGaVOyfDg36PByxvvH4rtlBL+UT9wNFM2F4ZeMGnPBNy+6ory9Mp3PDhSsK
JmrtqEeD0KOj8Q3d0knwE7BqLLbS17obTKmWJIvOXcFJe08bDiyWd7mVqNdc2iVgnMjX2AY51aEz
j5QwkOyiMRbEKqA057b1dxtpSpDw9sHxP2q5PbDViPfN5DACZmD6L8vHWqhTHZA6JEmW/k+b+XJI
FMCBtr0JHEn8fHu6fgaD9FM13cv/LuiogiaePjOfXTN8hCTAMMe6GORAbSgFWo9nTst2ssQJB2ca
pIGaoy1mJjiPdc7iscUmDmlu2h6OXqynvN/HdNVoFabfdAT/XD7tKfA1U8agScFbnHuQUesbKvvj
HJk5T0ZCmuzk6RZ/icaVVabr/HuHIxoLMIPoPqeBGsSHE+zEE0PHqhENJltvgnufRc0JijDz0cE8
GdQX5U8nezrD/SlTnf8Hs4iaYlkDwtJo7T1DSw5rFNZZtATdDBsaiJn0Qnns0jZqwfCGfVsCbdvY
+A+mlU0HkXh6dq7p/aOqr6WXQw6DJWUR+LCNgvFh3GAlV23T/7NWSGyzzFrhAOAjsPk7mlAlfXyc
JkMinPtcIl/lX22n61aZ4M5q76FF9j3s5UhAxO2hMLkc/K0n92irRI0z/9CkGXXFNjgsMc2dA5p4
cA/370h+ToVaT3HBgJKKsMPPBLw2ACCkFPstTk/1nq3thbp5NjEyL71EuEFOh6yI0/IVHAQ+D+3h
Hxc2UmhlZ2k+alh4vNzpNUNDwtDR+JvgYhT1zma2tag+zS9e4/dicOZvdDuzMKfnWO1KocN2H17s
fjdDf4As0hiRVh5KX36mL8rJygcJcaUmVUaubRqOGF8pWAuhkkuahzEsjcBL/XPYdfVLF0lOvns7
cHtegOac/dhgDmdkaSZ3yw3bQESUFJ8W4RmjQQb4vPvGpqmjgPdYnCZgQtnHZg35I0HW/TEaJnid
WLwD+KHTCC5MIPdTY4nxLunj7ysnozzBKmXcAq/M4faTXnVDvPSo0ysk4XZgm9+k508p5xC79Rg0
ISDd/Cst5xHJsasuHooftM5KmwsKjCSEj6y0jeAVRB5OQmu8GdnBQyHkg4l7m1q51TlU+K1gzUNT
JiuJtWQ6aaCtgVgqRni3OyLjawJPrdCoWQmb+RgDLQPI+sHYeUJUjkrHwa5mKLmYLSg3HVmcpkm8
Lb9CWANSulvWU/BSA4aRPKMSAHm1MvJx6SzI2l7CDbgc1bGkRhXLfXUfd6tEZdLvPMv/GpTo6oyq
oY29M+tSASJdoXLYMqlc35oVk7u0fR5MKTCvhe5LsooOhPzLahJLaAlRccva59NLbRwGUL36isbu
R0epS9Fhqn7fmpW2qiHhZKXsM7ZJz6zwvb8/SnBDVx1frPnAQqPCFrmx3ia56KXRrVhAszH1kovu
Hg6uHEVuselUWwV3paWP/h35YPr1+KE1BzJmzF3cz5mpbdKI6rYk/DkbcAiSlJDXpAl27gm0CssK
Tq4Kt6Yi9MXe83xgCEb43kUHJ0OMvTBJNl0q2PGNRyWw6RmqaOZkfA1P1IYyaMk6/6ZwwM94GvOB
/IQte5qH2Pzgj7ZTsLxJrvJO+4aUszJuwq4GKqKBJqw0L3fty0qIN0rFg4G8SbkFySZtJEWeTQ/T
dQvfwi16u0/qk6py8q78/Ua6ax4X5kwwijjnUwWgnhCIHBXb6SsLuaHjctxkROgjfYan7eFWwl3i
eoYZMdAIWwy6jyNkFszN6xsk1YuAx3OYfyPJS/86zf3DrO1cjBoCzb/WxYYLpg8vWUb6sY/ZL+gz
Tr9fpQ1FsVLyB+8FPQo3Kn3KmYAx4I57Q5z45U8ZVx475/v6vRkcig4yS+4touNvtD8yxwqriBG+
if25blOPMMU9c6oTOYj6ZdbFrhUQVF1WxaGA1ERAuwx+aqzImqyCWaENWLZ9ssO5uUHLJGBKOrAR
5fVflEOGeajGNhfCbztwQL1ywz8hsLsFkoR5tGGaa/wi0ZFxNoqArk3yjtXv0/a2j5HXkItFMxOh
CSK2tISZfWYC0SWit+whBv6AKQS/RKF171nqtkQRltcNEDJhK4Z1tNCt3zOtAjenu9wqW9LWpkNO
TV2b4rAPDlCivZ5i0ZK+/MWRUUHLyxQVzayaHHgVqhY04ad5S4nGX6H/EuyxPIZSO95pI71Ewx8X
xx5FZYR4aRAGvueHNgTYWj+fhNy95KEvgnXgYHb+wC3DdPD0wR1451I0ZWxn+a1pAoAA2Ds3RjjQ
fl6r7LvJbL0NGQJ3VsBsLuYlXtknMeiNdHN7PQVg+1nJK9JSZPK0HtMu5sRWZ0JMyQ8A3PEQUXDN
69QzKP6CpZww6cCLm4f+k2v4aK9Iy2KdHZLN06VcJNGU/qKQ7flYUX5PN0wkA1X+4Cdkb874JqYe
Cvh4MnxruUxh6/SxR+w27ixVUTGB/9/wVDBYWlcRsD9dFa9x4/F9RoBP257fGOlLwGnGndy3GMuH
Qre81YbTAXPxtp2lzG01aD4NUuOtaGTEv+RCMx8+bWNwUzmNjz60S2LmMsX06585HNkchrH5NwAW
L0vreR955+aWaKoittcXs48cFUFlzIrFiV+YYq/ls4g9rfrfiEgXWsR4xJJli4YzsulCSoEWNMpI
IBYbcphFNu0pwYEL0wc2TG3AlonA20Yu+DC4htJlR+BfK4XgsPg/gEpjBhXoQL4Fp8sEp++CqCld
kGWwMhtPWfOW7Ob960mjAZaviRCqhO9x7PDJNDtMOWsvuIZ6s3qwwX+HafcrjUFOLvkm3g2g+QJh
GmI7Wl5dKZAbNxbQy18+Q+cp6/Fjx3G/78M0bahG4hmPVw9NfBc8bVoJLpQH78MckeL5C0ZE3N5a
78S8tTy5rX/z7Y7MkUQLM9AiYGRZKpH/Je51zoYQ4uaU3Dkwxs9Lhu/us33L+iGR8b+N7ACqUt/i
al0UC7J3LWMlsInJw6OWJtngDVVnNNB7DRi/ESyR2aYl8GlVOjOr+jaTec1PwYTLMVM0S3pJN0/d
/Ym0JFciskWlAMDhSITUy7TJEkkYRorGU6JMvdRx8fB3ynjEdiZnCvt0eN6EfBUcgn3CQsfRSdI1
eX5u2MAu6Ug1gauadZ3p/nGeb3YkBP3GGBl2mioJR4eLu8UJjqiKHmH6dh1DfCMGGdefv7u0daqC
bDyYAI84heWRT+0t2gkJRyX9zAzDM2CYxUz9nGxEqY3vQSPgUi72pygZgSslLkh8Boy96G5h3OX3
It6hZsCujn7SXkF5rxIKUpLuMWqPSq0kfMRKdQ2m1M+66BsG3p/hOVvyKcb4nUfJjjGlyU3t+3/8
Eo5N1dH+PaKJY62VuU6GQ4Rt6owWMCHnA6KouHx8FvPWeUWMd5qTBR8vQshmOmccDdrTWXoiJhrq
VlefOqODu1EP0nLVA88xTNeqlGz17GAO4VfGbZjDWX7QseMGX4h65zrGuNNjMM2vya8TXxbnKIqd
vH2g5DgV0XzMbcQT0djc5+elgFvJ7cb0MWgeCN1XWnAfI9f+Jj5SLvhieVB6udee4yTs4ySwxGRU
UBdIXUDk+fhcE8YapWJ7c1aFW10CbG4D9Dr9ECQjZ16X0kM1VHbCbBdMMRmOZMGZ1lERkBieIfBg
K5U3v2XBmx3enCKYP+iXca/uLfOkB5/lmb13HkXaK9G5AqtLXlDqtNkyRzlldYBqvG/UDp9xjgNp
j9uG2JkARbuJ+EVVvccS0u0HyzjcN86h8Aes6j9GgfZE9qDr7nlfInEyeQ2a3hOq7gu6LBt4dbuP
pE084EK5wGiVriDAftBbiE5jnu+3e0HFWb6idw/pnVtMqE9kDs4RBTuUVgvN6oKzVO0lg03hBGWw
rqOLUFU6UJ7qJpPomdysRuwkO5CnwdYzdg0wNhT0L+1iTQjJfEmnS9iS+/vPh1v3C2vcxwCgU+c9
Itb3jk9C2KGNQ+qPKBy6y0LXpoVswSgZs9kzZBlld1aqjDYwuUsBUQVf33Q32epEQ/PO5OseQ68T
2HqpsBtt+aDDp0xTwABR+XKmq0bKZbgmWkdQWXeukQz6j3GKbFPLNMoqiWTE5yiHs1q5NgyHGMmO
0dpHcterDOdBabZwv6Qpl6pX2ABxfKRUeAjPaDXh0qs+qTDjr4mmI4CuoBMjsUglAwGknnNmYdYm
likOXbJIvWaHYHaCpB725pKSxd9p7eX2DB4RiXAp7c4DdSd2eukbaCV7AVv3m66YXEwIPj2X90by
7COWfCw2uMFn0vp6cjWC/XygXHHhXgaHONgJFduMyAKJ58kepNg3Oxl5ntz3gqxuqWmAXISFIhgV
9YLou/sJvHVbY0yuAV9CimpmPzdvj0PN3YWfVvdc9e4IHS+54tkzJMUy5WRzyD6ET1rHHo7BuO4q
fUMdO/SI7I7gpAtRmNK04xy7QoB/EwUq/g0VyP71IjB93e7tWBbkfrBb0qyWRBq0OkfRjBnGSVvT
8uaoTmFSDqhB2gNpiBOImvQbFfSapCE2VjhtqQRcsCJ8ULFxp34x8y45K8y0obw7B+MrQ96EmXKZ
DtOWLFlcBgYbYe1vYTUugFKjDLTpMnmIc7SIrBwBj2G+gkpKKqeRAs65vy/CmLnXteJkj608yUbv
AJ3YoU1c5Xu16QitjQIWIBc2Rs0j20qbYoFQR9XHgXoaSUSMZDdBtmBoKI/e0+DzpBqRsTRKABms
7VgHdJEOYhe7JAPcQUr4VcYl56b1XWRcKvJplJK8xwpHaGAkgfLf+ka8gYjrgEYwUm23vh0MVnKH
uI23LrsAZoO60g6+0NLpEZ5z8IkWJNpe79WZrrK9E1sGE5HYIfXudJMmJ1gl/Z+lZDzUe4J5/5vw
4YGFUKLhCpF9f8z4DtcYJ42X9ACHT0hJcoac596dFiwVyR7ruOxbsTfON/BusnKc9TTaBL+iUYPk
g5XohhOa9bPzPd6LKOauqK65LOVCBfLHv7TDhxd9cdByFKd8Rp81ZglNCQs8DVsH5A9Pdn9jpqar
hOEE9jJXHiUPnorXp0D1cuXI4oc3mdBnNXjjR73Eps3gH+oXocPkCZBtXV6MfCpPQbPGqAiqDPFE
6YjtNl5A+Og3XdkFf/fuJk9L44oS2J09OiDjIUZB2h9dKdcKTXCxDttwrSts5T677N/qhrrZZThS
h/fWzopnEQ0J/LKOdMdJ8KSd55ZAmDBVvLF0WGXW4TLYq89UoB3g5QavrJauhrSjVYWeXXYcFJvM
2f2AcdThD06O92lS6Pw5MP3n5RQLkTmGWbCGtjy4OYnw0ZsuydTFxtpVgsWdbOZp6rxgAuDgrTH3
fLOvAbA12kl0JBs77OV7JE0P/EWbNiC9B2FEUib6Piecj0dpmIjd0VQO2XYdPUgVHGq0doTpk6r8
yTshUqu93z0NsbZH9Z7kgY+qpeBrdwAHOFehjgR3H3zVSK7Z015LFHTWfmve6ITzdMS7sF/GVu0Q
Jx6iOQwUMedP9J9RJw58nHhxo7Mq2sSRWhOrj0ZZ+zwwcLTo+AMLb8lOkDDIgwR12k/KG6tBRDY6
GyF9DYzYbVerzo6KVsQC2eQ+VKrXf5TqxJufIyhC4qMALRvaLJYbB0HMNqUtU2+gg8P9bL/Y8df6
Hi8o1NxEJKisatMa4e/m0UC7PtWg4117XOzKYdcPzTlPjWnioJnZ4VsKdaSnDYaWOvXAlLJzZOBP
nkwOLeFwuV1mVOop636K+1LUpfs1A8LDwaNChJ4hUB5xa6dfN2u5Fo0cY6dl9BeO+5rrXTNODFfF
hL/MLSa29QINpsdB0ir9uhjyIWioxiDD9eemTpHyCtjvn12I5uZH6VO0ZgH+iqc7uL1xCoFlUMMT
StveE6xa0Qf3JWCvXh1+TwLbfZfJ1/1yZ1KDu1FZ4TS1K7Dug+4sR4MV2tPXJiW6epXTh6Ks0YyB
8QnEG3Wdp/3Xz/BSFFcSUGfEEw1xZHZxbIXOej4FcdEaN1E0sc9LzNW7b2GDnmyH1mrJITpNQuzG
almVWtL27fUFpAyI4x3RibUzQeefvSwLy32wDyN+mnvH5gV71Vti0n9GW0bc0VXhotd0qIkfKppc
SyR1tgl1OFJ6IoLCQmK/d39bcvZcZdM5qzJU+i+8Am9+ySC2T1E0wL9vxPunLPwZOSYsZxFVBlCs
ZyiID77EF4MUE8saJrrc6N/MJto3uDGbpPIqWLhQxNABCoRHOCWIaaIzbVU8SMKX/ksQw0kuH/73
y2GfssLURINQmRk+pECelExQST2RrS6PZ1AvlnP2+PGktXruGq9ZkaoXXqCbowOe0Y41634gFMrF
VEMZiL9YAt6LF/oBsEGUDyufN8QmeP5C8q3X5gmTBApzAlxJofKpEIPgNPMWy0sqL50EbnEYumnp
o7e13pmfL3R6RDTuFSKXJHoeeg8W/eM+OTg2hs/D0llimNRkjXBD1cCZjIRv1uF63nrJIDYUWeI7
wZyzxZ1f7vfpZ2YqKIQxp/C9od8YdkpiANHgkHrmYKAzS1mtbMz7RGnzKpal6BDyQnK/RtfyyGw0
oqcOwvSLWOXXjN1hL6PT5Jt63Uxn6tgspE3hyUlTev+yo2h6WFz6abgOnc9TdUDDogWrv/2B72k2
kDH53SSdkfBajEHJgwZ1b66QojRaNxB0Syg9Vp+94ji/m58XlmapAdYxn3RYg7dzIJ9mJfINWMnj
z9tGDoALNCBZR5C8HeFBEqaAUsQ6q71YRPmaHof7RQIqcovZWZqCBRRMmdPVuvXL94KqQPGp4NyQ
glsQ/m5YjTLv0Rk3bb5tP9Pg+GnYC4yrU+VVEvfexqSVdykG19zaKGWVzpStwbIpNwh/AX04jKsd
M4MzCdgm0rvIVuaqGhCdG9+lZuRhzh3dlToFv4UkyZ+T4vA6mQjtIgkjta0rQkmRQ6yXLiIzSSK8
NBy9x3LRAqeT7txB/HXNigWLIokBz/aeB6D9ORXkrx9QbGRA+6VR8SkGIxnk6OM0eTcm2dB1PVbX
qUZ7wC9F3z41GbHvQpLLXZNfE48+jgDINhTgplUKHksIKQZP66cWfjZ/bO7hkFZfwzvfcz+cC6hW
BqhP2YEKmXY/PQtjT8YfqsZGv2PpAkcKp2vi9t1Lcj7igQJmRqUTQVogsorkbgUj4KxGdAqJjRqq
3DxrbjsUcGSofmebFZP7XJSfCgS+Hb8CvfbF2rtEzr5j/Yjqm0Efn6oaJK3yH5T7jcDcepY70U5c
cM2e/11eUqM5kylpKySLvcWp8torZB0ZS2JPXqMx6LPpOmPyhUDgj0PqGRt6K5Bkr8+UahmTL7O9
g6MX0tTGjoA8a+b3VWHIlQnD7Rm/8uUtsSeMxwPraRlYs7aP9IrxA1j4A6X/BkDVffJB5lbq8kec
coOxnlF6TZPryyXxi4hHB+pYS5r1Wf4OkwQYZZOozsyyHtqwER+tQciPdSCYzFOAY8cRSupXENSV
o0NsFdFd72hM2RMP/SZTKDAAy+vQEbho/3ndaK/F1uGbuPdm6mzqTOmhEB3vUe9OdMUqGE43hF2G
qZ/Ftq+aWKMsrkuqkIfM6PyldSYGTr2azEjdl4pFxtAFIqZ2TL6gk9NrPhKb9BunhnMMQAqU78GR
KaV00x0ex+BO2ZeZKypaRdmRxjMp7CT2ODrFm+cA9GiO+g/VVfbZXlN8xtM+K+s/hUZGWG44SVJS
qOckvb6lmTHAd3mB4qYDPd+jz8DnBDlifZ344jr65cGGbz16al4wNk8EiFYM0MG+JzmJc1liOn4j
K7LQpQCUKpBlOi2vUY1XxVEvijWALJTZcUQU9M5z1STHBVc4JKtMEZTBe7g3/hj/x/XjGCAkCQv+
Y0Tcj7woaqEtryJBSiCHjcmCSJb3QeKIAq2UFT1bIWTT/pbQxLDG26I9epo9fw/Kk34Gy5J82Jqh
dGrk/LPuvNU7phRAb7VSSMrvOvHECaL9hAMxq1MCTp310eGVbJgEwIV0Lj6D/Yh+6SMgMJHRffKj
BKeakMG3gug1xo3fg1W/I0zzN9TvmsGlnx6AS8LXkNGgc67E9V+8xZ7OhWJ3udPfl1GK21Gn3b2X
Cf1WRtHf6QbRarQC75RqFfGTYaF2fmq1vqFQXfD9MZKZhCi+XpbrwpzMHFRTufPE/J3IHY5FYhvC
AeOts/wvv9n9S2eDH8uiKWPJi18N8YAHHG/KM/w5hEQZTzWbyqNWC+XCUscNjHbYGp4Ol8f0asq5
4YwgGZdgNpJW54dHUy3xb6sTJGYS+dJB1SuEQQR2yuYkM3tR5dOL9EUZORKEj/4aaopCQnSR1yRD
eoiHAvAhPcPT+TNHxbyb3HcxYv/rxwY/oKLm3EjEb6GQFePDF7IqIPmre2yxQXpiN7VgVClQnjf0
yi5/+n1xGso3Tykqi/FCx5wNJ2ngh8JVOQHLKCWsKPWARxROluA7ocxJil+AGm8GnNyGn/RhcyzH
8px/FW4jQEDBTYDLhmVm6fgTUG7QKMFCAlYbhNW2SlgVoqPNH36uYG7HEyoqneu42eWiCYlU597q
NtIJ6HIn3ZF23teWNn2kAwkzsh7QOCemm1m92YUD4fBikwhAeviC6m8Iw5zJYqBQzxOi5s17zELE
yTuDqj4VCAnhJSMvLoazmeO78NU0m6EwYcybBbNhlYWFmB/HVewzhRjehPFH5zL2S1dOzOU9uX3P
nKbI5yYyFY7V2eJspOuR5+yzWvJGqjaMGdcjj0uFt7LCQ4Kd5WTbQZIu/nkrjzBARq+PzteG+qiv
vECMXFp0eCAHuSlGOfbyx9Skg61UEsb1zJhn/liTd2gm1gFsMjNcqUgpUiMwom6t77UAB9nOYJYd
r92LYfi0DePzKMu8gghRjNWZNFtNGnQ+JlJBxMk2btLL+jwMNpG3fFD9eTQ9BY81bfYHrab4yl39
BUCUeL1HVy8EmsW9hBapkhOsrqpjTRZ5ZSHjCWjmDsThCuLHg6ZeRfpajJhTeR56vj5tvCCWNADy
6968/ySFy/uIHQinNvw2oq2x0qh+KYqHA2vOZJB3fkjepLJKaUy1p5aEQj7au6EP464y+nMUmH1H
e0gRjQLxUJT7nhuGlPyYMoLwWfh66q7NB0JrGrjl+9WoruAa2F3fkcWaY2PXOBlnWuNwGr+LQ2ud
0yY6qDE6jG8iaKjzmTmYmR1H8GsawvKfFtzX5wbTBlBy6pAVpiNTZaJt2L6pcMHI2Fv9PZh6EdpC
8MfgzdLqY+HdBcQgML9JsEooxAYdyAXCjOwHoMQuG4u7o/NHg26+mlFGEXhhHPnBGv9l9HplFDke
5DhzSCTilehWdn+QVabbCoV1Qp77VtvWQycZMCLMue+v+ABwjnBB3rUOzBJx+Nci5z1kPl6ni+so
Bg78/GSUd0WCjySXwNyFw9+IKmOEVNXc94m4ye+rIeBAjAdrSExGUOD4PLHYeViIEkVvQpcWRAu9
j/UxZB0eb+kVCJ9h8WsnhqJFj1qoKp+CMl8ZzMeEBYkhi0JoojjULaA37qdGXQfeG8HJcn8e6G60
7bSet1QUBBuZC+gecpDgAluOBcWo6vAkeZg0qM7lcWN+kebTi3mjPlguiN8CDhlLX2I7l0UuDhAF
OuI1H2ee+Xb29WpHf6UIwcv/eZ4RwGpPa5SKJ0yaULC2mBwiEywoWu6Gpr9aDMKp58PFG2H0X2Sz
k68X8ltYY/TGZQT1F0tzSGjpBFbVyAj7YzRHaA82Gj8iXg+cknOQ9pGzwe/U+uZ1AckfhjCN1GaO
9Tb47s8ad8GcpGwFShXzkWhoQa5QUMlmGEB2nLbetTXpoxddPcVEXpCz/sLthgAK4d9fmvLGoVl8
K/SHfmWvhb8audnXIVggXDIusUq17bMZDMuFSYA6oKBxBK9HAJUKUKrZu4ogyllASSY9fSmpAhXf
SSg8pcAPm/yOOPz0b7yPz/H8cq2dhXcDNdFPFpwRu9J64kPAguOj33LsLorXwWccg08cMSX+giYg
W4SMMS00C129dupvsTR3LcwvLiWwVULEi683zBKJnS0y3MKlkFNNvsfqc1+9t4El8tq2E6rGVHBE
eLt+szML05sURmYoTcEGyUA4BuYjr2XeLAqc373WD1hr9FFVfdAVkE6JDd1fQcZOm8l588RPmVBQ
O7nCOxt+BVywKowr8oXuMppLvysiATCyPfdmNZj7bEunwh+xZfd+J2W6HZN61gw6D5/UABVaTXTi
iqpIR2RPC+rWYETwucvH6H/uZI2ptWKwDcGzdcGAgE2j4iJ3upfx2aRfQ3xTe4KJFxUyo0WH4Gi+
TLSOv5KTWwVNyusZ3csfgq94nAOnXPHX1jAW4HpnV5OE8OODPeiuubf5NWWl+UW5aGjWGpj7AEHt
hkOqhl9JRpaSumUfRcvb9G9d7JDcSGfOTRfPrhrpsAM4FZtkrqafpvIyCQEXbtiOdEQbp7+J1l35
3/qVqXR1wcYAuIzGDrYpa+Z5+3ONndXFzMN6cPm458H/vGAwUEWCRowUu7ozieYe2+h1+oQSBL8U
p93/zHvrZgn/g4i/bwaEexd0dXFOx4ZNy5kWEfalAwQZvmkOs9eVfW+DD5Y+ndvJRmckd495/e7X
9jFo4/sFFY6UwbKUcQ0StXjNxEQYXXlF0umYGMBUL2ZPDFuMcaSLHEaZ0wjVvVWnoR3xUmHPHDD2
VSlTJtxbk+P91/i5LHEu6S/pDx9r/neFoExGccvLU76/rKKa3TvIQIEAzVQRV1peUE3lVO+ORm/m
2d+DBSqj6seBsEnKZ4wcigKxapl3zKcs166RbCTUaMOudX/3XkKNRJ03Az0I69Q+xNXj7WIibdo7
iKc9InpSf184BvPiTbdPP795nLfcAtlBZoQlG4MIkdsi3OCAdzCWEIvv7f2ErI22b1Nr45T+Kyk1
3r7XNTJKuyNCYh8XQpItdOyFzbWZPYi20WqkJdlkSanif5d3Yxewl07P6nQ14u87X5T1hHeZorYF
ZcdMnOdl+kW2oAkflDnZGgb5YYL07bGNjzridJS+KTK6My4kfB/fM4v8W0Mf/A2LAtvBNAl88ixg
XdjH923rL6wApOVUBr4qjpx2toHK4PaHzfJ3OaUsnO/w1H+GwNIvuJm8pME6XqeeyFZ/nONu/L19
T8+lSOYaOCuPwHvVM4CgGTtN+BqQ/TTADMlafMNovNM3tpBiM+ZwTBS6zUmfbA7enkhCy1kODUNa
3b/UlzubYQLeauxzYLe/RGTMJVutRoViVNE8EFqhXp65t9JEqQTE9WxZYFQBLUsa3WVIUj6iF3Nu
NtMtqY6960ZN7hgn/bTL3gr7YPhEhCf+MCPyRNbso/bVvvTrR7ICuIYYZPfEjK6BwaoZM/0NuzVO
SqJaLnVTlkLwqF8zM3p6jZDo1tNf+TutwwwHoDwMTZ+sha5BiUw5ow/c4Olf+s2TvseATIL/x2vw
58b8v+PWwXR9SHizjp3+uuRwkVmPTXiX+mDNE7TyyHYkUzuI63j2/IImjsgapLoQbPtGx2tuYrLF
STIn5S3YAuyc7220uNhbsi7rHMV1XAohRf/7u4/nIYKsf9DaZn1acgADB3k9nmGNYzbnWinb7s88
cmns9cNLmXgAUptPFxIax80eRj8GBgr+h+6w0lmNHc16DfJVhKtNrIVZGx3JQmrCdR5mMZmm9mAT
l/wsc1J08/R6UhmH3RYmcSgasZ3QXiBOL7vzTHgbhyBcAIwKym1hbNOcp3uvuzHC/bc7SoYbqETg
Kk/glToCr0zE42bqR1ys1qwrrYTpuqv7wfxvgt/BawwN9eh/Fv/ooIOgIeFAckLH6vxBgr/8nsQX
t9KTY3Y/IqJAbIGWaZgcNb9yEuZUGxYBSqhb5UIJZMjABaabbzy4SQJgQrHd6/XJ9VRvmdokLJLX
o0BBz2XUEdsPkNXwM0+pysGr2i4x7YrZlaT+eiYeybxzN8M1SFIxK9rJiv5KLTl7h0U3K5pjbnNZ
S7mmtwkWsmCV+46yZq76RvFEHXdZbHT5+3uZtjyd5ilbCFgjnLYKf6IFXIsZ/D0wya3LIgrvJQoE
cA1nNtRidmhW6oVCKpVrtYe2cQJktykRRaeMpwExTFvlAJMW6kMkCkobhk48STXM3r4FwHOQmsl7
6xAfIbJRs1G08jPQFbeQsag/PywtnxAbNhrfqxHnvtzeKhCttnbM58Si+4qxBBUrTHL3UdBPGU0B
/FDF10PYB+lzAc5PaVJvblOqy2Y0ZVoqeVgyGs+KwhSbz2R1R7EWM4t22GtP8Jw7c0QG4qXZ99YI
o+MJrTqVjs6qYBaOvlJa+sKWARohJa6OtBJRZjwQmnPkYFaKklhgfuY+LG1dLJZ2xEQF+7gun2hf
XXCVLNrDYbRvojT3li60JOym/H+rmDUfQpSUOSBaSkqeyLROWwVuN0PJeXsBJApKLlGRhUptFES3
cTsoKTEQ61IT3hq/a6fXgkScfIkgP5iAGIqExyBz7M2DkER7pDfglQAFQBPtb25br/CEo+ayehJe
jxVYt6Q1GfDs/GZ/DXKUqOTVn2/Tj+w279YvtSgL+C5qvAMSKExptWcaYrCFkwT7pVo2/4SumJFw
jU6R04TiH+703YFeKjBkNV39QdAk6XsT33FPKCt7+Qe02VFaDrMu7vH1sxCo7Ql9zpN9x1KEt3UB
8QoQRcowVhGOMaGco1P5aXgEENwP3QbolRIFBwXHdzZDkGV25g32seDy5rSFT4Y2ZuKudwNuSONw
lhyU4iXstqSHbQabPzIuds/AJc1VZ9W05UaKR02Z1SlwtWtP7D/0P9hNOy9fzih/a8MTtXMghJEz
EXWSh4gKNx+nyQRwB76sczF2IZfuNte+gJQbQRCvD5xmxBjzWycLHWnsd918iZh3nbcaHh3H0x/B
BzU4eKoFcPhsKjWA3lO1LUIm4iuZIVQ/+2wfvbYZg3vFp/m9zXdUHgjzN+RV3AvVQfgLR6cll0yK
ztKBtFq5HeYctR5Lfi6czsHqMjqlCgvJO/Frg8YeUuikj8CaGetQBG5YrGqUwUk86wj/dPF5pzdA
2Y57JHmFwgISEvY1pKlj4imZb3GlcJUT4ZdjxQFGm3flgTQ/YkCpstrEi8JM/zV+rhA6bmOsC8rW
Gu/g4p7WPAw4gbDjAU9+FMPMUy+2A6EkrZrKtMJiOhV1zVJXe9X8TDrtu+lHEPTF8wcvWEXSt5aZ
hL2TaNiGlcFK1D4sf7XEaXkKGaALLoSCpEXoQva6BsPx27SmTNcy0LYsS1ubAseXn9sV1phmTnw7
0LmaTo5GUoPHUaLUAFLIU9BW9bePk3+QUU+LiuiV9kcwFdy4F9a/CGHxFDu16MHmmPXhLIG6aRPC
+FEmbSeA+C1my0RMy7z9liHzdJqm8IksNWLaXLN5tKRBsKTbbJ+EfMW2QkzPrYopO3QacS0JLj96
LCDf9RWx/2IIcKE3x1VNCf38InY2oS6cLhsXCbKtPKT1I216cArgRXyRHtDYJ8aMMktnuPmphV4b
OHwyMRS/8D25dS44sYanmT0an0uPqs5PnWmu0PFKQCEx3wteBd3CFkcHDdJLfXk+cbGTatIgf1a/
BwFtrA+yW9k4ENv8GdyjQzfhmakVoXAbdigDJXCxtjUJaKwfw6/jGmj1TdoPrFxq1jZz7a7L10ID
xo3D2wfRqb/VPrI0C48Fou+Gb6RBPSQvZQOtyNFhL9N1EsqvEblUvuqtulsozUiWSbyQg6xWsSvp
1VqXlvo8gFyJhAFVETycVYNfYxt6njw/mprIQuQWOrNWf48vFHx4c68YYRrM1SingjPBA0MPAwGk
HOu5RYBTHpK5A190fHI0eFTfkO7hQNQ1CkTV9R9e6RZvjK2bGPwJdwErVZpOmLTLryZJ5yLUxoiy
kqRCmLwsQ83fF1qY1pFo9m+BGq1A6oespXVREfmFqQQAiXZWPKm1oF06GL0FCZTHIa+8fdB1zyrp
qPDmINVGyG0UBG0JdtMU2zdlaSdrm9WjTBcq8IWq/41jy1dHHZAwe7rbUYdsXT0wf8odg3XqClVL
t+hqzGLgNzUYy5WwrwxAprgfu3CYdM4tqWqf9SDJGWDCnSPjHzcLvgltY/w0GG/bYfTuZDVTEQ7N
UzyUdonyPjsoGVyHwEpZMxysM7gCnjnEkPF2TB75/BnexEY7IUry30tu5s4jaV3qLZeGhANql6aT
Y5WE7hnSKulzSzGH9gqmmXbPZnj2IImyYMLRQZL+xCENobB4EQKWVccMVAsizNV14NugbFehGLd8
mpm9Qkxgh9k4vY6lJaj7jf3o7ZGS7wv3YwnxKS+vVmfLPaf5BENuSLGnswIElzWHmAR1LUi0kPGD
2yDIx4QBbbA1/SnBTgPE/+aKtas6neqj2UikyR7bMtqqOHA2ImvwrMnouBLkt3lOGpFRK/HP1h8w
6UMA84hah2NaxkXs5eS8yt0bhZi1A0G/SMKLS/rnR1omz9zeK/oCIi6Vlx/Twx4187OvHk9U1J3u
1ZOAD/8LkPH5Vb53FYymi/wDw+AYmHCmWodw7SyDVUAFoQnIK4Jzx2kkQEiFSW7Iq/Gsj89yP9eT
HUOxtj5jXr0yPvcVrejjMzDdSaW6TgMNyUvI6clg2k2QbsTfMjATjtADXWEC3klZRuAMjC8hwbsC
EJMWfFyFT5neeItig3QF5N3W/mPii/nNncDthpvPfK00bxzTwfXvjM5wKpp4STIp0rPIF3OR7l5d
bGV9fGpTI+xgg0QJF/FEGAvuGVLVUi3KyHfviIB8my1u5KW4PFm7QlwutF5rKRNOUHOaWVVWxyDO
nix2a3zgG6tzB2AcLbCrDfYIhs7sAgF4GlQKAhKgZBHijZ1zc21TNTp2hdZPpnHAz0cggAdmm6Yh
ytAgbnGtspZ/jUc3g7hQIuBPF/j3A2O8yRsYjDjXKj2SMf3ipHnzW/+7QIv2mpnINH8XlmsMfPf2
0AoHKAZCEdeJndIZ6C2slk+1nlB+mLcSNOqgqXuErbqdIi+StqlW0ENVzToJcLA5T8fasOjcHGFt
w4WtPbovLX21kSYD7aMDlmOI5rukN1Y8FjBgWsdD/vtHrfDzwQvl03bpQGE6WiESONqeUfYgnI1U
F3jWBf5EZbiOcl09SpXbBaRzdTe4/Bz8D7R3EkfmZTfd84vzJ/GL71zJ28EehqG6kSJzRIZ0TPIy
Kk4QJnyNSOCDU+cgEegmxxJpEhaVwB+hZrkEMsdumNx+i/pmIUvWpMdMlNOgnvpiPTKKcwE6JECk
D+BwPfFmtb+WpjXJ2EAMbtx4BhWQih1QiiFU+WsZrzrfPO8n5MgapUffmKEECNDP9LD+2MJ39Mq2
6ap/z74x0VCTCqHiDPEmfCSkWoTvtxwQu8KPmZLCl9plVrOMf4UPa8XLhgsRbNr5F5FmR+MtG3sy
uvEtb3KTOZUpd3x650WpxeDzSuJpAb5YNUf2t4hdtjPxY7iOwcvE4UPBkbP0AD4WseLZ9Yr98fz+
7VbcNlcBToy6DCza5uDD7jIiqCAOZaEHiPyDjsOJg4OVeVBKEVZ09wJpy1Z+RmOhdCweSs4Rtvoq
P6gGNX84pZALKXb2fbJxL00fTrmTXGYoQnoxrtG3WuO/CumPzkNeoCB8dQhMdunYcYpskWNwc9Hr
38M1JuIae6ccPdJraWGCRw/CjNZ5jX3Tjpf0GVg75qSu1qlDL9b6tW08/PgSFeBpEmhuCe3JwzFW
ftw83iSqIpVLyAVUnOKyqrvTRyI7G9b0uh7ijHvaSynfoKNss6LRyaQJEfzF1jzJ/mAJDqSrJNI8
XwbFm2aRZB9bed9CAkGx8xN9/3PZIYy6avRcVsNYY8sGVqiP1CXFA1iJ78jwcc3joya6fXFDHREh
1lbhY8jzNS4w7AZhEVvCOFA7cdZXlrqKqBmSvc87wL2oG7Yth4BmuSTHxjnJL1OAQPEOOQZqXzq6
RfEzwzUtlN58pe5YhaYd/UGcGLzeSJeatglo6prPigtZHyQ7gsy9mk6KNglsnxW7K3bP/aTk+Zum
lzRQAbgtk57hfuOVKzzsskEsZVQtQHA5M0g0EI7kEh6thal0MrGJEP72I6HJ5BB7d6Fg5a4zT3kK
/IJBR5G+3WOEmpjSc/qPSRWX8nFRQm08/XKoXEFqCX6kRHt9w15mW8vswoLDNZHOmbe2dI3Ae4fs
X0rTEgJpFRwhWpRH1EWhii62fQDzPw+zTb+P3CTcsYGokkQBlCNnc+l23zPsEYSif1hZrSthniyP
sGc2XePFBPEAYV6QWnoeXrl8Sn8dRi52xd14CMFAP9Ps9x+PiyKuSJPz8MA7Nr7cKnaApElYS2qh
lmgRYVlgdYTzKXsqx+aejz+55+t1pjBl+5jt6QbVTdd3IHGDMHiKT3iiYiaCuy5W8IAlOH6XHyv7
h6RfOgMQoGY7I1gcmFiuuzM0OxRs7lsu3yqbvTdvv6wf/iU55akDldJVaxQcDOhCfX/dwFe/VMiK
25/EFbCpOgDqllo8CmffsIu0V10Qsi6igdtYO+niAiA0lPaTpx7yPMlrUV8lIy33LO+mkH+DoQgS
+O9XRA/VL4SeFip+YqLiS720W3xNnvVBPbX9S4QFYlXa3zSDshMFodlR6YpjH3h2tp1fHy8q/OaE
J+L6w0Dt2xsWO74eM2co0zC7gyf7A3Byz+Qzbt4203BUT+7pJxONkKTh5YW4i6T4tLJyfKJWpOYq
pxNpUjVUHPnPqQ8Cr3qMjCiu6sJDUaeJLxwxt/dI/Qw6uAFaRo/LKu6zvh9h4oeottELWTOpc1Ly
l9TsqtItTFkCLEuMQtdcS6LjoYT+haWVuYhx4GlciwcFBGZ/O3cMOz+ujcn6YSxSWYhPySzwdfIA
7jkVyZbvQ6RdV1m6db5iYdMiLXc/Ud0HbiKLeMBZZtlnji3jIizaULbY/JTHj3N23CAFl1BE7Klc
WL6fDg3cwaHQnkHkJRZmUDSUdQ02+zYhuujElAuxsqm9aSzQnpDpuYknL7rLIaG0VJrw/+Me0jx5
9VaC3ixzZlcYR16iXPkv18wLYBtRWS1G2CF3nAS82gslCel7YDDvsNE5SOmoDPJYXQqw9DTr2LuW
VKMwf8G6jUDYoBYOUnv4xBRQ3zmYMVL3TOZe9JXgqKImS0w+Zcy3XB0BAYivE2wzp/sWYfFlwU4Q
Wmczw2c9Y5N/X1li+EjhnBmmvBD1XN3gJD2zn87+CWcxQQfSKCP1hKSbd0/xg1ZVQQjHcDiBWBKd
v17rK3PmrOwcGnvhqwlFMy0KNywNGuW/odPJrTdh/n4pAbTZCt0wbSd7VRkRnM9Ere4XUtKd9+Cf
gj0yy+68n28bd3/jRpc7+ZebPI2zhRWG23dJuRh809oevAuWAyXX0Yvyx3ALO47um9X0IyKCaLqL
Ot8TNAYT/XGm44SdmGPSQpVKSeFImiV39EQKmS7XnVIROi6st7jxqcOJHCR42/NTMNT4pTmFw21H
iexMlIJ8SIGVNLYnbgNx1OUtsmlDVoEyuuj1ZVMiUk9KiYQOvjDrrx8BbFbgp6HSqPoEmi/TrUBD
YrabCoGVCA7ZacWA+RdFlcuRbUxLdn4AGKDEu3jJbuuCigzk+YjhfcrSQ9F/4il8x37nyM9ooyee
9ECxL5z8eor9kLQU/vpJUHIHezcyMASaUfoQ7LbsevdTDthQ8YrhXGxYwbjjEFO/2R0NEEloF2Kj
teRrFYlaXkjJJBQJDuQ1jXynET/KFCqY7Dc3YTQFj5wIWqY6Lgj8a0rohKB87u/eAxH9abdJI9KP
mf75uxeXt9eNqQEB6Bbp6ydeLppWRnIpowsJfblGj/3EGDPYUw1h/WGQIrgzddFy9XbJ2ip8hYDz
1Pz3jpu1TdQGZa7fmL+FGZr92NeD+20X9KfiW9tmWg/DWtc8ZbM4uwfT0wNXqUzinPDrZjH62BkQ
etrGNOOU7z7fI0pxnkGtgPeXD/a0C9Ks+j4viCP2v5h9U7Ppw6VueRILcVLchP9HM9/BzptpW6AA
kh0jNSKuuOiFi/fp7606JeCcB/qKU+ictTVCpUGg0nMWK5ii1f/gAC2aL6nb0dBA5yYuMxtjR4hY
cXK9pNXjf2s9R5x1B+in6DrgP8hJBsjvbxykLEWU7oDwbJfjdNLoqPNxVZbHGowqAQulLZIFzyCt
OCqkfPjNLsBgQ2n57oChNOFS+cXiQwyyXUPbBwHfSllByf6FvSWg7kkeI0Lkz7PwIoe6CqSYyWXn
Klp/6w5Bz68bZcjZ/ChfF0A6n9B1zRD7t2dbx/7t6RzY5QbvQUfO7B1fMtkDllAE3hMHBI1PsMm0
nCIdLfc3tmQQR5tJWxa/sDKjsD2bkYzG/aAepZLsIyEcMZSReUAL29g2QjKHoNXvNbes8GO2wRZY
VWsfC5umYuf2oNMsh8mFM5/ywRIlaAigVnTjjUO1k4xJ+beusfkR043kyhH+J3ViflZTBIM94ipu
c78mlZtOLVfgZs2qSZpPHAxDe4HkU2dlmhzvrmFMDMWWtehYX6ydq8Sj1lM3MRDlqw7du1gBTmSN
LI3OFqzGCU4m+RD3vVmZF8MutT4muIOsKcWZvotSY1NQFhoehiOt0Als559fF5wSmSHOdmulQKoH
v+/v2d21bJLwek7erhhOxsVs/PBHW/DKCSND5/VK/ln780BLbiJuIg0T4YZGzFrcjRbByXiT5cAK
hfkcIWxcEgJFjp1J/zYER5QzXj31yG2HmpbGwsu1ASOlTvNlBDDtB1w2So028AdKtD9IqfrH9I3I
qZM38uPe50KCrZp0a3sbQxjjM/ZLOo4HtM1TeESdYWCS5DacmViRXmvIm92GWRFQzileg+Eky0hJ
Um8tgY/cTdFKXVR5u+EDQRQ1pdKiWWx20bdMreg7pDYFGxX2dh5QwxzdfTxQ2T41JkBJaSPcC6v4
OIKqUqGfbJJXu71SEl3LD/5VMCvvcNOUdmvqFq+yah7KNEVr59cLS9BN2vE33IqT0u6NJ3zf5LY0
yVoHxe3OmuUAzOnIIppoADUsAIFj7OUkzYmGmVE3bP5RyRfqq9kG8S+jV2y0cdIJK4K9GUhJbdgS
VtC1ckmfyf/ewcTQ3yX6Y30MnbWR4Xpf0MEl+fqXCPXahLQjZHUItup4NQNypaiuJJ33F09ojqSz
/6IeBvTABshj3hWB9udn9b/mLqhY4HAz2l6rs1z6OfAmzcWheFYePns8v6oxj7N+TLq46GtuUhFj
/r7aMkMhBIKwKlFDBRoKRQpoDdlcHvhf4pPGVqfXduicp7+bp/mLStCPzwksXrm5LNbWcUwCsN58
A/iEKdLDvkTO+JZE8+u3S/AKG9J4H47qMvZKx/TGIa6n2faVcGcvjOmig3TtTY0OT+rqtu0rxqSo
tG/F5becHEtmMVD+zTdJz6/5dl6z01GKgfCyxQi0+vXgMfPSgJUPDYhTF/n6lHC+aaiPheLcSu4r
rfxpkfq9ykoJxf0fMaiQ3qwDMqMw9x3Y05wCPcsIaBZIvlBnVjXHnl2HyJqXTxuthNH+eE1oO9MH
4mTxh3Kvh7NocxhXinTiYlH1JOijtLtB0SAh+maA0kJnJDBR5pd4oWSDdaYSjxbl2Op5Wt2J08oB
tOn6t7ocmo8FLy/+9ozdyx76YOQeyB6C7U8bBpzfwqKysHWWe3pNrVoXLxAl6BoAotbZQ1p3HyqM
GA6YsEpvhnx6wgnkKLrFn0cY1q39RTVH+tfho+GB42pkJjo4437xlS/CAc3RM1FPbuXjLbhmvYQc
LAPKQ0yhqy5qJPBawjCbjvpSp+vH8on6y4Rw6yT84jJtARS3sARC/fZ5OFURyBqhRGi/qBzB7Io2
vmRIio6KB04Ke9aNjKhXsqYJVNnsZc9uqVmSFNTPcwgzJH8G4KkC5Ve1MWBQGDPfVYtyu1Dt9jY1
1BLTCbQBmfi1M7HNg+PqqqftDaVNd1+mmiFzUroD35wrjH2R2XFj+Ffpk8zykmOSJ/cGvKcPfnZs
Y0DkhkMnz+gjmAy4qfkgSSs2OuHsfdErXyV7zCplOxof4wIMjIsP8axPxHhKPZxQxRKplgTRqOMZ
kHjSIzpQXTzIujtKigW71NtQn48Vgwpeds2aPZKt6ZEvF8bth3Zdtr0tc5E0iDezJpCtiyGlXZ2C
yOwif1BxC0oZRt/yZPKYpCqFhmMHnIE8FFWzJAI/Mtoxlo3rKbS4aKpMWchmDOGWuxwGAv/3lRWr
07XxuLvKtbkhZ0wK/eTcnCV9N+smbK44XCNimoHwQk4lajFIH2H+WNPfAH6pxElGYxTEFE+vRWs4
UYlvpUZpIChmT4xhaIK5/7tvcDh8nhYVZq1Trj5kDmrsJXycEAeWLJek3pOUi4QMmsdtbIbaIO7f
OR8U4/GGCHQomE4Bcuz2vCAwLs3g2ikTNFXuoKFO/Y9tvNV1cSYDt+yKY9V1FBxrwZBm486zX0W9
I7jokjwTDG85c0gM37Ohd0zBBfhq+UundWYTmuDdYjURG1E1N0Qvn46emJGpl3Aqj6AjWaJliHp0
hSkO/uKt+RWIOp0ky7Y0aUd/RY6DwlXZPkjUvF/uh2k8zKZ7QO2lPbpbIzhjzpUS4BnCZjxXhcHR
qOqRoE6d9778MEf5o8lwAaY5eaxHOlodpA9myDvLfYmdMMI7JVA7KpD4l7V60aTQHHqy+vkgToQN
osjMaZBD/fmZFJAt4I40ZH0ujlh1qHdy8B4pTsaj55hve5pEvx6eWX+zBPRGTtdMQXZ9u3F/y3qN
Wm294a+Qcz/V/s76STTstMWL3vj2s4hrBNSDvuHEatObE+wjy5axCZnGLi3182ZNrtUmAfK1ufAR
94p9vxn8Lka17nfXY+/H28CNpaLSJTKWgThtGdUnM8bj5PuXdhPThLHeg4d1zH2qhKTkrZs7NmkR
+fZ4krkbHAtpYlcL1GGfXWkQw2zlhD/s9fqKEoWdcKj+JXkJQu9vO+H3V7IbUphyNQABMj9yJ5LD
doeOrKNEGqYQO0lsy0+92JHnX5Ie0zt5BYdnzNWSDe0JJSJiuTBucpwZdRyD3D8GBar33IfDggzF
Nu+56ETDebDwm+iD8gPfmd3DSkt4sCgra0cPIHzwQW8uLxi38qrD8hSi5p1/gOtHBALw/jb4pfJ2
cRKJQghBzL3LC31u3c6Lg0byjq5vjqizy8H6RVydD1DPzi4iJShQ0bL0mlIlEGBYV4jv9lJQDh76
Lt/ijqWAWLR+yCZH2JR4oxDUjlWSjUrCdtkfo9aC0NK6e92FkD7Cd6NeEFk1jtQdgmnsesT8fVsf
a8FL3MfjF7Dxf4zfc4eQ3/IhOxIz5Tv+5RssrKGrBZrTxAKbVB+QPGKhfz47Awls7VTaUJ+jszSc
nfAqDP4AxOnASIfnPPp9M7GUo7wHbZ1odn3Qn9B4fmDibRYRCJ4+REElPLixp5Y4E6z722ny+kgn
JY1AiOSP3ZrEJHs13KknZp0UuE+m48qdLj/2KS93ZEYcM3dXEv5rb0MbpMeKoi8efsWWG/v4UtCh
CyC9P4DD1Z8LgAC2yPZvc81Y77BEUv3RyYsh6z4EP0Mg30RQJ1tjRTmm37lRVgRxq+WNvQopTehD
5REK1lap+wf1ZYtPzYx8FdldmhT/SIWALZUbqTo6X0UdJPY/EDVBkuiHsxEY8PqCkJE3JahIvywV
Ii4FpBh0XA/MMT8PYdOhSpMP1ea5JbUtOkngGW9XVY5PwhxiyFN4T0TwQpHAebdlK5pZSacI1xSt
ZavWo0Ey4WwhYic/niHESeAnwnY24xNgvf+Sg9a7xGveDdMJZPxkOjinxkXg4ACinHzxmMSs8qK6
jBo/dG82hBRxmHxhTgBhbh+y53y8jH2xrY1LjBoVmiwS+W8PKw0Wwq0LwquOJaCSBx8K2pkomJmS
u9qBKg3es/8zeZISd/SAiZgb/sHDiIpMkELzNVEZCqPzhEXMimObinlxAQbKoE/GwWKmSwpjKc57
OXQ3HXaOzsEbF1GtR0LqQ0k59Y909Kfg5qSsbIrQN5hM/vH5Cem7qn3DvPnQwrNbQOsV7IkvvLLG
Bwn99Slpmz73f4bxUs2f/5OLfBc1XhtA6TMp1TreL1PDSSy6DXMlMaMkHkINqJaD97SFgn4zAgTD
WTnPPtbegU01jxzY7ZAo0nCYtjXbrs4IZXQBWaF/qbUNbMa741tZojDLT4qCk3cMqiAOgKMJ4n51
PBHZqA01eivyGWykHswtkiha0S+mYmCQS/jvurJzyY1TAkslmGTUEzp/StyjA3QJD1s+koZuU9dC
tJH9Ba+6dIm6JEWZLeHexbmwxfvBUm8l+LtRKQfxgoyAS4VsG1zCYvdqIPTJiaI/kHF2sDfCW+Vc
FuqNhDtlpy/3cfRmmGjTGCRYKo5dUCgiyXhjkGJOlaXf5UdssmiSQ+F6M4gupqFn5xO6NwzPISgi
U1W9JH8Cuhi4OGt7kDV8/D/VOhoxjvqM45uT+dpOZ/0uUb80q3Nh428Mg0BbRXu/HXl9qMSOcr99
vb6c8QJ0oohXeQGT5A4McZLdUHCadD9AI91Fk/PHhrBfFFwjFQVmqWt1mgVY/2an/pcjNPXtNMga
pYVIUp1q7oJGuUdcFYM98QwBM3cB8zCLOVrfh6wySJMzaHYi7+OUZ6HprtF13cJS0RdahPeZ+cnA
cjTe4Hl/A4zKXzLiimP+RMcGj5jLVCQIU0okC2vh8PxH11qMyo2QsTMJfnvTQaxOlMQQJI/7Omjb
XHnPnQeGkI2/a1IDBJrXZMjQxUTd927tQLKprsxvPkJoJNmLe8W6mmGAeSNzyMBfExn5bQVxXIsb
7NYRLBNLmLuX+NE3666+wbG3takmvg5AZxm7jt7vtZu3/6SMYn/Dy61hIpO9yw4CFVm5sSOy0b3Q
2gNGCngatNMaVueuxRBDs9qVJdXVWU9djouVqvntcEI2GCjBYEaT2AS8ZQloJDhoKauDFokNctR8
ZlrAw7rTY+pLuCqxqaPwRC/X9KnpztIn/EKBzqg1+KG5bDsTwwAGEDbvF5+K9x6CjXHk3SLm7iwZ
dOezwDw69ixocgKs6tinY3bx4Owg9wjaY16sD+TiDdFDt+M7Pg7p0P7PWj+PublxSEYVIASivn8T
pjrtY21HYupTzmKKItMshmBKQ0aa8qECHvcZqBHj4EiEAABVQrEFFV+N+/fzn31LX5oXVDoloHBI
UneVX6QA8MgE1Q1dkK2LCX+snLZydUtG9MQQ/3yxkSTQlzT8SJlPY8qmQpRNWBgm56M0LE3rmQVM
+lB/s/yK7sLZXkcvCO1KkYovmXkq/JL0dv6+fur7lJ+jpmqxdCK2+OdkBH340ntBX1owhToXyRcV
2ShefUB4b1p3dSADwv1IUzQfQ6/nmuNSIhYfhyQkXDvTjS2BDB3JJ91g/2I8gm7yyDwVLstQHeDP
Hp1J082KY6oPY/sKcoRtMqwqlSBpQYHUUQqnHkisKnIwh8d0Y1CLLNX2et5TW019pVp3kP3wBiYt
TUWw84/i9TimfZlAR8gWiTiXWRfQ5N72UGKEc0JrovGZo3xu8YBoxjOVIoWx9y7TFvyQ+vh2vPFX
S3jacad/ZNyCDbNKPs1XqyqaPBpLTY7I2CpII5lqPEHsTarafkyFysfF0+PMyPHrRXdpQpIIyuVE
JWCj1vcDyUv2cZ2maRsBliwAWhGywNltyvkhhIXUD99mvAj8Pwg+i0GL40XP2Gvq37GW7Y0IM/TP
xLxlp6X1w0UJ18LDMewnE0vnCuIdzoNmqUypPgkMX8IpE9Ifhdeqfl2XN+8KeIwUgHsqS39Qiztb
BO/TXTQDxrVAhMultsVqAWmdZJVamWR/yrls8N+mVj3iAbni3yg3J8HFrZftTgJ91lU9kxuKBMoe
45rHoV9Hp1ZZUxPdP4xjH6W2qFeAJHkT9JDPUkAYC99E447ShYjmX5ekSGZirHp1F9xcevbuXcvT
HDqvT9pnYMrW+r7rwJ8c65qf6jjBn5yH1Ra0VhtbSJ5hUZzzlgFM7hBplN5T9UzOhKVh92PqAouS
gstkyFIRnq6gvYqfjty3LKBL56nBMyzMdMQ4sW84zszs+dQ/DPvu6TTt/5qzOQT2MtVBZo7gccKN
TkH9LN5P832qYfxw9PbqSvLWoZuDe/akWvfcdvrQhff5sEBcuW2eeggELc8szdND0ai13SVjUCA9
JzT4yKN5gndFuY7XFwHULzLmYAfb5fezuCK3Y64ebqoZ0jKgt2tOldeaL7SMQL5zovWsGt7FXJpd
d6DsXAQI3oNXPh5xcEbwiboMcIQJ1E9JwGvNLXeIXYnaSIq3V2pHw92xxHMdpP4GH7b3jSf4n12u
TSns2sCIjpzpP4Ccafc5hVYZBFij+gNAb449zqYdCw2942rJoo22idkvdd853Lk69M+Wist4O8Ab
fU5ErTpqD7YTpgKC7oQkQwq0OzmpLH8glf8oY0bGYraWjdJa+LNGOCKgz/7BLu5d//qnYV0s8NfZ
cwqV0mhmiHZEvRWW6TqWGxnhaW4ykarRUZKeJ90n30TAy/jAsElc3PqRtB9RaGAa+rodN9TZFkJI
Zp+Y331ZQb3B8TDZL0CEShDKg7/EpIf1TAPlsvJFBzZyhr+1DVq3aCpTGkkzAGtBoEFaDzuhtKAt
JE4qJE0DPEGI3KjRFuJ7tgkPzSzs60Dd7H3r7IPVmaCP48FO8EFLHSGt/dJiXeFiyqjrgruh41UJ
ONaB35fwe0G8o/oCAnlzzpxIIafggL7yPINEf4xtJ1bzHitHktu1ehYw1urZMWhVjkGUZNlUWV1g
W5wr1X4cXpC22csIbT+RE3pv5zStHiOk1O5/LzImQv8he2Ph//245gvSDWbITsEgORJtYvhlFX0l
dp2uF0lIKZocR2kDkrHvCnV4k7+BG1p9IhkfudkuCIJXqHEdHxiCxaBX5rRuY3+ui8h1c2QaSvCR
VFiiM1hJNFYhagx0M9PMmXATxtOknYTk0mlDG7N1B0Tr88tcWpUj5kjrVBDdDr0mtXJHWTBzMIIH
tdzobRaiyV0hIAsbSLD8eogUxvrGNTXujq+/iFQCBO3RucB0qQAwj89nOsClwPYAdhIrdMQ7Pm9r
MckNre7uC1d6l1FojmEqUA4Z05PHIKyEbSZeT/pXoxKCV2tVdWQPysotnRMwFVSsY+iCquI4jYXr
pVR1o4s5tT2Gw7b0+Q1Dhw8mzVENEW9y8D2YqxRQ2ICC3chk8XL1Xx/XjQ0/8w2wnZ65rMphClMe
rGrhPF2tcSQl/CCmE2eZxSyT+x5pETz0xs+2KyGXAsp1bFSetb3HCAxv0z5HBzTKhYq1+nINpfuZ
wO5tlsYr6YLMRFicrHPekwdnPVZ+92A/nq0ExMGilL56xXUPY0tlxol32lh+vRJPrfbaMbHpohjF
yg7yy6PQNiHgez8+H/F+QJ5QQYJGup48jnuBeOy0YNNNoHmMR7pZmlyGfoiNj4oM498i7fITrhj5
nauW/64WbhQYXs3VhAlUXmYn2JIprvO0ks2U5ugZjT5qooENQgQn5ypAutdvLOJiFcvto6O2PKv1
aBg5uqrRjTJfVT3/SZlh4DC2YaM2oq+ohgVw471LJsdd/iexs5RU6v01Z/w4jKzMtXKJJuoLtfj5
OXvlK4+JY0PZG2AGbIG8QwbhGZ02w2MbizP2UxKR1MxYD3MfDs10L40uMGMMlj9jvEfumOYgMPsv
EtdOn8e6KmFosebpvRI9Mu5kR3FRfRz2vH5M78iGlcwXhJiFygdivSpXPOtthQo1ukCMPcNfDu8W
VVbjs1WdJWxCrUElEHTJsufmg+H36DkJqi1zI6exC/JJpseJlOZG5Z7vzMfmrXgIX60K0lIm659y
IwWGgx3hn3luwwwx0XHleCFj3XW3nCbavuEYvE0JihwZ4fILBnoyfd1JtqlxqjwN7MDraOgmWPij
9NCuVb6u3rQ9RAfWMv1E1YwfJyf/bwSr4OwmavLrG4zg5eXbHJv3P90KILcEtvqtBHGCevixP2k7
UPjPjzUwzFrYe5wdc73Y34RuaCmjKpQ/qwzo1HDhCbzDW0rfa7lTvjZ6qP5cEeXjmSqQ9vUFUWd3
rltWyS45Fl3PaAocrMwYxHwwtBINs3X/xj74MnGudkUcxKblKtPsSF0MCBfvNMrZflo1hJojMIr/
AaSw/9pm1Y3A8YnFsGYsFi8tJL5xXiC0ERJ18mztPUX4acrh7KUetwDGS/uucfeDojJisK4B4xA3
5f8UOTP7LydKHHF4yAOUaAXid+YLdp2IRrISkJ5Zih4POqRWRVbJZ45/gcfBDVuQsWJs527RtJkJ
gbkDGFlUS6vkril+Ab8TPILLG2ADAALg1/fX5x4qsr9RFM5+6SRd5aPwcqzjRzvWa8Ua7u26zjnp
P2ULoJtWmMrhXrPxfhOpBwsE0i+gJb6XFx2k1qtTmaLPzuJ7LgjBwuKO+q7+PuqLB/UMPZS9aZ/S
J8yWV8PeNRGGAaLqwhS3TcJ2HagGquYUT2Gs3vmekWWMW2hpDLGjnDbeTFWDjR0IrS2Yf5ash21m
s1K76D519KjaqN3tvoD14urIpk/bR6vv0ZI7qiPY41Bq3OoAkB7CBeJHydLkDsedLE/rhW/2aMpd
sglx86IbbwkA3ScK9XBJKilcyYn/iM2RkOt7bBT9lA0CZo81B+/oYWvn32FwXNgA+zSeed2CG3sD
Ty/g/TCyWx1GKTSfI46CTyRopsC25yX7gicKVJuwDW8LeqYAVtU7LzhfgLyqnoQajwdtw/X7pSNn
hxOwih8xLw5YW4RcoRJLE0Zi9rQNHUJFfVFRVywN1Qi5QCLXnuN3GnK+++liAvXEvpvAjTtub8pe
n9varsXgYfR3OLkihn4KrjoxnAyA7Yh63HUCd4WcunbEitMMp+Js9j+4NssG/M+c2poo7gQi8fKK
W+yTTN8Eq3aRgPb14cqLEEHXKmM2qKq3oWxHhIsuBcW/mUUU2WNECM/sYDoH9zxTaqY6o7tzc4Kb
FTle2j0UkE1HYalM4PZZ5X2WingL47JYcUXwH2MWWTSf0HxW7bLFt6RwJRFiH1leqJJoRKElUqe3
XahCJ8HoE+H/aXO/iiCJ8sUMNp0DClqCmA6W/M3/AsmKxkDDxoQynPgzIdsM9OckUQ9iEN42LDOI
hjBkNKcrc0JG+KhyZyy30i1UtVjpogKhxg/cKt1hUjcQi3jOfv0sh1ozn+uQHInykDNfhf6t++65
c7+UlouTsdXTjyJ9DYaHCUyC9ZDJdmpC1NCBrti5aDhykg/VJtI00F9RDtagmeOpRSdHt+03FDxV
MMFBj45Vkjy/Zrigh2qZHOq1OB4K4oXNdpmGvVmJ85tGyIP8fsLQDeBLVRH2UsV1Sir12nsKA4A2
KQet11I1Bos3idLoje8b2kavElCgr9OaRSX/doPxEe0aBvSFh4T4EU3ewOA2fuRTuagVutw/MHrz
6NtTs2yMCQbs2X0Bdk/ooNLawdRwXwpQMUsSNz1UJl1uML/NiIPEAoaDeExxhAZmCvacxmJHOhLG
o69ia/IDh+E0vhsvcDGrxUas0RXkP3tppGCvy2i/a21IX1P86UOIOM+JDTxlRtMhcXEO4l+cSd/p
KaGwF3njkqweHN7U5UqQUoeYlP9bJvcWqQjq+lhZRN24OQpL9qAMsTgoc056z/T+6yPtQJho3xB1
1LgSqbXxMIu1/pe+F2jVB0X7aZ9lbh0GLKsmBaY3edhtxDptpgZlpODcGleuNOsyaVy3JMPoIvGO
lVNXTzKZhaOUKWQEdko4e/VpMsAFbBNGl5IzOi8TSnmHscmdNRTYpSw4LLUWWJT6C5fn0bWlQADG
NStXS6VH4Az0aD5kr0Hsqtmf2ZEnFhqFfD3nlD9+CjOLJ+NCNi2FeNjzU14i1EYf2BLlHNBSdW3p
ldxffg0ffmHuNuO9rCPguLe64TupSsJ0+Q+5jM2K1OjysO41UmrChMCwIpw/0xetg+DhYaOOUim1
FdtGIzIZeKCN1QvaF2vZAv01kdv7pTmVtM1Epva1fvfElI1a4054JRbKuTWMa/cU/nf3cgWZF7Dj
oQVrYzo6f/piN3Wjrf8bgW0p3eXFHUeCPRXmXVj3TtK3WqOvZ8Cg01LyUuba7mp3k9CLfAjbX18S
LErLwhzB1c9LAUCH0A/8XxtlLLzTB1NvLm4ezbtuRACXTUOFWguFOVpM71apwYaumFqjC6sJQK/A
DeTXoJu10C31rVT/GBl7FeN65NXscLbgQmK201YIyjONLpX8JkbVISGstsbFj1mO9QAhxB3ZGmxn
MgvloXG6MTT2WhtRIXilIPkeDvS5a+AFv5LmYXQK2VvHmWs/W4ogdvLYwkjvh7skuuHOVjUGD1kW
ZjSywGQOCaMFfLeLDZHkzeI0xfyXjaRW/rIggVa+stumO5Wl1dYQTzkmIRez5hxLTtWc7Wlr93iY
02zj+lmQsLPkKGuwS9eBPM2FvVMLVO9cMjCXA8v56dzrw0Hc36Z2q9kauwtQ8apM5rcGFJ1HTL0E
7+9Fj4F0tzGMYvtA6LrCwUafKhGOKJMiEeRyp1CRlBvNBwDOM746+5jHbOfeBk3icyt8nzVbsgjU
MWAkMQ8759PER1tTSIZbF9i9+nCUr4573RNawFs4BGsjgsicTJRapJGOApx2iDP0RooZThj2VLfx
jDpddJn9xRMhvU3e0DejnGM7mQAZ0uKSyILmx0CBETGdOqsFGGcr4HnCxIhXBdq3cY2bu8Kvos8n
3qBkf4TXkyr9ygAlaCnUk1mWaGGijkasYq0Sma8nwCB0YOhjX+VUgCNmvFVsHzBThj6ZJVYO5QYA
Twlh5Rj6yKlMBxvQtx9WeWdZNBDCaweTADKcYJfeWWqCF4EeUUSVlKUZR92OfH0C3uRYcgHn0Dwf
XXBo8i6+iM3XlvRgNVDzDM3JWJNGu+L5iOjpFbS25I/MaJNAmQ1n7R3z21s3dR1wwHaSSJHcLJzI
+A39KCn4X7YseqweOTqXjJ9FTV/DdLIPHkNO3ejdnG8ebfKZNDGRVcY7xNZYnRK02/FPGW2uhKe+
v3jHHBcy3LtoyB48yN13g/Riyiap/CjrU2a4aIFImrDF8tG1iLKqwL55GN8bCFjjNd9D1eNRjtib
dOJVl3LCWHst4XVnY5d5k+TfnP+78Ugmpq+W292FrqRg9biykZlKesR48T07ZiGLg4q94EvuOKfn
MUe2LFJoVD6H6Vn49s7Y14QWPN/LDhQpu3bn4F6d5ee9gcMYKrj678nnPax39mVe4755j5WhK2dV
eWlEiDDDfpQxc5aazPS6PixUj9xpDyBwx1XzTKJm3XPITJd3J3lVs4eo23x54ckUxqtbgQh9my3f
7cpvXa9odF2v6Xh6rbPCLSOpFeQIHMho1C5RaohhJhEh5dvvG/7i1kZ9kaBjTC9YlehXV8LDscBp
Mx5DJmKVW3YM8dI0uMHLymM+n8FdZijzCUMLR/jKRwh7VdBwViQ5MY5grunARPaG4ZAyPil5rrhy
wvT0gUNQlxa8eT8rityXGFRAsLBT3pwAzo07oAC5RanaGqCzfSCG03KD/Js8qKD/unueuytNB/1T
Jn0w/oT62qihTaQrgLSDV/canzF/ehlQ5r4+56ddJR/V6jMhtaYD1FGwrt6MpGpI5doFRWmLvrmY
ROXs81dTs975e0UCjzvADRte5KMHFy8XEX+gNrz5CdPKp0+5BBN1cwocZNS7BU5YmHnfHDdSJiaG
PASJ3560F4jcZ6IaBdBvxCVNSGkYFJZVbJVbvtzlm3AApHv+lHRFbyycO6kVOiJANOwzg9qDa2br
MqNnuDCTprl77HFaqbF4u7YnK9IjTZiBHCoVJpn5wf5pITWb4CdLuscn8f+6xVRSE8PX2YN/ezOr
UVZy4lTDrRmgpL738pz9eKbGD0RhZHo8byWNiVADjeXn5PsGM4L7qEtrAf2Py5MLi4P+WjouPqtM
iaLaysrrrSw2Wb8xmqI2aSsQ8x5WA23wPlkhMe+fVDhpQfOXDR74r6DkuyB8R1TELkfUlHc4S0nt
kG3FlK2aad6K34Miy0nqFp3qmJGGy2UAq6k6M7TVyIxon8jYX4MI7dvbgD7r+njjmcYQHUoR4KL7
yxigfcyPQ5xPJelLec8bXJaJagYKczCi1xftnXygvFf19busATrfS9r/fVlDqZZDhW5kZaQ+usxB
Nb9Bx2rZ+lCHf4suVdNqkgb9tbesPVY1SYPXUyYoYMYaYjYoh+WLWKh5VWrdD2+WPMUoTZ0aNtDX
OWZ8GiARs4DaqZNJt8+/+PMICOrz/ioDvzBHS7ETLL02SmHb3rPwEAgBrnAF+j/uNfsip/crLqvI
BAP8HJws8ezyFLj8pxl1IiKV7HDXuIt1BzaYrX1vAtru53b4z5/bF7vBPFXsA9UZneSwifhvaeLQ
r3UuwNpJkyGk/62biHmhRPofX38aJL/G9Jf4tWeb66KOoMOcdfi9R8zfqfcdsT2iUFrS6HA43nRm
uLXMFpUAUKSiCPhgYGJ9oCdOeRe7ctcLs7RAHU0U/RvCXyvsnEHAyZ5e++VmMbrxEMqNu+Vap+OS
vWVlrExYv3C0sfRxNEm0YDrEcx/2+/97QtmbjR/kQ2c4cOZJ3X0pO0BPahyhdqYL474D452vsBXg
2/VOgZFiZPlA5xGMaRjdE7nXhRLdP3OsUWqJzBkWIrhhcbBTiBXwU8YCAIEJek+4KFocstg0oqyj
KmVVwYTSic3hgU8B1gdbAzeOBybe4BrtfTIj1J14CTvF9Gszekw9qmKw01HuVZ+iHmsbkfoJ2k2i
Gzgz8UNHcR/TEo3wYnOjMZQRRjfu/C7wJqg23SYsyoujF3LMDgTQw3yNd4S/wSHBbDtvI5Nh6ja6
wH4B+duUxZ6xC4xxud44kVVKBzlM6udjCQCrTfmoJRmuTSgYw/XpTudJHL0GqLXlOYVuy6Z/f7TQ
qfKEYI3fJdfys/y8hhAtaUBXRzblbCfRsC6GBoTQwmxD/mlTxDTutG09jzLVq51GdJaUPLVCkSe8
X4rp9/+9Q8WUITegYnJ7/c8Zv2m2gKzxOBZo8A65oryzl6FnvrMX+Obbj/h3k0J+I2SbgkMdq7vY
ceo1ZbUrSX5knYbHUBmPZ2vyb6eTlWLBVb2PGspiqnGWfO7o0T/OELxw8+tXWpE4liVYOKuLUrXt
+neLDIEb+Qh3l7WzcIsEs0k4oFFVZEU8Bf0xwqYzTUdbTGu8VBXxmoEgiutZTAYeJfnc+bjOtMcL
1CM3jqF7eGiTGY3EO3CO9TGuoOVLeNrcdSbpAAMtZwq8IiJANQSRexvPr5ashy/iXZa8uq8h8hGL
OW1WPrjWlEOuF2U2NI/ELlpIkmvXRHwWYQW5gFI2vdpXmARWOx8M9ZHY99WJEDWpg2yjgZ+SZO4r
bLQwnJaEth2RBOy8oRAe/hIZwfK8Ql2XDV6HnzsVo5sBCf4x25JPu0FfuaP4ofrGV1f/zzmG8eBX
8JK9o9sBA8FetX0WLZASfb8fgLpxxSEDW7Fw+Wb2gUEW/49hUeiGsxTcDKMqIY5p4MkdPjQ8+IpT
IidQuDCqam69ZtJVCqUqKVcdf/+JkcfX71xNBIa+SrlsrvGlhvnnPG0oNGRNFjVB2TRqztQTTDpR
YeRtPDXuv9KIf/gYMZZiCJX746drcbOoWdPJxMqG6JJmFFozytKLS0V/tdHuk7DXiyEEe1D869GL
0IVQLO6rQcs+P9CkbEuy+3ek4fGZpFAEI50mE2Tdv3ooXAeBeGACqrCLf4lsKn8KFmxoJqASE2eF
P5up/bu46+/VnGodG9FtUg3VtaJzTfhrLvQi9KtC3UFZH7RINxojylrFVuDmwzn2sAAT1BKURdOV
plVW0zrh0jgKFmBtWzN7cpENDlcHur7pTd2ae4OcyUljiqYxhNjuux+5hAR58ui1gAvyGcwleR1x
pcIE2LqfllMX8l/I0UEQ5f8PTKwO5cWvZeSJ+o5DvQN1EE4FPMA0qCkcsMpHUQL2ol7yso5J+qpJ
/a56aKIOSIR4W8kGKry0FXgI17zcgriZOLhOaEgJF9nzFnM32RO7YE9i2JLjSvsPiqrZREzPwip0
rm9v0ekDZEET4IvtxwiPvLvxJAJ9GjNRnlpTEL2JufO/A6KojML8Y6tiBQIQpaYH7E5hpfg+vaCW
xdSnernUPGmWhy8sOxKKZRNjJcxcCxRRunEGEeMMMx3zrD7nWVD+BSjpIlp1JPuZrcatI6Vdh0w5
HkRsCD6Li8eN73cvtsi13G45ltGaf8ynH5rcqVCxrRPuWYynoLQ2E++7Zlyps+lJ8Ed7SdUFhOdd
alhqy3aRCHkD4IshBeQhk4k4HOec7HCBWk9Hcn53QV88vStQwNFkeM6Y5Dm26vyRmgqEy4jJIP4r
3DX0GSwKrzCpUy5XLkRtcfw6FyZLoeRWN/aQFPdNzvTHHTsAgobaGmr1jmJdtx9bh8S4ojKrxIdu
FVaDulJ1IMBCHaHnPfMi93eX3OCmsx+wAoQ613p9QTmqRdT6dUBAb86RvqdUgVaA+7JdHs/VHDtg
5zOI4qTQiriFG1QezqsLTcKzbrL62vWZZ2d88FDrFbGsV0Ow9fOrf+D+Jm1tt/LS9Zq95fwbRXzw
qQDqgbZSgxLTmfFd5Adcu4k2OFhlFwINxPaSxP2frqJkl4uR9AK9+x2r7QvlrM9+vP/vIV5QFafy
kxnBakohNFG+71XaY1b2xZXcF43I2HmbRn/bsl05Z9Vc6TJn7o20ABWwe5tjhYmbC4qotKWMn0ql
dcIVcrZIwPMlfUi+VoOcX8ZVd4Bhl13lMsQ9xnSar8xu2Dq5xK9TOTE8t2gYXG5T0jhGAaE/2+0B
w6ISNyrc2hdXj9n9kdqp2DI0922lZgOajZr1ZudfsC8Ho6lqSS58BXLc2rBwZNXJeCMuPh1Ng5Wm
d8BZ5+V+vO9FvU10xLuBfwn96qv0uqiZv6cp3UBzytYl39tJgAPmx6QtVFH9tYSRaRCIHVmgvqiE
qQrRpa0t4LsO6LXhVncP4m3XW7OJoby0+nE7MeGGsCWNlQ5qaL55SbDfAov9Ky70auxm0R5OBfXH
n/uFGy8fJBdUJMiXFCp4f/wQ/ovxGT5rQkxaGGA2nSN2VGSm737LriMYeV+dPiFiYIz6twSw5Hbl
w/so2Nx0V+tq7zJI0bFQDiCT2ZrtRcafjYs3ZYbiHn608PefWRUIsZ0decum2xVtX5RchHPsZ08u
B0qaM568sGdlLGNGBdTsm+uEgn8Ry0TzoEU1lv4rOp3QlhNANiOKYE0sf2yGIvwFxpvZ9+lX/hZs
X5AjpqkqArjWAh6O0ucdos+KLNSyvOGSpN9wHYVfYs5Xo8waM5XqbzIF8ygNr0nhjdMmefC8Kgnl
grjdPmqLJxQAiK4xwcKFXG4Cgtyxb80vsVeWp0jTxHbQxacfF4+UCnXnNvolVy8Yp3bNOFlLwyph
BQflAe1OOpbk0rY2O/bJzkzH3yhKuhzGwILnaUoPIl6UqSAK4KSBjG05HrKw47tf2XF+THsgAGWE
XBMqm9C0PdzWWV5gIzREZ11RLP1nSmPi9qoD+fpNUBk4QDgW4a7kkC6s1DKbGGKFpayP4K48zjkB
VDtUnkcDq5biIiWTsFE34tJImg575giSRNLKN3e8qh9csMhDC+gXVJ9b5dHcicIwGMGsKYwdcBUF
tvnI65d5n33JszzP1TyX9qkVEoSEXryVJP7yG264Zm50+qEd7hxttxH1h64Il6tP/JhwIFOlf1IN
BqsR4HhPiadrPPRsNlakDmADh3KReqFuvOnIHhVjsxz8OlC024vQMuX6ZWN9oQtVgOd5aKo260vT
E67iyxtFdwzH+/GTUyIvUsxPsrEUpVOMB1UOBbNrcDZmionkSTcvQHHCZ7YhQgEopacsmrb0MO+6
MwgePneZM1qSDz5CldTHls77htTyFXZuUuA3a230xGZOdb0I5Vwxis9BvNdGL30cHyaZJqDXzxut
uEqhcqNXvgxTJLbiA4W6rLRoZpFeKcs6SKZEn2XqfUWxD1wnP4xZYTA6yV0cj5V77RpNIWv53zKu
KBiqUTC627bOuYoIFdKA2pnZrtxGFRNwzVACgRnPsNutK/FLLlPW5bdGhpT6fR2sNO8ZHvst3LWn
SOzQRZwEkLy6a74M4Fodpg1BrcR+vaZo3y0nMy/t5O4g9pe6pClnjGoLtH/CPY/Vg14KyntCOcCM
XXOiSAeZ1ywFQKe4/C2JffUV5h0wKW8mB7pCk5KgjMWKPkOvWVaRlTqALJj+o35Qhu6Mt62PjB0c
soUyjZ/nyJizDBMJYn5TMJqzbfFZyxFta02CQinYPuDGkZsqastia1SzBwxD7nVOgblkSrlISjia
/8lbTAaA5VHb+q+KjJpEPH/5RnlPUGDg4QkTbWX50ml0kkbCOALB5+BL1HwsF6Oc/nyZ1GOkGWzP
zUDZeq2CWKuMGRoWtWmk8jrEEMQQnJnScVOyELAIQQEnTdvj8Xy+OiX5on4W1W3iMlksI2UAdQOR
RuD2ChYjBfeSyNIGZXgTJF4YasABwrmf5kdClKPRbijN0fWkSVTT+nTLAUh9mKOtWo9zxEgw8r2a
plm3E6Zbne8H4sfNzn7nERkGu/mvCjeGAm6hNtyhcQSFc9kPbf4WeUM0CDHEIPhv0TZMo59Elbpa
eoxhcgJ1WDXDoJuHFEYi6tpboFmk1/E5jJJvinjlS9AEYb2qOtJ9EXdw7JXacNLYwQICMYUKc9rn
Q00CeQkExfxipkUO1YkaX9fkeRCtUyBE9ZUzOP5PWZLHRT2G39IMGAmx6GpnAFIKc0h2tERHHcYB
jwYxCY5eXUVhmkizxI7Muo28lM+bTWsSu/U+bNGD91qu6Q752YCEXL/XLJl8TnzkGl+/8ybLZI3f
5x9J90c6AoVHlcgl/sjBCfxFDPZjNHx4ll+tJACRKfsY/RcgeVZcncEqus4sfI5MjAnCt/ZTmKyY
hTTg/tTAuokymOoT9+rSaH3GVQ6PSvINBd4U6Hd1VA085zSVPeOy/jKQPLV4w63W75Ha+8qywOhH
5BfvXBPsahjzgc4yECY5FqIQp/n8PQ0VJ10HG9rMSOt8vMU5ewYLwGOAYNxuqposgmDu8MZBbGK5
Lwg9dELu55CyQ6NKOLNtHKWgjDOU5gQCbNxCZGcIJbzVOpxPoSB9WF80oiRdOu1vw9kr5GL57cvH
yd1BY6IKT9JFMNlq9MXvELxAvNRTPTLVw3kgvVnKuuvoxwsKx7KrWHGbnYcrOlDB8F6/BunxjpIe
QFSiSoLfbyWDU0bzlk2fenPh/kNuPJztXA+wb9n4tmwaZRWxE2NtbxC+1R+wtatIVyPzPG8HSqbj
SUeoiTibv7n2Ca4xr7KQb4ManUQeXn1WRUGrwR5VMTX3SulYB+niXPKbwNB5dlFWxG9yBePC8VSg
gT6ugOYuRtyvJTKl7VLhFUVbOCxOvhCGARhwqhlMReKiGTQb66QaOotDsEF5fHs/A9Mk1ltrxIC8
oXwxO71tfrJUs78vDtJ1OfsbdxTli8ioJBVdprHODbhKicKnrQKNJErWnE1rVGRPf/gFbKSyJQus
hAWckDruGv4zfK83sme8sKyv0PV+qqayRu+ZhNj7wDDEyZHbrB9yc3gQRFEnH3IP2jcX4ZDOCCa6
0UL53hkip9bl8jhMzTu/5UhoXitl8qXMjxojQNtKLiNU4sNtcfgeqMZqc52WE8P/3Ss3lMVKOMfJ
uYtMAA2WwZHIKbnNwsmmPVzdt5I2QJOfwhTf1q0cYblYgzRpT9QduPsxQhnAbnOXI93h1wVR4Cna
3LIeBBHoT6bpH6rD0a+I+K0aLsPQLe1/nFsE1Kzgp1REqkgjCgnmEB2hbxdRn2TQkL2VBijGacns
SGL9Ns58KTv/w4rdYx+eIGt29odD4aNm7zbOQOgA2F/RGSiUUojD6R3To4CbCJDguKYAI+uRYZ6q
D9Kfj2cY9SiRg7Qa/9sjJbmgS3CdZyynTsC78bzHSihgYkKcr3FSL9WvCDfk9iyrkb1cZ99rTxGZ
85rglukTjOahGwbJFcjxbWa5WV4iy1rnYADDGO07NyPcNr7fOHocfG+1w40OLfyE9X4O6KxlPGe9
NrYOSgileC+DwsAG6bj83VAWnzRSWM49/HGkk9oeLM0porLx1SPhF/3iL2b0f3/kOKKZrvz9n+Zb
olTKbXZdi5cjwhVAGZQL4WmphKcJiFi6LdtCNbkeVeCaKZMSwg1du1k96ek/J7ILssPCOuDjoujx
UBAhjK93YlSUFpbZ0R2i1z/xZt9/VibBY0ZobbjkVcH0qKQLyk0VCYqXNB6PV1u9UddO4IcSnPNx
PzKRkPCqccgkQ971QqUYdK19l4WR3mSbgWITum5K/kV0wHx33Y5Z/tEQgYM8hBa7VQco91cztJI0
lW1LqHmAfjBMShp4B+fYfaTZ8HrgEhGyz/JIwuCcby3nc6MDltMZ7lnR23gBGfkw73HOFJ5FfHR7
5UobFvNOhEpsGCV5X8Bxwxb+TCyBTx2ondOJEeZfk6WrDIdpxBp+vtiKlBfpoC03LiF1Lxuhybet
mhdacCjyZoCDM+fvulBixJpCeI27LnES4wehysZwhXLILdXR/0nuJPktBfCU3cea9CqkIZNmZ+ge
ASnkDLglvmIcTXwGjcsP1zgS1F+jYDTw1tCHK3AJxh0uUKGA26SrBpNA/KrjMAq8Thj0LHzFkDiF
AqmZujpZeGPTbti1+yB7LqjqVF1BKBRR6IeX87/LelhArtQr84oNHLd4gGia/hKgyBpK95AwLUW7
75F5ytFar7Z48fJi6rWBBfi0eKU2eL54/hlr157ohxZvraHY/tRzJiTKz9Nj5j8tDjVDbE/ElSkb
yIY5/B+ZIppW1WYRui4omEx/pXrL6tluqBpLd2poQQ8oZPMv6Rn6DWrJIWa1uKdTLqrZkN7HTEve
EUKuNavegPaVIMVdnVSJJmWuh7UrSuEYqu9wfbEpXD1ivL4kGLHJOdA6pQb8sXiT0yGKjKEvSCaf
m+2G3kUqQQdyhE9sD/+NnuvDfzltuNti0L60uuT29EZNhjyQHOlL9fJh4idQDBTDxbUIcPOEQ7Or
ZjcwnCw6odidmgLqJHSIo8vKxXl2qoYSrfsUEcxmB1c8ZFkIx9qwjOsTLk1f734aR4xahlf7hiTc
MSzg0Lp89mZue7VGl0dry3l7+9h0DKY41oqKNWDUjMrl6JV6wHSW0wRlxF4/1LyXo7c4BgNeMk5B
A7TRxq1dQm6yybaX9Z9EMelv0LFmsHrLjGccaMfpfn/PRzp39s/phhrKzuYEfBTpVm10GbMmdzK9
wY7ZDOiF4CrnMvvWHOMxmrsFvSo2e5p5BzmTRCXO7awJ7ZKrWTNgjlajbE2wrXWunbko9pyMSNnx
zeHbsFvcY5o8/kmNuYfADIeMk7bouQaxlQM4yutmHwnSIDeLrHWjQy2QsvdlrAkVAek+N0JQBiIA
4Eb0xDjMbez3STAjM4ZjMUXwxHcbMMhj1vqMkWFf9DghJ5xf5Cyig2L0eGYGrgwI1ydM2WcKJCNl
oBiU6/CSJCpUjw2Qrr0aw7tt7TjLkCk2fUYJXuL7KS8objX5Weladt00Ppd/YQsPqz6bgcb6+tqk
Pcaj9XwSGZIFRxnqiWPT9/Zd6NTZebFVPold1eELSFn2xID6YkRqahkG7jf21BTQL2S9KZp3LW+h
+HFkOeWQ+LDdG388JeBo0BZFFBZ69OdbBbi58EMatAJRACpV0PNEjg7pL7Owr/F6BHVdbTP8d2UD
G91FrxftVnE3D4tGimyI47hEzRY74Bfxy2rIOeQO9SmhD+B+lhinYa3YaKMka72PVYgj6FBFY1Wl
gpPmrSBWE9WGdDtY/Xxz2u6uSypJei8S1zdUAxdLcxjR/4EqoVqFMV0/8gKxXhygnOX7o1SNiN9b
E/3pbOmuOSRjn9AowBrqNWEWRl0YqwR3f0LD9fYMaoL0FFWddpZ2xNQrFK8RmygYi6aBAEMZWpyG
AK34t6gzIFV/LgPBqm5EC8tduWSgEL52q14mBJ2gLqza/nli4aXRUyjzwQk/TjGR5zJXahDpGVNO
QfQc58B7QfcSkNl2aZnO7crq5u/lssmoZBdADyx7DRkPYET5hBaiKr6jRgSiDUbGPYbZIJ7DNUuE
iwcfHgQOekunFAudkVcWlEl4rTsqg+L6So6GpYo6ogNGTV5o/+yLitSSomrraNB6UaoEYTNvd16T
3MWD3OH35d52Oh/LVG5DbxgILFdD4fwwvwv20EUqZiYhMzBNGzJakD11QGGZs+Bk81HVQZbAnzJI
3TkfrNf8GncVNfkVwM8vXZF+EAcZHdVcQU2xYDeaVqI7QWUCYRvQeNICNZ6KekMbr09QvNsGqezT
sfvYG31CbD+y2FYCAYmXdc4tcBx+VnixzYUAzW+L4gOyiVzQXo4pVAbKK1pGE3hCTJif4w+WanlN
1/I5CRFoUtg/i29Xzq/0uhWXFUvuNUiH9dCBB0eOBtjAZhljUT76y2RGVAB2LWjcwt7rYcGMm54e
bwCfnG6r0RkN+FDuaTx/avEHeHKhNiYVJK+K5EpGC9DukZrGUJ/Rl2rEl7WiypfxLdXGpKVMyvPd
O+0DbZirNaUzhoBmGUq3tgzW9raEHSrV+hINtFSM2enFJDWKpvOF659XezxzhfJhKsIF2UO3iv1y
k3ciGXhI3Iza0nWSt1/Z3hbdkOtJNr2AO3LFxnAeOVEfj++Ag3qhR59syCdwQqq5eLFa2Ftg66BT
pt648UZBEj4LJEDG+prJBGs1Oc8rWLGJJ4uTxTI/znprWUZ073H/B31Ce+1KPzE26QmofCTPwOYG
mygKQI3hAJYNDwaoxNmpskS8GWeqqodec5wRlomnU+GzvDaniM2DnWWSAeYx+Lv3czz2RO5/DPFG
DSJtj2OY10uMJcBWzRHhBapIb0oFYPIVC/7xwbxE+aN92oWo1xaciYTnjIctTx2hsD9v9n6RhxDq
pIzOMzfkZHH6QuiqCmOkCB5Km7BmIjzYW1xMSPDQDE8em8bmTRWPAkZ9RXjsbWxwgn7gkKcyWDr8
3gEAACqvijXcezM7p6x+yf1yaAdCilgLGDtLJzh181s1uxnifED+2ZIRsHStDk8umz4LY9nuDvyU
C8I/WsYBwNd6+L5vRPwZvcwvbsW43Re921kMTwSSa4luqxjgNIFsDR4N1RzV3NhC8tfjxs5PYX+y
kfBu1ed7otegXe/8sG2EHpCMRLIvcsNBVc2gZp/vVFO0fFL1UVxNGd6lKKsR7GBJegVSKUYmCvHi
w75lE+QAELCSLekkMc0YDnjiKTcJDuYGltLLUlWS82sCopfwmcsDSOvMnXkLoeEzgzFOptkHHnqU
RMyVij4dk7c3qUogc9LAurYF/N0TrxvMK+ZYkS50Z4X/D5mCntITaN1zclPM1JwLcZap4weTU4Iz
+ceHBm521YAnB2aAQVwgIz/1aoL5+BUvYoSSBSnnZ7NMu+mBiiYmGwpa+G8qoNmLxC76U/rRCP8J
TXZB4hq/jqXzbppj/UMHsibavBYH7/bEn9Tj4E9x5zmATq/JSz/FAk2L6GyesYKzSz1ACPsJGWw5
cvgZ+gt+uxnmY/yQ2rc/mBRNpijm7oUb848DMLdZlV8NrpKgUSTsOtDCULGiQxyIJSrgFrx1imG3
B1w7o63gh3Iqf10Ms/1LZtJQmk9vFD3ecfJl7b33GKitX8wDx5iJd57QQ/7V16l2BTItP5OSkFG3
hVLTU63UZqTX+9LCQYlsIDbFPql2MAEfoG7kQG7UsVZ8PUk3jaWTo8tAdPcjoKosm5C2ExWaBIKI
tQPV17oDlHeQbmMGO5wPt9tEROfR6cIeNwLR78Dofbzjloq6Dp4BG7bvQVSMVVOkm5IwKcIlRE4O
CDYHFQdnHURrAJKGMpAOT1bMs7ZUcfVnK4upR87H0s/R08eAKTb88Kee0MhMRJhlks1G19KstAVN
8iExEoddFOVENvPcoJuNs9MzGZLu4noA6SV6gPJXZN0Qpv0NFOdcSeBFDtUtm378SQkIon5AYE6m
1xQ6AFpk4oZ0iG3noa3ROGeXT8OjSNuu+GrckSRFQYcLNkRXE44NgZdMPM8nJJTrWUg+9vrWdE8M
2sVTgDbBbPfRcGpA/YbB1Fc4qZSTZQsz0KFCkvD6R96qlGbC70z41WaBihrSioLj9N4WorKHNs+B
Fd3QeG0b4JUDR19m9yDQ9YHrNBoeu28zhFD+Y0ycfXhspaVm4Vwoe3lDS/jh+h8BTxueo1CS/WAd
FqliKpM7M1hMxvpqzUfuJBQY3IDfPJ7hvyO7hZc0aczZGrHSaywHwZGR9qHFTF8jwMmy2nBu+uKu
t77ZiqxrEmoyks26Wq9iVtvDioAwlQXcMslk6J18BMUerkHC2TPRe8fRFtRtKirly8gwyUrKBcEy
cOFR0+tma9GVRGiCcMQ2NEAI8yhUsh8557AVb3AwyQCXXFbW1RUFEZGWJVdbWN6rb248C2rMt4Ay
nbXGqUKXjXSdKzNzev3MZRypFjc7ktnaYPElW3evzv+yB7DVx4GqfuVHLuZztZoORMXgSq4XkpVS
6UQEU3n++j6Cb50g2gcw1HKv1JJIH7tYTixPFKqjaXkaoqdnK0llSihmvcjHHm8VxKkcsHTweRvQ
qeubMkulbL+b+uZO9P1+H/nbaHvHiHfAgkfLYscREMO761iKsdhOgwglnNtwohCUbYofHElrB1LY
qlqmZqmf6eVbk8shJDu+iCFdmipw0dfRmtivkfc9CR6fUugTx/b8vRx0yn1ppi4x9fORaY6ejbGv
SrC4orZkyLOCWaYzj+Fq0xvQrmZS9tmr+Ab8wGLgtG/ugNdaa8L1TH9TJASkFiwPXwJwFLY4Cv7k
5I3R4O3iMwzVnDPXpDpJDR5/De83ob4nyXB2csRUYKDP7T8X9MXX8sl7e7EjE8+tugBnFThReNi/
f7iIDgy14m4eVVRvMMN1GzdhQNrT1oXULaB5R2o/1rt9kICkIJq9NSN/lH0eRz8L6baxlTbkuvRO
DRXu7/joWESyj58am0n7u3jtl0mDRPOdIwjPTqd4p8srTh/WlJJmafj9sN9Yf0bsYra8OyhEcC9n
7CYcaGNGUBJPbTqzAE50ZNnhF8up52jcfvvqSy6ePJDcaODPXhhljMjx+zSzJaukIcGxDh/5H0El
/Qv4P39fHJ+09qr0tdzY3ksm3gb4w2P1FJowwKBUTEdgftbDrc+wgLnI45Y/3Mw2FIb9dp3bX6YE
8OlI+6cFSdRMstsExodL37Oem+jpDQ0BbQzMUKm2Le+YuBCKChut7a1miLQS3TGkKu7fknIfv1O9
0M1z5eZYZ90Ix3oVWd6za4ioFDlM9pw9whNs6znfEuYV83/o6EvaN++IDl0grK3FGzWwkBNb5Y3L
x/DNbKDUnMsXCaPkRhWb/gOpS9X5Ead9SEkvD4H8LoKEA53ttxArOxfc/e0jQ1a8L96KcYk2o1fa
0/jf1/pYpejmQJerxNyhG4PJQbIkCzmdkTz61l8MZgssoXClFNZU+euynFFgJO2+ns/6duvc49wQ
77FWVfM0Rw3zlUbF5txCtgyQroCuzMfrwqyT0P32GA9wdg/WcC+ydGMsaV0IIaiSOfACkhbgwJ2t
emo3KvaP2S2QPfdlKNSj7i2hMeTsaU9EzuNXGlODlQZgsyLx3wAW/qavfQDX23y4CWNc9SCimNeh
P2hzXoKPkf9tjkzGAxvLrWLaoBVIfRLIIRUMmXL23MoPo+Rf9docvdmxKZhIyQuLjoNtgd77b6oy
XmnsIS8Lit1kauy7XfozGMtzGWkjcxL0OC9UuFLfSPLYj0glqWQw4fN9BIjgQIo9XAmJHA+fqz+U
8KChqlQ6RGIU+EUgK5Glbmq70YRtzvRUO0C9wygEZQscc1m/e7C8TDRJRS3LEVDOoCSIYDX7PqIn
9w3aM2IDzZEGTMs4ULe78UXwirpzALmtVmvRaWfBFG6KO8txken2T9QWYo9EPlbUfvZn640UcX6O
0wVDH64DdfRkhr1G3j3iGFYQ6Q3TPlUEm3s2cdX2tNjz7xayVLFTeugR6U4HAVhtao6uhrAz5BoL
LbKiwMqj+ecMkWf343Syg3dEGZ/z7u8DTAhok6Ed/x7qRZL3PharsNnNsaKhW11VtDyioDrhoZGr
salCwC6bZPYXcMePhAyVVD9ZlWL0/T3Qv2ZAWT1WLtOfTqKKpETVosvM8k3kZyT6R1QM1JJ0nlGZ
ay+X9aEkJW0CGSfUdlz1foJY6vRZHagTjh7JXNPibKp3PNar8bS8NrrZYY61ch29YfHzo+ZBPChr
yve5+X8aHHUVceL3scXfneuKfVPGaC+iBdTl7Ex9ZM2GtM0mjxFS/6QRDzGQVVbz2UNo3aLYPcpY
Ak4MQ4u1kcBjCMjq8znEPvBj2tRB8HvN73HSJRFyEPe7IHz3G1GEXTq9v6qdoKmOF9VbIaHfQtaK
M1sc9u9dt8P2y8UDfZADR6/5WkZZRWLuCKhAr7D/SHJIVz7I4OBD8ZWdJU9yxYkFPAm2tqI9A+O3
76zeRLRPa0XlcLMfUp5tCgFWCqFRjlPTeVoWn9v6JB0gA2Eq4bZZoQK3qVl47d2gTjL8TPo2EOdN
1IfJlSvQSJ3gMhF0Uurk4QLwmcOwWj/Mk2DIY4SYlk1ybStVaC70b+kCLRy8HMBQxo3zBBH1Fesx
9xkodIGge9gjqQq5Cpxa9Ca6fbLbaKr52haaUz+Xd38paObvADi8Kq2rLM2qphM9boolMNkF9ed+
X51+tHXJaKxKefis7PFFYUMGrjrjyaBfRNk/NKjwJNvNDxwAnfMn+cJSOJdQLvs7UeHtivCtlZPy
LwveHCBdYQPj8xDoNAAFo8MWcDjI4fBr4s/GwQ1iJn8kAh0qtK71zX/m3R6UjQjv0h2XV4AgLGGx
98NsdyjmqG3VW52D7TqQbjHm4jYm8a6wNnzmbBugXf5fCag3dKTFkb+2D0QZ8vJ+FwCvu6nhrLAk
i/mlDg4frZIKFO+Gh4JRboLMlLs25OEpVDmcS/5JOQiBAe82KQt3BP9+rWQj2VZyIqN5Y8Xz2KTz
wn7u5sfXkjNWu7j437Hq5cSky9ajszYw0xIeV/Vs8u4UbELR4WJmiMl4wOifhn4lbGTyOM+NJzwq
V50bcSQfXCZiDKrUel4Xt1zxVnsumwuMqGsOyT4olqx02CDuYSal09Q7JJVvVRnhmteQi1GVhR22
8AZrUtLW6NqAQ5ibHNQld3D3L5GiGABu7+kT4dEEVbnx2SXHEkP0QMANeDyAnyGNeLa99GXmA/q9
0D5OgjPVn5aG3QenVxpj79VDtEjaYLjBEFcypSPsOiXMMCMvbuRimJLdfwe8wvwrIOXEPsGMseFI
lMnPy/7E2o4yI9ZCzFM8SmhZKlmcwevZKgCS6C7H/aNMnAz5vio9eSO8d+/ryIDaOP3+pxkbfbNI
S0SuW+iU6XG+CFs15abnP3CjqZJUJxi2MwDoNxtxANec17VGUWxHdMnSKDS4de5bp+FzZgrhVzTf
sB1MgLGhAVkYfTBBJR4Tx6AijjflNvbKxxnI/EJWqW7Ruvnknqh8w2tj2xlVlFBbZCUvVpZh+VJU
thegXL2nzAcYSLi2lvzgT9djYpkMVgyakP20cmPyclrclHfWP28pmqtl4VIuaM9ZztnJRxbf0fRW
ym+4QNYAd+gvrpAg0I9Uyf0XLv72oY0pHQPTEu2qkFwkm3K6EyCrbJhfp08hxrqijg753Ocnce4L
aNiO+6qasIyiKzTGrEpUQyGYZNR1jwV29MehctDhs5OiS6fTfZSArOs5nkF8cunUVluVtOrv/VWS
9o3luVA+M9Fn/dCfQCWZ285Am0+c4exhrtv1nM8hhAmmAq8czhkqEqfjlAreQBfwCPNafG3nfnao
1Fh3wIwbU3XXyGofgkMojKqJzdQ+7RsDgSfwSpPDNfrOy0M7yJf1x0eLIN9uotTNvEMfn/iO6fsT
9Q83nsfFSBAQUn//f2lm03wPYxfn3hGEFw6j3L/CWUVNgrhtbdRfQKtdUq4C9a10Ro5AZCOCjjVE
DScJqLE+ScsPNBhZTPS4vC0YSaRG2K2GOinZKZIgNJK1e0uTjxvGRBVDuVeWYMUCRa44IY7ij3+v
+6YtKwv1V0AwSwVjiZaLfnjNp9/RMtAJ+XZWQnuXyka/98vuwGGKtiv8gh9cZWCAix7mbC1FnR7C
eRlMYU4jXXsD4z49p+lL6nRn3huXoKJF+u5g4t/dL5TDqjp11v5eMBFjbi40pYhgtqUC+EC+35F6
7nFj048GGCX/VMQx3JmuHC5LrC+JBg3lRVFtq9u2e1DCfIUUYzyvYNyDb6krrzpJ0l0m4PRH5928
KNbv+fd57otI0CvavrGxBy+4QSZLd+IPcdNeepIYUeiKm4MnotZlLDQfjaaIMM5/tcjoLUSLjXkm
6cKkQbMCMeuzZnInmQVd47swLERu0HD+ZHr4sYChstHnWXPZz43lrjKDGUZDHTNh6FXA7x6MPqus
p5rDO4iDMWN1j1jbjQNHgcO1iWghPMB/YA45TZrgX904Tvww0/rfufoY3nXj3wnpRUpjlKlwGFGs
ijE1Sc8RDzAU9gEv+J8OwLZGOIk/CtaURASS/tk7l9ATQ43wOwK1Dz8oOrLXFNn8qDM0IpKhgmsC
EF+dAFbfq0EpzYOAeBG3qzQHDbqmTMOmO6l3dhvF3CRbMAvrqZoaieg1aSGWwa7MXtqLDM4inBoO
5qz6MaD+48zBL2yCZE1Gi5E0CLN8T+LQmogXNz+TYvuhV77ZB7hk2gJnvZA1O9A7oKr5uXthvK1i
A4jpD8Aj1UAOi3HjSteAWp/9subJm3lw698eXm/UJVaysM0drlVWFp3tv0Y1gYW/u4a7yFLztMQj
jn4sokHBS8klbUOFX0jaeYMV+ePo/8pYbRzI73ghFyb9PZbV6vmtWTbQaVXaEPvP8YsjcOhN9gZ9
mWB9yqxXv5xgkrgbe0ErsPDcIOMGgRSnMMwBUw/SIc5mLoWN16MG3EzWJjmSXVMK/OdRNLQjOpUo
BKptkLBUnwsltXzpslxXUDBT7HOVAxWdY68xtZXbqxpBm9TFpejIuXc+6d1NCv8E+5f6TGpP4wHG
96xgz5gecpWSm66dNc0UnaJVD1UU+VJoRd634cntB8gavlclTqNKd9Mpf/NIGzPN27t/RV0/v4Fu
h3My1vghpyBEPvY5jXBT9Cv8XwhzvV2XpQiZxMpWT7hH8kopDhrtA3jL6nEA2dtNlRUpizJ77VSf
P+1ExfPhlGneuTDU50+zsPbss85p9ZhUsS7pVdy78TqqZ+m9RG/Z0bqeigO1e9jIYnfwky/i0NyB
ejOYJ4ORji1mTuIWcLyluOMuM50gDYvmpGSHcNA61P6PwmvyL1fcY49stpi8t2pMKt9o25zciDsz
IaYgBi96AeQKewdC++48BAb/Gq7Pfz/R/gaJ9ETdCHT5ierpl7V7Q+Izk2QA2D6A96K5GtjQzfiQ
/6qtG/c541eQ3otmEOcryy4g3aVj+jwLRC7R2nLfMwDk6f10BD2dZ1FH8pTzjVBD4SIs85oTaIEZ
/0KEpNAhQ/7yyxCmwWfPZLvpCx4yW7M5Syj76UcWvHQ5TQN9psrtY256EPHkq7w6ewTNweqO+lQt
N15N5iXcg/jXX5gRgR2yIsfqb+NJsF99A+Mc26qh+P1Go9XnlysUd8yMLrO1SIP8AzgYENLT5IPF
AdpSLGDyHwwtBwNLCoaqbthEAQWSF2/4dAxix9WL1FsO7f1brZBx9FhcaVWOdXbwaQhrz4/NVn/k
mUTbk7XFBBV8MPqY52et0OHvUBHDM2iJtGurUZ4LlWHAx2sYwio8YEDxAOrTUqsjQ7HgfIDe9vJX
RBKKkTfoSvRhyo4IIcuFM6X3SueTu/Mt2gqAYofTiSEhOqI8HuWWtY4p/E6CfzZlPbpKoIJNLS4P
Bv0jpENi9xKEKV/UbxYXBTgfhG9haiDA0KJpLbDCi17VQo/1zjF7grQc8ONh3ZU6m6I+N1YmipNG
HdJxUJ+RKFLo7s3RTxY5BszMjI6to0tpjEvBVJuSqg/viB4+sfC9T3erA7BQ1X6pBk7qTPvKVgP3
L9jCj9I3h+6hFur7JwwkRBqQxKGku5/dbP5M9AOVSlPI6GSCesDm0SMKb7fs5GQxVyBPj89BOjfL
alN3tWb6E9xCpXR7GLIiLJrh+sWnVz1PXA4bY2O6Ptv03+uKma44SbqNKrXJUZGb4/QZWWkz3q8x
Lm/4DKhKAZe9gjT1w7SDXJx8Q/sr/2bXaVFs6Ao6IUCf6tnYCrxeamhDjeQoq1+CNDpmGAzYfFzO
DABr/zZhqQ+CebiNmYE0f269Of0K8FHZjPcHZhFa95XXy0nr18sXuD4ngC8S7rEcdOAjthWvYZ/U
EbUskvFfcAHq1d623bgDIryRtx5Lhd6FftUBOP3iea4ug30MZjMZcZnW5yAU96zdpDILD7DXMYTN
5Ul7xIMcjZtsZGDf286hzqoXSg9TX2DnQW8MBAFe36a1ZzBdpHD6BypLxHn+/gAMqrVs/QPXapvn
SQi/eDcsjKXKLTA97KSYY/wNXm54w1Gy61ivrEKLaadcgwXbu0FOQIIGNlwx5Lu0h+dSdeKBavn9
kzsUasAJrM5NcQ8rj4Z3mkvoAhC+ldVpqr4a1QnLBpPv8gPFXUW/AnJITn3ZQv63YZZqJgdgClW8
qSBQZAsPAC0BPSo8xVOtzjSVhtLoYH5lDFlQcQ5p8GomJXn8wwUPBbJ+XlYvGUsi8SkrnanG0h7c
WAKOXH7wcK4OnO7ufVHTsnY9bujNRV5qo/yx50rZsmHdUt+rpGbEHsjy1bE4plaT5GNHCM0z9Oxi
EUQHg8f60Okxl8rUCdLu/FGpfDVNdqKMJ8OQ9hzOxCm4E+fkfyBEVxwCjRIL/BdTvchzRHioHX0f
ysqkPj7RXE1sPyiwN2hTLGB8YYn8ZuqTqLa/2+5sQnrNoEXZEcOhyjl937hawRxjOvwL1q5Qv+Ao
+ZUN297vLDz0iEsD1dZ9vtT3ACIyiDa9Byg7G/p6VUiXyfkKIL/PomfTsAje88kNAb8zSWNMk4II
M/wKZRUZgBdwQ9YxsqLIxuveN1YMeqKF3IzbBWJp4sbt7pHJla86GL3L6gFQTOT7T3ObzqvWPGjZ
7ytSRQTSz8sBxLW+DrRgf4tDSDe3zNBNSTbeoa4jfAT5BQZC5SWL27xUaBLbcA6iXBX80aR/tq2U
amzRyTiGvUxNqi16OMxwktWL+H5rSDJUv5nm4tagE8BqfTxNZsIP63H0ZDmvQBQuAMjpX8TO+FsS
swrDOouk/ouu6rxuJncMgMhdBASaY0mfo986tsoIljK2tGu2voWKEaDahg9/sPmOwx8hiV+QGqEl
gulTkc2Dc2Gme6E69GAtxKAX1+fnsFMN6qA1XBIZTK6dWO66UJdaYQJJlIqqCJZwFMa98uBzhSss
mQeily9dvFIlMAFYBP7H/0d9B8gMHd2Bot5fi2j6/dl8EVvrZHwlNWVYBpr9W/lEiT3WuzcPbe/l
3UlH/1uYPr1GdUlpwvJJWGpAz5QiEO0ZpgQsEzCIttjeTr8qwSMnnq17gT7gvAeo7tUitV4z/Duj
DpazHng1PgcWZsMXUfCbAeRzNRSqOpkU6gBLKTmtVFVWKgTopSFlSoyjwbOiOKylXjY/nLUekd/7
p+zqLYlkj6+4s9NG2qJGKwosnO2GOtdfUTWYIOQzMtXIAcWKfd9qWItujKScRSbtnxQpaDJuuk5v
jw1nwHNmM4t7HC6fCnoPsMlY9muP79slKqPvZO6J2B5FoBOpAUItkKxhOpLODhkatP+TsJrEgxjm
fS/O7A4tuSU848CU2zjJmu0R588k1mh29c2hcAGNcHXUnodcof3BGe5vnd7Zxkg+bNzDwjmYJ/fd
UpOKfdVT7r7YaWpap/hGHhbLdtsxlOa6ZWxa6/QFgtJZY9NzCDjWml+Dxh8uyz9r5fyJwV6zup+C
/IFwcJzY1qyrcamoF46uf6asJyxKs3r9zKbN/LsttPdArulwhRUnOB5j8e6tCpDTKhcvfo6fRCja
1Q38+x2UIXrrr3IQIOR9e5vdF5gvaz7dS9Agaug7B/mOk8FdWI7G3wvXGBWZgEKL2CWlJVPaFNx9
UJmtVMwjt64kd0lLgecA/X8lvf93xPqi+zt6zVj4A/2QqRNkgi63SKh4k9zMK7d0D9+7GjFhmUVH
7uTAON8v0Xg3lcv4bLlmueWB0BTSzOMAtKdd+XWeNZ5jWURyXK5E/sJWaM+hvvztwSduKxDCdlHt
pHWtsXrJaPC83UG5xzqyJVYqj2eJl3kCEUDM8cVzd3KuIYr77jehYrcK28e3ctWg7IIyziFyfwaQ
77f8l8wUAH25Gmg35pDN4yDmjwH0Qx1A0+KyaUy9kYBwg99IF9lkfGaSbbZ76gQo0IeMfs/78mcS
y6SNR3s1rAGNjHVtAQ7sz+h7jXFHQJ0goieSnWPzrMi8qx7NzRoZrbzKH6DT5MmWwuDlDOtueEco
LAzGKSx/Sj+KCzgkIr0Z5yokV2z13BJGjmqTtYI2/NzeDwi/+dRuU3wu8OeA8u4v7utR3F5aKRZA
3VHtrZ3xT481ppCrBj0EtiBXyzbRpOQz87cTKRDpABvEbSLp0SlzX8fgHA3+cSagc/3lgXTRf08e
edkzn85IOUSMl8ysFiIigk0tQsMo+JIYcRuSVWJthOoMGglGw34uoGgEiI5yAYdI7eTJd6w7o0ku
SgYPMpyZEtIMgkmnwGkasTSBhuDDE2EBs+j7zc34ZPMLx2F20/BYD5QwZCy+8eKMEHVM/Z1BepBQ
SkC5QI88lmsD8ins1iZiqV2lccfyq4IQ8e5OciFTLWbJm4GJ0MtMIxGuf5VLOPlq1uYMLUmdvA1i
wIaSRWRHwdd5F8nyH2Y/LvO1YB15JjebyQihhkjptba5lEmKoQsLRtWTToAwKcFbyNk2wchvHAsC
OdGlzTVnIU8To6sPe4KdEPVaShaGMMlr/83F0CGFRDsrRpJz+cb1GaSh8ZFg5BpKOiwdCaCP3Ihp
ZRUegCaJlkYvxgvB1iHbdqSG8OUx5CAlbWWPTpR6WimOVCD4fW49TmSTbUjH5x5sg79UY6dK1vDj
bscd11u0RLAkwTp3m43JATBE9+JkwUm5YCqrBDMdu51xR27kciWDHB5IPkAmLXJgTDQCsAY593++
dfRJVDBCpkyOM8sJn5vQh0czyAIo8uwCXxvVjk6DKfIDk/SLGbOMxrESx1TlRDO/Zhh5omBUulSt
WpXKbWeO+jhATVapKyQhhIOoBS53grHt4SjgZj4B5DO8Af2FzjG88jz0yKRnf2EZXZZ+9BpyKwM2
SE0/hai6oWELYgIQRZiJlsq6TqcKOVyKLvOMB5qbYsTe7ADBMXn4a/JkjZfxo7ouTgjZUMKlOEab
Vt83WDFs9BG7elW7m9dPePkgLeINjeg+wm2AyrHJiQbb2kwsjjMNtVbaqSTQ4KSeZHQdtywcrFNp
KoE0FDdcj7un9Q6eFs2imqhX4GjHovCYmP8ndLHYC0YVDvTM28gOQPDKZSlo/tIDymRR8MLQg4eZ
oDOfqnR1apjus8DYQBYJkD+SoOxgiNEcC46dETlH7pHBcA+hjeFqUaQpsXeCTuNTuaT1OnXLdaVC
bs598TBef+bm5xaDqb+93KGIG6vVM0zD8wtx+1SaWtvfqiWca1wiZfeqNGHAivQwblZrM+kY03lU
jNWqQHJXpk46dJ31IMoGK/cAOnraqSuLXM0n1pijUOvZkxmK7hn/d01xULhlnFyLgn0rBOODN5H/
PT+/agcjcTZviqwnkZkOCv/pN9+BtEQ/zOXi327pe0+7aL8boKQDNmaTX9JK/znhRYDJoI3k1eiZ
wmer7PkHqcwIzBBZCkwfOacdnTPPap25As8GGjttlr7EOrHek95BX+XeQwJIqtVKqJEb5T3Pttpl
7DXS53CEs94PtSB8ss27SCX+3CVu7ktrlGNCelLxSjA8Gaj3dE6980ffrmpuK5WweSQcrJK2jnnh
EpICn55AHfb7sG5PnC0FkVsx3+PYtY2ia5nK6CHeYMkqVkC6Of114FBvUCO+M9zmDSyff0LkKZ/6
5BKtL0s2Uc2A4z6noaYVgD0S6mtQVb5nPH8fyjmTlXUseVsjHReyD4crZU77b0LjZm3PEyzLJx0y
i2PcTNNV15B1DKoIUtVzoWXfwjKa1ZV8DuDnUE3N2TiQ+Yr+xeUEOH2VLG4xascndW4Q2rGgBBP3
TAYaplANY/VSSVrksBXrUJRL1pXC88Wow/uC1msGJBqCXtYhuYWbv5yn1LxfNhMuyCQpg8mjO1pD
hvMjshokomR87FJ+8pLx4KmxdPsTNKKVRF+fNraQLAQzptFI0ecSCXl1RnShqqlQ7ISrj1Wk50K4
7Uw5H91F79qRoH5Wwl0LIQ16oTBOo3aMeIIYWQCv1cBDn5GgK6GEYV0nAppBegBN6lny17VsMVR/
J4RY02xxc/vDDkjzZSwD21/bWUZe7h9AkzsAO8e604fSpQnFKjsYoiMgV7Q+FdxRVY9qY+4ckynt
OfHAFh16xlxs+UZBYBSFJOckQfDvvlf+mylQLTU2b+rzDjxm/hDP82gt6OBDXdkCGZgACtWiM1dJ
FjK5ul5iWf1GhE1mlkrPn+Pazor4nmpbT8u1IN2HshLmYKQrwakCCE7LobhYfKZZAk5JJT1c8pDL
r9Juwjox5Xjgaspc1kmOeqn6DwLUFrUnCOa3dcYLUH+HcKmWGoC0oc3TtFOnWYLkd1dz+TLYU8b6
RY9Z9RG98csAkpSFyjUsirSe2Y/tARJY8lrpjRwUTySw3t7zcFKcrU4EIz6HEH8ro8dLb8dsPieb
ykyNDBm2tnzhFhNmXehlie7a3N9uuLu9T9US/tG5OD+HXvveSWWvLQ3vYb812e0G6HYz6aXF+lO/
lLoJ4/V+YVPzRIL36jo/aVgoL4JnhbKju0gvKE1ob9FZQu7+JgkJsnoufDU0/uyWCfyv76aYURg0
JGAaMc62iRXxDArLjbnz5itL4DOkAozOUnsM1jQerCAzwl4PiUkoO2SB5MY31vE201BcpjbV+lh3
KzCwCeyhOVT4rwCEPjFc24Kp9YkC4SZ2FjAKXq8cks7X9+0BF3QKrQlbrsI/asdpeLFhoLEOgcFG
O0qNwrAPVR70RUzn+4VmADz9CzyLXzCNmy1oYweyjXZ8uOFecwWy+cnAZO5HOI01uImGNC8yRBBz
mJRV5dKxG++2iv0/RJv+VdGj7zolAQATMi9ikZ6Djibs/5g+P2vIT2ZE8NhM/wy6UUQ2O6sh5guT
S/9MX20RfB1R3k5bIB34VAqNiKun4USRGspIrWC1BoH73fJpNjhsSCqCTpQyM0rYam5yJO/r/wEg
yx3AdMW4wlYM/Gieg/vqtMBTdTeiQY5IlwszuyDWieEDcHlDxS0jc+iTHzm//+8vbyW5UV1Tdexp
Z9Uq1dGUh4+uzL+KPb8T8J6WJI/E125lvVLWvPfRArFSysMYwROM0riXwLopsrOMkwa3htDZp75r
1zYL0oKyEz9+Jo9uFPIM8Kq6FWH4XHTf2JzvrZHLy/xrQjH0OdWiBNgH1DcikKgUcp0yuq8bA9d7
X5SqP+JwI9p+Tz5ozHw4im7uvpyAZaiOsjTvp00N16JDY8uMDAyC0J7wPWZ2x5H3wafrfWiE8K/h
wZheQK+kOH7Bpfwbhc7XKchlUvxgDe8lNRbeKYX2JxlSdWBLc/B+oKW7tmfmtAuRfXLvu2ycebe7
CV19ghgtgyWbb9yPOLpRDY57Zkrei8fv1htA0TmaYqP4gcBrLQitDWt8TWaqyjQm0Pv0NNoy8smU
Z0E/NLj20rFS/bBoUJpAAlDZ9HkUCI2nfMYucjytoiMLoIR77Re6GX83urdvLX+5HYVZLyPmGH7F
oTT1ZBJyxCN4RrW8xekQ10M95esHRAhlEOXlVHitBSvWYnDewYYSXh1qKalkSxgXywOzia9XP201
ojUY5pU4j7af7OkEuDto8kW/bA49MAuA/QN0bKy63cXJyuCICit0Itvfc4ff8gX1Biu/rSPN2TTt
WHVUD3xwxCT36oj5nXUU1GAuWmhLBjXhKeKRUjMN5YtZmCvdVA5Ahz9XHbqP4TZCAhYRjZvLHd2o
IjnZzK9qO3etEZycvYgnGK2PcDKx6fUNC1bF3j232VfAY2JmwiIlS+FbKYcv7Obx9Z0FqmXGdkMa
J+qFEd36Wa3RPci0Cb37rUNQimclnEIleV/83nALZAWcW25Pnii+E7fkml8UqDt0hW8xL4VC9Fzk
IkGXEWzP6lPMQqr+F+aG14trhsgVIPOVUuk/lod2gHqO1y9pWbvjgtIPKOmw2Yjj2gcgYxj7Yi11
ccKuEwBlZM08yveXrPySn3lyGJfyjIRpRCPkIethqx03a7UHzDUtFsjSxxg+xzBe5jo0zpLcq/jn
iI3WkrnEygnMqCKiJWQ5WGjZSBQ/dFEQ4hMw6PNRvBFQwIhAfBWpvsq1LeBxI4wuF8icBYfCi3MK
slpgqlOp5F3ooJEG13HFxWljRufsC+ib19DKwFjy6MT+hKSiHxpSHOeIgeBIa38GrWQedCSuKIf/
C1V4+y09lGbovkmsOKfuQOHozJO9Pt09ueLeRcRR9A04DSOmKIMZt53W2dwq7xcRA3OxSLHRGfiB
MXEb/mYOBAt73gb/JYWT2axeiSzJ61Tz/cAuiLyaGOMim9D9N9TsAaxSUEQrXwGAHpSYrjggawR7
bcSRs3UuXavvzMYFXPc752RVeFiRK2s189a3YyVHcmZ1ywZZend0iqDrcC2OZoJhvuHHB1CLj/RO
2NvUpV8BmkvSlVYLUElXIr1dM2HF4ALXrr1rBpTb54GSy/q2y+mLH/6UPabG1hQOZfv9QTIphRxo
j/za2Oh8i9w4hmPSKP21kit2Ew6EbmZCOrkxIfADzpoUHWdxhCWmuypPuwFldrdXHiVhbfoUiKYi
NIAPbjs+1MlJOZ84NFTeeoopuSk0yAZqPUAKJYrs8mhRQERr1cKwg9RgFpCJUtQrvzaPdbhFHNJ0
g3sR5qfsTCT5AlUwCTqZ6yzGHgB+DpqciRn9lBUgPP0/fSrr/cqpPIjTu0URZ3pTuf4nHnwkcmAu
zeYEsDwBRUJABm5LVT3g/71MNMoMtj1zWY1MmLSWM3MThXy9X58Ge2wEE2XC4Z4SlV+geijE1CWT
jATwvhiBJ7nm9+C609PD3OSRlkk8OOFjozI1j+leNQzKxnGUHeTjGplluDCtc15RN9rNCaE606bw
vtnzdyqrQW9DZQEAu/JAt+PazxvL1kCqh090w0Xn8hSQAWXIrA12Zm+Kd1lLjUD+E7TUlPWvn8Lt
JmjqvfPaxX34kaU7/EsUJOmZO/QqllFFG7l2YdT1n6uSAGEF6K2aXLn+WciUl1OCbZtGagr4gHsV
E7wra9s8iVyEV76XqdqEjcWtY1IJF9bJ3VIxzb5ewoVIB0a9Rnk6gDq7wWPYkG4XwrNIBxVUAWDG
Xxj5QQNfv6iPLNLzzrj/kOscrLsKVL1XktmwSd3Jt9oA9ND+bwMNYwvDD/WP7bN7//5pn8yRAVOD
2ZcP2FGlzQ1cg5cpaKV6TDAjM2dTyiZjFenDKlzR+qgL7dmsedox4rJkUVDJMscFtUCJEMGBy9SS
7UfukXGKUaoCcTUTbsd2eE/VzEdenc1iljvWQ+o1+zA0GfEksLg171Ku9Wa2tr7T+rrEMXcaF9m5
Rlh3CfcY6nH/QRJdrQO1/c3NXJ21qC5u1RJc/uXOrn6DYUYq6noTKfTO7vQJak1w425S+MflNRfV
b2fHj7LGg32QVjQERbXCeFgp59MjmZr+t08PVKbRotm32UpApqEaWer6QrQ+a2v60YTDMMfgbj3M
oTvpY3Eg4nHxdNudMQGqQC42mEk62NDniGmw+j+dTyxlAf6FLR43Ga5XYYDDQdUpyakf2+Qiu+vv
Q6WJWhciiSY21RzVVQ9vye0jVynIQhOr2a8zLJDQbKNuCiZD/HdlYjLn/Iv/7wGYj0CdH+v6phXR
Dpz8SlurZ8vjGxE/PNSg87xxzMGNkJN+AebcurtE/NDe1frJKzTF/rmXyUoorM0Cnlb4ZDY7EIEE
CbnwwYNMoNuyW3wKtjeSo0QJoJm7WXiRp9TY+ZUbRUaPVDJWM/Ap2liLTzFeT1cPL6bNxXLISBSb
u6D2jN5SnhIz2UtMZN7IU1wlWTG5mOPta61jEc5KIQWhk2kP3NWkuwVrISaIfmfsSne1LawRlw8G
WcRmyb+aQGk2IZbuVsuW0xKhFh7lSrKRGNbM/AazMHBjLhjwVUTDXvXKz7uzMN1znmHZ7LastMat
/8bPQ8yTdcE3PbAfhzsvn3mSAumwbv/dGSNGb9VFyqn5q1o2rVzGeS4Ob6GDIxgFfAvnJhledVpK
pLhdrsxDfAEBDnXWE3wbYAcShZMo92e++NEarPmJJ6s/HPeH69BKmcHjEM0XlE5DkkGfXFbk981e
6/u/PdfBMDZ3kOyx8HY6AECJvKDTzg5dFnp0WwsWPKrgi1rizTauKXI95TcYL9rqIixywcZXBI/z
mEuyqhyAuhxLQa6NLQD56ts9fY/qGDzvLvueZ4MmSQl22ykeXHW+w7bUqLatxGQpLMqjzb6o9qZ9
CsRcbhxOY06ijTVnBNz5pIZkibZY9DECXaQnUcgFgHe6TRoDqaV6GCvGLzX9eK/3Zmfj9zNi93JE
S4GjC3wXAW++B2n73HWA6LZtbXsXgzf7mIOT7rmn/6BeVdDKTe0YZTM8axXh5RdQbEa/bKUtFfwj
5uXkS+Lr6GqV5T1IVksSkhDZ+L+k3Su/SzS5sBVNlyoHQqKQF7A3q17RoIy1OC/7++ft3jlO8GoJ
3V1ylllzOKKBtjFfNCLiE3lH+pFqRgiEnMSUhMOUqzZ4Z27/xzakKAEdkWvxrnmdUoar089pWn0j
iNG++T30Ax0Nr7fSFYGcmXeyceILkoT7P7vXkB5FaaoRbhRnJmcMxCBNhKCgOELPsZV2M7clzoXB
GrRvHQGSHLVkhwYbj3Sv4PcNg4LABb/PgkJtWH1u2FL0O8vlek59kYBIRgFOS09+eov8WaRMSAmI
hDR3x3UqtuNyS6Ed466qMFFkkKwq1tT66HzN4s0vgQW9861+BI3AHvhJwXjDDMvNIpOeKEfnOHSo
+7TPjs0TbRD6e2P5Yky2xxe3YSQFE5DzQ1ikyG9r6+zLPiD6MROMkjcqhBEbpSa9TCO5r7jP3Jun
+6SK05BXYL9pAcG/Mur2hMDOzOcMti34TvswRUz4Zt9DrDlFDc59XhWoj2gQfEbOSXauYBystJME
5jcJQM4+o1+qwy0S80k5DZb/ZZQJDuvjUjjUNolRhpwDAF88+q8x82ZnQYOJa3n78tcyjdGG5eCm
nbCPEpI/HGKClCXfwFHPesj9ikjwLfjtRfD3HT34zXAsf/plkBcnQIwYE0uwFh90EN7PQ/2P5M1t
eZjpRyBLpSeQcDnUPVM8nUBDHWuVKYEBnLrZqKEPoKuXtCQnY1BrMauaKox/WoJj/1ysvSfnb794
J126Q7EKdtdD0GnmRVbz9tb93ZiFbZvVIUj1ZSJfksndhx2ciIPWDgXUavKCZEJeVFUGCVmznFMC
aVCmTk6yDvCgqHo1uZk2TRzxtZPEUddnM5YhLbysVTnfsBVLJ1cM4kSSGPKhOTHZRcALsEZwuzsV
7dIxfxxDPAyXP/d76RuqUwteUr4DRAaDfoPIknk8626sFlbXRGaEnilD4wxRWUdjKvnNS0iW/Efg
4mkp3V5dJ3Hj9eK2r+WkyBd9X+gq8ED1dSTEYxrKAD3nlFNAlo7vG3zZ3OgKRQmVAM8oipK5fSAi
fjnwAqA3lJ7gLBLINPsih5j8zlF1QhyEEEjUvBltub8KExN9YrRmbo+ANRyb5Ev3JM5PewXH+od2
d2EGjdsm8kIavG8ajIKGRycKXXVj4Tr6u2kWOU3YWJi14wO4SvEACYuDhs6JtffTOa4yt4FjNvGo
xFEHowDVpiDiXKT56w5FIU/tY9vUzy+BnAVrh8YWqhEtD97EMeudA/YrHywZpRcGCfDFbfqAqvAu
BCJMsxAWEvED6/rN8sXan06DJ1POaMXtGXsSAr6z72oStcRuOPNK2QFzilb4M6JhbXQhnn9g4CYC
cpWLuSdidYunseimcJ3TRGPiHxFnP0R0tmupNiFOdaLLMBLYCzAFnwIktCwxG/S2pLsyFwdzLk0q
mGyYGRmB/iP4Bz33iHdgchyHJ0+Tpd0IOl4DbPaM9MCRDGVuNEX0OiiUzc+2NvWpE4+ru0yuSLHR
QyfYiUmk9yBDjGH3Keijsjo2qIsZofloKKiPDjJTZ3bEshrnF6P2UeNW5/nmgBt0Fxjk1L7Vt/x+
W8ywjYvkgS+lfCTKcw3kII6GIWOtiZfU1pzJLRvngxmQVluLbVMh2Z24zh4Sy2828qzP//W6tEmP
gRYp/IVEehMPeMvzoavjX1q/nJcJQqZwXr0hTVE4oNicN6tsqgMkvnD/m45LdTU3iq33zmnWg9Xo
d4X2X9lEFaZBL0irMC1Dgy0UTOPnRPndT05RDNWQ/zO3GHpDEA1np6FZDm7Ufx29MJXFXKTC6I5c
di4GcxHIowRCz2CXXZKevgiQaYNs3UO7I6f3b79kv4ETCKT9L2zZ3rWcC7VKIOrAohcuv7B2nwvp
e3Eg9bbIxiyCvePszfa6PWjHSkcO0YUPoGzdOHAg2zpAGGQp8+jl+HiiEpRDK5KG5uSwDydRsZYb
eaARekmAr7Jjt3egvGGNaNAsD97md2xwaxXAqb2+G13kswero+t3Z1R/qzEDiTGJxjbtjD7eS5dz
NjrEltdKZAa3znmgKFv6bH9xiodedxW+7uhD8/gA/9vkRGIDKAFWGZb2R1bN2M0/5JH9lFxfZ/8u
bP9Q5Kba+XxjH3vLzoHGm1gB9ZS+ZbHi+O4N4kzqJ7jFYO+Fy4V403LJVTACN8i39/mu4VoVFZTN
b07zC4G4RRo6Gr4JtaDUWNTYFNqp5MpUAUOuhmEFftLNKVR4fl2bOi3PKKX1Ptk8EOru0zMJLfaa
D3guDxr2XvuQnXxleZIM7jkwuc6g8yXYouiw9P3SMz2sNzMnjL0v7XanEv63vTvSmhRTvo6S1J4e
2jxeQNBl7CRH9JL8R1j267ilX9M4aj1jQgb78ugsVUBAeD8QSfqouLIIdTUFazDq3djl7kC+EwTZ
zT3yGbIU80wDSyjS36vlKe9CS5VwJwgJcX7pgtmGk4xYCrr2qzqj5b3QKZn5k2KzziorRSqIykE1
6r3y0hVmMjtgxLB4ffq8pdi6+JObau3lJgAGz0vgZbafFr3a4GelMgxHL8Zaq2hmqDHSHZZWcMe0
6i9MfWoX9cUBtZb2eNS+ntcufZJe6oC/XmRf0RjnPZsfix4NFpsVRPH3u0IJ74H0H5vXnyCPlFXV
PeA6lCiY0dZ5trc80vVzZPRA9uIR5/FEAzBBD9RB/2FIY7d+zlkvGCBM1dOwMgbNKwz9g1OFJpnA
LvkrnzOS8JtmhSuXlQvwkQ5Ec/x/2A6rltPJ/Aet68jnidYb7S+tXMij76CY8mFr+71fXPUIov3G
t/oxF6gVmAVcy++IWrplCnplZkLrSrSoiaaZXLPI58o4acJ/6NpyHVN2C5Mi4DoTa6++wAKMU1oJ
dtAAaJptRSIychUj5SMRXGJQhPWwaboZxbanuIXN5IdwsisyxB51uKXWNhALu2eX8WRfpKGOdmKh
C6pk3fannd0Gnyt8Y07BhNUdwbBW++Iy6rvlQBELgs82TerZfMi5WIQXx9ozFdubUurLev1ck8Sz
J9sUzzu4xHlOE+KuC3aMkH0CsHKhKLoKzRJgjs2gM1weQlQ03Uku/b8L9pVaBLXk93SlZTWAIsdx
Czv9rHoeKETYO+LSKWVO3iW52riJuXMOZnpVVUtGoEwM2wMjksCjK8L3Z8FvsIS88+salN0+1dDb
sdGDvKg3AnW08weAwJ+CCqzCpZgsHE/9csyX0GbpU28Lkok2Aj7DOpSOvTS7xO35Xcj208SK5/kj
RNJb8pJ8TRCYO3lAcCuIWJcrr90EQBn8q0f/ShBUQX5YYbQbiQyiR1R2T4WmNNchciwwVDfIihRW
oc11rzkf/jty7MfVgXG4IEUMSBWi9gmCzlt4AjnxIOqNr3a3cRW95X3GdIM2eox685JeI7C/QUD2
MUEIyZqIR/sbtJY/oxMInT0Tbnc7LTHXMlCf5VVjtVJPXdGZ8Sefs/CloEYllkD8JAnM5XFi8evK
Bvq6TPAbXh0QJ8X4o6VK8rCY2Taav6D9w2QHO2tps6kI0WNIwj4pPCmOaIZrlNvvjED+43k2LfIY
8Snjc4N1lFEB7uwRBOERtbB+Zk9I97JBFiCcWHp6hZbT9GEKBeDgnEpbZyGnoF5guAFad6NpKPzm
gHiUwZultR7HExb9FD5Bv3g0YoUpinVQR50Nfo6ucHUFKcimgwlWPwctEQtgcTpAk4GAQz8yGoiP
Z5KWznxjKgj/QudLaRpqUU76s3HnpabCcIyrt5s7//4P67XLO7eSr4Bv+nGjSN/2Zk7tyUF9wf2L
SnnjtQ08A8X6pSB3D9skOFnnST3SpupqWPRWLzBaFx6AGrwv8wlQWYjeztOchEv+yO/XWaYzT+vd
QV7Zvph9Jd+qjPzxGxK4G0cSyT55zfV1MPDRFjvV9+tPoxqWZvtYazJ4Te/KDfIIMtvlAH1b58II
/HBxphgz9rd3WHbsv024UFztiMOkA6+91+SsuPN5fheAmWutw5VC8JvpaXKBmmMVtQilhz0tOhEN
OYWUVRr9OELtWtk0+sQF0kLL5ELCikiGpJKrwYFaLcWVVh3pzQOxpDYkHgSlBo5U/SJWslLrsKK3
WtI2uQmkRjPOMYGbvQYIGbAetFpwKjNaT9oguDw93CoxUojl5f8y/Qvr1CbleE/XUQ8R0DHKQ4dq
6h45hUbqSWA849897Ta611IKZUfpt9vGLj9SdSa50m+RJIrdtlAzVOn2jvuMxhW+/Dvnu0q2mOoz
DqvN05kXxmmuQ6cuG/5c2xfWRg596pQo8UdVLku2haoZ34ynkFblerQfNeaiZa4bXBXMPIXusKGi
omEcSSdfqkPgrGx05dxYzwDx8sPUHJ5a6RTiTdgdcn7d6XW9n9vT0ykYtA0hBlBWbvDxdtd0aM0L
1LSel2QapWntQsjzTRiBg/hq/lnQSd6PATXiMW0IixFtdZNpP4457nISYFooxMBKHc/mJcfYfVTo
DEi9b3mk6VmY4FYFq4wxO7iD74C7lZ45pllM10T6QmwDAj7qVwxgSAzRiM8/C79lhDw01jAQOnW9
2LFHKr2bEU6l//uslCNtUhsD9sKNQYpDMbAgXUVMJMcavlZgvEUrVzUofnMw02YHE+b5GW3jajCq
6QF4ZYYiYvD9tcWpoXFrar2AvtyNpJK9+L0MeYq5yZH0k2YPhPbBcoCqnuQQG7mHEIXNIO5l3h2E
PIwhChbveffc7om3xFpbsilRS2W3gxXkhP5t72NkNHte19xWWjR2ih8dma9jwjDo275qa1jxVghz
zHrGWmmVCYH4wW63tOD8JkWEgzNV39uzy6BopDOHMEHU7dMzGJslVT2bKt7sJZZkbI/gofCg9qaZ
WQwR/wCw8SSOaH4RVD4p5Ctq0u5jri/twhyCyW4oEGtGx+gZFHSdB8yVKDIY2Ha15PIpZ+YFipbK
flCOuH/cy4+HPD4sg0pdMKltfo7j/aJdx1jfjImI7Ma5H29Z+rzLpxs32yg4dK2J73jDFprAnAh6
7FJ31k/q2xJjNUVKelk8KsnvHG6+f2hoYD+gl96sw4o34XDN6ecPxit2JK5e0wogvEBcLC16/YuQ
+86og7QJUHRcrmMy7wZu8FKbJfCzLpNoXp1xgUY9ywpeJvqmqkpfc4RWWQ8ft+XD327SvPzSkVnp
rbCS3+8leb0VbWk25Qsiw27CM9M7MF/sNEIBG4VheagRs9hAQGUHhisO/J/st2vRq7T2BOXF5j7V
JZfZDxNswhYgBYQ+en2R3D0EZ9KVJBm0GQ1ldOHoXNeKfcgWPFJ+B0cvMpsdFGvgrVwkD63uwy2L
GkHeeZLb/4MRQCKywBTfF5TCMgGA2tG4mDVnHpOnwXIHMzvGH7lDyTrFsEd7Aq9m99s7Z/EOOiH4
hTnKJ+QXAi1BqtTqyzxhCJA9Ptwr58svxLx3RLkHCst/mxNvvFKRQRm8qSJ+dqfiVoR6POVB7+ab
++eKsEsed+S9iLfdNi+HZB9i2nj0vnF20beC7lmlRmGV9Ez5U2xnTBppJD46U8LNPzz0u8SwMK8n
/X9H4jOepDHssgPTKE1uOBXIBSz05BR9/t5tN56YsVzogQjGZKq4pOOVHo5upbJa1K+5rIcswtCf
x0Lu7hQ58m9Y+nOslToI/p/OJM389qBUtoYw5KeUqYdJweYWNvPzYC/J0KhlzWSb8BXJyu5WAUsd
j0tJtJ05SiU5D/nh2LVU202qA00jqg4XGbJzM2to0cXPTVY7R/+166oUsE1trTA/yKfEGUTIJNIX
utrzEzt7c8KNjaKf+WSy9Tb+BX9wYoO693u7dlYO690013owXRJQqiiQgmlnmzjTcVDXxhP1NCuk
BcIdXKINhaAOqy3+p4YyqVA39fWjSbEmJmNs8gF9NJfiJ2IZhnHli0AwtM9qldoWGhnflrVUhgX4
tTm7l1qBSaNfSO89jgnEyAXGC5+JUSTsFghy4S/8/mPF3h/8C4z5zQ4XLJ4kdPlcYR2C0rJ8K/S1
sBqISbSC/Gb3a1nQtExDx4Cc0WIhi4HkodMlvV6e7nwTlHwMxsLFOuV68lq1SZvWK3QJzyeBdKg2
4wVl/yiiTHyiSk8LKni1MsVI6lWgZwViKVzW29rRKAPVK7OYchWgstBHKEwKHfCYjgPuYBoK7Qc1
4bli1pJQI8YvnhAxfj7p69Ossy7pZxAlLY3IacJmVf9IJHmr5gNp9/3e7tkidef/POuOfU3UxlGO
KNQeD7r1h376FsZQ+6Js1Bfo6gEEa0Mwb6pSCmL5iOH7B8qi1PH/UTj6inpzrYineAcxjJLfaNrH
El2MNljZVjjItKb6T3mVPqXe3l8Tt+kejDvXMfVB3tWbBgZ/JDxXuazF25olEmzrcWpzSjzk1xAO
T4EAaTnaqrLXHfnFTPzUvJQtRMQqn/SfyybltUpBe2OVgl0fng0qA9w+wGUA+vgithaIDwhlJcOl
EcFaKQvCxOpVYbfmBPcxDH+yi2+NnFnFVtDiUJTp6PmkIbkHd0ksCTQCSUh4JSokrtagpiJxyCyS
+TAYy4bEDfp94RQiDHlC9RM4E7PWmXib0wbE9qcqB/8gdhd/jS3IJmxjaoQazCzpyf9tM/xBlrW7
j3wc65F8q/KAv61ve4xEx1pC+qe4/CtqK+du78m0SnbZB1y2dBSWaiYHkbcNw2Kzsw/vFwdExJVi
xVqPX0zj4YDHHVMwieV0/j7nYVz8HAsRDZQUcv5KvijdZvYNagE65538R1STJ6/2ZCG58L7Omytb
DVgYMgzuVUtmaMcUzwypmh8R6mdggPz3LMSnn93yxvDHQTO2afG8xqHWvVB71aaQzi6SMXEUzqY+
WrKUeTugLumJWCg9Gc5e2XfQXo8xNY5CUcMGihlm+RfPEtCiq9qG0RFIiqKouEVTZvMOq1p1mslq
LACUIdDxalZEnwWlm/Fdw0HPRyHya9frOvdnRkg3x/hsoK66M/eqiob7x3wOXEG/PFcYidcgrVmH
wGnA0ZQJ/mOlOvASymubr+FbfP1LqbG5WPPrTRT6ZY4FGvld0ByVHK8vROtmG0PnmaLzy3ZSvr58
DgeP3/y1D4EDe7Hlcc27pb3Jh2ddTsCsOLjygNgYcHOgZ0eS7RwjasI6SxAtdr5e8ovh8743ZIxo
1ZSgCacepZSHGxmrGhvxg0CrrbMoXZmVgkLx1s0cb40xOWV7gSgIdUl5FD35L5V8tKchFiTCWuIP
NO237toYrIJWnPoN0HGnp9Vl3QpFURxzRM+hjxGyIGoqynh2sr49pniqwePOGaMUKQwWHpotcovS
dO39AqwkvBq9QU4fLWT0AAaafhc1c4MJ29J5SUvzwjSXb98phN7q+kfI6FqnSneSH8JhpYDucwFQ
xruiCfxyyFDtaMfkPyLbW4pddt5/XSeYPS/IBOkiXC47wQPjxev4Kgtn5UJx84/fxVw/y2Be5t5T
OrbR60iQjkc+b+FjTIJiWKmfJrqm25sitizeg3OGOYan+PQP9FAG3gJE5RcFL8r9cyRvpsQHe+AW
coLKchHCwMusKYP/T+24Qc+bxX7E398ONIvlPkDCVOc7MuTXSNBbNFKCyHoB4kWnG8VxseLx5XBT
DE+THXpKK92As3GKxm2IE2CcmhLQNnlr3oD2aFPSVNbwqfEcoueeN8wrTm2KiBiKWdDiB2BT2a3q
dXdMsmqOghTYsFxxtYUCs5KYZeRoPVrpN+6M0/3a11/2zdyosCJt02cxI1J1LdqYRsIGvwwTf1Jf
sj1Aao5miugPRkwNAUdLE8gvyxqXsAp24Sc30fTyuJqBOz90QftRlNjW+qigZFrlLptitpb1+aQ1
zx8fg9bQyHGEuKFlr874xPdhDgpGczOc0buVP/IRKrhoV/k1yQYwtX/jf1BnIsB5PqTwf2k/MYyM
d3KmOb3AnhCkUMLnhIk0fRah265t4Rb+dKNYj+fe1tzTiAwMwqmtJV1OtjlP5dkU1nRdi8TaZ+9c
xFCfLFNv0ISCVVQjIxcp1/eJyWhZ7uPOt3sH9MC6eGi3pZZbaUSvNtXbaCF2jrWoSwHhuWuYs+N+
ug1JzDORRke8EPin0XsPN6s5fKKa1YbkOeo6LT9+NWJiOQ4N7/OVKh4PZWJ1mM7J72o/OQsihxE5
11cmnpK/wr8xobSpJ7E21jcxP122pBkgOT0A0w5pYuYeTl3XvVNnu+gM5Dcl2NlnMAvLASkZhAsW
vU8XOtVnvn/ass2F2mSGP/v1FJbGeEcT8Rb9H4tYgR9XtyvXYDtKtCRJqNglMsrBYLLrOZ5f6wq2
Xn03nrss5cKDr7FDUnv+esAMllgaKjMHdjYNp1qjMRwfmm9yvgByrDdsKEkA9O39bTXTzCizcibo
KFy5FKcmUeLWVsgdqCnakr/flX7MQbSGeTI2hN9NwJV1Q353HdPjalgYVsJayc/fKI10R6fK2jcu
KUZqbFz945dDVIBmLorGMXBSlYWa1+wjGF2RZN8H7Sbu8I862Mkt77D1yAne2UaxdHChCYg1s8rB
0Tkj4k18agkizWtl1guOJALlRbhvjOpon2UVxc1I+bN4stj2YsQmQV0g4Q44SWtzZHSEVGc3jGGV
jkfFYIeaJJgHYyNOoW8WOh1rNLtTB+fdcEiV6uADwCm/0fY6QlPnlQaaXyqEzttKfnRl8bpfi893
sl7t4+DsR03MEeFwqAlZQKupWbniA0b0xKQ6uhUym/YJpobNl0V9nGc7GSHzcScBi5zeHqHtBGTU
pmZ8YJHdFV6yZ9Si6AJObKCcNo/p448dSpKXnSHKPWI+jhd49vrEPfoQmWqAP1xDzpwHXWTfmshs
N5qR5pOmHvsh9PAD/QhB2WCjPeKBarjE9NwH/hqQkpcFJFAs9f7+S5c4vysJ1wWONRt+jnEOeEYD
s7EqszWdjY80R863dZ7CBt2BC52jTbf61Z2GoI2RSHbfBRtcIyeGrRJ/Q/+UydvQSkE5WXOfiEMh
AmKMNpf8db9OJr0AjASK/q7l6aPG9NaDBydL4abrviBJ42BBc45ocbDeWo4k5CHQYkHxXcagJvcj
4X89gT1+0C10/d9c5KYWqJesepGX/2yQtg4ERt2V/sUlTO31dTJWwFBPKmaKhujkHb0K5XuI+tGA
KWLqejxHY3tiBbBdI+vZOvV/WKrZUtuOhwcYXCgljUwOWR8N17D9AUzrTxqEKiAuMPYorUd0abLG
+gT85BV8kPmZaG+M/R7pUUvi3SBjoNNFZelLoxlw6coUWYvum9X+zCDEBu3ievZhM5Dfu0ZHpHFI
KE9lCjzzSCI158AHlRuu8QEGn2gEiaJ3d+OnHudWcHYoaE+stlpUWqxQZZMYjZW3/bcAC6ke1RXj
1FH8jwvfjCTRvUD9QezuVk3WXYM1c87Gsw973qSxBRLEyzaLC2+PlE1uWtxO/zTyvhuuWgBPkNjI
94gJTHXQYUpLSAPHqHGHZQRmR/rvrQwHv70POlwTAcc8qD2nRFybqLkifBRmUVYU2XPS2wkIPFqE
w+fcnrtHbwQg9xPYP7krCEK7XiWzY6TOsYB+j8k2Mmb8MSxVYfvLuYtrPNrovnAgmv0jZJD1g9W7
nDpoK5EVPhTAiWAFBvkUJYgKAeZqi7ZXFB351bA76bcB0BCo2krlkzqRWMYnC9YcztmHKNn76iXY
G+93q6LvhDcJ+siiDqHmMsBuYGeitP5TeGgCOkKVcEW7VuAN0phZfmJJR0h1w0L/u8lzZc7qHVVi
2Rc/0CLbsuNBuM0ZQ9iFxJvARh18KvWFw6rhkjg7mxjy7IkB5kBLJnhHCMhgDw56iYPUDvHtz6Ft
oPScTvc+7Tpu9xCSyqsOfcfLRa+rxeUjbsdJWRwlzv4gAUHBBKe3+ixLpCnY8m4X7JpXN7e/KcP8
W/EBvgMOBVVSRoIZOju08XwAoTFl+sbuIZU6lT+B08SXMYmnYdi/j8xQz5wxTTSOUWjg2qyIXbg7
eA7SBTxtd1XL9oUEyJf+bINNhAy9NfvlUTJDn1QB01/vYt+MBMZ+eiJrkv9yYIQ4wwhNIzN70pYl
5TzmfXDmaTlTislEmEgs7RT7INvW9GrZhr2wy2Ectx0QCRY5CondSo4YIDAcQngNTWuoGw2NVBMo
YpwQUjhdnvOkMKbYqVHtvHo2kihBL7alGcGqs5fFnuKrbLfdSMX031yhbn5JLd3oOyVIuemM11Lq
OA2/tWKKUqwxVeuwbUfje3zyBcBF4pfPs0597G7x+yUVsenQO3gEpue/bCJbvx4LRsU8j+o/inhl
NCFb8KhLakL/h8BBdetx8rTfqGuk8MtTC0GLkst1xaP3cvNua/9aYV5uGAe9Il3FnwvvDRwelFtI
1sVQ1CRqVStcIunAKXnkxiHPfKf8EBzp/T5D4ZuMA3eP4yplc/xKgl69P3O3NYWgig2GQfHEuNUu
NmEfYULMgCmdlxpkR/zsYTUKI+Zsl8KrUs4uH/EcvXHOlOQmWu7YCm+TWKthqw9PnLlAqjpmOhdq
YrZJCAWZ+TH0feblyQFzqigS8QiRBDv3P/DtawrDXjrb7rLohYmRyOk48ycAzexbcmBgR2a20hLC
ggL+8qbZhupehgSIrX4ZzzjCY4UW60uZt5syZ6F+0oqu4UumnL8JkGB2MMT/+84Ms9pqvw19fBKs
aPcR2ZZ2SuLKIu9n/UKmgKOcpsvibdaVYiVLxN2od7SaHAg7dTXusg74iP2+YFOQE6E7IRnu4jcA
Q4Etb6vm/w5wNBRk3i5IyLy1lCjGDC6Cp969f4i6ndbVqQxef5C0OA4xhN1aigA7MrUD96w75WxD
oHE5YUVPcnUl3KLv+AtmQOhYZmoz6lzu0c4NyxbCQZeA8AZJMliBWVlMM77EWkzqXiyk53DXry3+
UyHUjsHXh9STdJO0tG2gXnAFZDHXR+LIqQM0s7hP5MuyvkZ/ro0dKGnVtg4oBflMZlddQPOlBLr0
0MLJwbHTi1+YIHTUeevwoPNWlvIj6WAsrU03QCPhfQqq2ZdqmGG6bLNfJp3AFZP6UItUk2fejqqW
nvQBEUbw72pdz7/Odp+CniR2gSu7X+EvrfWVB05NGdkcHdVaP4Tou4YLkH1dFoDVu5OmayxJjzY2
lSpcYa9TK6eLX8fZfIE8UiApRwfWfMIuH2oCzi4u+xUWgyAccEo12vE4riWxJTpuFTv8tmT18uIc
XY/NR8ICkkng7X8ZKAR41rAaF92YJY09PvX0fjPZ48g/o6lVYA7P05XXhe/zUpPc99xO+SRiJQEx
wRmKMduL3fUYCI8zuuLwSkiSVFoTTYME6bqT/oJSgkcF7ZIexzlwo9WgyMX6K46otsmQmlMWQ+wc
1T1dA5RJPRFjyQDz9AoPAcj/ff78bt/upgr67eWTqUnz3OTHPIu6BkiwCVfuCkyG810cxaz6ta4W
/u/ZF+C4OyQL062l6nBl0XaUZ7U2nu6yd2sy7Kg3cpbD9a6Cxw+ESkhCkFIzX1nWebUiB5gMdLXd
KspLnC8PbK6sJC1prbdnoyANTQLXAFROPQ0V6y11ozmGqvffbT1ttNwyhyH2cZFN5m5JlU21hBA/
ymZele/S4wqSQRe52vgkH+v0JIOi4YzoCwdbLW7KDYKsA5nk0DMwIB9N23tPraLVcva4ZscvKP5u
/p5OEUcCvCsvR+ZXSO9Le0zumevoUrkGYvSzsBg7YNUE2jmJ0vGPDYVBSoGk39iiKg3yT9G+ghv4
2ypFUBL9+61iJQqyFHJ4TcGYA3Epe7/Jvfk9e1fxuwdcFMJ4tPFp66apgNhA7YDKiXjCB3ctL547
jMoomfFHi+AdAX95FWuKvpN3Rp8nWpVW1AcZN/JdvKz1z7use4XxPkZ3KFUG6wvdYuU0ol4VqOzT
PvjYfA6jYOBpa4xaw+RC2VBv2gj+MgqgmfAcDIoUYGNYa+zOTZ2w8oLo4Anx6rOms90RuqDGS2AI
Z2zIdjMdd9vL1rCzRQ3M/sbSdEbanfzZrS2NdR0+aWtqZjHIwTw9oeKaKzvhwJCIx1gapg6U5mV2
q1srvfN/nJS3E2CrireIRbq6C8jJdNEuTggRebQvGDjQRQQk/ncBGvnvxHkCaMShod+kgZPwVG4q
eOBUdl9OBS656J6lP79TTCrbI7nrqLXXhA+fqJckPMl/U6jibtJC0xbJxQ67gs4e4UJfOxWnAzfq
fvhVnDMBERlv9W9bepC8zDRcoOuHp9POJT2ZatsBwAZYsWHLZg1U3iXKbyDMs+aMmZ3yngbMAmDS
ns16JtlERJWD7lVy9U8PnlKBMTgNMNg4inUQ/akPMlEtV4CfntdpA9JDwtSvJTnZc8cHMAtVA3Lf
9Z+0TuEvf4XMdnNEou3Z8o3sZIm25N6h4ZFQi/QeL6rOsQkda2nzM/ECC33PE9IvMZsuWq71+UVk
alqAIQ5gKTAI3957vXJ1aooeLNtumZ7VDqSNLWG27CynXUA7xls2tQnCAlnFxg8nljrlyLHloA3e
8QX4eIdwDBPgYy53c+Cc66d7ZYW35jt4qyep5Ea0FAbPt5Ttoe2G3BqwAzLBz7IN5Js0I0+Z8xDy
aaoo8aiRNfJoBFYJS8tyOoOKZiyKOon4h99Ln/IvyBtN/px95B7y2gzlusDEcp2KFCh3+7szXLPA
aH4175dKpolXa28nkvkehtfu+boEA2PbBqPcf7UB+UfTRbWDCV9IhLwM9FfrotN4OG9Ut9FVDyEk
4JvuJ6tvS28i8RshHtKpF4ztP6sBEd74+YQfReE0GIJ/I/4RJK1T9yuMlhko1Z1KxCrkaD/6pgpD
ST+mdqfwbDCWMyBcqT7xTrdG3uvYYUfk2olpokSJPM/ffWoBPS/wJ1IFwwTjp/b1YCURUx5Qe6w3
UnXUFxa5lVYMhmTnDzHSodzZzgp6bV4hyLK3SC8JI7DWWroh4D20JW3HbDOINxen/iXqr1dIFcey
ppU0PZ6ry47++4arfYs/Huweiuy1jt/BkxFH9geRlLQcVl6CNu7Sqga1EmPmz7At2Aff2jQQ19O8
es5+Ui0BtDldMuuVJiFdls2ffyHy2HbfOwylXaoJdu/IzGEddqw1a3FZ4CZYLeZKN1PEj99wXW6z
QaVK9hIeynD6IT7yyv9GH9X7QzT2TsDj9FpLQLwjNZcpUH9R0eVtU/xA6wS2mFKWBCp/el0buXxj
e35WpxEVK4L8VSBmetN4nC3qIE9jiHD2tD5D+OCeKM9A9ih2DsYCDjnJqHC8t4Ek3tc0a8v21VuH
TFUAD5j6xkIDOPjOX2kSF9e9py874EuffBVdHZeoHbesnW283bwqDIbgPhZ9UpgZgL8mtyCjgYZM
PzAQ8gPpJ21/sXt/3t1z//yxX62ft0p9FdqpEX0QoiMZ/YwwbmwJ7iUsYTpESTsbL3fykWLYgcWo
XD/Tx3oBwadQxXOccCh5NyT/mW0RfricJKuRetODwkhoypiAXmC+x90EWf1BFV4R/qOnSsOi8O0T
Nngnpq2M/tPFZ2EjITcuBGIUfxY2POgYamP2pLn/oEePg5j1Ec0u6X/h4vSY9f4lrH+0Umc1nmp1
n4+EjtiJw0iVUSFqcE7PCWcS94CO3v5E2d5+Ub6mlqhCY9QnUydy3oC4JQjePRwhXDtGkOzkxXaU
NkVAhAFBM6OAuFlUJ5xPE3dYx8Y9FWcgPSMyR9BCKSr6WjmNp0eFdO5tYofE4EoZwImta4yRoCg3
k6qEYXQfMbYYblDB+1Dv6JcSoe1RlSxf07BSyUdzi0EhB9orJnwGO7etWVd8R7B6VYS1KWo9PlaZ
krBuCx8y49fF4MVf+MT/SsdxzwRMidUlD9/iZaab1jMajf0pTXSJWt68TKJrK5d0+t7BNXuDP4FF
W43IZDVxDJsRHAsV5v7w74DU2jv5mDBc5HvFY6UPccOxpx215x+LceXaabLCeCfE5zEuZf+lcaZG
6PeWhHxs4Sx1lXVL0JKoVR95fRFnvV9jCn4fGtj5slt3yLZ4MbFGsFBvH1/qgCsFtdcI9y39eTMt
2Cgs61/ELpagKiKHV6DbCXfxbn6cMauPvEWV0USl+h56dbUe61URVuhjjKrBdVEaGoMm9QGdbSEI
jsAIQjjQCSOUAfaOipiHlniVu5RyhOIABnBT2eYQtFDE494k7xpBY73JGj2SGl/646MSG50XbLE2
PIyMaFKIiub+aRlvSH3MulECMaPRXwlruQEjJ+FhzYmJPZZeBLLG8h0VUNObvpEDp+Y+VcRzEeGs
9m3+/leqw+woVrFjR0ilPWP7CEDbpuyhbniRSLKJ/7ylZ5MT83b2aH0pWQcctF0XNksO51rtekIZ
FjzvV/m6Tloz/vzl+G0/jzSV25hg9V81Qec4sk7eRjEoRqdorPWexPFfarZY2wKD5tvl3sjPI3fG
cyqc3c3yJ6KSU4f5vSsf1N8GzLe/PyZ3ftnwmr/oz60cB8uDXUXl0jd2AhxV4l2lEHdWDmwNdKfY
jRKpKXvqjNAZOx7s/QFr8O08BSDIMbXablqz/MMvhLyNCf8NzEq6Bk5FpXa4Le130Ro6h5vwX+7o
YBqtiz2OojeM2fIhIwO87H2ZFBCwjoiC5we44sS8Pwd4WDFdSEMTtvGiFavjdeiB9mc2+hqBg87X
AWp5zREhos5hkpn7pGMwoa151+qspUqaxIktt1IviVmUPCMBPqzotrS5CbS4sVhK48aTF25gZ/Qx
Hw8PB5ndZly3ThMciu709+h1ZztwPspYSeNxPDL3OIPz5fIj/XB1D8F0Yo7Gk08wo7l0uQnFenFW
3sBuXu7CVR7CCC0Zm/I4oDBrCmtJ0QUGWzNvusZ8kXv8LHeKyWyzn6gtP/YWkT5+IVbdP6U9afim
l0tG3HOfjZHfOu8lqGfr/hK11dB7ClBipO3Ct3RhXoX+H/FjGqB+6ZhmrsJ36i4cRJYvB/JXdb4t
eSB67+i7qBCWHZgeUr76Jx1JBdUO+XaIhndZ63HDO0mS8czjaP4kzj+4/chpKS7A5eEHndsvrRq3
qX/wz+x8D3E2gVazaeoMo7kpn8UR3Hz9c3OWQPYM/pVqDf/KaKl8eQsBIdq4bg9bvf8k53m3Mfs0
Ev7lsverbI6RCYjZUbHiFXXFrtuTKIfY/yR3QtIXSc6nqnotwg/LE6cuZTOebzPNRjDeODpaiyYZ
Qdd6U65HLAEttf6bjseryyB+IzS6/Z0QTJclA3sGym/FAiCHWAs6XdlrkWg0PdGJ4GXm0hZda+kL
Y0txrQDdoX3t9Rm681rnjAm30PW+401iSyay4ApytgFD5AIsp4R0NMgryvCYv6hluMx1X0GxifNw
zk/6BewQ/yN+NXvQANkMeqT4qbnPqfmlNHnT/nyXAxcru98kiMsoiMzA6LNhzECNWWH3M/KlTGgW
O+wLSk9aKYEAPRoAde+hg0q7tMAECaYPe7Iv8L7HKAGtkv8u9hNygXLnXkXeCfOLqsPU9VNn0a/W
HMyDLFYAvk/e8pqx08MTPchFOAUpdeRVAQFmAoSLQHZNeNhthNvWHdA5b8lExyRTQ2aXwqW/txTW
ZUsZhOCGtLsfoYGNL7+JVLzFopar2G5PjDKWYw9dG9a4sr9O2RATQXZ0ddTE1cM4v/cVJFfwGqPH
r1U6+l10fjbCzY07FBF+qAYXPZXPFtpUrYvEyPBi25xGuoOyb+Xqrd+x4HcEk2UuUpldgA1owc97
73IdGb/7R1kq+Z28HSTpUJOvWJXn6zmeMF+q9KeLnJbpMeTeKv1NksN38iDfBC5R1MQc58gxsofc
Q031jSO/3rypzjzNt4jae9EvraVOmFYf8QWTM6gYslmk//iYPZ8r4EVBJxVpgaJGUFN2nYhqRk4S
Sbphmrb8fKskTVaWZIGfs7DE51j3gJQtUQCKz1SC6gvDNP5V3u/p/td1d1uv2rUIiqJk9KlcsFIY
B+IAwKxXsUMEFofAeZXgM+Ouni/oWPDdqYZRz3Ghx1eaYP22cXHVe1XGNNHn9yHKHygR0E4a2Igs
OzwY5wfbEUxdaPN62aT5Mo4e98+TEPT9J6espsLvMufB02W1zCjV8j4Hds42IC5BGienCBmI1FSW
di+kl/V0SbU0fJjADIfclWUtvpRpr6t7bW77PApzmXSowIW3X3LJ7kJ2iUUNLUbanHpCJ1j//qPI
39jGbJsadw2ng9CxgNlX1IOg9HFotvbtdbo5tC4AAcRTf/UGRAwmfw7CIoNNCo1P9ESAY1siUuZF
ZtQrr2KY4YygUgEihI1566/Ej4ectBPnyQ+kLyGaeHMn6YX4y8q4FgJ0cQeybQuyZ00IL2+302Kc
7sUs/NpPCBiLYlt1sZ8VHyq1BXdwnSb56zDzJ+k2Nft9YKwsbPf9S4C5j3LSM02CL5X+lyOFlYy/
aD9HcYmTdz8geP1dIFItUParlbQlG2cs5zUK5a1Rt0A9rzryfIfA0IcdYrEO43OMWKXXEyAy8ILp
Gx6kKXhFQIMdNb9XpsDlDflqWVjFp6uIUMHrAeRQARxNo3WG39CmndBUB4LYZB8i3nJcZzvfZYKV
QcmMV4cMkn8sH+E2oAsDRj0NZjwTWSqaCIsFUlQnJ3cWCXl1ZCbd3ECR+3DdQpO3O+2cEr/LB7gC
OrZb2wJFKg9NaevBoCE9SUFwDJ14WIjr8n71rSC6eZSeOiZQVprLjDYn94ge+K626Vui1CwMnDD7
oy5neSo3i7PaPn31hPjmSYhTGZEFC1sZ9fJP+kPJll26JV1bdnLeq3hDkJqtAAMWky49Qldyca+K
eDacyYhoZKKTMUOu6Yx+dU/6jt/p4tmdU4PioetVn8+/x+6H9vkPRCCXusvQgEPD4AqkeuoCOXhe
H3zDJ08+bVcZ8cqdTqZneFxSPAzMPfWFk/S+Cl1IRQmEjLWV43ZHxs+dwfdaVe9tarp7Bvf8B2Kn
puGWj61DX9tHzfRHZYI2WeQedcIELNIgFVhDgruh2PnmuIB+M0QSpNkaFSDTRqSUFGnKx6QyjD9/
VaBbDEkwtBB0DxFg+uD8F/ipVUvruOSBBP0dxgMUYUhf5We9uvD8+hPghoJQjATRmbcyxU3vtL7O
Jaq5LPHRVs4HMSwzMFuBSZjKY4buq9vaffZ05CxVsT5ZaXfpNNWUxSK4lqlrZEwVYLvGuBq5NGA7
FcAi3KyrGRpMB67AySn6rCNN58JxOGFF42WzgWM6TaNdyDUjqXBw6eE+wFfsLIJaoTXGKxnmPsi2
eEfHwQBOcYi+sqEUe4Z6tLw0cVjZX4q2baJJuR6NJWloT9N/otFjGrqST67pKohyBBnsZ3urxO3h
HohFe0/QrysrxM2rtucB+1E7vPoTdymU5dE5FmbmJnDy+Tc4rye0k/6+vVANM3HFYA3XB714NJ8x
67CxgmLzla6HiGuHWdWpoyPKBs93ysa9BAYIDJww9EmRrlZAj+PXigszZ0Qok4on+ggBSy3ga4uT
VQUWu43wrifBMFRTJD0Nu3lgq9+p+PjDs+Y4JMQ1f0m3kj5v9F9LqVSL50E/5qu0EaYTqKzAYNbR
xazf3Ds+vNG4dA+YvTtFNOLO5YYEBwYoY54g/Em0f0K0G+PVzWHfD8jZVC45XekzlLZMF/4m4HMq
anDTSoermzWStXudTE4UM3yhsT0bdShv37DK2ikyak8gW/kfBcvh/ifevPV1LmQ1NlKwA6Dcy/gm
CtTevUvTVWJClvXMS6ELQzYkwks4rmWYNS49LS5HQm/84797YMavd7CGqeZvbPkomoIe/g/qugFI
g699r9JiQNRzKqQGPlQzHIACDdkwMSd/h+MXG/NRcZ+zALUbUQHOSRULgC3rsPbAGUf+t3HI8bB2
HHbwsltlk2ZapJ4ze0Pm+/fxX80Nct/wzbDfBwcYMtjTv5OfnAV6RpN9jOYXXmhg87aYr8JWdlXL
Ts/o2NroWO/XDwYVQECAAdGivDb5YsOg3/CrIyQ84Tz8CdW+bxcAQhVZGmcAdWiKuLBvof6OM/ep
o2L2fqi2YRqx2OlroknrUaZRhr8v+qlzF1/kUBX3f4OXjZlsJm3NrvKJxEoHmYMZ0E5FcbMZjh7a
VWzrDzk76UbM5Cm72dInAI4jFeQmdfUd+D2HkWs/We7fmhctVoofaTusUxMqPx+AKxbpEUWxVokL
9CdKk32BvNw8v2eEZVXQ0yuZY0uSCrolBuR0tRgkIzGRJ2KNKy/q651H+LNnnX4l/3eb4cQEhsa8
tPw3UbuAPsaREPva5s7tgb7AiCPnyjPwgCpDvYmjZDLnGlbdH4uulXLKkN+K+ho+MbNZ67TksxtX
iUAa6G+4lbzMB1ij+aA97KmB/fpEEffsgU60G5vZJmQ1Bl1kqeA1JoT2HFu9cw7ftVDT2yzpEbnl
Tie31Pdf8KPSt27RgyQqgEhU86cs1349Xv4P4FS32+vYWoQIlCmyYb2LiByCsgTqfjPsk3qO8MQa
6HTAC8z8jMXLRMi1QLEPVuz0XEsy+RQmIooKFYARAFIKeQaKdHNvqHiy7CT+h6nTj7kwn41O4nHe
ga1vbKywmeKO65e0HPrNUSdNoe2sIv4x1/zyjUUO6yVIrPVduWLsnlIBLHfuELfkRZsiBSnd3AIj
EcrvjYEJDXs4dwJ6QNwSVOsYVLAgEKkrSxZIyWGroPNpc5VTCPubZmF7jrNrS8+/uQsWdVyPRgL6
0EhOf9XdLKlEMC6LkJY0c4LRtGpC7XsjG3neRRWOqigdOiEyqWjdOjJWj/4Nko6IrvlsMlE+IzEU
breKO9oi2eUjJf0mUhXDoF8DZzZWfOSWUU1pGhzd/b/QSbBc6ehrvKNVpgu6ly6qOz2f70fvyP69
J7mAjhgmmuvAWYhwjJny/+8UKaT4xGGPpDnSoFCvkGMM8O2OgU1FQPrD/0pnzUH3/MRGhuazw2Zk
wXAoXIl3f8F/oM02VsQtuVqtJjKhW+joVnyUFwe4y3A16nhZOpdUn1OslIEtgu4ywuYseownMoiR
kadnLNIuGk0Mm6u3TYwBdJ769xZEmTwtjpw+9gqYVI+ViSNlhfnGoMBc9FapzKcFz2eGen4D9eF2
FtXKq5iAJM09V6TH6DWuJT+fhlft2lvYG8zWybDQf+NV/NW+G+vdK0ofSQItaYCaEx0mbKpITuwX
KIDL3jRL00B8OnFiRz5J7LgUV3wQvXmM26F/Ap4ggWXe0l4bCYll2ZyHtZBh8q5srUwuEWSd97nS
SLTx61/o4Kesxn8fsdkais4BUzSWpMUFCgPHWIGzqHICa+Do50bFS2O0oU3pQHDO8MQnaVc3r0CK
0r9AYQ9qQjpZSRKhZeRWXPYm9/Gd/ljnecPS8wVr184ss+ozaX9C03XaGX6rTu5IGyzjzfpaqzR4
tfyeOfMw98kOtXwUlQcJOdkzwO45t744bynys6QqXowMWN/6L+hSMyAdiHO0CQvWb0n9P1vEaMTs
iBsv5MtKrAsRAa2utdw2rZp8qw+ryxDuLa/7GltjkgBX1UVkk2Diih/Ebnh/uuuY3zx03ymaCWEH
VPAgGbiLb2/rm/9obIz2DRY8J/a0TB3Y9WvOBqGAQYMJxwEBfZKlvRVoXLfcxt3yxyjDbVZJBR2G
DswqiN9zCs/DWbz7FQR+h51A2rh6xuftfekOXvOBVcfLOs4dxkBR2BLNx+KtxKEqB37ueJhR2kJr
eRZ6er24xYcePjwrjhg4Q4sBGWfuUEHCUD9cuNFK3wEdQge0NrxzARwMS6DsUO1PxE9JeJwnjnR9
97e0Pv5U5UXYzoX+mVfgrRphLJSCsXK9h86U1SUq8CI9ChevxJFVkoSsYiklRv7NRwbe81YLcSZu
nf2ZStSHiDNRzXw3j7a+8MxdosMvUoTRtDudwMM0TPMeENBWJZvJJmWX1UceAyuFN+RrU2ll9+jV
SM3N4Z1gqStJ0nPPCODedzwpVqVjqf6abU16ezJyGqpVleaLhIpxcqhhN79W6Bb1Ngz9gUOAc2cR
yiuB0BpDzTtXP5UkMnroGdEDBcFh1J99lct/tjf7tgb3U2XIF1fetFlwG3zv5DfXL4sCxDmRGRMJ
uUZQ0qPOfK43jd3X9bey7soMRmlUet4WsqJYBvHB09du36iWe5vZZac2ZulPi6DerPpK7HMYlP0n
Yjz9kNB21Ss+WSMze3liVUuEwVU+4ozT9ys2Xe4t9BmB3XLwqNqEQ4z/lD+IMLn8cgHdUibl9o7K
dqxJPFqjcIUBjy6GE6LSGSxXqD9zZq45nrHj+4/r63nj312BplC3nz7eHW6PoJ3N9iB+9rE62jPL
DSLd1yeelqjhkMLRvT3dMkiI7Z1Yld5MtLwPmKjRIyFapNZUAs/sMj/aWdTRJ2YOziNcD5HsydEI
uypJNy193iZl4y148qOkkm3mLb2MP1f1uKBjd4pGIXSNBTMjstl3VJcqXiGAHs7IEqt+RNxq+EcY
h5NyzPnqtW3I6TWuOi4ymOKoylpwp87R5rR2kV/RIzxiI1+r6EnsXLQAAJlMfH90gpwkozgl0Zco
wWGvBfugkKcCkxrTjq9oGJoLf9Tp4dV1ML047+ChJa1Q4oOOTAoPDpsEnVBlakOKASWPdwaaNC1S
zZh5WG2fYnZiq90BE4XxYGu7HmnFLnTsSlQxNL+DPTJsMHe942Ae+7C1ggq3p0hTGMBuPgj8e0iW
l7BnL6xAnA9T5yK/mw9Bwq4POq5yaZ+m9/kPSzHQzGPHZYb4bJv9xl5OQmRF2P3I+/jAIbOwzpN+
ZhyLpgA/Bp+gvx/dIrum0R08v/8voB53Wp/4Ospa7c8dERVGMJs37mDThJgakW9cBc9irGFVi3MD
H0jKNpiGvX0vItJKdcgtewWDXMlNCThtPbr5yZuLMVsZ3lgHCLMa34DC2endim6lh10ag+emsBFI
wWfmOTUB8bcv5kJlPE04AU9fowTDxAWHt2d6x+bLUg9YXE/j9E1MCjZ1vdtEnwx/KkEohsTVPiDQ
MZv2Ns6bqUXqXMBEEneo4nTnFTw28IV3vzoq9ggTPkWrTM0hd4ARKXptRMZ/luIPr+G7Igy26m1o
wTzz8cLg3Nqe2IHiWydOkDxd1K+7acSqndVi1JsSZSEFm3C2Gn1BaNSmTl4ioHfsmEL5PhzgwNHH
tPCSAKK66Hu6HzeG3JRntSxXNZA3KWmgP9GNOmPPcxkh1Z89I7uX0pJpuaMB9i5r/zBkWziAliED
tpmd/dlIZaYp5B4+MgeCxEw7plTqsORkWl6C1C3V1ygayI7IFMkhe3MUmmpdiDtkmUSNN3kBroBJ
CJQFybE2p1CLh2VoV3mUwS32jSzCu8dPr2bdvqEo5F4b3/uzZOKCDfqd/qEchNt/+JEsSSRo4uhG
q3atgr/asxPMnALpxF04qs8Fp54F7wsXFIe55YeW1Y2p2vtidVof+P/p8T8UpejvQnoVz9iLRmSs
BMpgQErrZbfIApgx3k6jC2i6HABtFP4sc9IHzbDkYm/eR673Yl6aMsO7dvP1UNBQAe1yHrLvUSX0
40ANCjYzaWZ4vec0OaY+RuWaj7OPNN2+UMq+2pJWZ9xjy2TR4Me2vpzOchu6flMv9rbNgcbHi7h2
H75od5SduZoUprObXJ2ct/AGZgy15Yzd7mmMbmb7PL/k01yv0joMaOJpL884seqCKgCR5nEKw6RE
np7/rLWEuObjaxPBDZ79iLHz4K6da+LluYsL86ndlCYQLU79RdY090Ws8HmTYHKpOebdzPFCcxs4
zEi1zBfr0PibMmFUx5Nkjn412e2Ft+vLrM8zinDrQtzJ6nsJZajX5W4G+1udnsseddemJizXMKFv
PG2ZUbV8qnIJkmIlq0fPCQqIuG97YLLkVbVTvs4r54jsjRBl+Ju5CeQCV5/4n3rPHHYVzzkq6HKm
kMSPQeP8Y4kPOoCvcg3wG82VpvJ+tr+mR4RKGyRkZUuiWyCrpNNubMoPJ5p//NCDD+zaTm2ihNnd
eI5ZQg/s9H9zz5GJjeKVtEojKcJEV2Y2P4x895rgAfttiMnZLPFeLIXt9wdmy1ywJrJ9gs9udEZ+
2dEwyKhld5Io1wXE4BKMO8ISPA4vSbBwu3nc6tNz/dQS/HEhpKmPIHyR0W6k2AIKY+Rucl9RE9V/
ntioqmL+F0vovOmLA49pqGy91/POIwvhlQd7YeBr+DGSdVejLpknH42tvICrBW0USrTZnWBs1/v8
5JQ0lKjTySX1f1LRzGrjzgQxSmT9qjqWPXAkBjzKfg7kKMpRzgYucjj8ZI9NLSjnhC2CKLc/FhJi
Ssv6uczkZEf/b8JWaULaralZxx7mH7PbS0TeuZtr17IYjLRiiumeJNvGVT5KQU1AALJ7pLfMbCez
kly2KWoguYtJz+YvX9uqj5CMB4RPXrZB1QG9d9SaodFEMGJ8eC0/xyCmX35vwEOLaGT1vHgrveaV
k8PBJnd1874xxBWUqqNlOTsFkAHDAxTmVAGZydqMpOWQqU7Z3ixik1kR3jtXAYIGl3xUCNwJCjY0
ulH+mBlpBDcRqnr2Y+auWWqvdDI9oQaCiCA7B3LY3ycmYIIlpyMUF1vaFD5SNdMI8KFXckCNmnku
jpUM2FSnU2gV5ru9zwHtwhMMmeE4DFSEbY+YJ/Kf8RfNkDjJND0/YaCFE9qld70L/PrRwBZLSrP5
XgAKV6f3TIKf7gddgk/ycWDzet2jyTtDIgTRJRHyXZHEqjYQL0hRSRCt5CoOO0GDNWUrxNbtM3WH
uKxeSxg6/K0Vov0l0Ee1yRqNd2fkhT3yXB56SsxczhKSGfsdVLGuXknwobYbcegnOB+iS8M0sJnE
ROAvYyWUhyIyd9tm1HJNxQxBnnV4M2vOWobEfrRa+Mta4xFENiM2v1MXoGFLWND/KlDQOG+fM7/A
Nb+1a3/VAf4muRw0XSrz3GiH0A6gX45qtk8wkjC7riY24TKkaan2coJAkLTtoegVdz0wHS1J+iYM
arWlK6qOnAJoWMHGyuKTtgZ15G6CMqaZSzB1oMOGeTp3An4/XRQsOGuREpXAm5htriEfTofGVgVN
VI4A72FwUUKQCGuA2TAR7H9QGHgMkTX4KMyZF7bVHOdo/7fkmGn7C31AV59P2cBgn7ljGRzek2H+
r5/HEgw735V1FgWvpG+ip8exK+F5RzlytuR6kf7XEKDu5FnmSjhtAI7wYuiPux54OlNsYoM9qnve
VBKobp9WhJ5XgyH2UOa6DQDqmQLe9mAnxs4WgeUM4ibEDCO2g5LEFgu3JBojvi6+1+pNXwOxTnN3
XzBX73d7c4pN2bVdkDHdmfElQZPW0WuO0fKynV25dA4MXLXmgccgHIQd5rr1eUxAjgfyYAy3Aqx6
DKLb/ZmSpA7RRa9ralaeOXu6ndLVzqNwCIzA8hu2FjJS3/GJKMCevkpkfavdOP57J+DZ0YhySw+W
FC4mNsLlpqTCcGPDtj9w44w04QFmYL5MKeu3JdqW1L0E2AJ1QMutsjqDQErOipJMQxVap1g2rRdX
fJrrYyOZs8bZEKHVQun4aOB+4A7kLk0F4xfYZN/sQCnP6K8MduriC4TqHrGf72v3v6qAjGBIlcRy
4GUv8DlcepfSP4l77pfyAxJyWlk4r5cS4ABZz5jiZ85tUXRj8lIHbeqAUB+/RR+qH4Azb8CF0lPu
W+BuCf/RmzgpyJfaVTuZhRA2I25V8yurIFP5EBsF5HbXNX+yPOQ2D3NkDpw0oteIn9ROjBvUao4X
I0RWpMqnfPZuutMWeEsCVKhrTERAr4PH9ri8y0SKcmG1cvLmL9p3JZf6Q5XtMfMeVMSpNZuWLiz8
vVteXKfo/4NZYnO03OCjaM+4PghkCsiwKb3yyORzzCqMcoeaPy0CMZX8r3dQZcZSw4krejq1pJ/O
u3+lT/iaqcTZ1HVaMOr+q19lHgObOAhlknQDz8XILyayp347KX0vHX3TI9SP7yconvJ6NRuSDiVQ
mmE9yAGYmjCk4Um1oj2+wvvA+KietNJiMPQrr22zkz+bZ8geJZ8JDP/XPkxvdGp6rvPZ/WekNqUU
K2owbZueDgE8tJ9q9VmnVLfDO/U2R9D1e66bvtUmT5/1XLj6iGBcmRg/OkhS4R3bRXD73x7Y7aeB
/pwNKQqzJs30hkqofk5djbHGdIBa0vwyxwc2OX2HKB4HtAMkER1xEdmCQePssMIoFeSKE+uHLS6n
fWFb3leQdE8j2cfv48pP68lkf9TiboTsyEn6Uj4fZ90pI4PU0p99hBV4JR5qBJrWwW1cyimSwS0z
Sq9M3CxgUUNng4OIwe/xYHZNYajEqLtzDPeadeZulBve7BUndp0jZ2jHrKmzh9lzV5WwPOz20abK
DZv8aITBqd3ab36W/RL9/J8O7xCgYpkd2WX5p7PIN0cQ7kp1QvqDCCzY4N2kbY/UZQ/5XDV29KLz
gixRJDqefXgJyyJMt20JAPBpuHlWLyTpfHISD6MWhudZPPTHNvLIwejxVkuTiTs3uv7Zija45/3z
Eykj4fs7skfbZ248k0Alia1P7tXm0Y3YPHzJP+qhPTJyVsJ9H8E82xsPakwoh2lwVbg2cxjo21w9
TcdWaq1cv0Ttc0SnnH0yiEfKdFBPbcypWY1bPpZLMukYdHTTkp19teOUp5j17s143LmwuhFNGuxl
oXlc9doa88KRybg3FuFq1Sa8BbN8eDmaXhK4a/Y/Bh09Y+HM/iQh2nfNUPY/nGriFATFx2Mxyh5j
XOjFwwjFK4rcb5zhHoNVzpLPj/8iRsknpSbMYf7YJCXEuRjk0quj/exXIOH3XUgGaqpFnIxeZtPx
W4WNI51A7wQ76KWE0hktu1+ObJM2R+qmErjRv9eURDvICXYNJ1RAUk2qqQ1uEz70s9obcw/VGaA1
XtlFoo6MCbEkW4I/qMYMp/Xd3WRQe0YdYu0xcGReKd5UF0Ikq2npjZ5ABl7i3umnhLbprhThaAyi
K/qJTEMPcEoMT//QtaTdphEIYY3HTwjL18XZ1JRHsA2kjsbXbJ4oLV5u1cBIIYoQF+e7MJH+1MwF
gC9kGS43atItJzZxLEpZGrNI5cAz5LKgp9VjV53y63952oAo1danoCumi8kjc5Xdy3RDqq1x8roN
mXdDkjTFHJdFuQrNZ91UoZWVIddjk//TWP9QDuwKSoeeaCXaaPEgnMXoEkJQhMgshRmizDWyks/i
JP/fkZGEFYzh0kAoUqjUHw3GdYfeiqzwRxRA163BIUmhH0Tc3WDoJeYsTIjs5Vw/li+FbDc2Ivam
YSUTh20SsFOv84sbcdPmNRqGeRI6puJ2Lqa29uDsAveyeVKlzv6BhTW+wtr3IbtH0cDYjQw0PE69
59QmIbrIYjJWL8L44LwEAjRwA9yHOE4NU0H93xjrMtY7jtpkw6Vr3cKs24eUKP/qgSlZjIaXYfnJ
B3DUzSNo9Om8Ryn+NH8agz+d9Mb7rObnJlWtF0gxIGFD+PeU83hl0TKMWOBPhxsDdSoaWZgwS5/B
JmU5iOB/MmmhDVyOhyomkeLzmTxQaxjbownk3SV0lxMcirVqBHrt5QDzfNPZIixEuIVJ11I/CIKv
AMwoA5fbiYSyevg0jA4M/2iLT/0XN8Af/mRlFuVyHab+xXcYZykG+jaZk1k5/brnvRp0aTPv2gna
YGtfsMOpxIBPxhc/csQ/kftG6xMJYi4VmmH6JzX46W30anmtIIghLMXrL6yMtcl2Dg7thySH3ISZ
kZAz3tZ2sN+TJrmj09efDkHqEUPABxoIsRcx/Qwucq6HTOwbB5wBX47FgNoiYzC/dZcsUeFb7BMm
g34EXS4OkMlDMw4ddhIcVHQTh8Euq8SnpwoMinpPOF9PlU3ukuu1QCLRT/4kJTy/EdDWDaTVz66n
rjlax1ZgRa3q4uVfa9QCagaDhzEF/Duj9C8izYocpCUTaxvYNhDUJcRLmVvGNt59lBZgzRWXiHe6
E1YVi+Tp/xFytlWrKWxd1i4EhLqx72SbXk2LNRyxJzBipJVgR/z61BoWqDiKwH1nmhHZ2fswdSkX
dD/m+QyVJjH0+lDNHmF1NmIMb5SJkJInnyPIWfWbCtWDXYmpy0g6aCGM19wAqIBdsO4iCBbkqZnv
kJmh7etJNAZe2hVxSAkxlbdPvcqo98DNzx8lLvv6NDtJXmPNpdht6Gfwpo64ab2p1LniiymXPfct
VVoRR4iZosGZcfk0m/l8dlJG1MdLESf0tr98Fha5Jx1rmhg8uy0NFQLe4nNR95CkL4ymYr6rjv3f
ljxbZkH7rkW+noptaM5edIL61tIoiFFbuEKORxyrCnrjgnA3Kts5Wa/5SDYXypw65BjVvPB29H7B
HcYhvaTQi9p327M6JNtEiPdfja5Y0ZpZAM6lt5OJcbjHhVl3HCE1D3RAJ9gP3A9PTzRl2CBJLfAv
yRi0FIabxwOJrdSk0NUGHfqQKWsmZ9EFNFe0rChTNwQ6SnkRkm55xzvwMzlI1wvGHbxSNGrRrpFZ
sl/Hdr9lNjBJ+YLh5Kp9qVxCWVhwgfRj7FZDd2RCs7yNDi4DJXkzkpL+luJeCFWZcfUpyXdfaDeI
0us7g43VbWv7eSNqKymgSiSbOZox8OkiT9xftvsJa/yBeTA3VoLVPHZy0MWPffxD3GAmNuln9W1/
RpGP/30TH4J/4ovz3nHU0109rc2QDP64UrhJIAgsR2VCpIYEk7nEFlqf+kyAK/PHgIdLvIEUcJ6c
mMQky68Uhz5JYC/uxn7UCML+JBtY8RaxS6j2nwmW0iKiiINd5qPL9uB95Iuua2fA2hspt06d16TZ
b2MBIiIz7C7f1eEv4KeX4P+GY4Yax5Mh8qZYz+fDakZqx3PeIMNkRy+oeMNzEiKs2+Cp0Suuim0V
CwTKSSTMOPPatEw8ErmZsFkJMlgTLesMoFL6O14ee8ZS/78zS1iFCTMbG5kopCFLGnY9Gcj4OfpR
TEFgmKNOTVpU9kZdwB3f3s4O4LxOkpYRPl2meqPeN2iwSLtYwtZKDwV2a1Y69P8XSlQaxa0v982t
QPHi/tDMzjSrDt+HjlEy4s4mxLG09S6QvHGduZrFLkZSHoRRb19ErAccPWg3C6CNb628oFLccozQ
rq6aeJgk1sCE+4pp0U8W5Ge4PrLURAnZPqWkUq2R+JEVKt80Bf9CBDdcfHd2sy/mYEYngUJxtiLs
fjEQ1Jc2YxXqoVUet7n8fFtd3En69gjkHs34SpDdrfBuJiYdyBz0N2TZ7dhbvrLRpuaYqLhpDPeO
KuBvycuKO24TfGmMhikB+3qctl2motVcUImWt6WaKj40261J/q+VL1oCpoAcFIZO2D+CjPcfPJtk
nwPRbIJvMUC+OG7AeYImRZSl0E0x4DDoUKg13DuYHoinwJZLNdafi8/HPuu49FYx2cEMwLFzXdT1
guu18FsQVbGjrMS0blUprHxM2d4h9NwqOO3kgWycTuuYbmTObW62stvbzhtZrzDb1c5iTMuJO3bX
3b/ZxC4jTyvodyOrka0NpeHOSCYByuwLnANqr5OCB1Pbw143ZrwbXgzSgF+X4AnoSbQy3P6Usty+
kvCu71/5GjEbfNAl9ceAAuDrHt4sROLhAF/DC62oFveKwvb5FKIpCkV/9GCigZTUHgjriezx4Aoq
BIT1QxgsMlEF0w0NgKxesSWzoLbas9ZwmqVmh2BS2eO/v2TX1FJ1ZolG5dt1JuCrgyKgzgm6ljnj
g0YFyITI5tCEImUM7aDKNbE47JxwDsnmtVtNfSu5cdEtLp7U1wNTp8GbaYD0W+wM35Wqb16MLdn5
b9P5DtoXekJeTAR/QG9lzSIEh1rTtNlLQobYTPSYo4fV9hJkG5e652FiC9Rl1rhsdpd6C8TrtRg1
trTMt2maT9ho7Jvmq9j0g/G+yMbpSFR6+5VQevKHciobLCm4AJuXoMyfkrF+pHYeqtklUSdpjAdd
97x3BS5y+WllrCS6ymfI6Dy8sWmEWTOMq0isjudH2iUnr5RikGm3SIytB6pRW8FeMZmnM0guKkd9
L6L7/sTlVZ9z0g+3436mbawqoWBznrr35yb4jzkuHVBaZm+fB9ziE3rOZIdQeh6Grh/RjiqUrRAs
jz67YkRwL+GXU4hzcnLOg7zuM/H9gp9ccidTnIcAlov5hlO5nG+y8Si0vEFdf7f9Bo1Q/+flh5zE
S3fAZom2vihD/OmgnzZsKcl/diuw3E+QEUyYXUax7DP8XOj5hV4I15NFq97B1jwBJ+BWLd1oJylj
GmizBMN64wie/C/hPKSF6qV//7Eqpres97o6031YRwU6VdBLa8t9Cyv1lkOLqeg0lXJ5oxOJ6R5a
q4CUqnyrjEJiGuQ45SWRxglPaj51zrQ6r2Nol+3CzRPVbrmQ0fmZsJ+N6rQg9sMb3k9dbFNEVdtY
i7tIDRr2xZRq11Usy0l40l4rRZTSimX9PYLCJ5jBcZxJAy8e7jK/sDDnDuvQTwyMaf0Z0VRcdaCQ
7VUndi/mgPlRMTiwmz/V/bZVng5oMeMViW0Chw7YBQvCRVSDAg0R/WKCjlLk0sV3Hw/PZBPeOxSA
ldFCIYa+O/5GX9iLLU44nc7kbsw/1jkMGbG3JPPRzNx1RRXkM9ssWULG4NBVJNDzKCbXpgnZ9fnp
B/3HOpM8K8rc9woYdAeNuUw87/vZbKuqXj/t9uk2fYGM5zOLotxZqHSSSWf18znvtCXLSJhstqoT
p6+NCpyBeN7T0Nt0f3oYw2+6jMblBvI819LLsp1304ILPz65XHaYn7D/uzBfpSWJ6rv10jrazl5b
9uL39/AdJifz8lp8hNPGfAnaylyVpYS9cMq8/LF/ZZx1z9I3cFZGucvMUZs56Euiy/JXTau1yE1l
ezhpN2rb5vqTzg90D+9SE8M8O+aDgxpuIrf+fqvR4WiLs7bsB6eorxpZMcaRqJdk9tAlxSTVWTEo
YDUXp+LN/v++dZSE6brJEwxsNQT2ZRNuz1cmmbRxKoIJvyiXosxZK/rHIYFWt3yCV3OVwYbkFilr
78jKwSe7SSmOkERFoQw0JbB/AWeN324nTsu6f2fqBmT/aBbj/EJtcJ0nNJHSFm5eCPzCH59z8Y1L
ahUTkCjORh9gyl2Cz4aEceruSLWiPIpym7VyqXgNIwnrksYizv/xlSU6taoBTieXA3vgUrehws1E
qeHo9zJ5vvYKNy+wlB29mARhcVCfitYzwhF5MWRPQCYaLLj0uYW4j1aMq8feMKBnCmVJbByP79MG
uFPwmppD0TUtb4JO+W5Z9RIODciVKhpyBgkByZSX6IHQZ27Zq3OkY2SGNUny5UGbCz/Yb5utYLb5
g1EAkR+5FN2L92qJRQNb+QrGSOYWqK5ywVh3g6K+fByVptk2k9GxdUZQ7E2IMefB/iv7YwDf66DK
ec6VO9pAJcoa3a2e+9GnYyvErJf1Yaz46LrubBc/rI368QfXL7CyuVAfOSqxhFpLu1Zojbp0P7V4
xQRmYXwhC/l/8f/CsdEwc4SepdM4JR0PN+R/5lD8QGx8L18yXiUksMXy+5/HVaSG547oXQGDCFQU
1nZLYreEtBiQQ/u9bR3o/z1+OL0IrRs20GnzF5MXZE7C2L9CttnHqMo+ahEULHJDu/mDgNhYDkzt
by8gxvV3TjfZ3HF1rDzWiMFOlrhSUKcK36gVh/uRUmR3iEG0NrRzO3yieRQ/ETdS1N+ey3OzZRoB
U3jgfO2MVuaCD4MXGx9skK+n/pmYrXAFygy8T/PJc9CTCy/VcnuoItMWcdIl+Y8RPbiGns+23b5H
uPlWidiqPalhXcWBAx6pHm6C3T5e1kpt4iI4/sgqkIDuQcfUwv7CQWJXBSgaBEBVg3SaLC9PIBAO
Jn16zxX7WQa2eQwxc7DH1dHGzmXmKoA+FHAk95OzfhEhjxuvQvRoix1tHj+CahXFVCK+mbS4/1dI
FKQn2EBiMtvYSZE9HkfaeSmjplCNdhCP5hF2pWmpoKj+Xz2c1E/QDXuUhqEJ3Y0P4ymB5NiZDb+M
8lLpPrhW+QoCWTPr2J6U2BJVA/u3fDxNEnEhp8ymsQ06l3PdMlPc/KH6cxH4tVX6RLI1KUuO6ifi
QlKkW0HR0g+ZIEQ77NcKzHxsBeYVGl3mam9I14UYaK6eMtQmY24GaX3sZzFT+AfLqKkmnI7y8Vsp
6d4MHZolpS3qcf+s+UMwj3aeQNJF5oMc+IhQdKpLLdgDm8jRP8rzC+rxbhVVV6a8G4ltT1xK4Kcj
V00lCBnla2GvVt2enlr+HuAMIIMPKj8iD3kVzGv1vVXxanRazlaVn6rMEKcbw5zJSYTuHWUFheiw
tEGPKmactmyhTFmwMj4nTW/99Gd7NFWSq/8zxD5UuIsklHKTOUIH8r0a3oyduEh/+dKp7DGKqNyv
qtiN3f/x2qFxiuQ3va2hq7CaRP3eGyA4C/P0oyPGBFepq7BXfrG4EAIsU7tcxWnZUoLtyIxdBLle
59epXGC7sy6qq6cIJ87nAzjBf/FAQiMDnU7y1kqET5Shh7GGx0RB76uD9XmWlyRshXKPj+du1GmU
OkC4jLcqMiS5PdAXmipUo5VQYmwqivrk0lOfaogz69PRrrV5C8SirRm/1tN9JlOtwjFCS8ZOlZIw
b8Jo/t+PZoVJ7+xf7VVuorSufIKzIJEU3wr7O+F/NNXOW6B6umBYTcy9NcTWnKCd3pvvxv+09FPY
z9uqILavMJKRKN9uiHtjsBJ1HdxL5mNIp0eeDVg0HL6RewVBn/+ggXfqXOTyPaxU6dBBplzuEBcz
KSHo1id4vHv7qNzZX5P3wN0NnWKvV+5Sd4ULtZ2mN7ofj//k1zwaY0tRtlX/3+J94x52EtbSM7Pz
GYCQTFLwe4YWyGjxrJzITjYc4Wyt/ixi0aRlj7ftSALz3oDrqMAqmKAOwHjFw9ToDphm7mlClh2G
Qo6Li4usWEMf9ffyx9GRECfv/k9+91o/IQTiFINRgP51BHZF5sCmGnAu3aQ1zics6ILEQEgJ6Mjb
FWI0aYlxrmjEDhRfBYfxLoToOO1AaEsL5klB5DwdrZ7yfVZfcHAMTkZRT0q6tlD5cpPOsOtqYedF
MfRX54W+nrTK1Qr4xhrtTSzCeISaHaVYXTjiy7TtboI/l5WyocsawYK+tyZoUpTomn67hcPjjc8f
//Ws4ERjVpTyMjVVEBLnpcYbP8agmpYxmXVDjJ2CtQfqKcchysl59GtmrFVkqgvUNQlAmtiKfXtL
XYk9fZHaeMtrtq6Z6umRN07ov6WQZBxjrniV+YeUazIbHnHPOYm7X9vjuU6M8aiGzWG/hBoJkZto
MbqZ0p8pTT+MEZSQ8RvK6IYZzuFPsvfRulBL3Sxuv0K92hj4AhYqqhkKRVvFnf1qU4CdijzT5eXn
o+B42icL7fvfGtjHD6cHMtfi/xheiyuXz6/5Wxq8BLPDMR6P4B7DvEEKA+vwC+gjTqnx4YgKAgrN
lx9vRvhsEArzZpcNYSBuSOt/ExKoUjL+8aoI9Z3F/LS97gXgKhjtxFZ3TnsnQxP4yiB6GpTSqstQ
qZI0qoa3401+/eV/QiOc0RYVQA6q8ETWZT9lT/lFrNflMXvnEhUw3Qu3ZgcFXPHcb6DHw1y4Nkce
aYcxTXybbREYkb7g477pf0XR7B7D+ognoDBRP6dohX6rEYAniVO1g0uNn6frI0Xmj+UkqJfCzw2n
76IcxuvvsLXaQQ8j2pylQA7PLKo14jhl8DeQiOUJQqPucp50higYPZsce6MeczJo2m4AdI1Uj3S1
Et/GG8J0WAq2sXRKaJn1R4OXNTWOSWNjd5OODK3VgkT91mSSzQXUevaizyMlVfw07xPfPSVIEdWf
467/XuWGq2X9rnUPc6Ll5zPitnLM1hn6WtO+mmzkPjEbX/IuTAegy0eDTBSypF50rJVek27+GAuK
apB17W1SiDzeGaEhFP7t5Z4Ow+a9HBwZlk8NmvUpgABTpeuGsCpuVbTkcO52x+D3KypjqExTEGPj
APHE8DXUqLjtgRljb9dNqupjWoq3gRUo6+eAe1WTgDRfFOBVU8gFb/k33R/O2UCQFQebshRhh6LB
N5uuLKpb6HUUkhVyKrfZ9i2BxKRQ+qW4Q4inQUATPvotiogCvllByzk5rW90toMtxGvFQYC1GL6D
cVh/MLYeS/nX0sWExPknHGzhEbXozYIDe0DpIf6CyX7gVgR4XZweKVrFCyCHnru037+l4IjdUP+i
TvykB4SOw/9z8BKGHHj+KUremXFrsKxYyjVXxEp/H68x56uRcztcBlhvsybtrPbHbPKUSr1BrKmv
FTPBiCRNXQS03rT2DRo7c2hwo0+G9Ko1NRWD6kMguJQFVJA++Q9zznOvFr11nrjBrxF0nGAQdc0f
rr3eo0zWP11eXYqEhUr+m9bKK+CTeTDAR2pBkLlnE+UAve6gz1tdKWNnP4l9mwuFzQUktub9cKMz
wa9sxPTG5AXRnmjnkrM1RNiIByCV15oBAhPumSEX+zGtBAq9gUcCiuf9RnYYPPxvEE9q/tqqcPV+
VXmP4w+YNLIqR8XZgYc3Qv1qrptrgbcDH8jdi3Lz723J332wyqMhAv4b/0D1ceXgywcr3h/uhqf3
50OHNyQ3jj3IDGbRmVfiXP8aWZp62ngIQsgbdFnIiPJ8ME2mE6Ty+r//AJDgI/fqsMwSGUj/kM0W
oSAIZVqkNtf/J8OETbqNqpOLVijNmKgkCvkZLJwv0V6Ln5fAs2+45Z0l/D1PnD/76XTLgoLcPd0a
F4sxnz136F3DddJOmvJ+qfmveDAyWgcTch3LLDrLGVZJaPLfXFDvusM6lt6IEETaLSjHTgHOJlpG
T2LIWA7If6ozH9p/WrBfBog5ORvTUnU5zukXf5p1vb7/dj1DMGx6Ez4+/4EakyjucpSf57DcOWWz
bxTduBQBgMGUuCHHS2HuWLjmVa5x+OOWWhrKH1ccIpm0XNEzRTn4QM6P6M6sN0yupt5ki74Iie0j
R5TFM/Vlmx4KPI3i0HrbrSRRNCmwVTv8w0/NwjTD+yGAgOtUcwwIOZ/iYxs1Z0mGJUtZPRncSluY
y6viGjXwc3ScEmanfeuCGEcjYCvirBtK2Tw/xm1FMmkpX0zEqtqnjiS3UJSgqQKDO5yOdwsMaoBM
D80xlhi4ZGiFOauESFHcQWnJVx9GqcZlhC27E27CFzmu/sw6IKBzL4sRzqNRy1r3/CSG5neWmc2k
W8nZ2NrksdSJqSSW+kd+VG6wovNdUZxLx3YPhQ/8moyHTM6+KPnYFTMlwmd5LDoUrM5Mos6U7R2L
xvzEI+X3vcioPaw1UrDWSfN4y1W/DyrZWUegMfMKURqzRvcQwQD7v3KfU8snAUaKT2s8kxaxCkF0
4cZK3rswS0M7Udha4mJ9lxmbT4Vue858yiRP+kT8Skvm2CC96By0odBo3hiyoP+MOtTtC8fKjhP6
XKtJjtDH6Hx8Pzrw4IR0fo0B9t53K8L3f2Uk1j0w2MVt6NZ+Wk6LJsBZgQdcyGWAHLb7jMnkuw3G
xd2rSyOc1edl9BvelmtFb2DHTPRsL40ILdkgSIo8IiZBdWY95n8DSoo4RA7cTob7Kpd4ikEk1YPK
iYGxKnlj0wocoppHHRy2wvyrtgVQ3S8qPrOSj7mi6uaU/eW3tP9P1zwE/ZFaSsUZKKifWii1lb69
kXF53LwWBYcpdp85JaMeg6iZXkcxJIXf1d/uIalDfbp9plnWCkEAq0K2FjZr8IdLLrXwOdeytNg+
hmhpn3GLzNDp1VLZTGHcmQKrQ9pkQnUXOOtVUr4MUTf66ZXfuqI3+4kUDZpK04n++Iklq2wQ7ZoP
614fWNpgdL6y8oTFRecMoEUPH9kIeY3sN9iGygjcXiEx2PW72HBVidoOSjrpKHY4++wuke5LH1BT
PEsIDf37BY+zCVYla+OWjv7trljqTUIeGGfH58zNkVQ1Nik5cHgv9oggnOUZid4Y1VKCblJ6fTYa
DDnzWu7WHrNXFBgOyy3OlCSQI82yOYBDUGDTB0oVuiS9q4rbjPMrYQ5N/dq9igF8L9OnwCoxmzOf
37fSAWv8+1eHjV3gobCpQZC4xgSPGqKO+txPQiomCWI8qogxiMnl/OuaZ+2UIFP0KYns6tZ3x2Eh
iDtCEpincYcVL0tW1IYeE/UsMuV5pDcg8wY5pYFd/fn0pt7ugKd/I2M1VMlSCkLoVQAl57tpLha4
+DCRcM7F9pxuw159O45cbi5nn1+DPZSpoWXFBmI/Jn1vQEAjNNLKBIy1w07CdpMAC6+3VQiMOAdh
oiXH94udIix+4Sv2DQ4Roa1zVF4OT2Dvqzvito01GfZKY5NPSJ9S+fIxWdNACz1zjHSIi2eUb5IF
d1o5dpb8k3z1C1P75widhUxUGc5kffLYxy3bp4PCCFYImIWy6SMXvKKkMi166Y7nCN1a5k90AkwP
G2KUOY4n/aK9Tst68CsGLo2raXqEv4lL1CX2uPpVcipuedq+R9XTUA93fviPyDvUNI3vI/RLNVSo
xxg1OpO6Aspc0PMAZgI/VNb3PCKsWSPBc1UUuklFrFsBCdpcGbZv6zLu2QKJ+0uYMTO9uyh84cd0
uoEOtBw/SnSpFGKWyXJTggTtHXVC6otPtPcqDcws9dz1sVTfJVq7y1g0ZhU6Dv3sYDhbUecIai2J
oG6HysjLtZB8yx0sh8kZDodON8yYLTgxSaPibNkzxO9vcSFcILc+4S8skzyTHsRJ238Bso7c7bMT
zIh83Zi0f+zzKyuzJdSQrvag9FqQVs9HSnBmi7j3Q6/JkJnlBmWim0zLnGD2lS5rzBbDtzWsbr2c
iL532PbNfjBELBg1Zpf1/pV65BY/Pd+QpaYy7QD9gJ2j7TSMAIB+eeXnjn2WP8mdc1lE4dJzxOTi
5HQ1vcDoEBMq0QP1yJ2uQ41YsnxXyudJDNh1pgwyuYPKySMW1sEgemjREWPyNu50icrGUAtvA6BG
/MldnOkp0R4mn4aC4b51SC1s9o8UYQ6IQDWZcy1q66dATBfo5Y1CK67iS7kyAsxfO44NtXtOJQlS
r32LnSpDF9JOmPbHiRvuO6xGJspNC5wWdRu882QsFGgJD0+0tbIfOO5ESzDV0pALkcNuhSQPyyef
R1gSqE3LR5L2ZcJat2cDO3O/x+wjnksmyZAXrnsBm9Hy/rR0PV2Mz7rD9RI6vA8+u4HOl9oSoATA
rA2u8yogfDPSd2qkVW5m5745ubjQZhBru9UJKJHb5SH8YK7/r+mVREGYL1YqnUh0Ho14h/a5ilX/
ctRWjgJ+ZO+HtVsYsL6t7kdy/9psoHZDujL0cK28/5ARSMrUAph0xgx52pXeLTzTKCEE+3FZvN+a
vKQ9Haaa6VlVr4W7tv3N3kc+djndM4ZlXVU4bzsmF6XMhI8TXv/zLKG1wotKbcDqSV2ThPESL0qm
TDzxy5CApcBSQ/hs3AymIuazpAExYi6EWDLBhfJYxR077d7zi5d1ABiTnFtmZizN9Mw/CgB9tyUI
JXQud35WarOXGy4BN+Bl+86vsEahGkUrL0HfiycqD0y3S/qAG3sbubhC+hp1ZO2u+SghJnE5ULfE
ccS9muqfvWP4NYsAdz7zYn/W4qzQWOZItXNAdAquhIjNIGvay5uwlh/gxjcGlGW0vNphnwRFNca4
SwmLbwcviX/eUaJQtjguLUZXtoT3m3Gz1/Q1DtFQuuR2N9A+LqBv/L6H3lDoYfNHBbPGXlmzaiOl
QMO4BVLjsXQcaNU/BOvmDtn+vzF0bXyE02vboodYvRYcGwrQWU1LvIN9mxaXkeBSVsrDaYXg4IQM
3HEctAYskR5L15ZQoqOAS3KUa8O47JneZo4JAK2EX/aKTpahoPaV9WwrbZxOSIRGZ7Ui59vx/axe
F5Wo+3BBJeNR4VCm/L2VbHB8pxtJpEFlBaWBUVRGAT2jr1Z6kvSf+hsBwX7Y4p6oT9DjVjlQY+fN
dIFdNm8heidvqTC1kmt5wTb6jwE8NlRKYhCa1dhenLYPSfcmwngUW78ybjoaZihY98Fr+2k2vflO
hyGtdMGR54gIJt9y4TR6TtktKZbznBsoA9OfyZoYVtTNX2fSK6kfUBfG2RLZNkW5OzGq5ACSGHLm
Xz3/HiIkV2jeUo6auMdMZJBz/3NCPw+lIBXzTvESQ2aJFYTQGQ4zANswcfzT+YjZrlWwihQ2PoRO
5nPXyRLb7TvKG9/oSJPc1hon+QYsdaxWac7adZ8H9aDY2VnCqWKcGtpc0BGcMtMfIhsOAKCbjuqs
YnWJU1IC2bxUWoEpV9G985oZiuj3TTVFa0RNqkWbUtfR4tkuKCswQNx0Q5Ri5CUloGIjBzJvnVw+
CL5J4LschZGRwblva3W2+vBM+kuhDi4XE97FRAp5Nl6jOKRW67JSISlEX9IA2qgiaL4ktgPeRLUn
yGzvcMlpD5sq1bGlUvMCf2lAyhFREivhkLdBYZnCkFy0/2O9PhyKsEfQs9TIrAdvE4fTw9y85QH5
8BkfHk8/LazTcLEKYtWEPDZcj2RLCyO1eIsCqPuZREcozfcXPf+a0XomSLXfTBSATVDH8BdAgEYY
GL0zj6BhdhDV2e29eMlT0piyGlh6Au/uILU8DZ8A1Ws9lJunxI4uGTm3Ascmwk1VW5ehk2FWnFhj
DcH5YORzYAUXsho8kx44VhR2OMY5jgvlmV0C3z5XDJ/NRwKq3tfIksZGuEDbeSVSsvjyD23wxsBe
kXORqeH4ZjPNpD63G4LN8Xof+SFc2wcPReCvK+hbi7XyuQNiphzObUIHLWSQ5IdbEjFHOXO9SmVX
ZZdXfMiphtpdcxoXK7CE1F7jx8PioMfFcYUvPQL4sn427fY2HZLgtmlm8MF199X74L/nYu+j48mP
+X3SosPEzlH9DnIp2+X5Zvok6CtBVkHkVflPbNbo8P5CJSwalvQCtrZGKg3tPi7D0497kretCqRf
o+PNsZVmuobawqVIAtzo3W+jpT7QLc9KE72Vkm4eyEFaRczBbHB3MROp6X9ehDMWpDfVGhEDzUC4
QzY2garPkdpPJRXQcos6CZI6l+ABkfzJMEDs4LnEZGS+VD+2vthcI7GMFPpL/d46tRG6KoiEGueG
gzf0xwR7u8LS12bDdyqYdSAgiZrVNZzQZFnaSKeG7omzYVmBFNA6JwwUmrosv68+uQhBuFQ/DuiZ
CHKIRx9Io4ZRbVsQOfpW8M4KPLt13+Vqwx20QH5aSC6rr8X7kE5j26XZT3U9z7rmsAbPEYTAiErI
JITuGRxlGfB6WgOlyMzaPuvqcPio5hRspyzRHgiplNOZX/sSbTMgNT5k+iyp5j+cVZY3UTxg4Qwl
3+wGINOItoQf5M3HtwpXCJBzQd8uAN0/s5Bmxe6yk2Xd8joYDbFyGtzaLmvDFqvpSPHkmU387OVh
BIB2zxocWWUD0HfmDFYSB5KCviJo/pBIQcfsHLHAXfVz7aPRfgAikZ+Iz9n3X/Z4DDsYV21JegPt
zkku6dXpkgwAhObpj9TX/mOPa7f24yHiNUIK3iYurtvR2NKNSR1GvH+WNDYHC4uSC1iQN/fj0Ryr
ZSXBDyZF5Vod1a2iq0wk86ZQ1zsZSwAYRDkM4Jv8m5Bz+96oNtQt8mijK/5E5pDlLQCualSR2wai
apVPi55x3DHkbu65CgTv6dvTnQwpSstb/+gD0zfViF8ueEmNewyOGrK7waIfwBEyQHo2NCgQG32X
8Nc8AEOHB2tAzNICEQR6JmzKSGOJ8qhWNi6w3g6Cb6ftsVnLIrRVxdX6dJsUAnVr320bEQ/rcvRg
2StLk8+2BI9Dvb32fLQaUVOGkvWtdH8kt6n/g4xpceK2dEFDjHmIcKJy/E3tUKQKgGNGjL1PmdVB
vmYWnzA5YbiwG67dWPCYfTCQbZBI5Dfh2JwAJRKATUofEHWMeZ1pajdmjBKZj9WKU6h03afs5BBk
lk08B6Ir9r9pAsH3O8TLfwf0oWzrHywkarFe6wL+mN5hGCFU2ep05Pt9nCSC8e2XAElwL+8TzN2g
tmn3WdfCLpUaJTqKzlJOm0GGAi0Tlr07NYQiK9u0ZyMLMaghw7H7oGQbYYiaea7By6FcREop95qd
kBJl0BI12D7V2ZjpajRRWxnimAm/IDbg/3yBTEpwws8NfzFzVYRLv2Rw0we4du/4T0KnFgUuRlb3
9vGviiGb1+vIh94ZilLf72+8HQ5SvxzhOgsV8JiLEK7DGc1cKgArpa0l8B43yKYpyDYk7sMwYplj
nU9HbJaPSG5kKoBIKualeZU/l49yTod8vSty9Cp7s/TCGSinnUgnBgMWZpPQnQXtU0LabYcQZ0ss
EYTd+/LKALj5mIxQ2H2H3js7XAhIc69q5qjzZ2ePhMnO5MmXAp7YjFSPqsbqdsPNBZzB4z+RSkT+
H9ieTu2r+kkoW1do4hgvSTa7is2xkq0yhaGIygWYZN1w2DSRSJSZGUS/EK5QDsvOCMcbJ/gEO/7q
GEbPKE6yg+qKjY5drMj5/3zdhjRTbxSkUWPff+KtBYjsaodLE6OS3k1wP6kz/i1B+3kHvwUWoIMq
NdfMvyH6YDFtuQcwpSwOxKLSWZxWVN4XF9LYhQXCbjqPf8qOsIVf0GhbeggCpfxQmRU8DT5RwjhX
6aSqMHGZpcrsCyZhvv1BqA9gSDy2G3CrBO3duMaK6RgZxulflI0tPU+eBF7YRKAV43oTBVlJNBzA
szeK7Lp09Tzz0RkFbdNiwwN0SXCIzu1/2kvAqj3TmXWSjhjuHXsMQCNBlOhryh9mAd3qTbfdGFAf
0PgZn7t332IHpxAH8yY5zztv87iFZJK/kgjKRFncnVP/eSDultCaVYg3I1+iOm5UB4OUD2BpFKVS
M53CuYYet0Pv4CPx6AMk/+OsRCKk1NYDKr0iRH0QIt/2AIhPMw0vEZrl1SbZnJQO/z6LeYNvyqbC
OidChh5InnCQtrXVSDP5RfXuNi8cpZzsOClmgdh9rkXslWF6PzmSPxGX3yl7aXPQ/Yt1DVEKl8Jk
RcWT/GyX4Qcxe020+XEIS9mQkwlXByWWExaXvKCR17j/fQKBPRgvDNcP7pCFCFGLzctKpDdIXOd5
SzdE3VQcpHUqQHmSP+5h7SLGmF/5VFJHAC0ZxRXIf1D5G2aCy/bbpnj+jGmF/dQ407AuXWP4yOD0
xE0aqerna3s9Xc3peA1GLR8dhzxI/GoePz00pBSshNIJDnaEET8tJvp5LixORLRPxaAkJ1aonqtE
uLyESs19XFpwY3CJgqKD9v2UE4zFZUZRjGSO30lS2Lh/HZCdt7l91NHZ35hZ6fSUl4Rg+7TUFU8b
qemnTdZLOkIVVUC1+iWzs/5Hy+nbWdQGvFPNsR+5gxNPbnzX8SxUjEhqQpYuXmZaJgQhmf+0UNrh
rK+vGyHPbNMF4WNSHNeeOHhuNasKE5KKNLD2WBMJOcxI8QtS3Q5HrJRErOSrH64F+mS/oxQuUS5W
ywe7a6SXVU38Ye8PO2YsB51XpBdB2mbrZ2Uk2Tsx/PFTuhHzZkfCwjcMZOYVZUa3Wc0EHvgSJ8hm
d0eF+d6sjB57cNavdZmddyP/oGK4xothxSYe2NM0enUcygK7voW1ogznSlfnCbG15+wZ0ZImpRae
Pvh/n3fBHin7iWgumfXWajagkQUfZujLVG927PYy1baj0Y8IJ+CZ0v/Fzqw8KPwAbZ24GtOfPUZy
NZHHISRJJaEL5n0fy2Z9eE3hV7qjqVwLpSqm9IMGqoFobxGJO8yw9l7tOUd8bKtvwPtV4uuZ27g5
9Yl9YxAdcFM4Rl5beb8/50AjWHTFaIF/1zcI60S5nHmUGX5MdYiQaryAIxgtY9Hq0pvd3173qXRf
CW8h/3l6K2O3dbJNVh14HV2qkaABtB+22ABGeH4GnuNlSCmnomo7YFI+5s04ipEfeWSYCz1XPb88
Mv4hLTuw/5srDgA9IxcFN/9JRSBqTY5zWl8FM28lEiWkpOWP6/f1YmQsbxe9N2y/Z2OE/SNp2ZSH
JP1GWZtGlV9s9NCnH1hzrJvrTwEyGqdHm5yoOQFeeNwpXD9OpIlTF1XmAUQoKjS+jKnc18/KlxKI
uogldybc2ogCnTE985Ij6ebB8V9wHxpaN2CK5Ut30SpGZghJH7FpjNcIhLfYd3xV1V2nGGs/1RvU
OQr8uxpttHBFjV+FzrmylF47DkRCQgVRPiNHsEfBAGPwxFRT+y4wigMqCWT+zcKR+y6QdnMPm3Xe
ZWsd7UouNCh8G9/Z9XlDdyQjcS4iTIcJkeIYIwOoAxGy1+mnof5Q/1zJn5r2ze7eIaGWHbamS/K/
8JYhpV4zP9vD4upm5dK8mm/81V/WNLwEjiONXCGpQofqRkj8Y5ASKfpg3Ju9/0Y5ygTT6U5H5ZMd
/QD3pqSyi/ClQCFnF9zFfrOtWgyx78Eor2Z1ZsbZM7g2qBBrqhNd9HpzxZ4fEhdNVJXEWnX3C4BW
+1p8eWB1AQA8T5strLlkTT4g8t4JkBCxcfuy2d1mFAui2Tb/0h61BW7b6g/91FP4VncLfZyfzIqF
2pWK01w/naEEJQV5imb1HUHf96dbbajJ98WZnz7D3kc0bc4/sWLsp89da8U7BJkDgkTm3ylOPHGD
z+JQ6nNSMr2qa6TQDCytC5ApSw8Fxv1yPfH6LdpypAX2qG6nHv7hp1e52nusSViwxq+P7GfyUfZ6
TzqggJofr3zVsHPMoopwJ4nGKKneEw/QlRBt7JVJ6JNs9WEAIsIVG3SSJGBVdG2Kmx0DTojeSWCW
WBRObfXHzMYwq/QOsyihBL+Co4UfCIdHs2I9FMK7Luvp2Hsv2H4WhUqcxqK7/s0LzdowA4WJ961b
H3cY8WVhkYzD3P6h2/S5UHjWgKbgpHffp7ZwJ/briZD5BTgHspVj5ccXZRfP8njHupJSjrEWSqDR
/GAhRwJBUrC7S/VG7Yx4UWWGRoOLzchN98fNA7ashOAuJI2el0w/NwQkSCOFvb7yyPjtFZGMluu4
HH75ZvkAQhPeuBUosgJeXNsUSZmu1PP9ufVJJ6S+n0upG/hWcWLiSKEDEysh1S8Mr41d2c/Ql2TK
8WJKK1BL1ytc3uY43rgbSi5lgRWet9i8LS52Wz8Y7fslgNR2ee0Q8PeixQk1Szlo5onfwIYwRLzF
o0MdlRAfsUFE+2fBPzkXScf4gO8RZ4JOFL2m5yoCRp4pQ/b9+Hd0E3f3z2Mce8ww9namqLr1nCi9
1Bs3qUjGJRQMSKBymjWFly/cPKSc8mLaB1j0G2CbVbz/8Z8diLdMwUSdlNLun8A5kvhpDMUnitXp
/L3VHjncrfD6AiJl3Zr6UP0hA5iCEfTRdyy71Zc7SGq9hgjuI0xoddBuMJegm0AavXbc5Cxb8LXD
Luy0qKBpHmsCkWQu81hnRICcPmdpsKejfaX497XcthaoNEGKIAqbVhjYMm+i9lc+VI7Um3GItpMO
+iubg7xFdhTr8JXEzMojRHgQx3Xduj6s6/QKs/PnSZtnmyhTn099qZG7rbjjGtjggQQLNLlfvyE1
tvr2dF9zS/xZ75I8BCcxYXjJZtIFjVNY9V2/KR/oY0/rqqSWBu8NEkFU+hqEo0bxDlT9+au/4EB0
b/wJYYj9IywOgAEtV0ZufXDYHHQMeAKf6msRfaHrXAm1E0dtUYKK35DaNIcldLczW559JsRlkcGb
lQOJ/NW8RT4HeUzBTPhF6S0hNXH5PkqHPeMczBKQUMsA4IZeE82k2LVRKyUntNYmvLuqb5eTs73C
rcYcqOSrsz9diFWHeSsUil+/43t8BIsyGUFVaJopuEAi4WUaOfBXWNT417GZXzOikgdtMCwvyzPs
qScQWn/vgiQqv/+Sb4K9NGf2FkISlUqN5gHq2lAOK4NvLhZ0hA5xGkRf7AeOZybzCerz0NN5rTcS
hT+aagHI3hNqVo34KtBW8QuGa1w8w3RPcnCbPq0xH64TFNOZFb6lTQAvgtnOtK3MmbyYgh/uBefe
QpSRkxIB0lQAm7jGrZ1HffrTe87i1bMP1UfAHaeet24aWUMYh+mGErYyThPxzpqsU4eccTPUb4lS
5/GfFtLTaKruBpZSZKdoaux4i2s5d1Rk4InEK6KIjX+ik+6DzfIZifqVqtcGsKA/zDdorlmfNzfb
9pad1PXjA/qnH4PWQ/U3ueb2fXk6q3AqdR0+QgSSIEifEP2koxIL83HU5VRznK1WAjY4VaX8oAI0
y2cd0iB60zeJbsX1BlIwYzVxwauDH6iGpyiSFTm1Ffw5KpmcU5n9yc+F+HnrNAYTTHVY/T/11qm9
cf8svEn0z5C/jsLespVgb5MNBV3FFznALgFgivuE6SPxPJDnNvan4Im6Awp+7p5vAy0uffp3TId5
8bCHjJ/esFHYt1eLYabNJH2Teo2rtAaKHL1qIGJeCPJ0CBbdE/9vxm0FtNpzdt40blymPQFw6Z8B
bWUiXtAUOrFwmS7aT2MXqYK+RBJcQF+5htLU94qTPw3wBHJjHgdDFUv9My7dWt+5+gCaZ0QMtgF4
WWk9+/qYmZ0fNw0jWxc8LIg0TPTUMqSMFYmZOEVNM+G03Fz4ncUuRSPAnn/PR3VvYM+WeaKI6DmG
hKA7sB9l4Wo3vvg3imQ5Sze3kdhCwvJqfarBIZdQAdZypy6DYjfem1vZx8U25wfe2DyRI9bzN6Ae
YuxRFSI2KEbGtD/PyMty3MjdkECk0omRWssvkx2xSQwVqRtYOxTXy5kndICoe7OuwRgPeiniVqoj
Tq8nLJJjLweGNuvcGKi6zntqYVKmpxZ+PNlznOaG41TJUi9elHv65+GBB68rI/UJ31RAATxwgRY/
OvkpxcyS9SbJ0QeaFVlsaafY71HkE/2aKGVRiyhnl97SXwfHT5VHeopOPu/ywgpJIpDiJmIEBA4b
TXK0naa5JG/NFv86HGbSgz8NsV8FPG7Ij3rYZDOaGJcsJcSX0a1QeNm5emp4WOSGb6c8EpzY6u7d
fnCsgibZCBSVukSsdlNjwAMh4Qeq1ggBc5Vt+L2u4oGZDOsnq5kSCjbn/RZTELORSEs/14h55PsW
6/XO65uTcBNKs0yUe60JMKrlq/3dncPhoo4FBPFEa+pRUdDB2efw10LwXh1lUdXUf5IHVEnHyf0j
J2j/cWSHdX7h9l0OwRfFPKApefO4LStKrVz96tWVGAhfJu1v0PZVtAmazI+Pb9UZNNvLMox+F3Eq
NvFpqRhtnc+AMUQAH6nuTdv8eIi9d9riSczwaP8e9K+qd/bRwpJ5IzyXvNcR13kw5Ul3L4lzE1u4
POLRyUhUAv01feT2OnuObB6qfidLoU2zg06ipC1P9HWAgNHUK0IoNnLeyh4j5zTeTRfP1YBupV7u
8YiWzJN0z/NiU/q7ZJ7S/56zz3wBmT5F0cOFf1rouS4G43XSENyhZFaOIMzdRYURqfKeNuGbrT9z
Gm883pQnJbehZ5LTOdU1Mw9meP+JfgjvETKDb+zHqFhiv651nss2IUZ5/wXXGc1gby+J304mit1Q
i54+Xyju9Kd8/egD7Y37T2DXVi2YjJ7FeuLVRPaji/HyQrOJ31G3R68uPx2Wf7JNbesw3Kg0TVRF
e3la8lRYtCE7h4OR07KfkAWYaIzy04sba6gRwL0QsDVn1CzvTST96tQAX/fliv8slShHOQtOHnXx
WjP9u9eHVFZYosA8tNPuxJXiQRyV+1791BnRUBaM//LAXHVVfjrDXXuAmMEqCn6G3bPJsdPDJtjL
pFedkfNBle8QGZjSlnJkukaOdhVDTob9Pr+DhdVaOokJCZ+i3VA3aqZqtU4RUImq26FaEVIb5Q8k
xec1Vt6PgAPMIj7KMXZl+cpMCg41MeYI3X/ndLMwD4BP/nT00P9UWh/oqohbCsO3f/iRMiz9hOhT
ghi3LO53LnIWu2yqr1LQT/lA63KfD2AikAX7NdvjHGB5rG/LkInPXkKgza2WbOEK9fvXZ6P8aSgs
0mp3iUAng/5IU1P7OgHbjUyu7Q6kQQH3H3VT9aelpbmQK0kWgtX53kgCqMCsDD08WA4JKQEeW8z7
vsBtpJKCerciiJbnV0GYns4LcyBIKO8oMY0Cb8UHzSdrFLthTnhqA7teXAEDXq9O8WynZWKJju7g
aMNNoMH5NRu/7npiphonqHuQMJmkJn2u+yxwEJaqtS/tfxOVOoIoOijByKI17xmam99UZV0U6xSj
IBJAvNDTpFFobSuw1qDeYCvRHnK9EwafzsEIfiIHsNFvBM63fvYWtEbjuJdlZjmFF0NwhThAOJAX
DmOqGXfwJH/asvoMbbCro/M0K0YE7GW41jjGHia7LeXdNYxw8lytXnKQ9Rkz2dBExYENlKVKhjRL
7yBJpb2LNY8ca/6A2LjuLH7BOzyNgYOtfuxPFyVLCpZZIhvgpqU44hEQJT/WsQjY2C7s++owUl/G
sCUZkuUV5aJuxVofWwSJhCd71HOcp/3+EAj95VBCOgiYbVZ+Arqw0nj5iI2nUzmqeOxEGwnWJB3H
1xcC/tPDKEF7AwOVzH+sbr6+7IgOR4AHegdibkIE0Df0d5f8gd6tw+RwimL+RIwSJJqpuFGriPUM
tHfDq1y343A03NL+dlQnFExednFw6CcANA8Z1sw8dkysxMLZQvo73wmtdK47YSVBa0OGLI1mQmSR
0KkzbsTWZeOhSp6LeuLmmE7ME8SaChbKpXUhQXQM2DOdQxMZUDrwVaiV+vZylZr13DUkNDi5/41w
53IHHIEknGGpJd4Zt/KiV6hmEMrbGLtHLAVvN8KD+6yaustrbizAPM0MjogLCcnerNQ2hw9zCPRv
B4QvB1ydB3bdeDf1gsFaH/Qh++Cwxhx6NoJXSwDYcViYny2EqvYgSfohbaZ2VQ2dWGuQDnAKFNqK
eDXGfHtjAK2bPRGNIN3/kIWOlV0FTomZul8CRijz6Jrr5SGGUUpeNfN/Z3SWrqheFNeZ2FD5k4Hj
Knr8HGluKLxMzydUZXZDqo+x21x+nZQwePHyTwB+9ec5+kMsDgUsVSF1Fctbs1zcHDhDnL4JkVHN
+DiEMqtEXC0w0/UHkvXbr6NwMO/8BoJaqnPEwzPbsBy4Xt1y/Z2Yq72sVLbXywlsclzjNwTlgRUI
9PkLrDAQ91evBDdz812PvroqdhuP5RJRG0aCHyYMToyIeBYrstEL7OP4mgaBGAgkcjl3Jnrig7Ao
EcMn9NKOM6GYTHskewtmK3c+SUG4/GDjQiLYj+Kr0ARuurvzptlzw29j16DQgoCmyQBadLmHPsJH
E5P9ZMpoRO959/rp0q9K1jnLviZQ4I/PViSAyeHk7efeTpasjrdlvfXHZ9QgDbZAwC0drvvQwfsN
zcMTS6NcgXAqNhUDozGXkKc2x4Z2uP/e9GF5Vs6czxrDmfk1fC8yr4lrwm+xbBkuK+srAgWwG+bj
elACnHYyIozmN2s/jCg2R4PYY1kOM3D81K71dMAIIfYplrjaiRnW7dH6KlEBRnDDKjYxCF3yqAxZ
kR54mnXoR1mA0RJA2tv+Tl/TY+aA6dKa5AzrHmNe2sCyRCqCOpAOejqnT9Rjaj5TiWBgWnyLP9rg
2F67BflqRGXnXCwAbZGLiXQOPSlPSF3SJhvRE/mk4CjKJP/iwDj9iwMwQDJ/eZznUr8QJJvxv3JI
eiPz1NHB/PoY7HVOpL+mKlFuJiuFmPYbJQm19DQuBp1gmqtlsZErYtB/UZf/YPURUD0RRCdPRGqo
4VKow3jfBNBFT0yiXhw/NmyAZE4PwpvTNJJYz21/ANN5nLQ5wSpch4aAowDJvdbrCAA1xrpIgIzs
4I+fb/EatnGHclw9P+av+yxuGWR6i5HlS9w/pt4qxdyg4N3cc/lGylow18S0xvsjojqn2BUZEYM3
vDzShH+SJq/xOckkcZ5Y5BqWQtbHUvXtWSq/JBhaXZCxEfqWvWlhAF3XSDXKYUfm7cUglfVipYIR
JyFLPawwGR0fTRJFDL88o7bgRokUDQDTM3ah/u4bYlIm7DoB9RXfBjVn8+HW9OSrAxPBHrX2dtUW
jUT0GgUOmDa5LC9ArKtH7+jNW2MsVwXMlOSYuLKbT9KS2GFXh88VBViUzLwPLn1zQ400V56JcYMN
wbNgzEUrioIRzr+h2UgFEycbiuWSyWcolwo8q8P8zYCNv4fSM9Lzsfm4jbwNqJVTYym8pIJD99iR
aF+6Ip0olfjE+p+QJhzT4bzuOf71DgpGqrKQulaDoYiZ0CqpEk1rCxl1/646PdrYikGSu5ZO+Y9R
E+P39R0LlzoM2I+i0CgDg3nsVkggAfTv2cIEZFcX3wSJD6DNmSTQ2CnSL3/t0tvax2EKbGqcwMI6
DrCednhQzG5oQKufHqGvOQWT27SRbocSEeJsGFrGtrAaFXsXCfjWAQuP7IUfmbEQaB6eRPNt591C
Hiyk7BukuMyDySwQqvr+88npi17MNU5gN3QtL4nbtwNnJ13uCiiQarmRkzFcwiIZbPKg6l9NfWxg
2R8NGge64w/LZ2bPeaQG7k1vlrTeA4s51GoADVLLkPRFfwf0UI4NQd52M/V2sK/wMMctHKAshWGP
DPiGxvkd0gIEqqkbvYPwXMmMR/IyIxrVhso9WZkWsbutUZ/zyUzMoar6wUHQIXd521cZ4N1KS9h2
d6BqRDFsvwFCXwav/D7yfrhnejaiaoOoCdBOixAvcuUkwxbCqEYuZzb2mhDFpNQQKuCXQpSH1Q6c
K/Ql7YuBx/TX5ztDUF0U8G01LYW2+700ntRkZ0180ZtiaFuipodQPTccZZYlcQVAiRRUcGuwsWKM
umfpoNwyxQrbPK+WKX/OSENiS89ExLac+B9uRkojchHP/zGIP+42HQupQgFrCbNBJUWbZb+4ZFAr
XoIMpMjQjaMomPHSxLa1sLXxhZKwAoQjSAPkcAyIvYFQgoAU35L6u63Xh/SFDT41LApGhNGbcG4z
0JT/tvKed0XnrAo/QMbWPmBcs2Qspa2nXjpr6T4K3wOH0htE56pvm9sZgxpY5y2aBGNgdR2M9Nhb
jNK3OPyruWfTUr2OrSy1HyyMXDwdOrkUDRcibMxvpjhvOIVvpoe/IZd1RGtvtl/mg33rXJuxfJ8l
gbrgZ2aaHwbxn+NEKcZEHeDj2/i2215EdpAoN0CbZdBVQekSzO1iRNgbDckNB9/SDL9sBjs7B0ip
+9qq+yp+Bu/1y9B/CSEicDuncTQR5DSwtdu3ekwRjAo9eZfb6cWQ2kbUACYMb7MYYVVecy+78N6Y
e6/OBNOhiC9CnAJO0BtHWUVa4LIaOuyknPXZMGF0gq3bj+64HW8zd9giN1fgnEPAn+wAB0pflLQ9
3Si23ZzTw/fK3SfnIgoUP5eywIpem+lH6Z0vTheE/LO1xWz2P1BBz8CC2IYjXXL/tRrpVGqe3aAh
vdYBE2CLq4hHHA4XiW/uhPOqZ0LwlMbpSncyiUoSTqCwQycPUaAKKFrOqjHk1+iLPQ24c8a5vxSl
Cu7onjqQmDSK7Ha/MSvOOSp/Kj9XonzzitzYmSbo+YS/NsSHSAXmA/14xEDL0e7uxNxogKh4gS5g
dCZzBwzLBdi7w++sJjfHU0IQx5ruw1PhEIstVVdHchBhmUZK5ca9G3Mo+UJnQpJe8yFwUf6oeysc
v0ZOd9fPweV8RV918DrcU3BFsJv5H91Bwp3Hq0ldOvVOgYxbaYZLC+k78Bd6GAtnADCU+5tdVbNM
1MItI8BOOBglmQkkYVUM3AKOc4ZSYJkoKLeGPVOr9RYSNhAVWSmAgMFJkNFDeojBV2JTioJ23XkM
4LgwbbE6/3FYvwOtKPfYtigiBdV81rRQPPPqcX5tlOI3TGtGIXq/WqjehgGP2WRObw3MDuCZGpyh
5kNhggaQBLYTXDjkc1CLnYjou7U22X1tEXP0GKmQ5y4/8IMxtcF+MiltQSSaXtpEoHE0nMs7+IpN
ti+BPZpNUvWWGCqpOQG0Ff1m97Gu4ao+ddAotrJTSIpy06teQozEhujZMOdjt8LSkvzSWeI9umOy
wDOahCoQ7D4xiRnExw/iVzPPrGQTF5pRlxlMyS55SiMXzDm9cHgY5I7CyZ0QLTP95UL07NXlpPe5
F8qWek4uu0aDWtwDO+JG2e39SCuI/pRn42cNisN29bWh5bD0BBLNZQUP8tDl1Th23CPlFyxjoswC
/eF60gp/doN9xzUAaGCfAv3jtkHcHZp6LA1zL5I0VhDfHbDBoUz27kOM6Y2xqVJl0P/tPxaxNeeZ
Q4qylpxc1t6C5Y+qrrHdgY0x0iZ0cenWSDoHKgL2agvEBLtJQvZ3sQbiqQdI7g9kUw0Jgh4POWxd
CaMMKs4h5zXelrBp1K0B1OhrACqJDZqrchZu5ZQk5azXBhEkmEFdi5Pj8MPZKqmJu5mhsnqYxJR+
tA74itscJivsYqR+PhP2oXMRJzlyE7aJXUu8h1TL176swksKTi22Dj/YW53rYf/+Mnjtd1COF2sG
r4JLScGwwbmMHZkq+AlQ7TreX9qo3OJoT28ht8X1cCMYeVptZSNogN5HtMHWHm2Kj/ePIYOBsttW
QxSXWN78kRrIa7Hc1GMVVjZdbmui3cVhnsfuMJHWTrMWRwFh7oDJEObfWU7PFOgH1vxm2U+Eqayd
zRTDx2wS/PCsmstJWCAWr7fK4C/mNTfsKKRQQ7spADCKzrbA1uREv8q28ya+ItRjae40VANVzXPj
rgCbBlgu1sqH+py9DMWZVFyC48Ypaq+40HbNPorPuLC1iCvJXUgtlKWlVJdMtYRF/XRKVeYjA7xd
rRymsunv5mQhjIA7oV7dkrK6M38X9zepzxIM29xL/xbq/Gx6mWFUZbhXyVwpCEZisXf34fVOEWg/
cM1gqBK4SdNL7Bfnsk0zvFBdFCt672DtzBaW6HxJj+d0dGvgaIyTdPcjtbcON7bd870njq+fr+HT
zlN12OeBfu8pJFAQY+S46TDSp3HKEU0IPVAvYlfKMYVUxUMcwZTbkwdyWi7UQu5tBk8K2egi0zFx
KJbuwG7AoRb+GB19JC9d2xZK+q9DYGkbkbXOInsSvcQj/4ObtdrMn0V/ltNQGzNUYs1Eu2DsKMX+
E49qBXr+4CROvTF4/1m0Ak7zXFk6qTyEPryJuDKgGpGELP5xXe8L/8+toLhTtuX5b0ZACqWYn0MD
FrIu/az3T/1Ddzqc2jjAEydQMQ9R8S2Gt7vSiDVZOaBGRrtoxxlXXYV5eKy0ioTp+689QQPMQEbh
fiQeg6Xi5TluFi1XN1HxL2GI9ivougUm/q0RRMrTg4X4+iLl5fYW/yda2FrZKsf2s1+ANiuJ+OWp
qY8uxUS6L+ceABChIK3lYFqCvmU8DsTOOIYqo65j8Mqixgs5jX5kiBq6OqTxADMtIe6dy0DuY6tM
LpuiCEj/qUkjsASHweru3iRouOCfIN13nru9Gl+988YrXSZ8sHyH0dtGKq4Beh2dTKZy0ybsmZ+T
JvOhlJ7p+flzqLrhiCHArGySvVwN8/p1d+S+8vq2TJfZGgdRcOK3Z+MHoWIE2dZGyXHIP1OyRlkL
ymzRo1sIPJzqWMhLtW7U/ZJqS7i8o+xlqRjzsUW2+1e7Wit90zsSrfvBRFmkF8Qtn+hmTvvGsWfv
stjZin5KmxuVr+rALW4dvrhnAtmZPBrYEmnBxQfSBEvQoyEYu6QWqU+RGDF/O+7mCz10ZE3sRgIL
1EXQ3O0qKB851XVB0xCNDfM4hWynICZXiq79HDuHq70Ud1oyQQ4HbjjOLs2lC9RswJnEx+eX8RLz
Ru46NqgIYm8Dr0Zg8nFrOS41fzzKBNzng6t+XSZP0Q/X1sH/eAW0fPSDnhHIp+8T5wFc4qw115Cm
RaeYLJ+0zOGiqdxLUUXpnafuqbfZ9gCKOSfCOG7FjyDIxQM7dLFWUQYhVcr3GL9AKRSMbeLYYBhR
AdSCxKtbYP1VvGZbTfQEIuUucAK9c1ApMojgFY9jzYUJ5aH///kQdWaekiIXY8VSyXyOp/zjB7B5
t0T8H19Qy9dwkGGR10UMDmMOjPjZWxb3YRxr7drGL1aT611lORnASJHw6kW/JOoZvlMHdUDujg3U
9XUGiVCtsXULLHaaVCOH7E8jUUFEAF56Z0YPb8rP5Tc05bKbwRIQvL2Hx3e94NPxKaHcm5bJV9Bm
xOKh3m/OYkeSEl3ltFtOyf9rKMhNN8aDPPCRgw+kRJ8AR+ez8YIM3sokppe8vcs/4S2Df/0yAI5l
xQS2lZrOofE0Urefn720RKRniOm43vTQKxwSnqyvKBrKvd2WYUOvG8rWyHWUAMNtKOVxScarXqmO
oqMrn2BsamffvLLbxlLFZU5xPktZmmXubQz6+01DzJuy6FxwRwdNS5dKvV+2qFAna0F1I68GZUWf
GUc22RjZZZ2Mr+IQm8e/l3fY0Fqc9iNBAExh1A2nE1+fqXPYC8S6FTDQttcqDOH8f0Ln1penNpUB
ZL6uTASI+AJpS/TuIw+gi6c4kn8kMj0urJ95BFlDkFXSEggi/eORJFUrO1wgVKo5AKPxoEGajbbO
glqROdOcasWn+QlRNdq4d5sRB509inCgtoQ9oQ41pYTp8mzPgpDvXgwsihpo+Ei4eC12QFdPuUq8
6yRQSOOiTaxuZ112Y4Pe7fa6aCM4UIsTAWORgsXXvy6SAdujbGEt74KFBEbBwXE7RtS8CHs1dVPM
1JyOyECU9IwVv5C705pyWZ3Nj0fQXr5TWrQXGS9nFdhJnx0/DVbqn+8qsPYc8v4Dt/WoQcbcZI5X
rR6nf/SR2LceycnK3y1kEOf8GM88lemtNxbnDmoR3So8+V48BK6gQ8r0sOHMOLIFcof9oYdI49N9
60N7f8+mbwx4DMuaY3LRv7UWdpcqqPjuSpvqNv+nmdN5GiFKCJvUYhSJuoth393O+637eFYvYgJR
20TUUW37zlVcywnhFh2y10M9Jc94IWUFkKwn3OhJaRs1cS5pnz0clUkM9Nw78P335Pxvc2hcoogE
vGU1b3G0FG2dNSliSUspVSUMU+NG4QSSOwMlNx8l2UZg4Uv8l1++2oUKboX+b98NgvfSMQxbvvsR
HXNi8PuToj5qTpODqEDql8rgkyDlnIV2Kfpq5rVy3SWK9vEygAz+ZviHea9TU0XA1Uyf0Y2wa4ps
P7Y/QDMMPNtbfYp4AQ5to2QGv8Zbj860FE8Z/jIREgeLSdKH4k0eXeSeGjHyi4q644WIMSeh4IQl
NI6UtpIsGbPlYD6DI3Ny78YP+N8TT3pFwtXYi41vINkgUKfXREjmOrf7Rh8IKynGlOby1s7ardB9
oPR/9MShxLHgIiK8noBkV3hEnUnuNrfmlYMDowHmP86KCyZZGVoLZqBImb6+0Xkb4Gse5+YKUC0r
ynoRiP2WFjmiZWWZcrWIy/xo+HkqpQUNU1ZTL9Z+rFChHFswu476Rwu9uVOaPV8RHxVwVM1WGwbD
AO+YSepiCyofob9E/cmB1y5HnZaQcSeT6HnOWgOFK12VnCSWwJHHai4rK5NaABUxms9igZA6WK4K
MAQn0SNn3jAEpRPrZyO6uLdFz4KNZjkMjguOL0gyGTpPppSTckJ7lL6gTo/wv08LrXMvY+kLX31c
tkjpAQgnxgTpsU2xU7RZHM9Fu6qm++p68KT7sefM4KQnI5+AaIJO4FwdVeqLvR8lcUISvod+tSQr
QyZrLzJfPKTYo1AD8647hkV2Je+ol+VYhdeZEMHsIuKG9tRSipxz86fA8KRa1gm+G82z7NqUq+64
iOFgbwarR9e9hZoBtif9A8TUQLnlhusST98rp4JQ2zuYFzraO6jB4KZkbZ7iD9fijNYszLjnJf6y
V7QVUPd9cXixC8Js042Ac6GZZ67di6SE6Wvmgfb/IdCEDSaLIpXGI0O7PyTh49ctJL44oepIJe31
UfZxjJcdte1/pxqdxcfg3f2iQI2l/GPd0XGIV72pgdPVlTvvRfy8d0G7pXIY4wNn8620m+RgNK4Q
yQekVIkZlTSkK1QBDQAaJny7m7lqI0n1D+sY9rvF9/Tt0lpzMKNg9JioFiUKPFYt3feilxX8LDdY
ZbANEGc9IiSgLbz6/rPZkTkp/DewHjDObQ9xDP6nlGPaAwVbU5Dpn0rkBb0Lkg95qLhNgt+3gzfq
YthYDK58iHwAH0gcmJbbwucNqofvcXkHIgpEDN1uK/t7JiKAsszErIkYaOySg4f4OOWoi/mn0ZOx
IeZdPY8QF8hmiqdkOS/0vPWAgct4F3OM+80aSDNqNUCbS6j3GY/Abo7LPDcLoswn/bg9rj+LGml2
j1llxS7qbUwCa8NpBoWNdZehGTfCJrpqLFhfjJXcknrZPOVncEInX7Gq7VCtAiIJwvQNWsxxaWAY
XxCe2MT6CXIE2vMmmVSfm7B2WNuNpN+s2wk9zCWtEJ35hLm3k/PS4h4Kq65Cc+HUlrq/8C8XELL4
JcxwiA/bYYjLww9OuaSfXzl26O61/4sUGNbqjVc5aIMNfkqfEvCPhWVRYIn9WObls65e0WtvttDa
BQCQSm1GO5v25wq28sFiRyAf6sGtt0QNwRAsrC+rmLJgeJHaCAGFoLhwAHlqs1P/bihcp9Oo9/Dh
Jhm31h4xmdxaypiML3fvqLh2wGaYPvueJO9qgK/YIXdH/jzxT4j2mIrKQYrTD0QKh/z5EfN0UOXY
8zXOmYZ3S11PRVzH/vJjlR8awzQG3PVQl8fkuNrSDEastm0spt/eRTSe6hMyokOgper9XTps6JO/
dcKZUTRPjvfNy2jQw2NvaMzeLRcJ/1Odj+fEhaS/b39W+48vSiHlQgGMWJDyKL1MBt+zlN/8lAjD
TLQok7ok3yf5hKSKAVABm3fAf+d2Wta/BT2lLDunb3r7D0y2/ZwPI/7rOoeF3Bl7Ealf5mmP6Kkf
X972DNUWI/+b7QqouH0S034FshJbJSxkPF2i7Fbn9lBo+rFv45aPXUiRVQocv2uY4VYNiWZ9kMEM
i8FzupyAaaoCyVeU1SsqBZaqBWbqdrF3p1j6bICWiii7XipH5EFegDbe3UZCf0Ck8+ATwq7A4WQI
z8akfPJQAByD/nQSkYApp9mnxP7pcxsGb3/l+S7GQzJrQ4YaK/1gBtUIDrbkkvRSF9kg84v1vGqW
BHmxTHy5MYCNs+t1TPygtWTfVIgKtsHwInOaXVNgKSJo2ESe0EJy/16BAr/99U0R9friNkLDed7G
Q4LgTaxdwxKIfL3Yh0t4CyXRJhAbutZhbovY3BJgqetVDK72QXOTX72EBCE4+riiUX9IJYX98p/t
8T8GDgKJ2aoGR2WkWNRL6Ay6ghMea7PT8oymVlBrLklD3V7vFjMFbSU1UfC1ouZvqchHBdrRqAHL
ISOosfRdF8Joj1pwBd4xP1i2V7x4GNkQYs789k2Tsorg6+t6t9cmEPO1sb4Ve604PBlhKXfiE6ty
Sk+/wpWhgQKzcmTTeYq4ITHhtfC8Tlv4s5JtbHpl98EkHo0HaP99myTAj9VzuJ6osXKNa3vfT+bO
1atyh+F5gpmUvPztRi9KVPkN5N2AKyBWa+bBstLG/gfy8OIob1kTNiwhJa+A5UhQDn5N++ja9Qa4
W8c2j9UwxvrpAiTXtEom+/pUiIg45Ong+6THCTUXQE2u0lwiZE7eAokGAk9LXM6NkPQJxY0U0qMb
pVTg+yniPEp8rY7sxCcsC8QXxllVvwUu9JACuQtEWGYfYHVWRvk7aiKCsQbg0ewr06mmWBURmWBC
1Xz7X84218aN3zCV6QUeVGagnjBtnPTetzilJujLeydMwOJQPtlXGwlAFcg78o2r/70JxUE3/rP/
Qq50sP+1Kk0U07XSEOKZN2Xv+cT8i+IQDIowSgBlDxGHzCcCMzT7R7rHUk7YY7U5An1Xs1GCJbyO
afIS+SxrpCSlNCsG7kOxGX1KF1FTPNJnYAhn+NRdykUZmWYTdgtroBtm5ZE23RAlr4NMdAM9zOdI
lk1R+AyDWYuxS5XVJ+j74ccGibxQj3HGWnZVKM+1hkdOxnmywMlE/f11fe42GjyVPLhoB/z3z2QU
xT5U6cxpQYPDyJ/bhASQLcyXoQSfPEN35eXrkNLB9tbzsMJY/vR85aLX9UB4f6jkT59SHfbEjn/r
JYMk5uRCWbueEJ8oeUftsxP4kxTzUgNPj4XU/6jAZRjBl7NrZAIW9j6udMeycN3D27NqMSOMd3Cr
iy7HNfzYwZV4agr4M+nEtgwOHuyq4O7KQoAIypUF2Um2aN5dq2A168qR4EnKpnOURBhHg/EOP5K2
j2HJqptGp56c7AcVinfwVVLjIff+5vACLOnBcVoMpGJyTBT7lK+WNSkhCKD+SmK1lY1K7Cm2YU8V
Z/J+lExjm33MoBT+p3HfpYH2y6L01GEBWazUmjI9+4Syhc/i5E9QtZtrs8eETvSTfSvyxWqfJCaW
6ohXaiYyDOBu6us+/Apttg0wgQzDWSPbZ3bV+3AMD5AY/U/EIfqU8p6zIDMxc5iUhK8VTpkFbbBj
vAF3dMiUoAyXzq3D11dpbxFXxlDsyelXV5uHyhiWNd3ePcjxVg6WKk+Y1LYHxzy6/CKubeNWH9Tn
3cqXplX34QHKy2RD+ThY6PdNbpEC9KhgV/Qb5TVbr0pfGvDUYLe9b1+X2NXYCJL3XmrouiDZs3mu
9eODBSrH6r2GxsYLKzA2iBsKzPOLF6ubLk4tJqRrWclc7jSBodnx0GNa2Hi1/YzfgGu+Rme90cgN
UC5KyiQGVHXR1JLG95dk7SjJNsMCQgILYQCf7g0ubg+eahQ09YEp4FScQt2v5ViLM1UhjALqREfw
WyWkiLFzFvOIcXzKN40PsmKNXGelWUghyb2Y1gJOz459w3qsxBmDstQV8dKPDeC3pg5RnWcp3z2h
sf7tRghbqTHQUr9mOeIc7Ue2rpXWVBBUgaeiG9lX2h8HJAheP0nrz6NKbmEjVUd1C5ZW4uJncW6Y
9ZVnovgj4Fe+RDOtV9dEmKARaxY8BW8+Lw6PhOjRIOj4dCaIP6I6AMDROEamz3PZrUb8QvCwF83/
PYZcq2yYFDPPmeqTYi+UZRDEVT3o/z3GTy5A5URvjC5QgE5begq5k48W2uzavWmnVC4MPcvKQz5y
vBZH6nmnQi6qjPfMlZhnDDGOJ7Yd2eWml2Sd+clZ5LNWFnyYjENKR5qVNhCnUxfkrskirDKAWAJP
UiRZZBHyj35H6SGj5aGGrs+gF5vfzL4v6K0ji38X5kkGNM6/jOeUFPGVQhhNJzYNkSymvquXVGQe
apkxKGjtpunE2RLbSmQr9PfeOMcqHhxU122WVLC/dMnCbFMWSE7mA6iIaOXCcvx3E5JNDYpO2EYN
9YMFLbvwXCQJqIzLWEtxtz7kdx1YVe8jLPdY602u019Pt5+VmccL9eHRian9R0vdr/adV59YlAlC
TIEdU/C9ii2oXHVjPMo2Eqn33hpPhmxRrY6gcRj5bOkgdck8Fm8LvVnNuEDVH/2hSTvYKk+MLGCH
3sP7UhxJ8sNg9HTapdiqihImWaKBB3k6p0rzAl/KBVoAldlVuII6tmaObIScepyZLvOIfme9K3+e
zwaZYPhdxK39k0cvP16cL6tjB3FRQFv/ekHGjmMFKw1OjIuBR9R3Oho+FvJ70t3VYwt7P2FRz4mT
xi9r7XWb+7DCnnEN+nMH6dpg/L7KFWdLmYeYQEd4VltKXBIDGtCwGnqXWjaLbgM3L6m7yDC5qULc
bOjfbWc7cvwPAhVEiAzjyUq+bzoaXo6DtAq9bCbW3Dh3yDqffzN8UDMn637q6BritIJvFHnQDFUc
W+pIYtT+iehhevajSCRdjwh7fdFGE4fh2m/ZDaAPoY5RjqNIVh90hWPT8cWcikAn+60CXyl/wN1H
D+NzScvt3K1DwC7MEFwpu+Lc6PVes6Wiq5k0gwJEfvDGZhnPSeHjEH88pgwTb++HzVKHsTDTll0d
lSX44Sy1Lgi7QDqSBgjUrVvWjmdV/BZ9BDMGiynyeTZ49jpaIqoXgu05vScr87J9+9TVl2QauWjk
QR9dgi2AqCX9TlUvzwkOm4gfJqo7mLi09VXulbNKjd6vJ5r6jUAodBZoMSrR1rWPzgVVcxmBFhN9
WD4JAbp7kCjoPvEigxXglaULs5WN5vk7uQURWMEFtZPNwOv7da+aCYp0lb/kon9rj62sQpsG5OoF
DGf3NM/iIULBPn+4xugBF7DwtAizFhLIk3PImuZJNcYvwQejdDu0cjcm2tvam4eDOuw82v1KMl/H
5OUxECYJrAN6q1/zh94Z2BPw5RyluX4zYg00tj3LSj1eQwkgRluHsypIrEptfn5CLXZ+q2ALhbg/
lSdJy6TCtNHp76GG31bulTpDx95R4rqMQwERCB0bO2sDMjUeFJD6+FrQPds2/JYEWiITf5DhHf9L
ng1poM+Ec4ia1Nkj04xRXBsJ591hIdyQZJPj7ztUqPlU5pGLHmA+wm/pQP79hqXWOiEsgSdktvYN
C84XT6RKtqECCQcxtd5JRBbVbBr1XvqDgCBC+whlnnRb3hKcqivBtIzFDWQqAqdoXAyJC0NeoBL1
w9tdg1Nq/kzgEr2qrC542/+3AVy8J/17TdhKhbi1yYuYqGfQtxdNR77ANtnS+a3rjmv85bh/k6ka
6gMmSXrdbFXLCDh3sO5AnI/Nr7oHC0TvTOdo6EyYDqZ9KBX3oXO+65rXTC7zP+Fts0w9vBhvZ/sX
WFt0HSxhtz5/izaioyDXDPtW69ZrfYut4HEOXHxi0dR8KN9FUttCUB3yN22vDPOEeJSgI9hxaQxg
tyGuKDYGz9SpXNLA5uLHnrS2iqv3JoLuTldBoDFwriCK0Na++7XLkyNB5CE36S2OXp2cN18JuWtC
3eLVd2bCsJGDBRTPlhkdua2Vquv0MqsAiGWeuQle++k3Lfeu+428f6A1BP+zv3rnZ7C9B0tqji2j
mPYX5wOoxheOcWwRemDRcgRAwYEUEyN6pqUd49Ymoc/cfUbU/EhZ7l0KsPwAFCiZ53NAdx8UoZsO
yGxHcRx4ajVUNX8LSVXO09+599FmlNO7Y1pOa89G4YbeT86KO+40zmryKXHL5lZABng5UztTn42m
YNDN4bl4RpSI9aR0SqrmJjqvPgqtdP59OiKGwHk+8cDGYJbuGIxrihnS1Lxlhm3b9JQfhQ6bm0RG
XKf25vz3/6Ds+Qcc9y6z5KKdgVvpiSRzEjKrWA+gxAGzC0x/tizboOBxMmZbLfjMgaYKSrjSFaOX
2UoyA8g90o3m9h61gRupy8ULIVMgBjLv++1GwdsxZSYPhN+OxA6yYSvhRjq2/KhgSpqtB/XfCDYB
BGkCErMLFDCaDMtt3S4BrLzG68uX6SjtqFau9NH7/4y1ITCpVCikFWEggIvn+EFe1ifgK/jlDVq7
Bql9gSIUIC1onuZLeI4fD3ZHFyRQwPxCsNpdMyfbQ0XmnChZnCNP2ZodZi7RXF/Kc331XULRHBG7
fTHbdEiMXPtmf9QZLL4M0aTBAW5tzox4Jg6ZhO4NNtKAbje1wNBs/Ai5VfMT1typrSYI2QoRQmCh
Sa/AAf5Vhtar7kfvdqzuawxCSfehWxaO7768MjtXwGhCeA8ahhkVr1o7My2Cwglciwb83QNSAGJ+
Pki7Tx0U7tn/xrcpATdjlrCxRXyoKIaFML+9Nr3rCM0FmqfGrbHmNb2fQ0fwvpvp5LZThVerQnyN
+9kKp2NV29jbiPIAQCQ/I/n85jN1vnTKlsQ7lwfyRxdW1NkXzQKL67qvBUFS2bS85I80W9KB6l32
2I3nYOVwh8v5zXonUXNWd6yYjvOxiKk61acXWEISM9z+o2YMTX7DSVLdUec/YN26NHPGL8Gq/8yd
WN6GHKvlkJBG1W1dVunMosEOuBIzNbQxlpPhUF6Dj3NieC599N2PWH1TBtIMRmPEBvlWuTwdvlIB
GgXZY+IWYwt8j9W1tQUnIJ1l7K2L77Ir4+KnHJ88x9xPvWHVjRYtrFXwN9hq3njXxUH1dnziAgJl
6gTps7rRqMuBAnGc9MtJqYstxEeoUP9TrAyfa70n/MPvHw24TRKl/g+kjjBzQTOk1/+sIt/M2vs3
DIkgjXv0Cr+P5N1mi47NI5bVsaXHkgI5eJOwkH54Brscoet1XPFzAVJn3AreNWoV+OE1FaOni7X8
cnAT91c3kf98+TeJH2kyL9CG53ZGKSfy1kYJH3LyZjx3HfMk7JxvPq4o5UYFm0fjoGHAWz9T9dqo
JfaBd4XuzT3lnC80/xyIl6yAgOpSe1QpthNswBZm0WdAJCNcF7ZgaBziIweeMFMhEc+T9yJmQWb8
WELbInLew5lPtBHCzwIVSoW9irCQ2QUdVDcEop4eXFjWZhb+FevjvFtERfkm15Ap9v/y5/1BRF+0
be0TrS+vwYkD2psuZ0iDRsmxnlnpLsTJBGvhPEJO++V8ai7Y+mdjo76Mr8tL3SD2aL2DuHjyL9yR
nf+wWb9hnCOmclRdZBcBtJ1MpQI+ast9SrwlrVQ/yn7IIcE0S6BKZ3vtrDQ3LD54sOZysXZxbeL5
OVfVJeyUcpUbDI0vgfhl6CwqFjL89X31SzoFfAl4oWszskJol0EMv38+hNUWAbMbECJ8eEjuOQX5
AB2Je1qz50UEv/V5omu98V9z/ExlULbycELPo88J9MrPJPgSUtmCt6mzdM4UG5URFxyfzaw/3V50
SMq8FCS9ZPhdlkaaCCO3JriKotuy9k/m7gT6ElfAB20oZHgMKP1cEtwLFFWOTIZAEta0lF7Mf0ZV
lXuKKuSWnyW+QEzqWeaKaGqm20C07cPCw8KMeO1LFJGUJ9d5MSP1qLIJxWSdii8P0XMiLWVrMiEt
7nvqN8JqQ11ba/edBAt8WFUTEI6g7YJQfuV0+2cfBQ8pMTGwhwHMcfZtGQXKnLDNwi5aT+gxBDRr
f6m8e+j5eZ4Ep+PpYIoyMCDknMDRif2+zXlPB/9GT1+KqbMOBF8GQGISQyiEVgCrJyL7vwqBEqdS
eCEPM7xP6sDa87n0nAdHC7Abh/bPbAx36sojBuKvmgM76C8E9rYnW8oygIIGoy5SfLx8w/ajYNbc
hmffq3dh4qSTO6Sp1o1VUOoIpNeHtW17Kx5Lb8XtxZD+4HJi1J7DKj2YBAb0MfS/AKvSCpgXDSiw
FRxV8pYW8EowqZbl46TP+9d1bMU5ap67FIovljqC8eLGyKjXmiLVJkDMNmPzrHhkA3awiOezeUM1
wdVQ8GAOkmNqzmZbIz8FPQkV5XRNt0icWSOQxtaeXNel5lZJmr4NyZ0aCMdohjFH1xAAbuhebFRJ
SN+S3Ajtd5LnUdissKSqi77I0OBocxLjWUsFkUabwIFojoty9x/u22mZnlZMCfZvfBSF86Y2HTSW
NtuiHdNNvih7J9HmYfp3xCK4xHxRADPJwUWjTIY/Qyb9A0bYKWBEQBUURxvoDgpmSs4jBqgRrUwv
ISAn5C/oQtQdjJ9PbZ7pjAZqoGBL9LUj4P2RTaCzlhNeLEJlOxLxV61JM7NBgeuv7PBvNEzyBPyG
SdrvoX/zfj47tldg/lcGfiPQ3h3n2yUwdxULR3MAvRfBf/8SJWr7NW5R5KJLFdWnFhSGwD+PTT8f
Bx2ACAczbpG2/YcXyZlk/FeHyBtbWUw9fcgS4vMxDKr1p+j3roe5cpbwQoAdlO5v89uT05LTuqfX
1Otp2PrjUD3v2idUz9tlP3argrBCLXn7CUnJB91r7nfMV4HdTJePqfs4UWEIoF00lfHhAl+AU2sZ
33ZSZqxpwF8viydOO4RhB/UGiVLws4c6fR8/SJU/zWAg93soy6xRRzWSiMV2L4+9eEYAVNtYxi0j
PhGZWuQzmt9NmkwZY5N37cTU4wBr723V07ksXRoNb6Vnv4BHWB+KJrTZkTItW11BnBwLcsmFWM+M
lu4O9Gto/qWmSw/Q/NBd7TYoCeE9HoFyq32lPp/BAP52brdlroHNHRvLJMnqaPH+F9Rq8qpBLUF5
a/5pmsnFhN9EE4xqkKWqvJ/8i/uscme/GJkkGKlTCS7UNpZrroDcKYVoNg7eUYZ6Y3zt3TNZmXoi
1rNDx2F/+mkOG2xtBJuB3yUfNbMEnWlLhBeeE59svDbxFSLiFf6+hWuPCMBUSH8X1ZHrAfGVSME3
M1eywMIJokKAvljXfaJMavXjQOy4Pd6gWvFtQ027/CIjIGFa7zrR9zxs0AnJMWDIhZgpS6TveFfP
wYrOd0HxY1E8N5rMLSAXMUhdC4se37nelbrj9yNrsyQxWMQKH1hRsT8/yVKWWIqYjerfY9pm+exi
1JyKWDquwUP+CjMDJiq4etQc/vHi5UcDyCKX3/cCzHk0OBhrMb6fgLqpICEXC0sC9ubUp2o9b0Yv
95I69kn/YwpNJhf5APElCxpc8AD/v8IBDWN3S6qibc2wdDjpr7PFbpbNTvv/0oLCf/6oxWSRR8h7
mJAfW3gyiJpoTcnNcn08EWgYVYI0qjNwQJmXjNzV5I8OwWIepLu+QnRR8cENuQADkgYHj+LK9Rxf
lmXpMgOTn4gYXo2axMetfsOyma9K7pSg0DLOwfnBZQrMJz/G/gcWi8rHsLk1k+X+h/jtgA661Vum
6YIvQwszBfwp1ro4ZL2zA+MEqzXKInytIE77SE4GJ08rcRGW4PmsKEXYLHm9eExvBdmmwHjTHJux
b3it9mB2M1yO6+Gv3lVZMGLkUyF781IGV6VbXou3VCi9DGSVw4LJsrQIi8tU56TP5t7HNn/BCumF
sswsTLsm32nI/L+5FF7ro0fhM51vNWrbcBCzedm+O0A3k3yDHyaIHNPqJjQOy/8SazZyrRi3urM6
qnASzGANdExxDhNAA5Xf8amhw7CP7uTfr0Um0iAv4yglQSPajYBd82NHDuWYC9qiiCsgO10tdh1h
+0qlYAapePuMSISSVuh1jMmX/gw3emmjmzo+9UbgZV2+J/oftsnU22ZfNC0QoX1V3uzOU0UeuWe0
6WNgBBu4ATFgpydwOU+PhmlzVVWOY4y9TJWh7oVrLTj6yYBnA9QrUyoA7sXiP4xzjfDry8v5ESNc
KngikVt8dGbRKi3rC9WB77oNX4LJo9DeYsnKRSYbII9u+gJD3Vx6tdNALVyYP47FGJvlT/2WvGtl
xGyCM6F4HCnQ8kPw0e7mHNIOqFc19Q3Ew5YSIV+UyuXHAJq9PD6Xd/rkFeDuZWtM7aRyHMEIcmFy
z9fK2HyQD0QkOLHJAf/crl+Mc/J0d/RvJMnU09LEUGRlVJpav9/22fsfp/RMhUP9qNtm596C0aD9
ekzYfxnqKbRjzs9/bIF5uP7Rt05n+nVu8dsRhotYv0lKBfed0GJ+NfARe13kbqnip/GAac4FDd1/
xT8p7Vr6lsYo1Yjma/Fre+ah7S83v2BqrIlyQZNWNwUWKLJP57WfLLzTU8dzuolxAVc2/gN+YNVP
KzlcTFWxr6+1nw1ICOXMg0ZiCysKPXBIN4tzyrYwwuguM4TthC7EmRJmRyFPX9HgKnbUGTbeJzlH
2I/93fvFrsULMm/AWLl4wRjCJMrY27ZxKdexpBVAXnTYw9ERWzMKC/w/tiRny4Xyth3SmR0X5RjP
WvEi/Xfg8KRkRRScEg3bibL6tRpY2IwNVLHTaME/RwjA7Fo5Kc9H1vVgTdn1aED5/TI9v2bZltuA
bPilOeopA/3+6i1SZ0wiCgbKajygdQ4Givnm1FlVHCi5S4dNmQbv03xVluqUtfFXGKHwwbQswNSO
tuNM0RAX0Z0Sv2Fke4O2k1mXEX1Yj9vseJNRFmvOQNtpOM0pHLLwLKIxx8sueetbkR/R4L7F+Jb+
oOa3OGU/9ZanAbjRbFhwBCgApYJoHw/npIEvlCw3vgpYCd+eFFsTbJUXRYqKcCGnu8FdMm2LV7o5
gTSNyHm+YjE6ka4vSGpL7pSoHfn8PqzqcmzY3Tj6RaKw5V0gj1ps9z3OwQjVxau6X7Qp0e9dePe4
61yqw/1t21cVYimHh3WKYic8JfWgH8pK/w1VzN7PNIHNsVzakyFuj2NK00EyQQt3MnrvtEd1PRAD
LojHpIQSZhbVh8EKH7wwZighZaPSAXA9c9aeM9CdFx9kxRXGPw2WYhCUCvHRgbQ65PJXZZFi+nCL
/2JrNiKvfCD6J8bFp+PVH5ezmCLeOKEk2mFCq0yNgq9lhVy5xeOl0P2L/FLqRP3975kxpHaPGLtH
qEniy5A9efjyemyJqpYjPotGuo97IZgiaquRKnpafu/q/UvJcT4OR19yhD1LoCVgXqAhtKxYLbpv
eAVFja64FFjWQznU20AYp3OnlE/KGXzint71pt44kN3G/Xvco6EXQMYFaQBS1VoVqUW6Kx0pq42q
2dJouJTdXIGJblHQDfb2i5TrFjXoi2V5KD/dMcTIz6qakH3S9Q3uQCONlsjJej6P45QOVs++vBrq
N5Aq2VhuPYPpy/N5W5t4vMwhxNcqw8FW7nrMeggbt4He1t+/35WV/RonN5TFimQ4OBv8ioyB0MpO
zk/O/gNODBVzUe28VdkbC8z/LOv/vLhte2xJFz/kLsY5/qI/oMO0Aig2A8FyN8a3CAx9XWxhDVwB
1eMuAgaHBCMgeW5g6By6Qc5t0ZPr230X4y/lqnm2U23fkW5tGQei3InhXe+XGbo6xPBHAMLRHWtc
rrjI5kldylEkd1IVcxtiEpOPyxWVFsNUBfn7ze2TYx+5zAPLgeoziqxwZ7WnXJa+9vVajgmus+GM
iG1/PRRUbOr3BerDaOOyGg5gIolrQNRJFut/qawLS2FOEyS1RDepUuzwgoSA+XUZUPZogsaQRIIr
U7mqokEglqxwl9thLfqYUhOc/FD3zqDfU9EEM737XQ3OQIy0e2B4j7mUThLzbfYxLs1NuInm3zw0
kP6dFP6lSeVEA13sUnuBMhb0CHDZsjGRtPoPoJdiKLDOxBxmtmpcauRlvIUQAkXy1rpGTkGKQDeM
Ned2tZJgTJcvuo3TyDEE392+CVMzvoX5APPB+NOz9yj/FyVFrTQSP12/EXLZfwT7oMtJceSB2MgB
TQie7cbzUSSsoGIxC3iiMZc5jkkLvXNTkOJWZTh33Jh3fxrmJ2Y66rQmA5+Pe42mJa8xqesnq1lP
Tx+TLlqwCFmR6LCu6/q7/sPsug/lBgU/Ia3lgS/XgFAGXKsniYpACIjP/gat8Kp+IiLh5L9JVjSH
l6CBrok1IXT5H6pskAzrvn8UNFYSt4iHMYQtSRVzblVvgJtF+PyETGGQcjQKQpnewzxOI5VNZAhd
hmQ9RyhX4mLqLgaSfQOBRMZeKoAfLptQS6HIvSyH5XlaM+sqWNBdeZVk7OPgxR+wTrB0cCZKYTts
VarvU2h2bXTDjN0joGNG+yDl2UBeIUA3Ms/1nRiC5xsByObtMVBrvh+DBVpXuMpkyXqxg5L+LgnD
+rnw3Q1HMPAjphvj06CmxFU9o0CwEXyZQSFGcg6cmr/CtG30DS9e0kdelpF+ai7oD1UDJAca0Jcy
vxLXkkSB3rdafnd5XnJ4zss1oo/93nLe5Tv7Iy3wnmn6Hxi38jLDDePAJK0oqy9ec+YBg7trfKms
wXYk2IvLPJFzmT3Sxv3sUTGpCCVM/Z6176iR7XN+8UrXviHuIQTAllAaUCjYGrwcFkDD69dgw4Qm
m/22X5BzNzuOre1eM9/Q+fdmOMF7TTIUBf6+FwbdXaa2nGEV4lgjjBU0bUGIZ3dgB8uHAERia3Hr
qwuaSVa+PZ0qFl648NATloP1rgHiMpp88b6/JEJ923Sc+dTphOnbV/nVWqiN2FoNrqqD1iuTdhEy
rDg3Z6+YURT6yCqM3tuQxH+m/0hM+OaDCfmNBdDhBy947OKSDDUCaYfTKHgjm+iMQLijbYZzRD5L
YIJckatEJ/W7TekDhiNxfu672ftfp+/IaWSydGkYQb9Yc7KtyD0UgD6KvnsXRs/b79cI5Fzx/I0E
ndtoB45/2V4e608zZ7JOGQheC67mfJhhlH2BcV3bEcsH3L5qIQhUaMCkU9pD7mVJ0mwYYYsRQgPT
RSdh8woYzG80r3v/Uqq6cTvUbc8/A8gMjx5EgO1iY8Nl2AKk32UVseiHUFCuVeZz2c8IGzIaXPPt
B+HAhcyBj3cy2sh+q171UG7cgOovRyEsc6fiDdRA4tgRIS45KFgjXOhLzpehWjxCt79rlFcL06VJ
Cca8zc1HS2ZXzNKH21KpCQEng1JLaerUuU/qWQIix41AshbGbHwdpmtwefxxb/4Mfxu5ln31JbkC
Ifqb4oNh1ZYtzc0MhAxSwag0xjo+4zPvTceXrpc47yeuIwztnNq5P70VddiThjigERXh4l0o5WPH
6NsBOzk7UwzQGw993T8IpfaWzrOlQcoB2ZGuzaAPycKEIDahG3XkaN6TCk19JjQ0VhyzjzN3s08i
ujznT3VdL3oRqzKbxfKs0o2N1wcbHItVZueW5pGWGLE5ssENT0eEITg9qZ9R3ygS0fVv0dEYyhqb
uAhq8blb6pf3UNQNcv14nr065g3RC5NqcFpgJJul1oyc8HQ1Dw5PnzEd/1wdEUM4ibYl9GhjYDsE
GdF63PIVxFgdlYuJQ2TbvmRAYfTFXh8npnZuy8/8eaOjYDrm5JsP+E92AbwmC69l+DuD5MAb/On+
STGTM31qxYeI2shYQ54l6vc0lexuNhslXIrZ/gav8kTYoluWJq5RsnPmp0k2grJqtNNUefa4aSDI
s0njG3nOUQWR+N3aa2F9PjCVgRAs8zOODkG5g0BU3K07tWAmxA3ZX8dQBY28V5UEUh2n6W0txD2P
2mXHt5Wy7Yj1PokdieVroVaWpGpHRwct1EVS3Yol/K8CV8iZhx8LQovuUUJWG/Xa6w1/ORBOSZ5K
GLaXfsa5cZ4nhOZCOzE8uE9R+c3b0qaApvx+ThFxchwLxVwRUSZ/FakKVL0UlVCCFDthfoXIAoAw
nEbXE+FYP+9yiPUoV0cbev1ocQ3vXj7N+9ACTW3IVl7oWF1EsrQygVuTi0/qz/I3dY9/ok1DJssz
MicSnPqUCN4fE5eFIV/KEod8MOfYUApaRJZgIl8DtNGVJgHP5LbUmUSejDFlAr317yQljUL5Eqla
IErmQQdlU4/kq1G7/BByPFa0zYc0akpNGiQ7h8Pr9Z7BIwEJPcKs91gEvCm51hfizLrqGsN6m7PJ
/PbkIZINYXDrvlZjehkL5oJPx0Av/oFFdfUcSYgFwfnn+qUJDYeYEoXXw60BHTELvHzq2kESR3j9
GvrleRHY8V3LhH4Ybho5g9N4QQUib9yvpA/W1iVwH53x03gXvskNREvtTFSXyL+Crc89IRB3/WYL
F+o6DCOEyLlzw9Q8ZW3o45pWdgwA2iHiWLcRbb1jULXv/dZcSPmJfX3DblqfAWa6CH2ymM0pRn0Y
hL9yUGZ1vdFRm+elGiJnlmTaysuEZNu926bl399Q3S4wN3j9UkbWKepFUl/Gvhf8jQ7UL/JQyzUX
Qx8lBYT2qjwaSsSpsVhc9r+Obsg4KcIAUp7Vhe3Iofq8RKjTD+3q7Fu+m6w58M4yvrIfuaSrxdOK
1yw1jCfcMQyoNcVRfswx32BGqUXC47UgVj+/xpVkTzkeg1sdBcWmegG0JLgcrz+ensUXqu7kezyQ
FSbce/sDorWwCcIAubPqT08Of3v4Xo/k4Uo3FWRkZWubEyTBoZi/zcIUQx2iYQP7wj97axmpN+8A
Do5V0ErvM+jEMFserqpZhSiEOYdaiROgagP63eACSlXJnG3zyybohlM+vs1DAfd5IEUso0fYU+6Q
qG8od6BC95f9WWXHbcTg09BcxePwhwsf+j5tiEIjtp6zQ21QupgCp6nmLVk+yLYFXSv0ZKvhSDLY
+AiikUx8ieC9U8xBPTBGvfhD+w8O0qEcHyAebGcTysLzBYcBb/07ekfsPzNWJhQ12VkiOC8SkPip
W7SgbHJ0bOYMdJmco4amLE1uJN+yJY7winSVpIRmD6Hq1fMS1DtJOIXr2qg22Zz/EP5/6qtSJupA
URkDf4UFqJCwLszp7NnH6JqtikUCCs4VJqfmouHBIudBJzahjlOODlsHsQk3h46J40NgnpWHn7/2
JHIwiQt3TW1Xd0N1MB2+GWiKhtWkSr7+zvLLCS+x4tBN3HIJajoUW8D4GU4fwIwJdvYEKnG80i6Q
kzWzYKF49ZuBXz6hdYbAp0KJwJ+IUY/3OmF5WVWN4fdOYS2Tf7uHLVQhGgs7gYG8KaqQrdTc0Z0w
irsrjEJ6eDshRisOXwbs8G3/vzzGXR5xqnY+0KnFQ+fIUqJok5s+SWd/Qj7mbmNz/OAziS1Q7iCR
28AQ5Ka1DVx75QFbMz43WwpU4LlFTFh6iOfYb/91WIbAD5zn+j565QGS9q3x7z8sSrgBz1AYgL5W
dKZd5S0owkKIWK4eRugPyIEcFwOTD5S8nEoEVM/V2uf2fgYGWeW98fq9WgY4Llew2ATGi7FMz74P
8BaGOAQfu9HvvfabWcNB3ow5DztVxHkUq/0iMqVt9dYLG7KHwjXs9Uw9wreupAEQQpQ01IV9ZYn9
7SzStW2vsobmAUzdZqmmFSzW9JepNKsbSlMM46kztt5Mj3EXDEnoxr3cir99ND07KpmKg7MvMITm
lYLcOdWB0CCfuY22iJT3OXTv7DKetO3EkmJGYBcUFB7/I1ySqa2Jf658iLBB1AunpQ9Fyx+B4OhT
Yrv9/kZQcvRuBR0WNkA/LKug/hoo+b8Q0nBlKDMHSlOrVqzEpM6PUPf7ki/7x/b6BqFqxdvIA1vr
wqc2+f/9F4NUaiscz9C+liRV3GRzYoMbjHYSeFsq6N/7sjTkcOxlCij7hH7ceIyP0JWxtz5sJv76
BZHkwGAqdyTO+ypeHitjgHNzeYOTTNhIdvjD/3dUY8nQ7pVlueDI88+gvS3+lh3fSXC3sHRWUF29
C2FNpSY94SOIo7iI3fOGnD3mE4d7GbpbYXnfieOGzdsn+XFBhe8xGgHBOQzFS19+LFU0yHN5tpUP
dpTCHqpdQ1FdGyl0WPSDwrvv55+WUsR1SOnx+iJSrGOhdkhP1hv4cXJZBTYr7hlKtM/AjFXXTJWF
5RtiqPeEy8VAm2uQ4nuqans/2wwhIm+If+ZJLNcHmsSKVquX2+pYqPCp1oKezD/GCOVidI4UWlFZ
x92Jj1edlnd+5MPmTMNxVkxMjvOjK4tcZRU5dUuUxvJkQg3pdNeAwBd9lzsSrpet4TUPX6uTpeHg
Zdtn/HGJKEbeHAjVIG22iA6mGBEn5TuYVRUo28HNVimVkYOEyy070k/thiyfpnvaUG3bq06C9HJP
928LA3d0KJg4IW7J+wDk/6uZSPm/un1YuaVxllBnUJRFBQvQyAbtH2lk+Dy66iIQikBbZAAiyZQ8
R+DtWB4NOqyYvOa0SkEX7etf/fAdxeJ/5jO3v+bFgshWaPFwQEn1oy4kylXmuRHhonex15fiTR9X
Z9Lhm2ugkzRtnhFPLmUpK4nr9RTvwdG5uRftb/hW1xKoturN2HHGdFUdfKPrsp6QfTy/W+K6S8wm
Ks5coutYmPoinH3mbFUMqqEk55iUFQOZ580i88fT17A1pjReowfGNPwG+EyK3FwiELjT/AV+9FEd
Ina/dUiNtJjspy4KNEd3lf/y74kZ8KisNOaEaB8NHschs1zMgVUWS6mX+i4wEBZIaVAfwisN4K2v
pndt3TJMms9AZF8fD+t2nI6hZc0Bjbp5UsGWKye7ZLUZu1CPyY+6nYNiCoMs+ttM8NC5U87JXtx/
oVEsHqOmg5bsGtNlY20w4XqxcikEprQIONt1Kd/KeysJFXBsW9eXqaG60lD3p+vBqKGc64AZr2VF
s+QNtpjr9KpR/AhKBYYfAVPvm6aUv0qg8AXp2A/SIBXQNThIiQhIcjKyz5S3XsslAFCmigW/awK1
Rh8xe+W63XGleYHG9pu6aR9ntRvrix9d2QvxGgcEfBjhEcN+/apNhGqQssc769jMBuBrtA1mwqSp
xLLLM+0oxjhbcppr1vSs+dvvjh39ge4haT0GZFhhEhZU3kSnBLiOXc/k0wG3pB0D3ifEGZId7nNo
f1RPavsYVWXRUDgK1XUbKrQHwSX8dVSDeYN8dCX8dDE0Wzxzgk6yIWzt0BO+l0uiFwhOomc0NrYj
zq6Y0wndMwpgnTySx+Ux3z5yF3RZZtBDUqRpb4UReeC9PvMD2SF3Qs/VMZLPAlOlGG9+e1+cPNG/
ivrGuP+D1U4eDYXu6t3j8QOOfwooB21sU8Fi9i/jT+CjsdqrEaNxoeU6rz3+/cPJpTWIh1VGXJFX
om8/0xMM0B/2KJqam/03KbPWyR6bCu7R4I2BQ/PU41qS52gUP2Bgpd56RA1Ehv5sCRT3gx7kdsdm
5FELEIB23Lm9KbEtDwXQBVFqe0s0VA733mA3WzXUrkkZsIVolW3NoeJIkPKtenOUzr4t0C/NG4YI
q0YmoTg51oBZ6/sc79h7XKJp2WKJGSZNOf8JvxoEf091JLjocYIufi62j06Tjnw64uHBukr0IkjI
4uSiRKg5t7FMM4FIZPQrJFoATobITa9fvwke8QVShOi5v5lnNpjs0a52C+UxEVfxqosef0qDftWc
9+oqBUelySOu4oaiL5kCoaWxjdnL9zp1pNTTlvxhve9GYwIKE0o/NQ2AgCIReyDeKY5HuFgIv2Oq
SB5a7Mvrg742+xK09mku5LNAOJND+BNDxTjX+FyM7U9P31HUsbkn+Ri/3/Xe075/DywaCduPIaQk
wZMJKla1FcYEEvaIiczgRkl9WbFvp1G3T9EfFliOxNdGylkVQ5K8LsUeWyqtMpB4bmN6qaqMbX3c
IaYAwyuU0kgqIWfILPhNkyIEfH7GlOs2Hj8QYLT8dSjqgiOiU0OxAz+MulVrNfG4xFvNxSmVn0bs
BlGKwrG6u1MtaFI7lZM5LhWVy15YpkvBz1UBzyZ8Lgp8NuxNn+UTXSljGst+Iy/hd/F5I9jle5Wz
D17xAuS4uQn/F/p80a/z42az9T2MZnS8kAWQkz/zP7sFnWn/6XKtOksmv1vmrXiqivj+CwXH7Rtx
7Je6iRFjq8MyngFSQhCAM0mu4186K1JXmcB8Zp+LsCCKGPVHFTdkB11INhEhPdVT7b+X3nb0IAu0
yM9YbU0zbkdhkwMnpx7+bhx2ZpFqlHizwpv2oK78yDKGV4vvCtkzhnc9dJwaS/aJYjqReI94CaQ0
iwNnSIKhSINWlwRbJSiA04JcnmWpD3WQKzp1L0iVuhJjR8x+3tLsm3Z/zRDl5AOGiKDg/zMFgQL1
YbihG6b549DxUxMkf5/bkPZN0obbN4BWUnqCH0AzclQpUzGThmOySrxWn6TS1nvmfZEACnz/SRc2
dMCQvz65949M2u3md3HqE1IB+tgP+R2iNNVLSFtc9bKZxT+mKJqvkyyo3VttyvC0zngprGAen5nm
5+POMNpXfYFSUeEOVmvByku5YiIm8QMchKN/G6WUtOx77/JOAXFgjePhdFjHzLWosnpeyhCHHMwP
jFj20gIDp6+6wYhc3TSCXxJ1UMfl8ttjmhSf5FdOSt1ORQa6usYSL/m8uFrFSl5wsIXmIpxIWT+b
3QEVmIYJyInhxcVvF6MfPmRvJE2Tkyz97Py0oYXWg3tW64/nWYsEdIN5AEb0XdLJxVi6oxa5bxjL
Q7oiOZWU3wUsL2R+wlGLVoCsoaJ8+rm5JiEiaVAooWLiP6qTfHh0uz1uXcrXIIkmshp2/yzPBvSs
aIqYLtys1i54wx99cdG4ckCZr/OfGBS1v4yo1Hk6j2GyUQX3CiWx44xHQ+aegqg3T+irYutzxKxX
B+ojUhbigsZ5co3G92O5duIPJiwdTAvfl6orFc2aOCtTgAr9zTf+tDMsI45Vd/usDyh9h/2emyWu
kVfgPrdPPK76LNtvYIO5XFpTH2NiWVkS+v6tcDrvqdXxZHSQGVTbzE7WwM2czQhP7kczPvRKBR9p
Ys9mAw7yoZFlmzHMYEPmJTTf7EOQwV0tbLZzu2xP0g9VT4fa7gUwEkET8yfaHwlmVnp6iz6z07TG
XtMtC27FJLVexnhW3aqyrmW9+6o65pmY8furnu3a4imcgzyJ4t9AxBq+olGT1qIPCrutUDPoC8Lp
U2TpNkP/FBpYzjvmXsG0ZBUvQkTRcBrNr0TtZIP3ry4vNVGevCTkbjDn5eddMse4+LF1wHrShIvl
HDhK0LWwRsKUJA3/c712u2HS9mCt8wUIdAKLjEaxb4zOW46GLs/lhM0PfxarF9xyOQZIPYr0aTv2
bCUsPxzuENgVgs5locWCj8CGtQEAKCso+6iv0+eyWq8uoI5Ip400VzsZjt2jtURtgvAK3k/ZPGwF
S5zROplp0O/ZqY03bUbO7x0AQFYr3AkDl6w/SfGYIWeTNUqo0wqgmxulU0Pm3llwSO4lvCc2/ymM
3tMTQsShipn1Huvqvc/Ebp7cXIkfpWbqhtChyujBNrUoulZGx2hCiiER0caPpChYQO3uH2gA29ZG
w8fyBbbfFNIW2ahVQIQ+I1eC4r++gDxH8gQUWVZOQot4NGWAu2PY6vfkVSpot2EkZBFPUZ1SSExg
2sJEgyFz22fSlYzhUA7RA131CCwz9szALdjwmHTPOCfd2KZFwmepy1Q/V901UIeuEQf8lcje2+Io
KUS1O4RHpU2hAcYe9TaM8kcQB4zSVHdyXfeVYo6kMjvyQg0gH8udTLdhvSUOAk3gx+2FRggWjyOY
/FraypatM7QT9c8z+M97vRYr8Wz7IhVrQTiC5WFexnRzYFoAaZzBopp8bkMbFGjWVXxcyBRp7kUd
AL2VCebWss93vd0e+P0CjsQRlS2hhPS9u7FV3cfUvFz/SJCyVeJuOhh2P5OL53vb1nKxqI+oV7ju
++bBsAY50p4Wf66xW5kyViztpf2oZKf0pWU1vOIAP4/lSAzM0nTr5gMhOOWYrhr91JaE6s+dOWUw
4CYQrnIhbR3N3vG/uKck74BiBYRSTdt7kfpy+bI9mvzeKf5HtnD8zS+iwk9c9Ty1TL4rw/4s+OC8
OkqIe5WN8jWMkjsppwaz3mu9sC3KjfRZLEhXlcQrl6dXGtU6gWowxYRNPuC+r7H+Y6sMfPadAR6X
liM/NSPOCn4orvcZbd+AtAyd9P1lAjNQMUTut905wbfpMtKbiA9HR2R8CeLvDiqblvtD/kZngDpf
qjbGxPYWohY3NGjzZZHG/OMqosBuCl9LOdsbH424q4Lg1ei+K6LYe5ArQKgfeC6p1FLaaiBO8lLO
wfTTYjXtuS645X0I8JdyI5WoLctJ3zlDW174HZNoXPnuKUU0JIlXCikEjegwwhrXI5PITLZkhWA6
3TZqXCd2i+eGys2KVZMcROsOkLxfaxtcJlvE2wIDT7cCiwJNCA/rb4tP+TEGZswuQPbfqR+Yu+0k
a/VVyEG4LJ1/cMT8g1fU4GEgL7Rxzfv/sreEQNQLFkk0SvWF4cXDTItozxyDLWy9enUxT8RQVGb0
oLb5uXI/B9GtBX6ZosL9zDXNc018SIiTElgIxso80MWWQSDH3T+gxHfHzEz4Gsz6a+woCVbvN04c
GDU/yEHaFXfuGvPDOHM3tX3Xl9FWHLenTiwL53wN7lb8jij1QyT0kt7uZajCZW6gOUWnMNHwCBd2
gE6fhY5mshnIFTbCOhFpEXUDxuyFWraOwZXh2Wke75AbpyVlEP5OUum78lm1YTrCJNWTOeATOz7A
Qm/pnnvDkqS8wIoORkGHd5bQau+ek4RlftSaWwv1MCzCwpR9C9KHZibHOByKDgkBg159zUntPZBT
21w0W+3WoT6Q9mq32tRFeqJFV3wJnRPEl1lvFPrhmWSZDuDjR0SOpzciITDnHqLQVINQc4KnemL2
8BFnqf60WMU10Pf9bL58qj9oyUHu+wCX3y5dYYGieicFSFchugtxskhuvZFKYRdoSDFQjUfVs1xk
l8h88Tws3sPRDnHoeHBHILrvNOcpbQVhHntf+mmPfPqMy0ipHGPjOv+mOWXdOlTnMcopLt9+nKjV
YhtteWK2KMrhVrTtcOfcKJ3V7Dp59sXNXwCPKlyw9rF0ImKa4Ig0SiMCcsdc1E4pgx1fjpNJrg6f
dLL8lv5LFB+J3hWE7jG0pW4tanqCkDrXujArkp2h8/PZkk7wfKEtQgvwtisHkcpdt8qmYs0N5SgR
J8vObcPc5AkWLfnpreo0bPPsyyPMLbouXX0qaOLmhIwWHRKx9ePyPLKWySggav8by3QQNIGNfggR
6IGXGKV6R5OOxs9rudZkhLSC6SF4q+1dFVIheBK8pbmDBBjLY02E3iHHKpwF7GDDnf5OCCt09YFf
5M6W7RYWJIvNKZIIS1SJ5OAImND+dQXtNNkvQ9JMlZFWbpMe4bbz5gqtA3Bm+1GrZkt0FHBOczeM
X4WW1qmWCbpcwzx5JAe812e4d3phS6/xzZnrsNcwMSIJKWp3rjxB3DYRjijnRFwoi/cD2P6fN/fb
i1A4awg09e/w4gH+nCgjsJ45TvriMYfV3jC5pJ46oOREpBpxjusTSQiLTGCw1wNlG3Y0klEyAiDd
OtjcOuBXjdsYAZ6OKDRStKnutdBT8ZNv1AIkIK8PYnViVrHv9Uo3ck1Qc4vmM7I3cUblCXzA0mXA
2YX9sNIOq3wqjPjPcAj2Ko71tFJs7fwktE139xK8yXhSg39YLuPXStIizGub+1plsVTMbrXKQ0xx
qrAqMOqUflxC089iFCytZwz7TAZ4vuwxFJ38kyVkYIzkA5oq5TkYWN7Na9UU0CuG5pV3VgNKNgXj
3K6jjTguoAraFZmSX+CSVFdRMfIgQnW6L0O3mMFbtFRl/VDfC/KbqUp039efJZ1HMxsL/tf4NTwP
bqewcsyejmWnjMnFn2MBVjCkcIegKOIfSqZ8jwrmnrZ6mn0Jwk6sPq28z+yHepZBwT3ilW4Zk9xp
ViTXBpk9fVmJ3jJ4wJc8zH+a2J3RfqmNN/xoH3x5BCecn6LDP9KXhrTy7zJH1e0udh24Mudx5ttf
CP0hgIPvvl3L1O2Ew0ufcxjZaCKioxb689owEdJCUJ8Z5KonZg2LRv3RdnzjMBkwpDMfxItNVtd8
q4vZlvAfvi4IMNwAi05vZW8UNVfVMXmKqT4cbVrNBGeZnbkqGGhNNm6pLLcyHvZcHPEBNCQo+ijk
KpsXxN/XooJR2bscaltiCBxNTStT9BiDUqrCo9uRlivV2FdBeL2D6Kwwyg1p2hXimkPFup1cwKpd
R1ez8gCXkCagMit3o1t9g/nBTBzWTe/jrZ9RwnB05sY05MlC7gxqbdU3PFRqRk5N6pavJUYLSko/
T9AGmrKVC95735mgi1xAs4zyIHeKhnt7hc0IAe8tnBK5Mu54BKZwmbm4BiBoX/dSHJTj4ithOj9N
4JkHot8LULkZoJAUXjkgeDXUiOnSvjWcIS2EdTNVFEYt95GWJOAQB3QShw3PniVHVdmHlpFG4Wl2
zunRfZR/jZSXoYjCo34+wjuDEwjdISGHbqbeh0IpLPDYHbz7MyJ2zk6H+XYRlY5bLuE1gtamnFEZ
FlkDdBEWBdqPS954DsqZtcNXtbox3KHmgAfgJUD8DITcmjjt4JeEZLgcZuS7Gxv8n31ZS5DnBBDk
Pf1iNmrEAaTCGeRudSCbqY9pGFHNOM5s3xdzrsbgFA2rE1Xz4nudxaC2GlgeREDxmWTm4h5bW4Vm
mn8ZN3bbiCXMvw3Fp6VoSGxJYmEga0PjlG8xjhtqlSskKsmJdDhnqXZZSPbdhwlXeBKvtq4D3pY/
JS4FoPQ7pUAPdr1OsXMr4/MHGibkTFCdi/r9JdYxECVUUiEHEuHNiIJhY/TERvmbg9LYoi2fQL2Y
jsw2rk9zz+LQ5OC8URa/ArlexPQjX2epheLOQCPV39VdZYhKtnLvX5U88ZiQcU9g55cnY+/B2Mli
KQ36YH/bfjqEaUrbJS2SPFfALXiAdOAA1J7usxINUWQw4az1UxcCBt8DPJ1aMhmHvFyEm2D0q2VJ
2RWm4kKw52zwQGc5GXcsf2AxsENgoetoKL6jHyxvO1aCZffjD2z+pK9lW9Mtb73XXlYCVDYezYZm
d8KlDLHetDC1bmK1s8eAAo81fbUkbCsmnNrGpRPciueQuE2K0TrkkxMkQmsLrhVapQDZQz+ONob2
3ODSEG4MwyMJ4bTTMR8TtZnfk+O7D+jkT4gzTC2zevpUOj21M73jqUr+I1ZAmQgbQ6ugjebPVhRF
FE31q2K4jIRE+16+vmdvcliLhNoUSFsSTgEFlO4a1mNNtiKi6I2dPO7UvXkWUnP8jMo7H6Pn8AHj
l3grsmWiRy2+bV6++ANmkkDP1znzWx63fza7DOMcTgz3Pzzg6eLxi5lZ5S4hfGM5bmrG7/vwt1Eh
fZUht03YC2QM/VH+3Tn2TbE+p0oepjjombUzNq7GN+70n97cp8cJR4Estc7uv0dKHI0pfVKJGTBf
+lOT5rkK6AJSTxGBflbqPeUo+Td3WMKEl7rYeiaeonttJ2DVBVg/SRSCwkkNrXLPoMKyNXc1Mvcv
GdZbovjKrGVzd9ZB/IeKJlm4hNTCPuHELKs6PJpCbOhwEc9KNmIdZQfb3Yky3qy3z7t8YSGhzBHk
RFsjBmJ5BfgZCmy5rvfG+tZvhg8ArPHB3QE0RFIxzFfRrrgjmiawKSgGe2fR1NPx8bjm6RrhB5tl
YeBXRavAlizdiCyTyXSpiUTVVX2hOeym2xvfgyCusXt/MRZ2xLsJFYaFY8xkBn9Bfm8xEKcFMP7j
mE0mml2EfDBSOWy/b2bPKoVdEqr0t8oc+v0h5SBg7OaB1BMhZmhA9QzkfTvpbI3XSaZcWh+0qChY
eqg8AajWDs1o3JXcIZkV9xwM3aXmPXn0Vg06u35j4jzaDpTDxmAAeWAPEihhHnfcNYqZpS589cJi
2Njlbeav+JCEDg7qdv+WuaGkEPcyZE3D/QZJO4e40GNXXjBdztc4K23xxaunTjfnBCyS7L6XKQ/+
JooI9OJzJC3FvW6U2eX7EtAuQ3gr1NQyvarcuj8BshXQ9TrvIi5BkvSdRAjdTbpSLFQMy/s/HvzR
M7J+QCFqyzjpW7H4dKoZPoH+yS+FHlOaWocd6IlSOmykdWRpdf70keuraJW6dNW1SXxpdgYzN4o4
Aey2h3aiPDFW+N/1z3dGmnP2B/Wj3vsSOdpcpPy6+S3kTMpZ+mHLdwOWJldTVkxMdG/s+lV22MHL
2a1Cg7/WPgwP8xJejUrOdLviuFjvkfXfPfwGcAOuN2VpYu3Za5wwuDdE2jeKlNxhOYMwWdX2SInX
2uiPbtoAo7OhCs7mc/m/cGrwjcZNtGVuix62FTmoFoOkH7k0mHwxaOGbACK5aGZcodflv1kN2lAR
L3m5amNn+5zCQHJ+qruo1lWLLkVBWjspK0YXwPqU8qhNWTNJD0uvdkcvDSZ+ZAHUgnYZUZZckXU8
fIJj+BL48kUjnU3CWeyyYjwcIinFcMLodJsbQH7ayw84mCz/72L22nteP2Blzz3kw2iMiYIMVTMj
X+zlx+Qo0vRAlwmNs3+H5fe7u81SBVWSD1X+B7K/RlCo7gW053Ixc9ROTQ20BccJZVEoUMdB7ZNs
YQYh75P3aBSKQ+vqGTXeYAaEl8nFuKBuG6ZWfKrcxtvkzy2rlrSpvrK0AcV/swAt5Ls2iGfVvgyX
CK0EYYd2DdgE0lU7TCe+eCOobO0P8bUu3KD2fgKGazCXKOZ28vSR24JRgIQMzSa9MECQ6Vc2Ukjm
hNrhufwSNE4J0/KSrcxOzwCiwEBcf5KOaPrjtgDpyMQJLinFNak1aJ8ta9U9PXUgrqRK8ppFAh4m
IxABjks6tejn+rnEMmg0rP9o7VknZEXgJMKs4shAoD+phGQKVqs+LrT8FlLJbzT27SViLrsbNdLE
et4gAY/dbpRVT9dZLR1YnHq/pQAqaC+o9IF+Rg0JRM0IzksL1+KwlPq6WUSCK+AlTldNprC0/dIC
PBqronGwBRSzHXDauXF12W/7LEzefqsy2qPvtDW1tcNMgkGGHj3XtAKWJ/WHzb9rczJ3JHMWylMH
4CpnH+X8ssvK2LkdIHU6VDhBXKzAmAP0s7MElYa59YNjZFNrSc6DvXoOTlO/h+Ln+XyUVBU5jEsQ
Foz8e+wcvMuncQDokemtdVv5xLSNUfJ8oN2xWIe0ayUpfTkBs+NaGKflAsVpf91IkLt4vVJa8JW9
esj+udZMuzbAazot7hkH2iygA1kxdzM8uibgCZtGDHGTWbyN6XzZe5FjC17JoHxsszDaEFsvU1AY
dc5OBNErNq24lIQSFvXLF9NEu8HgAi1BMzDowe+aDCQWniBCysnFsBX5x1LCO7tu/ryJjKrD15z2
JyEfjCX/Tjy3VMaEz9atItXmoTXNyA70BsEf51WDKExNJzl0N2uVhWueV3YtI5hCq5nkjfl8s1Kt
kcHJpUX2Lf36M4TUtLYY8HaouS2JhEWSunuUrIy0kU3QkfFOkiNnSiOLf5w/dqp4emAhj65UcMSB
1gJsi1FLfYjQC63VbeXyUDfziKTOp6BrCTWZJMKZcFSfGu96csGTJ7R7sJfJtR1YTZ14ByBaV8aH
Q4TXf8gr/DlMt7MzakT/ZjnQW+VY/v3f4HFzZuRhMZrxGXC9lVGHwh1G+sT4dcFwAuRtkQbgiJnq
Dnn89qu7AZzk9q8mNGY88jN1AwS58rl/nn76bVu/GkLAZEQfq1keld5qBFkTfDI2KOKsz4E92o8Y
N9bQFeDByeA6sTMQMhMVgf6tWtonVxFvVR+pymyTZrkSGO7SBzjlh3/TLMXX3R8aR83M91Ye8SNe
0IGnc4eeYIfsP8RHaBFlbh/Ikp6fJRsJeHrQB9qqUFcVvx5Z9RohsK9Do1eddws1aRONmsF3J2y0
iz3AdahimK7eZxVFEPtPoErh9aRpfoL0fOslS447hYoMPOy3mVR6DVANFOD6iE/kaAETGOA1fk7h
IQaShMVQiLHizEbH3HCxh3NwByRkzM/0ZK2Yl1Bdt0Cc4ago8JeOR16NZjft6z5SqnBI7bE0uDZd
ZXtzKf7J6Ezd4HvOHWfZVxfI3kUBOfeNk+f11YwQHpk2Mmv5C23aNw6BcKd+YLfimitpWTljXLNG
IEh/yUePwTUDNvRUlJklmPYMLzuYxhgGzo7sOjTSaH2dWTBoXYxI7fMI5ZuC08PmXknIuV7wqDTL
dSmaDXDh67IILwSpcOWFudWyFKGhFggbFPH7dE1ORAC4/8vcELLOS5Jv9QM7p4AWNT9A/Iu7OZFv
MUgSp8ilqI4olm74b41GNbnaksQQoAnnEy4KiiCJ9A35QkL+L5r4OSMAgBAqQUF74vyFCyXgGt/K
uygf5SCYUiHD8U0hR8bddi0n+E3gJDkEWEyD3B4z5AMocyAHfnEFRWpeaCOnwNkbNlitPTjKGjRV
ubkazodPMY3EJUZy6P1YqKtMhDJbaabVR57rrQs/g1RYWurgtqXQgnURflCrd07zbnsrpPprvfr8
M6vTBerhjpKqaHvf8ri9fr+KwcK2oOTNk7u87/uSZ51w6DiwBxMcFNvy3ECuWBOIc67Zc4lp1URQ
Yqq4NdBM6tFlXtk2lN18QMOhrIYVLwyCHn/8yZH1UOBlbq73J7m8UVd06N1IeiuuZ/Q6IsjSspNQ
RZlxjIJoUEQe8Ss+s2fI42HKfAPoNR+MjWZpxJ+2X4HIWZA/GeWEl/4IuFTUEskAmHKKAr2Sy2D1
YDbMeXLJHf+C3lUItMX/a5p2bMrrOvt/JPbKdBHwaz0zkW+slKiIhlfqPGHDN5M+wrji2Zngx3q0
SqcYiJlkQhZ2siTIgxo3CXtstD0aFxrQFxOByXi4OUVetaWIhezChYmEr9MTxet/vb1JvDHsX2/D
/U5EEp5aQJ7ECu3CfPP6eaa0Ysk2BNP0Bm9j/olQzhTCWUwfRoeVpxP+JjLOid7bVeLSOIPW6uN8
Dc54Tz4CMhJPRhZR66/VGaYUSifXkkS4UQEVG3iqBWXl3cm9AMRmMNDwS1cmeQwiCJZoW8RRRWPO
KDNE2M5aYhl6Sxj8JfsIxyyD7nv8VK87ppFF24uEZhvODSZFjMUYY4ri8JVkeGof27FqMiKU6ZlJ
qEamfkngiolUGa9JLNNT2/idH1zDYNOoZ4YBzb+51HeipJKfNKBdSOmAkky05XN4RAACVC0swotu
p9nRXP3JR51eq4d41Hr/WcgkeipDNjgDGiO0CY2QvKIzgsB9UtMZ6eeI98/Yu70CEUpMwGD6NC7y
7dODwUO+z2FL7TRwHkyqX4vN5JCkjs3mlLkkTDNDnVEo2HO0681+3GapTrjJnv7BrGN5PiYgJsVp
9i8BoF+bmcvU1T4foMdjYR9Mppl3RPWnv9m0eucBQPwxX7URzYFP1PNI4RUXtyX6jl5CsPGxC922
VTHYguBqzhvvGsykpP4fJP/5x6M3UG/FySNI439OihWHySubnNvrOWWpOkmDe195XjyoYhmK6ucr
DcvmfwOv4G19zwiD4LxxF+V1e/4PLhf3gARglx/a9WEHa1r9XvGh0QB3yo/nCEzkpRDKkxoqO7vf
OwmZ+cOZGcJGeLQ0fGbEiexJfVsLyQPQjPz2+Ac1TbHAafHGnqSCPrP+ogYd3dq9gSBbWYb2FVm8
zWdv0D9lnEYxuAh2Z7sqcD6MiutuQsRORQuG1ng/gmB/BEiJ5zD7/9ikiCzqaRuP419TspZ3VbMe
m87CHz3CeZ10+sXqJlaKd9TWcJANhAOGSZb3dt/9jzw/efq1Gf1QmQPrVZ+0G1gtw2IIsKCJDDGU
6vNgLlR3drganTH+xLhQV2pJlKkdiu6rrW+uZAlixomqIYwJYn+8aqu+xktDoiCiFrOfCbq+JR4I
m/LofmjL+P4VRa5uj5vZj1lFDpTXnMGTdGlsvl14DSmb/22TylvmlSJdHi5Y7zSniGi2pW0LBzKT
dZEtbGhg022fc00WzyQOLp81ZYZ0LZAy9XUe+G8LIWJPxNxYUpBpwoFToTviRB02FGr8NBl1/EWl
/B06X1UEuofp1olnBiYCcpHO9qlrrzIVvwXjAil9dNCZwwkVKgzcn9FNL5onmbKKOs0w4ZITAMne
HDYdb8zhnMM5m4JB+ldN5GuDMLanTA1DZaifZU4u1yTAZjn2eNvCADPLusEZEXN6CGUftOOL2oip
KrQAhQJ/p0dfJPCQfqUAsoRolZfO70NDB9ZdcdF9zxWXPf9A5fEYhUv/upoSnk/vlGRNLPvDtkxW
f58FXggSSLpcasxILYlrWaMjexEfryt0H4FflJvmOHyMIVqNYxto3K1UFitXE4b+EoILan/3o64Z
12+bu1wXAdaTKYXpwZs6jN84hpWFHu59MCZJmdunfKes22qgcVlXR2SrOHVCKLq6oe4tQLtsozfl
I/qlhz4Q9TgRIx2s1tt3C0WTdcwgpx/mqY2W8fS8Ha9HfGAybxxK2Cv4wnZf8OJilMVI12S7gYIj
/4Zh9CkdvrlITYWeVlFcYuAfOGl97AvKFiqvcDwa848LIw3N5TOmF6AL2f3h4qcxvvLO7EbDpWBN
W+HGIv6DW6Y5WGPMQTwDBUqQjCfshN5E2xrACERzD2RJ5FaVXf2kdlQW9N+CHdWwLrZSSo3a/HQF
v8KbOwzxs6Z4A3HgjILXH5+EpVX8vvjtZCNvva0tX5DhFmP0nzacbujHwdBfRZG+ibgqtaXB64Lp
84+it0nrHLMdxCwFRBz7LUT54XdwggZ1yq6UYtP1Oy8SX5UntpkkS4r6boCULl+sCNNl0fzUemOs
HMFCX2YrJxtKTcmKiIN9HzWDDWO/xANQE170h7MsXA8XrRyMlTuACpNDJLjU0GyxEHm1btNPz65Z
18sVXlACCFecPQ42ysbJFPcM1Td5FhGymfYSG7kffrDxC0z8pJObUJI67ZN8BDHJPhfIhfKfrO+T
EDXFxLv/v7UG2p8aq9NRuhjzlw9NCRqB3GYGXl/IRbmXkRLTzvj+C4wqOQ3UtfCjOqqB7NIyaO8s
iPkBvljvqSvK+gZSvoNi45wkQaDP77INKeLy5KAYeSPgOgcJv7HVKJ3Ev1yA26wYG7/6az5jH+/5
p9MmnM8jhpT5enZPEF0d3UjwpQ7eJMrSy1OdrVQiS/IFl+OHfDAmNhTpWFNXLJT/1H5fQMO67GvF
UP0bE1Rs9wgHh/cukpevkhVU/wc2rMbqEeeev+JnT3Ls9CvLpOoUP/dGFx+g7ehkRbjvR4fcgY8N
OU/iTkkumdzWmLe1x5QUEpbzKdWf7Dgc0hjrvg/CkDiqbpL572AB29nDLym9f0GqDjsg2soyUGsw
Qwv5fV5QiHPcBUTcdeYxq6/vZRYpqpU8/nN8jnTFF3eCEqdD1v7n2TwDBHEkS59ZiEDINpDtYsKX
fokTDmf/k7XfIE3ZPOraXM/fTCsHSMNc4v0gos0pln1I0OdBsWriCWj3eqokALsYveDJ7jR0qjQk
/yumYoYj/qYi+TOfLPT35HOEoz3wHwCk2Z8MasfxEWJ5SnGkKy5RK+gZRDUj5E9WkHFx055sLQwa
oLaM+buT8M48lFkkTbzXNUGlLxlDkhAzTQMPN77taoP93e4EK4ZNKjzMh7y6C6uG1HLjXWax2OP8
YwzRCIzmDswbaSdrwOK5pp7N/bqGNarduMgpfcS9gzJ8JtvQV1eubaJsnfpawHK8I5YvilASNhv/
8Zns74sKoNZ8FU3E4SXU2zCqu1+i59kL2nxPqJKfbusbRQEVe15X1opYSU8NylqvbPjeTj+yfcxC
XMlf+vUn4Dc1ee65FYi3Um+P7hNqOKsfNlZLQOAFw5Ceb2fvPgmKfpLEOrbGun/X8aFGyh833xJ1
o/rp6Hm4m+B4bFs7vax7Xqmc1Zmo/Mc7LXk8EhtSPocxDPx/CDmgDfe1C/NCnlorYPAxwsUzSfCZ
Y3/6zUDBksCTH8SH6O9T5uJNrkGqHXags3PZu5/qUmlBkTef7invX7AsSPGAsdXDT0rhxXTqPGNv
NYXH3btyTonV/kqtJwUi5RhSChSKaHdMyNqVg5uX5NbNTqyR9/ljmMR8QxcrFcOBwReiM6Rij1K+
jMd1KtRNNMnhKlUs0RRhG8lpQ3pANf7jG2NeKTMs547JRWmO68wlCaIosGZCjqKMLxT+zRYtcw+b
fyUJqSLQXWE++ol6FjAuYT50lPnLFb3za37O9K3oJFvKQiV4YW1nuouLQSEJhElWnR8XhvIBeats
yaYBXJi0oeo+0y49VgPhXuWrYK+CcN/MJHrAZK3R8/S/Xc4l8FvQ3sPLxvtOQWwFoHvGB9ruUH9d
voO3gDs2yXwqjec2jtrQL2WU/ROkhO5sjU0CuKMKrE8oeTQAwjXE3tHS7RWVycKbrD2fdO1JfYV9
YBsEBQrb3hxyP6v0OX7F0Lu8BmF5csCYWZmpqo5zf0phc9LtaqrR8FNDmQKaxydXxn2r+DQ1/Ni7
vEiPoliSmRzt3sWxh1wysrAmdY8VrsIoDIOY8WS7ngqlKZh0WTe4DcLkP0kjbl6Ave1C32EmGEqC
4Yj9B+5pNeLtcsAPfGroUbvqiVweWoI7N8Uh60tESljtBa/7WX9bOMjcW3LYn7LG3pjJaFDc/VrT
/Wl/g5n/Jxpom9Tj6G1OTuMB/6cVWd7BSYKJpl3sL/lsMfoDIgZcHKscH304/S7u0tI4XPV2Zycq
p4Wc9t0iyFmpGewrAC8gd0dvWeW8HlJQu1KABzZCmd7aS9zsLR/JhRGcffqLnCfnGA8Wl23BTNFb
rau2j60SPlLh6h/WmfzGrTU6otW0b1hEUzIeLksr3bMoy8Vbsxmwi/jXjizMR1W2FFgikb2FxQeE
sV4+j37U+NGNzTiBxo+t4w2SLxti9jKx+r+PIP2WNuUqTw1aTy8qPTmZpf3DrFN2/04BmoYvbyaq
ZsjAmA/Qo7gXL1RQOE+16ydWnryhtIkpV/AIsaoKGSJc3+NDcY1DAsTWdNJnmw6RTP8CYL5f6/db
lzghubHusPy89jSIzZJj8JHKSX84P5rvJYnb46BsB/CEMLEELPxgKaFRH7z7paQ8Y6YD/0kksLZ1
mCEg5tlKU6xwVqGFOrnYtHSEVVMGYXFn3FtwXW3ZxhAfZA7FwtpCzGdMWGkI6AQWnAXlpAgP9TJE
zrqthQRp5g3fGf3iQqn+up9L8cCisudyo3q49iAEKfHsPgoP26Z5UCad4VLAN0xf1wXJvi3syCQj
7jhrlXa5Zf5LgILidMwakxAlyv55dMRhIqy2fLyLSNcBu99sqt1EdOu/CYXxFlI0pdAQvA6dxM0q
BlQm07OU1E8YIoGw4S5Y/3W4JmiHUurqKfa1rdENUsz/oJ2qUsXuJJxD1weskuGcz9XA7emG/auP
kWPouBfsL3qW/wj8ZQ99sNmfSX06noP2Fo+LoJ8atGTeCFMpgAYD1cPiro3ELjfS6CUnmaTYaeSi
HJJubMM9agugUnM2ra26t7waRob0ngF5ny3UVhc1aTZL7BDIrkzejibgp8G2v6mbzilngCpzjGNK
B1GzzDU/uBgHeqkBuRI6vn14O6gtqekxkQY1Ik8FUwBqeG5Rd5sMFOCVChkQdjBaRCFI6ijdTvB5
plUW6L/Jpi0NyWg2L6ZJzPElHvPG4foVHGZNUZQqtJYj0QGXH3+5BDYAWTTRcbz1cVZ7oE1lh0Ze
qDMz0rrGNspgaBYYejOZvfMUlRtjOsYT2IuPLukuLIx6iLPHL/F0pjbzo+PVxpilqE102/nXC9g4
9aQqh9t5L1xg1KwjBpLosIiwnfW7tLYW6R5lY8l8egweP0Jb022HSxiFWhtX4YWNWLqdfu7pYaWB
Y9OQJceSJrlDr4GTHl+ZcF0sAkmKU5Z7CHjikcr4Ai8IpfDpymLwgW6MTkRKm29/4vTURdkyi0u4
NfRhencaij5ZC7h2g9XvXl9NL46atE38EOsfnAfj/VqZwTt/UWdyj9Z1usADIuqEhIZUaCAJmUpL
qqVC+EJUFHMsx8cYCzAbkCtFX8xSZYShDU8SWJgQMB/C7NmYQ2P3Q6J7qbRSFN8wMpKLFsRaT7nn
MCAd4fYIADsw1Gp0M6O1+oaoGsK1HovFvP456w28bGEUGqgbxknxU2vckqaY0WyLeuXVo1jLkth5
EK9teB1WMqSAUs4/S/8t6oEE323UhpfniZGFMFua6VEIk4r9DW0rZPPMIod8Zo6wIe6OwCJyydoL
BfS2MOyMXCfcPWd7UI9faLHFOyxNchzTuNaNIWvUd/fZs2Z3FTRajxdBcOyQ7knG+zbM3dGsVd0+
AWllKnu46dYk+7s4D+JK4VZwbs/pz1FxpDof65bwjVrBjPpHNJ3cKYFiXP/rY1m25oHRskRkWp/k
oTk2nYnArQxqftDN5stqpKzItFoDAl2mdELt/3jvm66LMhq5T4obQZc+Sai+8DbwvZ94AaHeNr4w
fTit68PMnh5G5PpR76/nlHJENBiM0ukTDwcEQqVm9o0QTV3+uTqnxbXmri2OWKVLVfH3BDIr0VTX
UMrwfIl4UtxPKNi/STpsLbLWq2G6cnTH2szKtyLqtLciGe4lRr6iSSLt7ixZiJtxtOyU/ssHWEWC
RKHlg2IFBiGIIJXg3Y9l7ctaN/GfSowpjS3dbMKuHSsxMTLWiE6S5c78qCgJcW/nShxHIiNS/lH0
7FUkWU63TI4K6dlTKUTyN0Ivje/51Heyw/BAWWRz8Ir/bSFmQR4+5tVjvExFApOmj0rVUrmEXWnP
Opo5UtreHa8dl+No7D8Q3AnLiK9DFrrmXzri8Bjvh0Y3NOAxu9UVZVmqj/ljVIfCYt19vr1fOgbp
kYfoW8LrgUOEVlO5DScWiOrVaUUYirBzVeOdwhWBRra1ac0R3UND/bh5/us/NI2cuxLWDI0ZkOFG
hSTYfvOMJPtkPIj6Eq5d7xuPJQT5mCiBQuSiOpQahIck+P60N8X+Tiv9ckN4g9HJE/6ZmTKXU2hE
cXYtpB4VhKaQOXJGOwoPds2x7ee+ulBEGEEnxuukuVVBP3wO3HaP66U67LjJ7CCBuUdm2wv2S1DN
LreygQU76DfkRvzSr9TdwEyoCoIWoRSkBYd0NYJ7KLSrVIUEM3eX5yz4c+XAdpIEcefGJrpBOOml
6QV6c66o/yA9YyX0/Lg37IMF1QuilGQsbjjMyVOeKz0k8mn6Vpyz8TyGhEKKqgnHH0JhxXE17B43
oOtKxKEKkJhyWw7UTPJJkeMTwyrHKgKNXhycKHnAShmIbbj1wODoEV6eOIFKTEZgshz+WmyLX21M
Dwv2wE3tbqsOjld1X7jT2PaGqt073/c3bIjJynrStkCTclgP+LVqRYRwzlVK54WbCQr7k0LbEi4z
qmyy6gIKjK55EchU+Wdyy1Grj4Ab+0Dd43ZUlGmtyuOmir0Hy5+ZIoBdOcG/8m3rhWuZoTkZNHq2
UAuHcW9tahxqdU6QicrrQrhd96i4L1rtyNVyeJT7qP/wMulQewrF1Rbm/ujw2siumfc4zjF2h6Hc
W0p0VIY92qZ8iT0DTYjiZhHVMlKppD9+mkKTTj3BMdgeRK8GT+9UmRsdzeSUTjnffTjcvJBCgcpv
b2pnls5pmS6YOR8U3tU4ura2jrOCtm3WAFEGgnPO9I2UdbgQpcRSqnIJq8F2Pj4R6wcbjQ+HaagK
t6W8YtrITMLf9lyvQTkKOCvlr83SOOcwIxXJ/+yr4EMy6Cc+p+85egsG+KpRhNuKB7Uq4fx3ZUSR
+fxYDoC96KaO+i/O72rWpMT7iPsW7DYD3D7hCbdz4kUdmmntwk2vqMCj5nA3KTnRF0pde0KCmas2
U0eMB9wX3LqVjJixBxfbYaHInmSD6aMwq09anNUrEFjUFyDRXw+O6hlMran/8NXP7T2QikPt6GFP
hCYStGC7kKtLmB3ETycIal172sJdqmk6kHG0vmH8X7aJ6J+ArPXdGXTjDnp7/YiN7cIauf2MmX6n
7hIsMmM/URZxhvlnYYKZ5FnZU+D8Hk0V09XB3U8H824CxKwH1Hu/OZC/NkFQzATsbbGeolWVBzaX
rriJvFiRstwbKPIxNDxr6wZ3EJAvgS1+j59EbbUVrzVLV+cyCPJruJJZ9eAbMTcsi3fsKOPRC2oe
ZJ0aK9yFXT8AU5A/Xz1WW4k1QBkHKV/K0yxVhHpwWGEYk7CGX3ujGZHlAu8mZBgbJdLVrHpRHuA6
zri+/pKwRf1lwtMvECweOEqnWHXk4jgzBdJgP2LzZFyfjm8yZE74ERcttCvHsdCpi6S7YWreZmmQ
YlgfTmMPiTEQdio6uqxfXPGVWLA77DKgHIfkFxW31mEuCQmLHJUD4LHdOc1EzowH9qWmjCGQxkh5
CjFZl9vfilYgjkvr+OG5TMVjBGjdXax1+pVH6lMP2xN6Q5JDFEIy3lUfS1LfE5q22JcQOtI7ECxS
ZHvxVMy0INWai74Du0cPfP1F/7bOkm2PC+JXMkSK/lcBgGbm29ywlW1mzfW6WbSekIHLmJg9kyYY
pMkjHmp+KohYU55M1rm7RKqQgHGiYobTlj4bJJuJjF1zTq5iOOwMhVac+W6+Sar/rk+z2eDfzx79
q9FoEKL5ua1Dr24L9lyYnIr6AlCsOADlv5wqxJni12fLTGFcTQkEn73jQCO0Oaj2NVWftfQ3i+fh
Ewv0q2OhF1kEXLyW4Gk/QE8xWfNnYsSI6e5WsUdwiR/R518ZETpAZAjBgmkhALnFjNJDgtQfgCJq
X/PT2hj8NZO6vP7WDHlxvk67L9DZMN5i6YChUDG7HpUPlUek+ayX/W6yPIE=
`protect end_protected
